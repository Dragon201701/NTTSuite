
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.v 
module mgc_rem(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_b-1:0] z;  
   reg  [width_b-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  rem_s(a,b,z);
	else
          rem_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> ../td_ccore_solutions/modulo_7c916ad59326b02df02b1a80099f3e2761bb_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Mon Aug  2 16:56:58 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    modulo_core
// ------------------------------------------------------------------


module modulo_core (
  base_rsc_dat, m_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [63:0] base_rsc_dat;
  input [63:0] m_rsc_dat;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [63:0] base_rsci_idat;
  wire [63:0] m_rsci_idat;
  reg [63:0] return_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire [64:0] rem_12_cmp_z;
  wire [64:0] rem_12_cmp_1_z;
  wire [64:0] rem_12_cmp_2_z;
  wire [64:0] rem_12_cmp_3_z;
  wire [64:0] rem_12_cmp_4_z;
  wire [64:0] rem_12_cmp_5_z;
  wire [64:0] rem_12_cmp_6_z;
  wire [64:0] rem_12_cmp_7_z;
  wire [64:0] rem_12_cmp_8_z;
  wire [64:0] rem_12_cmp_9_z;
  wire [64:0] rem_12_cmp_10_z;
  wire [64:0] rem_12_cmp_11_z;
  reg [63:0] rem_12_cmp_b_63_0;
  reg [63:0] rem_12_cmp_1_b_63_0;
  reg [63:0] rem_12_cmp_2_b_63_0;
  reg [63:0] rem_12_cmp_3_b_63_0;
  reg [63:0] rem_12_cmp_4_b_63_0;
  reg [63:0] rem_12_cmp_5_b_63_0;
  reg [63:0] rem_12_cmp_6_b_63_0;
  reg [63:0] rem_12_cmp_7_b_63_0;
  reg [63:0] rem_12_cmp_8_b_63_0;
  reg [63:0] rem_12_cmp_9_b_63_0;
  reg [63:0] rem_12_cmp_10_b_63_0;
  reg [63:0] rem_12_cmp_11_b_63_0;
  reg [63:0] rem_12_cmp_a_63_0;
  reg [63:0] rem_12_cmp_1_a_63_0;
  reg [63:0] rem_12_cmp_2_a_63_0;
  reg [63:0] rem_12_cmp_3_a_63_0;
  reg [63:0] rem_12_cmp_4_a_63_0;
  reg [63:0] rem_12_cmp_5_a_63_0;
  reg [63:0] rem_12_cmp_6_a_63_0;
  reg [63:0] rem_12_cmp_7_a_63_0;
  reg [63:0] rem_12_cmp_8_a_63_0;
  reg [63:0] rem_12_cmp_9_a_63_0;
  reg [63:0] rem_12_cmp_10_a_63_0;
  reg [63:0] rem_12_cmp_11_a_63_0;
  wire [1:0] COMP_LOOP_acc_tmp;
  wire [2:0] nl_COMP_LOOP_acc_tmp;
  wire [3:0] COMP_LOOP_acc_1_tmp;
  wire [4:0] nl_COMP_LOOP_acc_1_tmp;
  wire and_dcpl_1;
  wire and_dcpl_2;
  wire and_dcpl_3;
  wire and_dcpl_4;
  wire and_dcpl_6;
  wire and_dcpl_8;
  wire and_dcpl_9;
  wire and_dcpl_11;
  wire and_dcpl_13;
  wire and_dcpl_18;
  wire and_dcpl_23;
  wire and_dcpl_28;
  wire and_dcpl_29;
  wire and_dcpl_30;
  wire and_dcpl_31;
  wire and_dcpl_33;
  wire and_dcpl_35;
  wire and_dcpl_36;
  wire and_dcpl_38;
  wire and_dcpl_40;
  wire and_dcpl_45;
  wire and_dcpl_50;
  wire and_dcpl_55;
  wire and_dcpl_56;
  wire and_dcpl_57;
  wire and_dcpl_58;
  wire and_dcpl_60;
  wire and_dcpl_62;
  wire and_dcpl_63;
  wire and_dcpl_65;
  wire and_dcpl_67;
  wire and_dcpl_72;
  wire and_dcpl_77;
  wire and_dcpl_82;
  wire and_dcpl_83;
  wire and_dcpl_84;
  wire and_dcpl_85;
  wire and_dcpl_87;
  wire and_dcpl_89;
  wire and_dcpl_90;
  wire and_dcpl_92;
  wire and_dcpl_94;
  wire and_dcpl_99;
  wire and_dcpl_104;
  wire and_dcpl_109;
  wire and_dcpl_110;
  wire and_dcpl_111;
  wire and_dcpl_112;
  wire and_dcpl_114;
  wire and_dcpl_115;
  wire and_dcpl_117;
  wire and_dcpl_119;
  wire and_dcpl_121;
  wire and_dcpl_126;
  wire and_dcpl_129;
  wire and_dcpl_136;
  wire and_dcpl_137;
  wire and_dcpl_138;
  wire and_dcpl_139;
  wire and_dcpl_141;
  wire and_dcpl_143;
  wire and_dcpl_144;
  wire and_dcpl_146;
  wire and_dcpl_148;
  wire and_dcpl_153;
  wire and_dcpl_158;
  wire and_dcpl_163;
  wire and_dcpl_164;
  wire and_dcpl_165;
  wire and_dcpl_166;
  wire and_dcpl_168;
  wire and_dcpl_170;
  wire and_dcpl_171;
  wire and_dcpl_173;
  wire and_dcpl_175;
  wire and_dcpl_180;
  wire and_dcpl_185;
  wire and_dcpl_190;
  wire and_dcpl_191;
  wire and_dcpl_192;
  wire and_dcpl_193;
  wire and_dcpl_195;
  wire and_dcpl_197;
  wire and_dcpl_198;
  wire and_dcpl_200;
  wire and_dcpl_202;
  wire and_dcpl_207;
  wire and_dcpl_212;
  wire and_dcpl_217;
  wire and_dcpl_218;
  wire and_dcpl_219;
  wire and_dcpl_220;
  wire and_dcpl_222;
  wire and_dcpl_224;
  wire and_dcpl_225;
  wire and_dcpl_227;
  wire and_dcpl_229;
  wire and_dcpl_234;
  wire and_dcpl_239;
  wire and_dcpl_244;
  wire and_dcpl_245;
  wire and_dcpl_246;
  wire and_dcpl_247;
  wire and_dcpl_249;
  wire and_dcpl_251;
  wire and_dcpl_252;
  wire and_dcpl_254;
  wire and_dcpl_256;
  wire and_dcpl_261;
  wire and_dcpl_266;
  wire and_dcpl_271;
  wire and_dcpl_272;
  wire and_dcpl_274;
  wire and_dcpl_276;
  wire and_dcpl_278;
  wire and_dcpl_280;
  wire and_dcpl_285;
  wire and_dcpl_291;
  wire and_dcpl_292;
  wire and_dcpl_293;
  wire and_dcpl_294;
  wire and_dcpl_295;
  wire and_dcpl_296;
  wire and_dcpl_298;
  wire not_tmp_54;
  wire or_tmp_2;
  wire and_dcpl_300;
  wire and_dcpl_301;
  wire and_dcpl_302;
  wire and_dcpl_304;
  wire and_tmp;
  wire and_dcpl_306;
  wire and_dcpl_307;
  wire and_dcpl_308;
  wire and_dcpl_310;
  wire and_tmp_2;
  wire and_dcpl_312;
  wire and_dcpl_313;
  wire and_dcpl_314;
  wire and_dcpl_316;
  wire and_tmp_5;
  wire and_dcpl_318;
  wire and_tmp_9;
  wire and_dcpl_324;
  wire and_tmp_13;
  wire and_dcpl_330;
  wire mux_tmp_19;
  wire and_tmp_17;
  wire and_dcpl_336;
  wire mux_tmp_22;
  wire mux_tmp_23;
  wire and_tmp_21;
  wire and_dcpl_342;
  wire mux_tmp_26;
  wire mux_tmp_27;
  wire mux_tmp_28;
  wire and_tmp_25;
  wire and_dcpl_348;
  wire and_tmp_35;
  wire and_dcpl_355;
  wire and_dcpl_356;
  wire and_dcpl_358;
  wire or_tmp_80;
  wire and_dcpl_360;
  wire and_dcpl_362;
  wire mux_tmp_32;
  wire and_dcpl_364;
  wire and_dcpl_366;
  wire mux_tmp_34;
  wire mux_tmp_35;
  wire and_dcpl_368;
  wire and_dcpl_370;
  wire mux_tmp_37;
  wire mux_tmp_38;
  wire mux_tmp_39;
  wire and_dcpl_372;
  wire mux_tmp_41;
  wire mux_tmp_42;
  wire mux_tmp_43;
  wire mux_tmp_44;
  wire and_dcpl_376;
  wire mux_tmp_46;
  wire mux_tmp_47;
  wire mux_tmp_48;
  wire mux_tmp_49;
  wire mux_tmp_50;
  wire and_dcpl_379;
  wire mux_tmp_52;
  wire mux_tmp_53;
  wire mux_tmp_54;
  wire mux_tmp_55;
  wire mux_tmp_56;
  wire mux_tmp_57;
  wire and_dcpl_382;
  wire mux_tmp_59;
  wire mux_tmp_60;
  wire mux_tmp_61;
  wire mux_tmp_62;
  wire mux_tmp_63;
  wire mux_tmp_64;
  wire mux_tmp_65;
  wire and_dcpl_385;
  wire mux_tmp_67;
  wire mux_tmp_68;
  wire mux_tmp_69;
  wire mux_tmp_70;
  wire mux_tmp_71;
  wire mux_tmp_72;
  wire mux_tmp_73;
  wire mux_tmp_74;
  wire and_dcpl_388;
  wire and_tmp_44;
  wire mux_tmp_76;
  wire and_dcpl_393;
  wire and_dcpl_394;
  wire and_dcpl_395;
  wire or_tmp_185;
  wire and_dcpl_397;
  wire and_dcpl_398;
  wire and_tmp_45;
  wire and_dcpl_400;
  wire and_dcpl_401;
  wire and_tmp_47;
  wire and_dcpl_403;
  wire and_dcpl_404;
  wire and_tmp_50;
  wire and_dcpl_406;
  wire and_tmp_54;
  wire and_dcpl_409;
  wire and_tmp_58;
  wire and_dcpl_413;
  wire mux_tmp_84;
  wire and_tmp_62;
  wire and_dcpl_417;
  wire mux_tmp_87;
  wire mux_tmp_88;
  wire and_tmp_66;
  wire and_dcpl_421;
  wire mux_tmp_91;
  wire mux_tmp_92;
  wire mux_tmp_93;
  wire and_tmp_70;
  wire and_dcpl_425;
  wire and_tmp_80;
  wire and_dcpl_430;
  wire and_dcpl_431;
  wire or_tmp_263;
  wire and_dcpl_433;
  wire mux_tmp_97;
  wire and_dcpl_435;
  wire mux_tmp_99;
  wire mux_tmp_100;
  wire and_dcpl_437;
  wire mux_tmp_102;
  wire mux_tmp_103;
  wire mux_tmp_104;
  wire and_dcpl_439;
  wire mux_tmp_106;
  wire mux_tmp_107;
  wire mux_tmp_108;
  wire mux_tmp_109;
  wire and_dcpl_442;
  wire mux_tmp_111;
  wire mux_tmp_112;
  wire mux_tmp_113;
  wire mux_tmp_114;
  wire mux_tmp_115;
  wire and_dcpl_445;
  wire mux_tmp_117;
  wire mux_tmp_118;
  wire mux_tmp_119;
  wire mux_tmp_120;
  wire mux_tmp_121;
  wire mux_tmp_122;
  wire and_dcpl_448;
  wire mux_tmp_124;
  wire mux_tmp_125;
  wire mux_tmp_126;
  wire mux_tmp_127;
  wire mux_tmp_128;
  wire mux_tmp_129;
  wire mux_tmp_130;
  wire and_dcpl_451;
  wire mux_tmp_132;
  wire mux_tmp_133;
  wire mux_tmp_134;
  wire mux_tmp_135;
  wire mux_tmp_136;
  wire mux_tmp_137;
  wire mux_tmp_138;
  wire mux_tmp_139;
  wire and_dcpl_454;
  wire and_tmp_89;
  wire mux_tmp_141;
  wire and_dcpl_460;
  wire and_dcpl_461;
  wire and_dcpl_462;
  wire and_dcpl_463;
  wire not_tmp_332;
  wire or_tmp_368;
  wire and_dcpl_465;
  wire and_dcpl_466;
  wire and_dcpl_467;
  wire and_tmp_90;
  wire and_dcpl_469;
  wire and_dcpl_470;
  wire and_dcpl_471;
  wire and_tmp_92;
  wire and_dcpl_473;
  wire and_dcpl_474;
  wire and_dcpl_475;
  wire and_tmp_95;
  wire and_dcpl_477;
  wire and_tmp_99;
  wire and_dcpl_480;
  wire and_tmp_103;
  wire and_dcpl_483;
  wire mux_tmp_149;
  wire and_tmp_107;
  wire and_dcpl_486;
  wire mux_tmp_152;
  wire mux_tmp_153;
  wire and_tmp_111;
  wire and_dcpl_489;
  wire mux_tmp_156;
  wire mux_tmp_157;
  wire mux_tmp_158;
  wire and_tmp_115;
  wire and_dcpl_492;
  wire and_tmp_125;
  wire and_dcpl_498;
  wire or_tmp_446;
  wire and_dcpl_500;
  wire mux_tmp_162;
  wire and_dcpl_502;
  wire mux_tmp_164;
  wire mux_tmp_165;
  wire and_dcpl_504;
  wire mux_tmp_167;
  wire mux_tmp_168;
  wire mux_tmp_169;
  wire and_dcpl_506;
  wire mux_tmp_171;
  wire mux_tmp_172;
  wire mux_tmp_173;
  wire mux_tmp_174;
  wire and_dcpl_508;
  wire mux_tmp_176;
  wire mux_tmp_177;
  wire mux_tmp_178;
  wire mux_tmp_179;
  wire mux_tmp_180;
  wire and_dcpl_510;
  wire mux_tmp_182;
  wire mux_tmp_183;
  wire mux_tmp_184;
  wire mux_tmp_185;
  wire mux_tmp_186;
  wire mux_tmp_187;
  wire and_dcpl_512;
  wire mux_tmp_189;
  wire mux_tmp_190;
  wire mux_tmp_191;
  wire mux_tmp_192;
  wire mux_tmp_193;
  wire mux_tmp_194;
  wire mux_tmp_195;
  wire and_dcpl_514;
  wire mux_tmp_197;
  wire mux_tmp_198;
  wire mux_tmp_199;
  wire mux_tmp_200;
  wire mux_tmp_201;
  wire mux_tmp_202;
  wire mux_tmp_203;
  wire mux_tmp_204;
  wire and_dcpl_516;
  wire and_tmp_134;
  wire mux_tmp_206;
  wire and_dcpl_520;
  wire and_dcpl_521;
  wire or_tmp_551;
  wire and_dcpl_523;
  wire and_dcpl_524;
  wire and_tmp_135;
  wire and_dcpl_526;
  wire and_dcpl_527;
  wire and_tmp_137;
  wire and_dcpl_529;
  wire and_dcpl_530;
  wire and_tmp_140;
  wire and_dcpl_532;
  wire and_tmp_144;
  wire and_dcpl_534;
  wire and_tmp_148;
  wire and_dcpl_536;
  wire mux_tmp_214;
  wire and_tmp_152;
  wire and_dcpl_538;
  wire mux_tmp_217;
  wire mux_tmp_218;
  wire and_tmp_156;
  wire and_dcpl_540;
  wire mux_tmp_221;
  wire mux_tmp_222;
  wire mux_tmp_223;
  wire and_tmp_160;
  wire and_dcpl_542;
  wire and_tmp_170;
  wire and_dcpl_546;
  wire or_tmp_629;
  wire and_dcpl_548;
  wire mux_tmp_227;
  wire and_dcpl_550;
  wire mux_tmp_229;
  wire mux_tmp_230;
  wire and_dcpl_552;
  wire mux_tmp_232;
  wire mux_tmp_233;
  wire mux_tmp_234;
  wire and_dcpl_554;
  wire mux_tmp_236;
  wire mux_tmp_237;
  wire mux_tmp_238;
  wire mux_tmp_239;
  wire and_dcpl_556;
  wire mux_tmp_241;
  wire mux_tmp_242;
  wire mux_tmp_243;
  wire mux_tmp_244;
  wire mux_tmp_245;
  wire and_dcpl_558;
  wire mux_tmp_247;
  wire mux_tmp_248;
  wire mux_tmp_249;
  wire mux_tmp_250;
  wire mux_tmp_251;
  wire mux_tmp_252;
  wire and_dcpl_560;
  wire mux_tmp_254;
  wire mux_tmp_255;
  wire mux_tmp_256;
  wire mux_tmp_257;
  wire mux_tmp_258;
  wire mux_tmp_259;
  wire mux_tmp_260;
  wire and_dcpl_562;
  wire mux_tmp_262;
  wire mux_tmp_263;
  wire mux_tmp_264;
  wire mux_tmp_265;
  wire mux_tmp_266;
  wire mux_tmp_267;
  wire mux_tmp_268;
  wire mux_tmp_269;
  wire and_dcpl_564;
  wire and_tmp_179;
  wire mux_tmp_271;
  wire and_dcpl_568;
  wire and_dcpl_569;
  wire and_dcpl_570;
  wire and_dcpl_571;
  wire or_tmp_733;
  wire and_dcpl_573;
  wire and_dcpl_574;
  wire and_dcpl_575;
  wire and_tmp_180;
  wire and_dcpl_577;
  wire and_dcpl_578;
  wire and_dcpl_579;
  wire and_tmp_182;
  wire and_dcpl_581;
  wire and_dcpl_582;
  wire and_dcpl_583;
  wire and_tmp_185;
  wire and_dcpl_585;
  wire and_tmp_189;
  wire and_dcpl_589;
  wire and_tmp_193;
  wire and_dcpl_593;
  wire mux_tmp_279;
  wire and_tmp_197;
  wire and_dcpl_597;
  wire mux_tmp_282;
  wire mux_tmp_283;
  wire and_tmp_201;
  wire and_dcpl_601;
  wire mux_tmp_286;
  wire mux_tmp_287;
  wire mux_tmp_288;
  wire and_tmp_205;
  wire and_dcpl_605;
  wire or_tmp_808;
  wire mux_tmp_291;
  wire mux_tmp_292;
  wire mux_tmp_293;
  wire mux_tmp_294;
  wire mux_tmp_295;
  wire mux_tmp_296;
  wire mux_tmp_297;
  wire mux_tmp_298;
  wire and_tmp_206;
  wire and_dcpl_610;
  wire or_tmp_820;
  wire and_dcpl_612;
  wire mux_tmp_301;
  wire and_dcpl_614;
  wire mux_tmp_303;
  wire mux_tmp_304;
  wire and_dcpl_616;
  wire mux_tmp_306;
  wire mux_tmp_307;
  wire mux_tmp_308;
  wire and_dcpl_618;
  wire mux_tmp_310;
  wire mux_tmp_311;
  wire mux_tmp_312;
  wire mux_tmp_313;
  wire and_dcpl_622;
  wire mux_tmp_315;
  wire mux_tmp_316;
  wire mux_tmp_317;
  wire mux_tmp_318;
  wire mux_tmp_319;
  wire and_dcpl_625;
  wire mux_tmp_321;
  wire mux_tmp_322;
  wire mux_tmp_323;
  wire mux_tmp_324;
  wire mux_tmp_325;
  wire mux_tmp_326;
  wire and_dcpl_628;
  wire mux_tmp_328;
  wire mux_tmp_329;
  wire mux_tmp_330;
  wire mux_tmp_331;
  wire mux_tmp_332;
  wire mux_tmp_333;
  wire mux_tmp_334;
  wire and_dcpl_631;
  wire mux_tmp_336;
  wire mux_tmp_337;
  wire mux_tmp_338;
  wire mux_tmp_339;
  wire mux_tmp_340;
  wire mux_tmp_341;
  wire mux_tmp_342;
  wire mux_tmp_343;
  wire and_dcpl_634;
  wire or_tmp_921;
  wire mux_tmp_345;
  wire mux_tmp_346;
  wire mux_tmp_347;
  wire mux_tmp_348;
  wire mux_tmp_349;
  wire mux_tmp_350;
  wire mux_tmp_351;
  wire mux_tmp_352;
  wire mux_tmp_353;
  wire mux_tmp_354;
  wire and_dcpl_638;
  wire and_dcpl_639;
  wire or_tmp_934;
  wire and_dcpl_641;
  wire and_dcpl_642;
  wire and_tmp_207;
  wire and_dcpl_644;
  wire and_dcpl_645;
  wire and_tmp_209;
  wire and_dcpl_647;
  wire and_dcpl_648;
  wire and_tmp_212;
  wire and_dcpl_650;
  wire and_tmp_216;
  wire and_dcpl_653;
  wire and_tmp_220;
  wire and_dcpl_657;
  wire mux_tmp_362;
  wire and_tmp_224;
  wire and_dcpl_661;
  wire mux_tmp_365;
  wire mux_tmp_366;
  wire and_tmp_228;
  wire and_dcpl_665;
  wire mux_tmp_369;
  wire mux_tmp_370;
  wire mux_tmp_371;
  wire and_tmp_232;
  wire and_dcpl_669;
  wire or_tmp_1009;
  wire mux_tmp_374;
  wire mux_tmp_375;
  wire mux_tmp_376;
  wire mux_tmp_377;
  wire mux_tmp_378;
  wire mux_tmp_379;
  wire mux_tmp_380;
  wire mux_tmp_381;
  wire and_tmp_233;
  wire and_dcpl_673;
  wire or_tmp_1021;
  wire and_dcpl_675;
  wire mux_tmp_384;
  wire and_dcpl_677;
  wire mux_tmp_386;
  wire mux_tmp_387;
  wire and_dcpl_679;
  wire mux_tmp_389;
  wire mux_tmp_390;
  wire mux_tmp_391;
  wire and_dcpl_681;
  wire mux_tmp_393;
  wire mux_tmp_394;
  wire mux_tmp_395;
  wire mux_tmp_396;
  wire and_dcpl_684;
  wire mux_tmp_398;
  wire mux_tmp_399;
  wire mux_tmp_400;
  wire mux_tmp_401;
  wire mux_tmp_402;
  wire and_dcpl_687;
  wire mux_tmp_404;
  wire mux_tmp_405;
  wire mux_tmp_406;
  wire mux_tmp_407;
  wire mux_tmp_408;
  wire mux_tmp_409;
  wire and_dcpl_690;
  wire mux_tmp_411;
  wire mux_tmp_412;
  wire mux_tmp_413;
  wire mux_tmp_414;
  wire mux_tmp_415;
  wire mux_tmp_416;
  wire mux_tmp_417;
  wire and_dcpl_693;
  wire mux_tmp_419;
  wire mux_tmp_420;
  wire mux_tmp_421;
  wire mux_tmp_422;
  wire mux_tmp_423;
  wire mux_tmp_424;
  wire mux_tmp_425;
  wire mux_tmp_426;
  wire and_dcpl_696;
  wire or_tmp_1122;
  wire mux_tmp_428;
  wire mux_tmp_429;
  wire mux_tmp_430;
  wire mux_tmp_431;
  wire mux_tmp_432;
  wire mux_tmp_433;
  wire mux_tmp_434;
  wire mux_tmp_435;
  wire mux_tmp_436;
  wire mux_tmp_437;
  reg [1:0] rem_12cyc_st_10_1_0;
  reg [1:0] rem_12cyc_st_10_3_2;
  reg [1:0] rem_12cyc_st_9_1_0;
  reg [1:0] rem_12cyc_st_9_3_2;
  reg [1:0] rem_12cyc_st_8_1_0;
  reg [1:0] rem_12cyc_st_8_3_2;
  reg [1:0] rem_12cyc_st_7_1_0;
  reg [1:0] rem_12cyc_st_7_3_2;
  reg [1:0] rem_12cyc_st_6_1_0;
  reg [1:0] rem_12cyc_st_6_3_2;
  reg [1:0] rem_12cyc_st_5_1_0;
  reg [1:0] rem_12cyc_st_5_3_2;
  reg [1:0] rem_12cyc_st_4_1_0;
  reg [1:0] rem_12cyc_st_4_3_2;
  reg [1:0] rem_12cyc_st_3_1_0;
  reg [1:0] rem_12cyc_st_3_3_2;
  reg [1:0] rem_12cyc_st_2_1_0;
  reg [1:0] rem_12cyc_st_2_3_2;
  reg [1:0] rem_12cyc_1_0;
  reg [1:0] rem_12cyc_3_2;
  reg [1:0] rem_12cyc_st_12_3_2;
  reg [63:0] result_sva_duc;
  reg [1:0] rem_12cyc_st_12_1_0;
  reg COMP_LOOP_asn_itm_12;
  reg main_stage_0_13;
  reg main_stage_0_3;
  reg COMP_LOOP_asn_itm_1;
  reg main_stage_0_2;
  reg main_stage_0_4;
  reg COMP_LOOP_asn_itm_2;
  reg main_stage_0_5;
  reg COMP_LOOP_asn_itm_3;
  reg main_stage_0_6;
  reg COMP_LOOP_asn_itm_4;
  reg COMP_LOOP_asn_itm_5;
  reg main_stage_0_8;
  reg COMP_LOOP_asn_itm_7;
  reg main_stage_0_9;
  reg COMP_LOOP_asn_itm_8;
  reg main_stage_0_10;
  reg COMP_LOOP_asn_itm_9;
  reg main_stage_0_7;
  reg COMP_LOOP_asn_itm_6;
  reg main_stage_0_11;
  reg COMP_LOOP_asn_itm_10;
  wire COMP_LOOP_and_cse;
  wire COMP_LOOP_and_2_cse;
  wire COMP_LOOP_and_4_cse;
  wire COMP_LOOP_and_6_cse;
  wire COMP_LOOP_and_8_cse;
  wire COMP_LOOP_and_10_cse;
  wire COMP_LOOP_and_12_cse;
  wire COMP_LOOP_and_14_cse;
  wire COMP_LOOP_and_16_cse;
  wire COMP_LOOP_and_18_cse;
  wire COMP_LOOP_and_20_cse;
  wire COMP_LOOP_and_22_cse;
  wire COMP_LOOP_and_24_cse;
  wire or_1_cse;
  wire or_6_cse;
  wire or_10_cse;
  wire or_15_cse;
  wire or_21_cse;
  wire or_28_cse;
  wire or_37_cse;
  wire or_48_cse;
  wire or_83_cse;
  wire nand_276_cse;
  wire or_88_cse;
  wire nand_274_cse;
  wire or_93_cse;
  wire nand_271_cse;
  wire or_100_cse;
  wire nand_267_cse;
  wire or_109_cse;
  wire or_120_cse;
  wire or_133_cse;
  wire or_148_cse;
  wire or_190_cse;
  wire or_195_cse;
  wire or_199_cse;
  wire or_204_cse;
  wire or_210_cse;
  wire or_217_cse;
  wire or_226_cse;
  wire or_237_cse;
  wire or_270_cse;
  wire or_275_cse;
  wire or_280_cse;
  wire or_287_cse;
  wire or_296_cse;
  wire or_307_cse;
  wire or_320_cse;
  wire or_335_cse;
  wire nand_281_cse;
  wire or_377_cse;
  wire or_382_cse;
  wire or_386_cse;
  wire or_391_cse;
  wire or_397_cse;
  wire nand_215_cse;
  wire or_404_cse;
  wire nand_212_cse;
  wire or_413_cse;
  wire nand_208_cse;
  wire or_424_cse;
  wire or_458_cse;
  wire or_463_cse;
  wire nand_198_cse;
  wire or_468_cse;
  wire or_475_cse;
  wire nand_189_cse;
  wire or_484_cse;
  wire or_495_cse;
  wire or_508_cse;
  wire nand_203_cse;
  wire or_523_cse;
  wire nand_250_cse;
  wire or_564_cse;
  wire or_569_cse;
  wire or_573_cse;
  wire or_578_cse;
  wire or_584_cse;
  wire or_591_cse;
  wire or_600_cse;
  wire or_611_cse;
  wire or_643_cse;
  wire or_648_cse;
  wire or_653_cse;
  wire or_660_cse;
  wire or_669_cse;
  wire or_680_cse;
  wire or_693_cse;
  wire or_708_cse;
  wire or_748_cse;
  wire or_753_cse;
  wire or_757_cse;
  wire or_762_cse;
  wire or_768_cse;
  wire or_775_cse;
  wire or_784_cse;
  wire or_795_cse;
  wire or_837_cse;
  wire nand_84_cse;
  wire or_842_cse;
  wire or_847_cse;
  wire nand_79_cse;
  wire or_854_cse;
  wire or_863_cse;
  wire or_874_cse;
  wire or_887_cse;
  wire or_902_cse;
  wire or_952_cse;
  wire or_957_cse;
  wire or_961_cse;
  wire or_966_cse;
  wire or_972_cse;
  wire or_979_cse;
  wire or_988_cse;
  wire or_999_cse;
  wire nand_57_cse;
  wire or_1045_cse;
  wire or_1050_cse;
  wire or_1057_cse;
  wire or_1066_cse;
  wire nand_36_cse;
  wire nand_29_cse;
  wire nand_21_cse;
  wire nand_222_cse;
  wire nand_223_cse;
  reg main_stage_0_12;
  reg [63:0] m_buf_sva_1;
  reg [63:0] m_buf_sva_2;
  reg [63:0] m_buf_sva_3;
  reg [63:0] m_buf_sva_4;
  reg [63:0] m_buf_sva_5;
  reg [63:0] m_buf_sva_6;
  reg [63:0] m_buf_sva_7;
  reg [63:0] m_buf_sva_8;
  reg [63:0] m_buf_sva_9;
  reg [63:0] m_buf_sva_10;
  reg [63:0] m_buf_sva_11;
  reg [63:0] m_buf_sva_12;
  reg COMP_LOOP_asn_itm_11;
  reg [63:0] mut_2_63_0;
  reg [63:0] mut_3_63_0;
  reg [63:0] mut_4_63_0;
  reg [63:0] mut_5_63_0;
  reg [63:0] mut_6_63_0;
  reg [63:0] mut_7_63_0;
  reg [63:0] mut_8_63_0;
  reg [63:0] mut_9_63_0;
  reg [63:0] mut_10_63_0;
  reg [63:0] mut_11_63_0;
  reg [63:0] mut_1_2_63_0;
  reg [63:0] mut_1_3_63_0;
  reg [63:0] mut_1_4_63_0;
  reg [63:0] mut_1_5_63_0;
  reg [63:0] mut_1_6_63_0;
  reg [63:0] mut_1_7_63_0;
  reg [63:0] mut_1_8_63_0;
  reg [63:0] mut_1_9_63_0;
  reg [63:0] mut_1_10_63_0;
  reg [63:0] mut_1_11_63_0;
  reg [63:0] mut_2_2_63_0;
  reg [63:0] mut_2_3_63_0;
  reg [63:0] mut_2_4_63_0;
  reg [63:0] mut_2_5_63_0;
  reg [63:0] mut_2_6_63_0;
  reg [63:0] mut_2_7_63_0;
  reg [63:0] mut_2_8_63_0;
  reg [63:0] mut_2_9_63_0;
  reg [63:0] mut_2_10_63_0;
  reg [63:0] mut_2_11_63_0;
  reg [63:0] mut_3_2_63_0;
  reg [63:0] mut_3_3_63_0;
  reg [63:0] mut_3_4_63_0;
  reg [63:0] mut_3_5_63_0;
  reg [63:0] mut_3_6_63_0;
  reg [63:0] mut_3_7_63_0;
  reg [63:0] mut_3_8_63_0;
  reg [63:0] mut_3_9_63_0;
  reg [63:0] mut_3_10_63_0;
  reg [63:0] mut_3_11_63_0;
  reg [63:0] mut_4_2_63_0;
  reg [63:0] mut_4_3_63_0;
  reg [63:0] mut_4_4_63_0;
  reg [63:0] mut_4_5_63_0;
  reg [63:0] mut_4_6_63_0;
  reg [63:0] mut_4_7_63_0;
  reg [63:0] mut_4_8_63_0;
  reg [63:0] mut_4_9_63_0;
  reg [63:0] mut_4_10_63_0;
  reg [63:0] mut_4_11_63_0;
  reg [63:0] mut_5_2_63_0;
  reg [63:0] mut_5_3_63_0;
  reg [63:0] mut_5_4_63_0;
  reg [63:0] mut_5_5_63_0;
  reg [63:0] mut_5_6_63_0;
  reg [63:0] mut_5_7_63_0;
  reg [63:0] mut_5_8_63_0;
  reg [63:0] mut_5_9_63_0;
  reg [63:0] mut_5_10_63_0;
  reg [63:0] mut_5_11_63_0;
  reg [63:0] mut_6_2_63_0;
  reg [63:0] mut_6_3_63_0;
  reg [63:0] mut_6_4_63_0;
  reg [63:0] mut_6_5_63_0;
  reg [63:0] mut_6_6_63_0;
  reg [63:0] mut_6_7_63_0;
  reg [63:0] mut_6_8_63_0;
  reg [63:0] mut_6_9_63_0;
  reg [63:0] mut_6_10_63_0;
  reg [63:0] mut_6_11_63_0;
  reg [63:0] mut_7_2_63_0;
  reg [63:0] mut_7_3_63_0;
  reg [63:0] mut_7_4_63_0;
  reg [63:0] mut_7_5_63_0;
  reg [63:0] mut_7_6_63_0;
  reg [63:0] mut_7_7_63_0;
  reg [63:0] mut_7_8_63_0;
  reg [63:0] mut_7_9_63_0;
  reg [63:0] mut_7_10_63_0;
  reg [63:0] mut_7_11_63_0;
  reg [63:0] mut_8_2_63_0;
  reg [63:0] mut_8_3_63_0;
  reg [63:0] mut_8_4_63_0;
  reg [63:0] mut_8_5_63_0;
  reg [63:0] mut_8_6_63_0;
  reg [63:0] mut_8_7_63_0;
  reg [63:0] mut_8_8_63_0;
  reg [63:0] mut_8_9_63_0;
  reg [63:0] mut_8_10_63_0;
  reg [63:0] mut_8_11_63_0;
  reg [63:0] mut_9_2_63_0;
  reg [63:0] mut_9_3_63_0;
  reg [63:0] mut_9_4_63_0;
  reg [63:0] mut_9_5_63_0;
  reg [63:0] mut_9_6_63_0;
  reg [63:0] mut_9_7_63_0;
  reg [63:0] mut_9_8_63_0;
  reg [63:0] mut_9_9_63_0;
  reg [63:0] mut_9_10_63_0;
  reg [63:0] mut_9_11_63_0;
  reg [63:0] mut_10_2_63_0;
  reg [63:0] mut_10_3_63_0;
  reg [63:0] mut_10_4_63_0;
  reg [63:0] mut_10_5_63_0;
  reg [63:0] mut_10_6_63_0;
  reg [63:0] mut_10_7_63_0;
  reg [63:0] mut_10_8_63_0;
  reg [63:0] mut_10_9_63_0;
  reg [63:0] mut_10_10_63_0;
  reg [63:0] mut_10_11_63_0;
  reg [63:0] mut_11_2_63_0;
  reg [63:0] mut_11_3_63_0;
  reg [63:0] mut_11_4_63_0;
  reg [63:0] mut_11_5_63_0;
  reg [63:0] mut_11_6_63_0;
  reg [63:0] mut_11_7_63_0;
  reg [63:0] mut_11_8_63_0;
  reg [63:0] mut_11_9_63_0;
  reg [63:0] mut_11_10_63_0;
  reg [63:0] mut_11_11_63_0;
  reg [63:0] mut_12_2_63_0;
  reg [63:0] mut_12_3_63_0;
  reg [63:0] mut_12_4_63_0;
  reg [63:0] mut_12_5_63_0;
  reg [63:0] mut_12_6_63_0;
  reg [63:0] mut_12_7_63_0;
  reg [63:0] mut_12_8_63_0;
  reg [63:0] mut_12_9_63_0;
  reg [63:0] mut_12_10_63_0;
  reg [63:0] mut_12_11_63_0;
  reg [63:0] mut_13_2_63_0;
  reg [63:0] mut_13_3_63_0;
  reg [63:0] mut_13_4_63_0;
  reg [63:0] mut_13_5_63_0;
  reg [63:0] mut_13_6_63_0;
  reg [63:0] mut_13_7_63_0;
  reg [63:0] mut_13_8_63_0;
  reg [63:0] mut_13_9_63_0;
  reg [63:0] mut_13_10_63_0;
  reg [63:0] mut_13_11_63_0;
  reg [63:0] mut_14_2_63_0;
  reg [63:0] mut_14_3_63_0;
  reg [63:0] mut_14_4_63_0;
  reg [63:0] mut_14_5_63_0;
  reg [63:0] mut_14_6_63_0;
  reg [63:0] mut_14_7_63_0;
  reg [63:0] mut_14_8_63_0;
  reg [63:0] mut_14_9_63_0;
  reg [63:0] mut_14_10_63_0;
  reg [63:0] mut_14_11_63_0;
  reg [63:0] mut_15_2_63_0;
  reg [63:0] mut_15_3_63_0;
  reg [63:0] mut_15_4_63_0;
  reg [63:0] mut_15_5_63_0;
  reg [63:0] mut_15_6_63_0;
  reg [63:0] mut_15_7_63_0;
  reg [63:0] mut_15_8_63_0;
  reg [63:0] mut_15_9_63_0;
  reg [63:0] mut_15_10_63_0;
  reg [63:0] mut_15_11_63_0;
  reg [63:0] mut_16_2_63_0;
  reg [63:0] mut_16_3_63_0;
  reg [63:0] mut_16_4_63_0;
  reg [63:0] mut_16_5_63_0;
  reg [63:0] mut_16_6_63_0;
  reg [63:0] mut_16_7_63_0;
  reg [63:0] mut_16_8_63_0;
  reg [63:0] mut_16_9_63_0;
  reg [63:0] mut_16_10_63_0;
  reg [63:0] mut_16_11_63_0;
  reg [63:0] mut_17_2_63_0;
  reg [63:0] mut_17_3_63_0;
  reg [63:0] mut_17_4_63_0;
  reg [63:0] mut_17_5_63_0;
  reg [63:0] mut_17_6_63_0;
  reg [63:0] mut_17_7_63_0;
  reg [63:0] mut_17_8_63_0;
  reg [63:0] mut_17_9_63_0;
  reg [63:0] mut_17_10_63_0;
  reg [63:0] mut_17_11_63_0;
  reg [63:0] mut_18_2_63_0;
  reg [63:0] mut_18_3_63_0;
  reg [63:0] mut_18_4_63_0;
  reg [63:0] mut_18_5_63_0;
  reg [63:0] mut_18_6_63_0;
  reg [63:0] mut_18_7_63_0;
  reg [63:0] mut_18_8_63_0;
  reg [63:0] mut_18_9_63_0;
  reg [63:0] mut_18_10_63_0;
  reg [63:0] mut_18_11_63_0;
  reg [63:0] mut_19_2_63_0;
  reg [63:0] mut_19_3_63_0;
  reg [63:0] mut_19_4_63_0;
  reg [63:0] mut_19_5_63_0;
  reg [63:0] mut_19_6_63_0;
  reg [63:0] mut_19_7_63_0;
  reg [63:0] mut_19_8_63_0;
  reg [63:0] mut_19_9_63_0;
  reg [63:0] mut_19_10_63_0;
  reg [63:0] mut_19_11_63_0;
  reg [63:0] mut_20_2_63_0;
  reg [63:0] mut_20_3_63_0;
  reg [63:0] mut_20_4_63_0;
  reg [63:0] mut_20_5_63_0;
  reg [63:0] mut_20_6_63_0;
  reg [63:0] mut_20_7_63_0;
  reg [63:0] mut_20_8_63_0;
  reg [63:0] mut_20_9_63_0;
  reg [63:0] mut_20_10_63_0;
  reg [63:0] mut_20_11_63_0;
  reg [63:0] mut_21_2_63_0;
  reg [63:0] mut_21_3_63_0;
  reg [63:0] mut_21_4_63_0;
  reg [63:0] mut_21_5_63_0;
  reg [63:0] mut_21_6_63_0;
  reg [63:0] mut_21_7_63_0;
  reg [63:0] mut_21_8_63_0;
  reg [63:0] mut_21_9_63_0;
  reg [63:0] mut_21_10_63_0;
  reg [63:0] mut_21_11_63_0;
  reg [63:0] mut_22_2_63_0;
  reg [63:0] mut_22_3_63_0;
  reg [63:0] mut_22_4_63_0;
  reg [63:0] mut_22_5_63_0;
  reg [63:0] mut_22_6_63_0;
  reg [63:0] mut_22_7_63_0;
  reg [63:0] mut_22_8_63_0;
  reg [63:0] mut_22_9_63_0;
  reg [63:0] mut_22_10_63_0;
  reg [63:0] mut_22_11_63_0;
  reg [63:0] mut_23_2_63_0;
  reg [63:0] mut_23_3_63_0;
  reg [63:0] mut_23_4_63_0;
  reg [63:0] mut_23_5_63_0;
  reg [63:0] mut_23_6_63_0;
  reg [63:0] mut_23_7_63_0;
  reg [63:0] mut_23_8_63_0;
  reg [63:0] mut_23_9_63_0;
  reg [63:0] mut_23_10_63_0;
  reg [63:0] mut_23_11_63_0;
  reg [1:0] rem_12cyc_st_11_3_2;
  reg [1:0] rem_12cyc_st_11_1_0;
  wire [63:0] result_sva_duc_mx0;
  wire COMP_LOOP_and_26_cse;
  wire COMP_LOOP_and_28_cse;
  wire COMP_LOOP_and_30_cse;
  wire COMP_LOOP_and_32_cse;
  wire COMP_LOOP_and_34_cse;
  wire COMP_LOOP_and_36_cse;
  wire COMP_LOOP_and_38_cse;
  wire COMP_LOOP_and_40_cse;
  wire COMP_LOOP_and_42_cse;
  wire COMP_LOOP_and_44_cse;
  wire COMP_LOOP_and_46_cse;
  wire COMP_LOOP_and_48_cse;
  wire COMP_LOOP_and_50_cse;
  wire COMP_LOOP_and_52_cse;
  wire COMP_LOOP_and_54_cse;
  wire COMP_LOOP_and_56_cse;
  wire COMP_LOOP_and_58_cse;
  wire COMP_LOOP_and_60_cse;
  wire COMP_LOOP_and_62_cse;
  wire COMP_LOOP_and_64_cse;
  wire COMP_LOOP_and_66_cse;
  wire COMP_LOOP_and_68_cse;
  wire COMP_LOOP_and_70_cse;
  wire COMP_LOOP_and_72_cse;
  wire COMP_LOOP_and_74_cse;
  wire COMP_LOOP_and_76_cse;
  wire COMP_LOOP_and_78_cse;
  wire COMP_LOOP_and_80_cse;
  wire COMP_LOOP_and_82_cse;
  wire COMP_LOOP_and_84_cse;
  wire COMP_LOOP_and_86_cse;
  wire COMP_LOOP_and_88_cse;
  wire COMP_LOOP_and_90_cse;
  wire COMP_LOOP_and_92_cse;
  wire COMP_LOOP_and_94_cse;
  wire COMP_LOOP_and_96_cse;
  wire COMP_LOOP_and_98_cse;
  wire COMP_LOOP_and_100_cse;
  wire COMP_LOOP_and_102_cse;
  wire COMP_LOOP_and_104_cse;
  wire COMP_LOOP_and_106_cse;
  wire COMP_LOOP_and_108_cse;
  wire COMP_LOOP_and_110_cse;
  wire COMP_LOOP_and_112_cse;
  wire COMP_LOOP_and_114_cse;
  wire COMP_LOOP_and_116_cse;
  wire COMP_LOOP_and_118_cse;
  wire COMP_LOOP_and_120_cse;
  wire COMP_LOOP_and_122_cse;
  wire COMP_LOOP_and_124_cse;
  wire COMP_LOOP_and_126_cse;
  wire COMP_LOOP_and_128_cse;
  wire COMP_LOOP_and_130_cse;
  wire COMP_LOOP_and_132_cse;
  wire COMP_LOOP_and_134_cse;
  wire COMP_LOOP_and_136_cse;
  wire COMP_LOOP_and_138_cse;
  wire COMP_LOOP_and_140_cse;
  wire COMP_LOOP_and_142_cse;
  wire COMP_LOOP_and_144_cse;
  wire COMP_LOOP_and_146_cse;
  wire COMP_LOOP_and_148_cse;
  wire COMP_LOOP_and_150_cse;
  wire COMP_LOOP_and_152_cse;
  wire COMP_LOOP_and_154_cse;
  wire COMP_LOOP_and_156_cse;
  wire COMP_LOOP_and_158_cse;
  wire COMP_LOOP_and_160_cse;
  wire COMP_LOOP_and_162_cse;
  wire COMP_LOOP_and_164_cse;
  wire COMP_LOOP_and_166_cse;
  wire COMP_LOOP_and_168_cse;
  wire COMP_LOOP_and_170_cse;
  wire COMP_LOOP_and_172_cse;
  wire COMP_LOOP_and_174_cse;
  wire COMP_LOOP_and_176_cse;
  wire COMP_LOOP_and_178_cse;
  wire COMP_LOOP_and_180_cse;
  wire COMP_LOOP_and_182_cse;
  wire COMP_LOOP_and_184_cse;
  wire COMP_LOOP_and_186_cse;
  wire COMP_LOOP_and_188_cse;
  wire COMP_LOOP_and_190_cse;
  wire COMP_LOOP_and_192_cse;
  wire COMP_LOOP_and_194_cse;
  wire COMP_LOOP_and_196_cse;
  wire COMP_LOOP_and_198_cse;
  wire COMP_LOOP_and_200_cse;
  wire COMP_LOOP_and_202_cse;
  wire COMP_LOOP_and_204_cse;
  wire COMP_LOOP_and_206_cse;
  wire COMP_LOOP_and_208_cse;
  wire COMP_LOOP_and_210_cse;
  wire COMP_LOOP_and_212_cse;
  wire COMP_LOOP_and_214_cse;
  wire COMP_LOOP_and_216_cse;
  wire COMP_LOOP_and_218_cse;
  wire COMP_LOOP_and_220_cse;
  wire COMP_LOOP_and_222_cse;
  wire COMP_LOOP_and_224_cse;
  wire COMP_LOOP_and_226_cse;
  wire COMP_LOOP_and_228_cse;
  wire COMP_LOOP_and_230_cse;
  wire COMP_LOOP_and_232_cse;
  wire COMP_LOOP_and_234_cse;
  wire COMP_LOOP_and_236_cse;
  wire COMP_LOOP_and_238_cse;
  wire COMP_LOOP_and_240_cse;
  wire COMP_LOOP_and_242_cse;
  wire COMP_LOOP_and_244_cse;
  wire COMP_LOOP_and_246_cse;
  wire COMP_LOOP_and_248_cse;
  wire COMP_LOOP_and_250_cse;
  wire COMP_LOOP_and_252_cse;
  wire COMP_LOOP_and_254_cse;
  wire COMP_LOOP_and_256_cse;
  wire COMP_LOOP_and_258_cse;
  wire COMP_LOOP_and_260_cse;
  wire COMP_LOOP_and_262_cse;
  wire COMP_LOOP_and_264_cse;
  wire COMP_LOOP_and_266_cse;
  wire COMP_LOOP_and_268_cse;
  wire COMP_LOOP_and_270_cse;
  wire COMP_LOOP_and_272_cse;
  wire COMP_LOOP_and_274_cse;
  wire COMP_LOOP_and_276_cse;
  wire COMP_LOOP_and_278_cse;
  wire COMP_LOOP_and_280_cse;
  wire COMP_LOOP_and_282_cse;
  wire COMP_LOOP_and_284_cse;
  wire COMP_LOOP_and_286_cse;

  wire[63:0] qelse_acc_nl;
  wire[64:0] nl_qelse_acc_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] mux_7_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] mux_3_nl;
  wire[0:0] mux_2_nl;
  wire[0:0] mux_1_nl;
  wire[0:0] mux_nl;
  wire[0:0] and_273_nl;
  wire[0:0] and_275_nl;
  wire[0:0] and_277_nl;
  wire[0:0] and_279_nl;
  wire[0:0] and_281_nl;
  wire[0:0] and_282_nl;
  wire[0:0] and_283_nl;
  wire[0:0] and_284_nl;
  wire[0:0] and_286_nl;
  wire[0:0] and_287_nl;
  wire[0:0] and_288_nl;
  wire[0:0] and_289_nl;
  wire[0:0] and_290_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_xor_nl;
  wire[0:0] COMP_LOOP_nor_nl;
  wire[0:0] mux_12_nl;
  wire[0:0] nor_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] nor_516_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] nor_515_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] nor_514_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] nor_513_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] nor_511_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] nor_512_nl;
  wire[0:0] nor_508_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] nor_509_nl;
  wire[0:0] mux_21_nl;
  wire[0:0] nor_510_nl;
  wire[0:0] nor_504_nl;
  wire[0:0] nor_505_nl;
  wire[0:0] mux_24_nl;
  wire[0:0] nor_506_nl;
  wire[0:0] mux_25_nl;
  wire[0:0] nor_507_nl;
  wire[0:0] nor_499_nl;
  wire[0:0] or_61_nl;
  wire[0:0] nor_500_nl;
  wire[0:0] nor_501_nl;
  wire[0:0] mux_29_nl;
  wire[0:0] nor_502_nl;
  wire[0:0] mux_30_nl;
  wire[0:0] nor_503_nl;
  wire[0:0] mux_31_nl;
  wire[0:0] nor_498_nl;
  wire[0:0] and_1168_nl;
  wire[0:0] mux_33_nl;
  wire[0:0] nor_497_nl;
  wire[0:0] and_1166_nl;
  wire[0:0] and_1167_nl;
  wire[0:0] mux_36_nl;
  wire[0:0] nor_496_nl;
  wire[0:0] and_1163_nl;
  wire[0:0] and_1164_nl;
  wire[0:0] and_1165_nl;
  wire[0:0] mux_40_nl;
  wire[0:0] nor_495_nl;
  wire[0:0] and_1159_nl;
  wire[0:0] and_1160_nl;
  wire[0:0] and_1161_nl;
  wire[0:0] and_1162_nl;
  wire[0:0] mux_45_nl;
  wire[0:0] nor_494_nl;
  wire[0:0] nor_492_nl;
  wire[0:0] and_1155_nl;
  wire[0:0] and_1156_nl;
  wire[0:0] and_1157_nl;
  wire[0:0] and_1158_nl;
  wire[0:0] mux_51_nl;
  wire[0:0] nor_493_nl;
  wire[0:0] nor_489_nl;
  wire[0:0] nor_490_nl;
  wire[0:0] and_1151_nl;
  wire[0:0] and_1152_nl;
  wire[0:0] and_1153_nl;
  wire[0:0] and_1154_nl;
  wire[0:0] mux_58_nl;
  wire[0:0] nor_491_nl;
  wire[0:0] nor_485_nl;
  wire[0:0] nor_486_nl;
  wire[0:0] nor_487_nl;
  wire[0:0] and_1147_nl;
  wire[0:0] and_1148_nl;
  wire[0:0] and_1149_nl;
  wire[0:0] and_1150_nl;
  wire[0:0] mux_66_nl;
  wire[0:0] nor_488_nl;
  wire[0:0] nor_480_nl;
  wire[0:0] or_165_nl;
  wire[0:0] nor_481_nl;
  wire[0:0] nor_482_nl;
  wire[0:0] nor_483_nl;
  wire[0:0] and_1143_nl;
  wire[0:0] and_1144_nl;
  wire[0:0] and_1145_nl;
  wire[0:0] and_1146_nl;
  wire[0:0] mux_75_nl;
  wire[0:0] nor_484_nl;
  wire[0:0] nor_479_nl;
  wire[0:0] or_175_nl;
  wire[0:0] mux_77_nl;
  wire[0:0] nor_478_nl;
  wire[0:0] mux_78_nl;
  wire[0:0] nor_477_nl;
  wire[0:0] mux_79_nl;
  wire[0:0] nor_476_nl;
  wire[0:0] mux_80_nl;
  wire[0:0] nor_475_nl;
  wire[0:0] mux_81_nl;
  wire[0:0] nor_474_nl;
  wire[0:0] mux_82_nl;
  wire[0:0] nor_472_nl;
  wire[0:0] mux_83_nl;
  wire[0:0] nor_473_nl;
  wire[0:0] nor_469_nl;
  wire[0:0] mux_85_nl;
  wire[0:0] nor_470_nl;
  wire[0:0] mux_86_nl;
  wire[0:0] nor_471_nl;
  wire[0:0] nor_465_nl;
  wire[0:0] nor_466_nl;
  wire[0:0] mux_89_nl;
  wire[0:0] nor_467_nl;
  wire[0:0] mux_90_nl;
  wire[0:0] nor_468_nl;
  wire[0:0] nor_460_nl;
  wire[0:0] or_250_nl;
  wire[0:0] nor_461_nl;
  wire[0:0] nor_462_nl;
  wire[0:0] mux_94_nl;
  wire[0:0] nor_463_nl;
  wire[0:0] mux_95_nl;
  wire[0:0] nor_464_nl;
  wire[0:0] mux_96_nl;
  wire[0:0] nor_459_nl;
  wire[0:0] and_1142_nl;
  wire[0:0] mux_98_nl;
  wire[0:0] nor_458_nl;
  wire[0:0] and_1140_nl;
  wire[0:0] and_1141_nl;
  wire[0:0] mux_101_nl;
  wire[0:0] nor_457_nl;
  wire[0:0] and_1137_nl;
  wire[0:0] and_1138_nl;
  wire[0:0] and_1139_nl;
  wire[0:0] mux_105_nl;
  wire[0:0] nor_456_nl;
  wire[0:0] and_1133_nl;
  wire[0:0] and_1134_nl;
  wire[0:0] and_1135_nl;
  wire[0:0] and_1136_nl;
  wire[0:0] mux_110_nl;
  wire[0:0] nor_455_nl;
  wire[0:0] nor_453_nl;
  wire[0:0] and_1129_nl;
  wire[0:0] and_1130_nl;
  wire[0:0] and_1131_nl;
  wire[0:0] and_1132_nl;
  wire[0:0] mux_116_nl;
  wire[0:0] nor_454_nl;
  wire[0:0] nor_450_nl;
  wire[0:0] nor_451_nl;
  wire[0:0] and_1125_nl;
  wire[0:0] and_1126_nl;
  wire[0:0] and_1127_nl;
  wire[0:0] and_1128_nl;
  wire[0:0] mux_123_nl;
  wire[0:0] nor_452_nl;
  wire[0:0] nor_446_nl;
  wire[0:0] nor_447_nl;
  wire[0:0] nor_448_nl;
  wire[0:0] and_1121_nl;
  wire[0:0] and_1122_nl;
  wire[0:0] and_1123_nl;
  wire[0:0] and_1124_nl;
  wire[0:0] mux_131_nl;
  wire[0:0] nor_449_nl;
  wire[0:0] nor_441_nl;
  wire[0:0] or_352_nl;
  wire[0:0] nor_442_nl;
  wire[0:0] nor_443_nl;
  wire[0:0] nor_444_nl;
  wire[0:0] and_1117_nl;
  wire[0:0] and_1118_nl;
  wire[0:0] and_1119_nl;
  wire[0:0] and_1120_nl;
  wire[0:0] mux_140_nl;
  wire[0:0] nor_445_nl;
  wire[0:0] and_1116_nl;
  wire[0:0] or_362_nl;
  wire[0:0] mux_142_nl;
  wire[0:0] and_1172_nl;
  wire[0:0] mux_143_nl;
  wire[0:0] and_1114_nl;
  wire[0:0] mux_144_nl;
  wire[0:0] and_1113_nl;
  wire[0:0] mux_145_nl;
  wire[0:0] and_1112_nl;
  wire[0:0] mux_146_nl;
  wire[0:0] and_1111_nl;
  wire[0:0] mux_147_nl;
  wire[0:0] and_1109_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] and_1110_nl;
  wire[0:0] and_1106_nl;
  wire[0:0] mux_150_nl;
  wire[0:0] and_1107_nl;
  wire[0:0] mux_151_nl;
  wire[0:0] and_1108_nl;
  wire[0:0] and_1102_nl;
  wire[0:0] and_1103_nl;
  wire[0:0] mux_154_nl;
  wire[0:0] and_1104_nl;
  wire[0:0] mux_155_nl;
  wire[0:0] and_1105_nl;
  wire[0:0] and_1097_nl;
  wire[0:0] or_437_nl;
  wire[0:0] and_1098_nl;
  wire[0:0] and_1099_nl;
  wire[0:0] mux_159_nl;
  wire[0:0] and_1100_nl;
  wire[0:0] mux_160_nl;
  wire[0:0] and_1101_nl;
  wire[0:0] mux_161_nl;
  wire[0:0] and_1171_nl;
  wire[0:0] and_1094_nl;
  wire[0:0] mux_163_nl;
  wire[0:0] and_1095_nl;
  wire[0:0] and_1091_nl;
  wire[0:0] and_1092_nl;
  wire[0:0] mux_166_nl;
  wire[0:0] and_1093_nl;
  wire[0:0] and_1087_nl;
  wire[0:0] and_1088_nl;
  wire[0:0] and_1089_nl;
  wire[0:0] mux_170_nl;
  wire[0:0] and_1090_nl;
  wire[0:0] and_1082_nl;
  wire[0:0] and_1083_nl;
  wire[0:0] and_1084_nl;
  wire[0:0] and_1085_nl;
  wire[0:0] mux_175_nl;
  wire[0:0] and_1086_nl;
  wire[0:0] and_1076_nl;
  wire[0:0] and_1077_nl;
  wire[0:0] and_1078_nl;
  wire[0:0] and_1079_nl;
  wire[0:0] and_1080_nl;
  wire[0:0] mux_181_nl;
  wire[0:0] and_1081_nl;
  wire[0:0] and_1069_nl;
  wire[0:0] and_1070_nl;
  wire[0:0] and_1071_nl;
  wire[0:0] and_1072_nl;
  wire[0:0] and_1073_nl;
  wire[0:0] and_1074_nl;
  wire[0:0] mux_188_nl;
  wire[0:0] and_1075_nl;
  wire[0:0] and_1061_nl;
  wire[0:0] and_1062_nl;
  wire[0:0] and_1063_nl;
  wire[0:0] and_1064_nl;
  wire[0:0] and_1065_nl;
  wire[0:0] and_1066_nl;
  wire[0:0] and_1067_nl;
  wire[0:0] mux_196_nl;
  wire[0:0] and_1068_nl;
  wire[0:0] and_1052_nl;
  wire[0:0] or_540_nl;
  wire[0:0] and_1053_nl;
  wire[0:0] and_1054_nl;
  wire[0:0] and_1055_nl;
  wire[0:0] and_1056_nl;
  wire[0:0] and_1057_nl;
  wire[0:0] and_1058_nl;
  wire[0:0] and_1059_nl;
  wire[0:0] mux_205_nl;
  wire[0:0] and_1060_nl;
  wire[0:0] nor_438_nl;
  wire[0:0] or_550_nl;
  wire[0:0] mux_207_nl;
  wire[0:0] and_1170_nl;
  wire[0:0] mux_208_nl;
  wire[0:0] and_1050_nl;
  wire[0:0] mux_209_nl;
  wire[0:0] and_1049_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] and_1048_nl;
  wire[0:0] mux_211_nl;
  wire[0:0] and_1047_nl;
  wire[0:0] mux_212_nl;
  wire[0:0] and_1045_nl;
  wire[0:0] mux_213_nl;
  wire[0:0] and_1046_nl;
  wire[0:0] and_1042_nl;
  wire[0:0] mux_215_nl;
  wire[0:0] and_1043_nl;
  wire[0:0] mux_216_nl;
  wire[0:0] and_1044_nl;
  wire[0:0] and_1038_nl;
  wire[0:0] and_1039_nl;
  wire[0:0] mux_219_nl;
  wire[0:0] and_1040_nl;
  wire[0:0] mux_220_nl;
  wire[0:0] and_1041_nl;
  wire[0:0] and_1033_nl;
  wire[0:0] or_624_nl;
  wire[0:0] and_1034_nl;
  wire[0:0] and_1035_nl;
  wire[0:0] mux_224_nl;
  wire[0:0] and_1036_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] and_1037_nl;
  wire[0:0] mux_226_nl;
  wire[0:0] and_1169_nl;
  wire[0:0] and_1030_nl;
  wire[0:0] mux_228_nl;
  wire[0:0] and_1031_nl;
  wire[0:0] and_1027_nl;
  wire[0:0] and_1028_nl;
  wire[0:0] mux_231_nl;
  wire[0:0] and_1029_nl;
  wire[0:0] and_1023_nl;
  wire[0:0] and_1024_nl;
  wire[0:0] and_1025_nl;
  wire[0:0] mux_235_nl;
  wire[0:0] and_1026_nl;
  wire[0:0] and_1018_nl;
  wire[0:0] and_1019_nl;
  wire[0:0] and_1020_nl;
  wire[0:0] and_1021_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] and_1022_nl;
  wire[0:0] and_1012_nl;
  wire[0:0] and_1013_nl;
  wire[0:0] and_1014_nl;
  wire[0:0] and_1015_nl;
  wire[0:0] and_1016_nl;
  wire[0:0] mux_246_nl;
  wire[0:0] and_1017_nl;
  wire[0:0] and_1005_nl;
  wire[0:0] and_1006_nl;
  wire[0:0] and_1007_nl;
  wire[0:0] and_1008_nl;
  wire[0:0] and_1009_nl;
  wire[0:0] and_1010_nl;
  wire[0:0] mux_253_nl;
  wire[0:0] and_1011_nl;
  wire[0:0] and_997_nl;
  wire[0:0] and_998_nl;
  wire[0:0] and_999_nl;
  wire[0:0] and_1000_nl;
  wire[0:0] and_1001_nl;
  wire[0:0] and_1002_nl;
  wire[0:0] and_1003_nl;
  wire[0:0] mux_261_nl;
  wire[0:0] and_1004_nl;
  wire[0:0] and_988_nl;
  wire[0:0] or_725_nl;
  wire[0:0] and_989_nl;
  wire[0:0] and_990_nl;
  wire[0:0] and_991_nl;
  wire[0:0] and_992_nl;
  wire[0:0] and_993_nl;
  wire[0:0] and_994_nl;
  wire[0:0] and_995_nl;
  wire[0:0] mux_270_nl;
  wire[0:0] and_996_nl;
  wire[0:0] and_987_nl;
  wire[0:0] or_735_nl;
  wire[0:0] mux_272_nl;
  wire[0:0] nor_435_nl;
  wire[0:0] mux_273_nl;
  wire[0:0] nor_434_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] nor_433_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] nor_432_nl;
  wire[0:0] mux_276_nl;
  wire[0:0] nor_431_nl;
  wire[0:0] mux_277_nl;
  wire[0:0] nor_429_nl;
  wire[0:0] mux_278_nl;
  wire[0:0] nor_430_nl;
  wire[0:0] nor_426_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] nor_427_nl;
  wire[0:0] mux_281_nl;
  wire[0:0] nor_428_nl;
  wire[0:0] nor_422_nl;
  wire[0:0] nor_423_nl;
  wire[0:0] mux_284_nl;
  wire[0:0] nor_424_nl;
  wire[0:0] mux_285_nl;
  wire[0:0] nor_425_nl;
  wire[0:0] nor_417_nl;
  wire[0:0] or_808_nl;
  wire[0:0] nor_418_nl;
  wire[0:0] nor_419_nl;
  wire[0:0] mux_289_nl;
  wire[0:0] nor_420_nl;
  wire[0:0] mux_290_nl;
  wire[0:0] nor_421_nl;
  wire[0:0] nor_408_nl;
  wire[0:0] or_823_nl;
  wire[0:0] nor_409_nl;
  wire[0:0] or_822_nl;
  wire[0:0] nor_410_nl;
  wire[0:0] or_821_nl;
  wire[0:0] nor_411_nl;
  wire[0:0] or_820_nl;
  wire[0:0] nor_412_nl;
  wire[0:0] or_819_nl;
  wire[0:0] nor_413_nl;
  wire[0:0] or_818_nl;
  wire[0:0] nor_414_nl;
  wire[0:0] or_817_nl;
  wire[0:0] nor_415_nl;
  wire[0:0] or_816_nl;
  wire[0:0] mux_299_nl;
  wire[0:0] nor_416_nl;
  wire[0:0] or_815_nl;
  wire[0:0] mux_300_nl;
  wire[0:0] nor_407_nl;
  wire[0:0] and_986_nl;
  wire[0:0] mux_302_nl;
  wire[0:0] nor_406_nl;
  wire[0:0] and_984_nl;
  wire[0:0] and_985_nl;
  wire[0:0] mux_305_nl;
  wire[0:0] nor_405_nl;
  wire[0:0] and_981_nl;
  wire[0:0] and_982_nl;
  wire[0:0] and_983_nl;
  wire[0:0] mux_309_nl;
  wire[0:0] nor_404_nl;
  wire[0:0] and_977_nl;
  wire[0:0] and_978_nl;
  wire[0:0] and_979_nl;
  wire[0:0] and_980_nl;
  wire[0:0] mux_314_nl;
  wire[0:0] nor_403_nl;
  wire[0:0] nor_401_nl;
  wire[0:0] and_973_nl;
  wire[0:0] and_974_nl;
  wire[0:0] and_975_nl;
  wire[0:0] and_976_nl;
  wire[0:0] mux_320_nl;
  wire[0:0] nor_402_nl;
  wire[0:0] nor_398_nl;
  wire[0:0] nor_399_nl;
  wire[0:0] and_969_nl;
  wire[0:0] and_970_nl;
  wire[0:0] and_971_nl;
  wire[0:0] and_972_nl;
  wire[0:0] mux_327_nl;
  wire[0:0] nor_400_nl;
  wire[0:0] nor_394_nl;
  wire[0:0] nor_395_nl;
  wire[0:0] nor_396_nl;
  wire[0:0] and_965_nl;
  wire[0:0] and_966_nl;
  wire[0:0] and_967_nl;
  wire[0:0] and_968_nl;
  wire[0:0] mux_335_nl;
  wire[0:0] nor_397_nl;
  wire[0:0] nor_389_nl;
  wire[0:0] or_919_nl;
  wire[0:0] nor_390_nl;
  wire[0:0] nor_391_nl;
  wire[0:0] nor_392_nl;
  wire[0:0] and_961_nl;
  wire[0:0] and_962_nl;
  wire[0:0] and_963_nl;
  wire[0:0] and_964_nl;
  wire[0:0] mux_344_nl;
  wire[0:0] nor_393_nl;
  wire[0:0] nor_379_nl;
  wire[0:0] or_938_nl;
  wire[0:0] nor_380_nl;
  wire[0:0] or_937_nl;
  wire[0:0] nor_381_nl;
  wire[0:0] or_936_nl;
  wire[0:0] nor_382_nl;
  wire[0:0] or_935_nl;
  wire[0:0] nor_383_nl;
  wire[0:0] or_934_nl;
  wire[0:0] nor_384_nl;
  wire[0:0] or_933_nl;
  wire[0:0] nor_385_nl;
  wire[0:0] or_932_nl;
  wire[0:0] nor_386_nl;
  wire[0:0] or_931_nl;
  wire[0:0] nor_387_nl;
  wire[0:0] or_930_nl;
  wire[0:0] nor_388_nl;
  wire[0:0] or_929_nl;
  wire[0:0] mux_355_nl;
  wire[0:0] nor_378_nl;
  wire[0:0] mux_356_nl;
  wire[0:0] nor_377_nl;
  wire[0:0] mux_357_nl;
  wire[0:0] nor_376_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] nor_375_nl;
  wire[0:0] mux_359_nl;
  wire[0:0] nor_374_nl;
  wire[0:0] mux_360_nl;
  wire[0:0] nor_372_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] nor_373_nl;
  wire[0:0] nor_369_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] nor_370_nl;
  wire[0:0] mux_364_nl;
  wire[0:0] nor_371_nl;
  wire[0:0] nor_365_nl;
  wire[0:0] nor_366_nl;
  wire[0:0] mux_367_nl;
  wire[0:0] nor_367_nl;
  wire[0:0] mux_368_nl;
  wire[0:0] nor_368_nl;
  wire[0:0] nor_360_nl;
  wire[0:0] or_1012_nl;
  wire[0:0] nor_361_nl;
  wire[0:0] nor_362_nl;
  wire[0:0] mux_372_nl;
  wire[0:0] nor_363_nl;
  wire[0:0] mux_373_nl;
  wire[0:0] nor_364_nl;
  wire[0:0] nor_351_nl;
  wire[0:0] or_1027_nl;
  wire[0:0] nor_352_nl;
  wire[0:0] or_1026_nl;
  wire[0:0] nor_353_nl;
  wire[0:0] or_1025_nl;
  wire[0:0] nor_354_nl;
  wire[0:0] or_1024_nl;
  wire[0:0] nor_355_nl;
  wire[0:0] or_1023_nl;
  wire[0:0] nor_356_nl;
  wire[0:0] or_1022_nl;
  wire[0:0] nor_357_nl;
  wire[0:0] or_1021_nl;
  wire[0:0] nor_358_nl;
  wire[0:0] or_1020_nl;
  wire[0:0] mux_382_nl;
  wire[0:0] nor_359_nl;
  wire[0:0] or_1019_nl;
  wire[0:0] mux_383_nl;
  wire[0:0] nor_350_nl;
  wire[0:0] and_960_nl;
  wire[0:0] mux_385_nl;
  wire[0:0] nor_349_nl;
  wire[0:0] and_958_nl;
  wire[0:0] and_959_nl;
  wire[0:0] mux_388_nl;
  wire[0:0] nor_348_nl;
  wire[0:0] and_955_nl;
  wire[0:0] and_956_nl;
  wire[0:0] and_957_nl;
  wire[0:0] mux_392_nl;
  wire[0:0] nor_347_nl;
  wire[0:0] and_951_nl;
  wire[0:0] and_952_nl;
  wire[0:0] and_953_nl;
  wire[0:0] and_954_nl;
  wire[0:0] mux_397_nl;
  wire[0:0] nor_346_nl;
  wire[0:0] nor_344_nl;
  wire[0:0] and_947_nl;
  wire[0:0] and_948_nl;
  wire[0:0] and_949_nl;
  wire[0:0] and_950_nl;
  wire[0:0] mux_403_nl;
  wire[0:0] nor_345_nl;
  wire[0:0] nor_341_nl;
  wire[0:0] nor_342_nl;
  wire[0:0] and_943_nl;
  wire[0:0] and_944_nl;
  wire[0:0] and_945_nl;
  wire[0:0] and_946_nl;
  wire[0:0] mux_410_nl;
  wire[0:0] nor_343_nl;
  wire[0:0] nor_337_nl;
  wire[0:0] nor_338_nl;
  wire[0:0] nor_339_nl;
  wire[0:0] and_939_nl;
  wire[0:0] and_940_nl;
  wire[0:0] and_941_nl;
  wire[0:0] and_942_nl;
  wire[0:0] mux_418_nl;
  wire[0:0] nor_340_nl;
  wire[0:0] nor_332_nl;
  wire[0:0] nand_12_nl;
  wire[0:0] nor_333_nl;
  wire[0:0] nor_334_nl;
  wire[0:0] nor_335_nl;
  wire[0:0] and_935_nl;
  wire[0:0] and_936_nl;
  wire[0:0] and_937_nl;
  wire[0:0] and_938_nl;
  wire[0:0] mux_427_nl;
  wire[0:0] nor_336_nl;
  wire[0:0] nor_323_nl;
  wire[0:0] nand_1_nl;
  wire[0:0] nor_324_nl;
  wire[0:0] nand_2_nl;
  wire[0:0] nor_325_nl;
  wire[0:0] nand_3_nl;
  wire[0:0] nor_326_nl;
  wire[0:0] nand_4_nl;
  wire[0:0] nor_327_nl;
  wire[0:0] nand_5_nl;
  wire[0:0] nor_328_nl;
  wire[0:0] nand_6_nl;
  wire[0:0] nor_329_nl;
  wire[0:0] nand_7_nl;
  wire[0:0] nor_330_nl;
  wire[0:0] nand_8_nl;
  wire[0:0] nor_331_nl;
  wire[0:0] nand_9_nl;
  wire[0:0] and_934_nl;
  wire[0:0] nand_11_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [64:0] nl_rem_12_cmp_a;
  assign nl_rem_12_cmp_a = {{1{rem_12_cmp_a_63_0[63]}}, rem_12_cmp_a_63_0};
  wire [64:0] nl_rem_12_cmp_b;
  assign nl_rem_12_cmp_b = {1'b0 , rem_12_cmp_b_63_0};
  wire [64:0] nl_rem_12_cmp_1_a;
  assign nl_rem_12_cmp_1_a = {{1{rem_12_cmp_1_a_63_0[63]}}, rem_12_cmp_1_a_63_0};
  wire [64:0] nl_rem_12_cmp_1_b;
  assign nl_rem_12_cmp_1_b = {1'b0 , rem_12_cmp_1_b_63_0};
  wire [64:0] nl_rem_12_cmp_2_a;
  assign nl_rem_12_cmp_2_a = {{1{rem_12_cmp_2_a_63_0[63]}}, rem_12_cmp_2_a_63_0};
  wire [64:0] nl_rem_12_cmp_2_b;
  assign nl_rem_12_cmp_2_b = {1'b0 , rem_12_cmp_2_b_63_0};
  wire [64:0] nl_rem_12_cmp_3_a;
  assign nl_rem_12_cmp_3_a = {{1{rem_12_cmp_3_a_63_0[63]}}, rem_12_cmp_3_a_63_0};
  wire [64:0] nl_rem_12_cmp_3_b;
  assign nl_rem_12_cmp_3_b = {1'b0 , rem_12_cmp_3_b_63_0};
  wire [64:0] nl_rem_12_cmp_4_a;
  assign nl_rem_12_cmp_4_a = {{1{rem_12_cmp_4_a_63_0[63]}}, rem_12_cmp_4_a_63_0};
  wire [64:0] nl_rem_12_cmp_4_b;
  assign nl_rem_12_cmp_4_b = {1'b0 , rem_12_cmp_4_b_63_0};
  wire [64:0] nl_rem_12_cmp_5_a;
  assign nl_rem_12_cmp_5_a = {{1{rem_12_cmp_5_a_63_0[63]}}, rem_12_cmp_5_a_63_0};
  wire [64:0] nl_rem_12_cmp_5_b;
  assign nl_rem_12_cmp_5_b = {1'b0 , rem_12_cmp_5_b_63_0};
  wire [64:0] nl_rem_12_cmp_6_a;
  assign nl_rem_12_cmp_6_a = {{1{rem_12_cmp_6_a_63_0[63]}}, rem_12_cmp_6_a_63_0};
  wire [64:0] nl_rem_12_cmp_6_b;
  assign nl_rem_12_cmp_6_b = {1'b0 , rem_12_cmp_6_b_63_0};
  wire [64:0] nl_rem_12_cmp_7_a;
  assign nl_rem_12_cmp_7_a = {{1{rem_12_cmp_7_a_63_0[63]}}, rem_12_cmp_7_a_63_0};
  wire [64:0] nl_rem_12_cmp_7_b;
  assign nl_rem_12_cmp_7_b = {1'b0 , rem_12_cmp_7_b_63_0};
  wire [64:0] nl_rem_12_cmp_8_a;
  assign nl_rem_12_cmp_8_a = {{1{rem_12_cmp_8_a_63_0[63]}}, rem_12_cmp_8_a_63_0};
  wire [64:0] nl_rem_12_cmp_8_b;
  assign nl_rem_12_cmp_8_b = {1'b0 , rem_12_cmp_8_b_63_0};
  wire [64:0] nl_rem_12_cmp_9_a;
  assign nl_rem_12_cmp_9_a = {{1{rem_12_cmp_9_a_63_0[63]}}, rem_12_cmp_9_a_63_0};
  wire [64:0] nl_rem_12_cmp_9_b;
  assign nl_rem_12_cmp_9_b = {1'b0 , rem_12_cmp_9_b_63_0};
  wire [64:0] nl_rem_12_cmp_10_a;
  assign nl_rem_12_cmp_10_a = {{1{rem_12_cmp_10_a_63_0[63]}}, rem_12_cmp_10_a_63_0};
  wire [64:0] nl_rem_12_cmp_10_b;
  assign nl_rem_12_cmp_10_b = {1'b0 , rem_12_cmp_10_b_63_0};
  wire [64:0] nl_rem_12_cmp_11_a;
  assign nl_rem_12_cmp_11_a = {{1{rem_12_cmp_11_a_63_0[63]}}, rem_12_cmp_11_a_63_0};
  wire [64:0] nl_rem_12_cmp_11_b;
  assign nl_rem_12_cmp_11_b = {1'b0 , rem_12_cmp_11_b_63_0};
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd64)) base_rsci (
      .dat(base_rsc_dat),
      .idat(base_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd3),
  .width(32'sd64)) return_rsci (
      .d(return_rsci_d),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd8),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_12_cmp (
      .a(nl_rem_12_cmp_a[64:0]),
      .b(nl_rem_12_cmp_b[64:0]),
      .z(rem_12_cmp_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_12_cmp_1 (
      .a(nl_rem_12_cmp_1_a[64:0]),
      .b(nl_rem_12_cmp_1_b[64:0]),
      .z(rem_12_cmp_1_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_12_cmp_2 (
      .a(nl_rem_12_cmp_2_a[64:0]),
      .b(nl_rem_12_cmp_2_b[64:0]),
      .z(rem_12_cmp_2_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_12_cmp_3 (
      .a(nl_rem_12_cmp_3_a[64:0]),
      .b(nl_rem_12_cmp_3_b[64:0]),
      .z(rem_12_cmp_3_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_12_cmp_4 (
      .a(nl_rem_12_cmp_4_a[64:0]),
      .b(nl_rem_12_cmp_4_b[64:0]),
      .z(rem_12_cmp_4_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_12_cmp_5 (
      .a(nl_rem_12_cmp_5_a[64:0]),
      .b(nl_rem_12_cmp_5_b[64:0]),
      .z(rem_12_cmp_5_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_12_cmp_6 (
      .a(nl_rem_12_cmp_6_a[64:0]),
      .b(nl_rem_12_cmp_6_b[64:0]),
      .z(rem_12_cmp_6_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_12_cmp_7 (
      .a(nl_rem_12_cmp_7_a[64:0]),
      .b(nl_rem_12_cmp_7_b[64:0]),
      .z(rem_12_cmp_7_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_12_cmp_8 (
      .a(nl_rem_12_cmp_8_a[64:0]),
      .b(nl_rem_12_cmp_8_b[64:0]),
      .z(rem_12_cmp_8_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_12_cmp_9 (
      .a(nl_rem_12_cmp_9_a[64:0]),
      .b(nl_rem_12_cmp_9_b[64:0]),
      .z(rem_12_cmp_9_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_12_cmp_10 (
      .a(nl_rem_12_cmp_10_a[64:0]),
      .b(nl_rem_12_cmp_10_b[64:0]),
      .z(rem_12_cmp_10_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_12_cmp_11 (
      .a(nl_rem_12_cmp_11_a[64:0]),
      .b(nl_rem_12_cmp_11_b[64:0]),
      .z(rem_12_cmp_11_z)
    );
  assign COMP_LOOP_and_26_cse = ccs_ccore_en & main_stage_0_12 & COMP_LOOP_asn_itm_11;
  assign COMP_LOOP_and_cse = ccs_ccore_en & (and_dcpl_294 | and_dcpl_300 | and_dcpl_306
      | and_dcpl_312 | and_dcpl_318 | and_dcpl_324 | and_dcpl_330 | and_dcpl_336
      | and_dcpl_342 | and_dcpl_348 | and_tmp_35);
  assign COMP_LOOP_and_2_cse = ccs_ccore_en & (and_dcpl_356 | and_dcpl_360 | and_dcpl_364
      | and_dcpl_368 | and_dcpl_372 | and_dcpl_376 | and_dcpl_379 | and_dcpl_382
      | and_dcpl_385 | and_dcpl_388 | mux_tmp_76);
  assign COMP_LOOP_and_4_cse = ccs_ccore_en & (and_dcpl_394 | and_dcpl_397 | and_dcpl_400
      | and_dcpl_403 | and_dcpl_406 | and_dcpl_409 | and_dcpl_413 | and_dcpl_417
      | and_dcpl_421 | and_dcpl_425 | and_tmp_80);
  assign COMP_LOOP_and_6_cse = ccs_ccore_en & (and_dcpl_431 | and_dcpl_433 | and_dcpl_435
      | and_dcpl_437 | and_dcpl_439 | and_dcpl_442 | and_dcpl_445 | and_dcpl_448
      | and_dcpl_451 | and_dcpl_454 | mux_tmp_141);
  assign COMP_LOOP_and_8_cse = ccs_ccore_en & (and_dcpl_461 | and_dcpl_465 | and_dcpl_469
      | and_dcpl_473 | and_dcpl_477 | and_dcpl_480 | and_dcpl_483 | and_dcpl_486
      | and_dcpl_489 | and_dcpl_492 | and_tmp_125);
  assign COMP_LOOP_and_10_cse = ccs_ccore_en & (and_dcpl_498 | and_dcpl_500 | and_dcpl_502
      | and_dcpl_504 | and_dcpl_506 | and_dcpl_508 | and_dcpl_510 | and_dcpl_512
      | and_dcpl_514 | and_dcpl_516 | mux_tmp_206);
  assign COMP_LOOP_and_12_cse = ccs_ccore_en & (and_dcpl_520 | and_dcpl_523 | and_dcpl_526
      | and_dcpl_529 | and_dcpl_532 | and_dcpl_534 | and_dcpl_536 | and_dcpl_538
      | and_dcpl_540 | and_dcpl_542 | and_tmp_170);
  assign COMP_LOOP_and_14_cse = ccs_ccore_en & (and_dcpl_546 | and_dcpl_548 | and_dcpl_550
      | and_dcpl_552 | and_dcpl_554 | and_dcpl_556 | and_dcpl_558 | and_dcpl_560
      | and_dcpl_562 | and_dcpl_564 | mux_tmp_271);
  assign COMP_LOOP_and_16_cse = ccs_ccore_en & (and_dcpl_569 | and_dcpl_573 | and_dcpl_577
      | and_dcpl_581 | and_dcpl_585 | and_dcpl_589 | and_dcpl_593 | and_dcpl_597
      | and_dcpl_601 | and_dcpl_605 | and_tmp_206);
  assign COMP_LOOP_and_18_cse = ccs_ccore_en & (and_dcpl_610 | and_dcpl_612 | and_dcpl_614
      | and_dcpl_616 | and_dcpl_618 | and_dcpl_622 | and_dcpl_625 | and_dcpl_628
      | and_dcpl_631 | and_dcpl_634 | mux_tmp_354);
  assign COMP_LOOP_and_20_cse = ccs_ccore_en & (and_dcpl_638 | and_dcpl_641 | and_dcpl_644
      | and_dcpl_647 | and_dcpl_650 | and_dcpl_653 | and_dcpl_657 | and_dcpl_661
      | and_dcpl_665 | and_dcpl_669 | and_tmp_233);
  assign COMP_LOOP_and_22_cse = ccs_ccore_en & (and_dcpl_673 | and_dcpl_675 | and_dcpl_677
      | and_dcpl_679 | and_dcpl_681 | and_dcpl_684 | and_dcpl_687 | and_dcpl_690
      | and_dcpl_693 | and_dcpl_696 | mux_tmp_437);
  assign COMP_LOOP_and_28_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_2;
  assign COMP_LOOP_and_30_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_6;
  assign COMP_LOOP_and_32_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_9;
  assign COMP_LOOP_and_34_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_11;
  assign COMP_LOOP_and_36_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_2;
  assign COMP_LOOP_and_38_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_6;
  assign COMP_LOOP_and_40_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_9;
  assign COMP_LOOP_and_42_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_11;
  assign COMP_LOOP_and_44_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_18 & (~ (rem_12cyc_st_10_1_0[0]));
  assign COMP_LOOP_and_46_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_18 & (rem_12cyc_st_10_1_0[0]);
  assign COMP_LOOP_and_48_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_23 & (~ (rem_12cyc_st_10_1_0[0]));
  assign COMP_LOOP_and_50_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_23 & (rem_12cyc_st_10_1_0[0]);
  assign COMP_LOOP_and_52_cse = ccs_ccore_en & and_dcpl_3;
  assign COMP_LOOP_and_54_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_29;
  assign COMP_LOOP_and_56_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_33;
  assign COMP_LOOP_and_58_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_36;
  assign COMP_LOOP_and_60_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_38;
  assign COMP_LOOP_and_62_cse = ccs_ccore_en & and_dcpl_40 & and_dcpl_29;
  assign COMP_LOOP_and_64_cse = ccs_ccore_en & and_dcpl_40 & and_dcpl_33;
  assign COMP_LOOP_and_66_cse = ccs_ccore_en & and_dcpl_40 & and_dcpl_36;
  assign COMP_LOOP_and_68_cse = ccs_ccore_en & and_dcpl_40 & and_dcpl_38;
  assign COMP_LOOP_and_70_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_45 & (~ (rem_12cyc_st_9_1_0[0]));
  assign COMP_LOOP_and_72_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_45 & (rem_12cyc_st_9_1_0[0]);
  assign COMP_LOOP_and_74_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_50 & (~ (rem_12cyc_st_9_1_0[0]));
  assign COMP_LOOP_and_76_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_50 & (rem_12cyc_st_9_1_0[0]);
  assign COMP_LOOP_and_78_cse = ccs_ccore_en & and_dcpl_30;
  assign COMP_LOOP_and_80_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_56;
  assign COMP_LOOP_and_82_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_60;
  assign COMP_LOOP_and_84_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_63;
  assign COMP_LOOP_and_86_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_65;
  assign COMP_LOOP_and_88_cse = ccs_ccore_en & and_dcpl_67 & and_dcpl_56;
  assign COMP_LOOP_and_90_cse = ccs_ccore_en & and_dcpl_67 & and_dcpl_60;
  assign COMP_LOOP_and_92_cse = ccs_ccore_en & and_dcpl_67 & and_dcpl_63;
  assign COMP_LOOP_and_94_cse = ccs_ccore_en & and_dcpl_67 & and_dcpl_65;
  assign COMP_LOOP_and_96_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_72 & (~ (rem_12cyc_st_8_1_0[0]));
  assign COMP_LOOP_and_98_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_72 & (rem_12cyc_st_8_1_0[0]);
  assign COMP_LOOP_and_100_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_77 & (~ (rem_12cyc_st_8_1_0[0]));
  assign COMP_LOOP_and_102_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_77 & (rem_12cyc_st_8_1_0[0]);
  assign COMP_LOOP_and_104_cse = ccs_ccore_en & and_dcpl_57;
  assign COMP_LOOP_and_106_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_83;
  assign COMP_LOOP_and_108_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_87;
  assign COMP_LOOP_and_110_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_90;
  assign COMP_LOOP_and_112_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_92;
  assign COMP_LOOP_and_114_cse = ccs_ccore_en & and_dcpl_94 & and_dcpl_83;
  assign COMP_LOOP_and_116_cse = ccs_ccore_en & and_dcpl_94 & and_dcpl_87;
  assign COMP_LOOP_and_118_cse = ccs_ccore_en & and_dcpl_94 & and_dcpl_90;
  assign COMP_LOOP_and_120_cse = ccs_ccore_en & and_dcpl_94 & and_dcpl_92;
  assign COMP_LOOP_and_122_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_99 & (~ (rem_12cyc_st_7_1_0[0]));
  assign COMP_LOOP_and_124_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_99 & (rem_12cyc_st_7_1_0[0]);
  assign COMP_LOOP_and_126_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_104 & (~ (rem_12cyc_st_7_1_0[0]));
  assign COMP_LOOP_and_128_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_104 & (rem_12cyc_st_7_1_0[0]);
  assign COMP_LOOP_and_130_cse = ccs_ccore_en & and_dcpl_84;
  assign COMP_LOOP_and_132_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_110;
  assign COMP_LOOP_and_134_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_115;
  assign COMP_LOOP_and_136_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_117;
  assign COMP_LOOP_and_138_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_119;
  assign COMP_LOOP_and_140_cse = ccs_ccore_en & and_dcpl_121 & and_dcpl_110;
  assign COMP_LOOP_and_142_cse = ccs_ccore_en & and_dcpl_121 & and_dcpl_115;
  assign COMP_LOOP_and_144_cse = ccs_ccore_en & and_dcpl_121 & and_dcpl_117;
  assign COMP_LOOP_and_146_cse = ccs_ccore_en & and_dcpl_121 & and_dcpl_119;
  assign COMP_LOOP_and_148_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_126 & (~
      (rem_12cyc_st_6_1_0[1]));
  assign COMP_LOOP_and_150_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_129 & (~
      (rem_12cyc_st_6_1_0[1]));
  assign COMP_LOOP_and_152_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_126 & (rem_12cyc_st_6_1_0[1]);
  assign COMP_LOOP_and_154_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_129 & (rem_12cyc_st_6_1_0[1]);
  assign COMP_LOOP_and_156_cse = ccs_ccore_en & and_dcpl_111;
  assign COMP_LOOP_and_158_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_137;
  assign COMP_LOOP_and_160_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_141;
  assign COMP_LOOP_and_162_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_144;
  assign COMP_LOOP_and_164_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_146;
  assign COMP_LOOP_and_166_cse = ccs_ccore_en & and_dcpl_148 & and_dcpl_137;
  assign COMP_LOOP_and_168_cse = ccs_ccore_en & and_dcpl_148 & and_dcpl_141;
  assign COMP_LOOP_and_170_cse = ccs_ccore_en & and_dcpl_148 & and_dcpl_144;
  assign COMP_LOOP_and_172_cse = ccs_ccore_en & and_dcpl_148 & and_dcpl_146;
  assign COMP_LOOP_and_174_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_153 & (~
      (rem_12cyc_st_5_1_0[0]));
  assign COMP_LOOP_and_176_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_153 & (rem_12cyc_st_5_1_0[0]);
  assign COMP_LOOP_and_178_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_158 & (~
      (rem_12cyc_st_5_1_0[0]));
  assign COMP_LOOP_and_180_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_158 & (rem_12cyc_st_5_1_0[0]);
  assign COMP_LOOP_and_182_cse = ccs_ccore_en & and_dcpl_138;
  assign COMP_LOOP_and_184_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_164;
  assign COMP_LOOP_and_186_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_168;
  assign COMP_LOOP_and_188_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_171;
  assign COMP_LOOP_and_190_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_173;
  assign COMP_LOOP_and_192_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_175 & (~
      (rem_12cyc_st_4_1_0[0]));
  assign COMP_LOOP_and_194_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_175 & (rem_12cyc_st_4_1_0[0]);
  assign COMP_LOOP_and_196_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_180 & (~
      (rem_12cyc_st_4_1_0[0]));
  assign COMP_LOOP_and_198_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_180 & (rem_12cyc_st_4_1_0[0]);
  assign COMP_LOOP_and_200_cse = ccs_ccore_en & and_dcpl_185 & and_dcpl_164;
  assign COMP_LOOP_and_202_cse = ccs_ccore_en & and_dcpl_185 & and_dcpl_168;
  assign COMP_LOOP_and_204_cse = ccs_ccore_en & and_dcpl_185 & and_dcpl_171;
  assign COMP_LOOP_and_206_cse = ccs_ccore_en & and_dcpl_185 & and_dcpl_173;
  assign COMP_LOOP_and_208_cse = ccs_ccore_en & and_dcpl_165;
  assign COMP_LOOP_and_210_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_191;
  assign COMP_LOOP_and_212_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_195;
  assign COMP_LOOP_and_214_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_198;
  assign COMP_LOOP_and_216_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_200;
  assign COMP_LOOP_and_218_cse = ccs_ccore_en & and_dcpl_202 & and_dcpl_191;
  assign COMP_LOOP_and_220_cse = ccs_ccore_en & and_dcpl_202 & and_dcpl_195;
  assign COMP_LOOP_and_222_cse = ccs_ccore_en & and_dcpl_202 & and_dcpl_198;
  assign COMP_LOOP_and_224_cse = ccs_ccore_en & and_dcpl_202 & and_dcpl_200;
  assign COMP_LOOP_and_226_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_207 & (~
      (rem_12cyc_st_3_1_0[0]));
  assign COMP_LOOP_and_228_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_207 & (rem_12cyc_st_3_1_0[0]);
  assign COMP_LOOP_and_230_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_212 & (~
      (rem_12cyc_st_3_1_0[0]));
  assign COMP_LOOP_and_232_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_212 & (rem_12cyc_st_3_1_0[0]);
  assign COMP_LOOP_and_234_cse = ccs_ccore_en & and_dcpl_192;
  assign COMP_LOOP_and_236_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_218;
  assign COMP_LOOP_and_238_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_222;
  assign COMP_LOOP_and_240_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_225;
  assign COMP_LOOP_and_242_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_227;
  assign COMP_LOOP_and_244_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_229 & (~
      (rem_12cyc_st_2_1_0[0]));
  assign COMP_LOOP_and_246_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_229 & (rem_12cyc_st_2_1_0[0]);
  assign COMP_LOOP_and_248_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_234 & (~
      (rem_12cyc_st_2_1_0[0]));
  assign COMP_LOOP_and_250_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_234 & (rem_12cyc_st_2_1_0[0]);
  assign COMP_LOOP_and_252_cse = ccs_ccore_en & and_dcpl_239 & and_dcpl_218;
  assign COMP_LOOP_and_254_cse = ccs_ccore_en & and_dcpl_239 & and_dcpl_222;
  assign COMP_LOOP_and_256_cse = ccs_ccore_en & and_dcpl_239 & and_dcpl_225;
  assign COMP_LOOP_and_258_cse = ccs_ccore_en & and_dcpl_239 & and_dcpl_227;
  assign COMP_LOOP_and_260_cse = ccs_ccore_en & and_dcpl_219;
  assign COMP_LOOP_and_262_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_245;
  assign COMP_LOOP_and_264_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_249;
  assign COMP_LOOP_and_266_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_252;
  assign COMP_LOOP_and_268_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_254;
  assign COMP_LOOP_and_270_cse = ccs_ccore_en & and_dcpl_256 & and_dcpl_245;
  assign COMP_LOOP_and_272_cse = ccs_ccore_en & and_dcpl_256 & and_dcpl_249;
  assign COMP_LOOP_and_274_cse = ccs_ccore_en & and_dcpl_256 & and_dcpl_252;
  assign COMP_LOOP_and_276_cse = ccs_ccore_en & and_dcpl_256 & and_dcpl_254;
  assign COMP_LOOP_and_278_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_261 & (~
      (rem_12cyc_1_0[0]));
  assign COMP_LOOP_and_280_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_261 & (rem_12cyc_1_0[0]);
  assign COMP_LOOP_and_282_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_266 & (~
      (rem_12cyc_1_0[0]));
  assign COMP_LOOP_and_284_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_266 & (rem_12cyc_1_0[0]);
  assign COMP_LOOP_and_286_cse = ccs_ccore_en & and_dcpl_246;
  assign COMP_LOOP_and_24_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  assign and_273_nl = and_dcpl_272 & and_dcpl_271;
  assign and_275_nl = and_dcpl_272 & and_dcpl_274;
  assign and_277_nl = and_dcpl_272 & and_dcpl_276;
  assign and_279_nl = and_dcpl_272 & and_dcpl_278;
  assign and_281_nl = and_dcpl_280 & and_dcpl_271;
  assign and_282_nl = and_dcpl_280 & and_dcpl_274;
  assign and_283_nl = and_dcpl_280 & and_dcpl_276;
  assign and_284_nl = and_dcpl_280 & and_dcpl_278;
  assign and_286_nl = and_dcpl_285 & and_dcpl_271;
  assign and_287_nl = and_dcpl_285 & and_dcpl_274;
  assign and_288_nl = and_dcpl_285 & and_dcpl_276;
  assign and_289_nl = and_dcpl_285 & and_dcpl_278;
  assign and_290_nl = (rem_12cyc_st_12_3_2==2'b11);
  assign result_sva_duc_mx0 = MUX1HOT_v_64_13_2((rem_12_cmp_1_z[63:0]), (rem_12_cmp_2_z[63:0]),
      (rem_12_cmp_3_z[63:0]), (rem_12_cmp_4_z[63:0]), (rem_12_cmp_5_z[63:0]), (rem_12_cmp_6_z[63:0]),
      (rem_12_cmp_7_z[63:0]), (rem_12_cmp_8_z[63:0]), (rem_12_cmp_9_z[63:0]), (rem_12_cmp_10_z[63:0]),
      (rem_12_cmp_11_z[63:0]), (rem_12_cmp_z[63:0]), result_sva_duc, {and_273_nl
      , and_275_nl , and_277_nl , and_279_nl , and_281_nl , and_282_nl , and_283_nl
      , and_284_nl , and_286_nl , and_287_nl , and_288_nl , and_289_nl , and_290_nl});
  assign nl_COMP_LOOP_acc_1_tmp = ({rem_12cyc_3_2 , rem_12cyc_1_0}) + 4'b0001;
  assign COMP_LOOP_acc_1_tmp = nl_COMP_LOOP_acc_1_tmp[3:0];
  assign COMP_LOOP_COMP_LOOP_xor_nl = (COMP_LOOP_acc_1_tmp[2]) ^ (COMP_LOOP_acc_1_tmp[3]);
  assign COMP_LOOP_nor_nl = ~((COMP_LOOP_acc_1_tmp[3:2]!=2'b10));
  assign nl_COMP_LOOP_acc_tmp = conv_u2u_1_2(COMP_LOOP_COMP_LOOP_xor_nl) + conv_u2u_1_2(COMP_LOOP_nor_nl);
  assign COMP_LOOP_acc_tmp = nl_COMP_LOOP_acc_tmp[1:0];
  assign and_dcpl_1 = ~((rem_12cyc_st_10_3_2[1]) | (rem_12cyc_st_10_1_0[1]));
  assign and_dcpl_2 = and_dcpl_1 & (~ (rem_12cyc_st_10_1_0[0]));
  assign and_dcpl_3 = main_stage_0_11 & COMP_LOOP_asn_itm_10;
  assign and_dcpl_4 = and_dcpl_3 & (~ (rem_12cyc_st_10_3_2[0]));
  assign and_dcpl_6 = and_dcpl_1 & (rem_12cyc_st_10_1_0[0]);
  assign and_dcpl_8 = (~ (rem_12cyc_st_10_3_2[1])) & (rem_12cyc_st_10_1_0[1]);
  assign and_dcpl_9 = and_dcpl_8 & (~ (rem_12cyc_st_10_1_0[0]));
  assign and_dcpl_11 = and_dcpl_8 & (rem_12cyc_st_10_1_0[0]);
  assign and_dcpl_13 = and_dcpl_3 & (rem_12cyc_st_10_3_2[0]);
  assign and_dcpl_18 = (rem_12cyc_st_10_3_2[1]) & (~ (rem_12cyc_st_10_1_0[1]));
  assign and_dcpl_23 = (rem_12cyc_st_10_3_2[1]) & (rem_12cyc_st_10_1_0[1]);
  assign and_dcpl_28 = ~((rem_12cyc_st_9_3_2[1]) | (rem_12cyc_st_9_1_0[1]));
  assign and_dcpl_29 = and_dcpl_28 & (~ (rem_12cyc_st_9_1_0[0]));
  assign and_dcpl_30 = main_stage_0_10 & COMP_LOOP_asn_itm_9;
  assign and_dcpl_31 = and_dcpl_30 & (~ (rem_12cyc_st_9_3_2[0]));
  assign and_dcpl_33 = and_dcpl_28 & (rem_12cyc_st_9_1_0[0]);
  assign and_dcpl_35 = (~ (rem_12cyc_st_9_3_2[1])) & (rem_12cyc_st_9_1_0[1]);
  assign and_dcpl_36 = and_dcpl_35 & (~ (rem_12cyc_st_9_1_0[0]));
  assign and_dcpl_38 = and_dcpl_35 & (rem_12cyc_st_9_1_0[0]);
  assign and_dcpl_40 = and_dcpl_30 & (rem_12cyc_st_9_3_2[0]);
  assign and_dcpl_45 = (rem_12cyc_st_9_3_2[1]) & (~ (rem_12cyc_st_9_1_0[1]));
  assign and_dcpl_50 = (rem_12cyc_st_9_3_2[1]) & (rem_12cyc_st_9_1_0[1]);
  assign and_dcpl_55 = ~((rem_12cyc_st_8_3_2[1]) | (rem_12cyc_st_8_1_0[1]));
  assign and_dcpl_56 = and_dcpl_55 & (~ (rem_12cyc_st_8_1_0[0]));
  assign and_dcpl_57 = main_stage_0_9 & COMP_LOOP_asn_itm_8;
  assign and_dcpl_58 = and_dcpl_57 & (~ (rem_12cyc_st_8_3_2[0]));
  assign and_dcpl_60 = and_dcpl_55 & (rem_12cyc_st_8_1_0[0]);
  assign and_dcpl_62 = (~ (rem_12cyc_st_8_3_2[1])) & (rem_12cyc_st_8_1_0[1]);
  assign and_dcpl_63 = and_dcpl_62 & (~ (rem_12cyc_st_8_1_0[0]));
  assign and_dcpl_65 = and_dcpl_62 & (rem_12cyc_st_8_1_0[0]);
  assign and_dcpl_67 = and_dcpl_57 & (rem_12cyc_st_8_3_2[0]);
  assign and_dcpl_72 = (rem_12cyc_st_8_3_2[1]) & (~ (rem_12cyc_st_8_1_0[1]));
  assign and_dcpl_77 = (rem_12cyc_st_8_3_2[1]) & (rem_12cyc_st_8_1_0[1]);
  assign and_dcpl_82 = ~((rem_12cyc_st_7_3_2[1]) | (rem_12cyc_st_7_1_0[1]));
  assign and_dcpl_83 = and_dcpl_82 & (~ (rem_12cyc_st_7_1_0[0]));
  assign and_dcpl_84 = main_stage_0_8 & COMP_LOOP_asn_itm_7;
  assign and_dcpl_85 = and_dcpl_84 & (~ (rem_12cyc_st_7_3_2[0]));
  assign and_dcpl_87 = and_dcpl_82 & (rem_12cyc_st_7_1_0[0]);
  assign and_dcpl_89 = (~ (rem_12cyc_st_7_3_2[1])) & (rem_12cyc_st_7_1_0[1]);
  assign and_dcpl_90 = and_dcpl_89 & (~ (rem_12cyc_st_7_1_0[0]));
  assign and_dcpl_92 = and_dcpl_89 & (rem_12cyc_st_7_1_0[0]);
  assign and_dcpl_94 = and_dcpl_84 & (rem_12cyc_st_7_3_2[0]);
  assign and_dcpl_99 = (rem_12cyc_st_7_3_2[1]) & (~ (rem_12cyc_st_7_1_0[1]));
  assign and_dcpl_104 = (rem_12cyc_st_7_3_2[1]) & (rem_12cyc_st_7_1_0[1]);
  assign and_dcpl_109 = ~((rem_12cyc_st_6_3_2[1]) | (rem_12cyc_st_6_1_0[0]));
  assign and_dcpl_110 = and_dcpl_109 & (~ (rem_12cyc_st_6_1_0[1]));
  assign and_dcpl_111 = main_stage_0_7 & COMP_LOOP_asn_itm_6;
  assign and_dcpl_112 = and_dcpl_111 & (~ (rem_12cyc_st_6_3_2[0]));
  assign and_dcpl_114 = (~ (rem_12cyc_st_6_3_2[1])) & (rem_12cyc_st_6_1_0[0]);
  assign and_dcpl_115 = and_dcpl_114 & (~ (rem_12cyc_st_6_1_0[1]));
  assign and_dcpl_117 = and_dcpl_109 & (rem_12cyc_st_6_1_0[1]);
  assign and_dcpl_119 = and_dcpl_114 & (rem_12cyc_st_6_1_0[1]);
  assign and_dcpl_121 = and_dcpl_111 & (rem_12cyc_st_6_3_2[0]);
  assign and_dcpl_126 = (rem_12cyc_st_6_3_2[1]) & (~ (rem_12cyc_st_6_1_0[0]));
  assign and_dcpl_129 = (rem_12cyc_st_6_3_2[1]) & (rem_12cyc_st_6_1_0[0]);
  assign and_dcpl_136 = ~((rem_12cyc_st_5_3_2[1]) | (rem_12cyc_st_5_1_0[1]));
  assign and_dcpl_137 = and_dcpl_136 & (~ (rem_12cyc_st_5_1_0[0]));
  assign and_dcpl_138 = main_stage_0_6 & COMP_LOOP_asn_itm_5;
  assign and_dcpl_139 = and_dcpl_138 & (~ (rem_12cyc_st_5_3_2[0]));
  assign and_dcpl_141 = and_dcpl_136 & (rem_12cyc_st_5_1_0[0]);
  assign and_dcpl_143 = (~ (rem_12cyc_st_5_3_2[1])) & (rem_12cyc_st_5_1_0[1]);
  assign and_dcpl_144 = and_dcpl_143 & (~ (rem_12cyc_st_5_1_0[0]));
  assign and_dcpl_146 = and_dcpl_143 & (rem_12cyc_st_5_1_0[0]);
  assign and_dcpl_148 = and_dcpl_138 & (rem_12cyc_st_5_3_2[0]);
  assign and_dcpl_153 = (rem_12cyc_st_5_3_2[1]) & (~ (rem_12cyc_st_5_1_0[1]));
  assign and_dcpl_158 = (rem_12cyc_st_5_3_2[1]) & (rem_12cyc_st_5_1_0[1]);
  assign and_dcpl_163 = ~((rem_12cyc_st_4_3_2[0]) | (rem_12cyc_st_4_1_0[1]));
  assign and_dcpl_164 = and_dcpl_163 & (~ (rem_12cyc_st_4_1_0[0]));
  assign and_dcpl_165 = main_stage_0_5 & COMP_LOOP_asn_itm_4;
  assign and_dcpl_166 = and_dcpl_165 & (~ (rem_12cyc_st_4_3_2[1]));
  assign and_dcpl_168 = and_dcpl_163 & (rem_12cyc_st_4_1_0[0]);
  assign and_dcpl_170 = (~ (rem_12cyc_st_4_3_2[0])) & (rem_12cyc_st_4_1_0[1]);
  assign and_dcpl_171 = and_dcpl_170 & (~ (rem_12cyc_st_4_1_0[0]));
  assign and_dcpl_173 = and_dcpl_170 & (rem_12cyc_st_4_1_0[0]);
  assign and_dcpl_175 = (rem_12cyc_st_4_3_2[0]) & (~ (rem_12cyc_st_4_1_0[1]));
  assign and_dcpl_180 = (rem_12cyc_st_4_3_2[0]) & (rem_12cyc_st_4_1_0[1]);
  assign and_dcpl_185 = and_dcpl_165 & (rem_12cyc_st_4_3_2[1]);
  assign and_dcpl_190 = ~((rem_12cyc_st_3_3_2[1]) | (rem_12cyc_st_3_1_0[1]));
  assign and_dcpl_191 = and_dcpl_190 & (~ (rem_12cyc_st_3_1_0[0]));
  assign and_dcpl_192 = main_stage_0_4 & COMP_LOOP_asn_itm_3;
  assign and_dcpl_193 = and_dcpl_192 & (~ (rem_12cyc_st_3_3_2[0]));
  assign and_dcpl_195 = and_dcpl_190 & (rem_12cyc_st_3_1_0[0]);
  assign and_dcpl_197 = (~ (rem_12cyc_st_3_3_2[1])) & (rem_12cyc_st_3_1_0[1]);
  assign and_dcpl_198 = and_dcpl_197 & (~ (rem_12cyc_st_3_1_0[0]));
  assign and_dcpl_200 = and_dcpl_197 & (rem_12cyc_st_3_1_0[0]);
  assign and_dcpl_202 = and_dcpl_192 & (rem_12cyc_st_3_3_2[0]);
  assign and_dcpl_207 = (rem_12cyc_st_3_3_2[1]) & (~ (rem_12cyc_st_3_1_0[1]));
  assign and_dcpl_212 = (rem_12cyc_st_3_3_2[1]) & (rem_12cyc_st_3_1_0[1]);
  assign and_dcpl_217 = ~((rem_12cyc_st_2_3_2[0]) | (rem_12cyc_st_2_1_0[1]));
  assign and_dcpl_218 = and_dcpl_217 & (~ (rem_12cyc_st_2_1_0[0]));
  assign and_dcpl_219 = main_stage_0_3 & COMP_LOOP_asn_itm_2;
  assign and_dcpl_220 = and_dcpl_219 & (~ (rem_12cyc_st_2_3_2[1]));
  assign and_dcpl_222 = and_dcpl_217 & (rem_12cyc_st_2_1_0[0]);
  assign and_dcpl_224 = (~ (rem_12cyc_st_2_3_2[0])) & (rem_12cyc_st_2_1_0[1]);
  assign and_dcpl_225 = and_dcpl_224 & (~ (rem_12cyc_st_2_1_0[0]));
  assign and_dcpl_227 = and_dcpl_224 & (rem_12cyc_st_2_1_0[0]);
  assign and_dcpl_229 = (rem_12cyc_st_2_3_2[0]) & (~ (rem_12cyc_st_2_1_0[1]));
  assign and_dcpl_234 = (rem_12cyc_st_2_3_2[0]) & (rem_12cyc_st_2_1_0[1]);
  assign and_dcpl_239 = and_dcpl_219 & (rem_12cyc_st_2_3_2[1]);
  assign and_dcpl_244 = ~((rem_12cyc_3_2[1]) | (rem_12cyc_1_0[1]));
  assign and_dcpl_245 = and_dcpl_244 & (~ (rem_12cyc_1_0[0]));
  assign and_dcpl_246 = main_stage_0_2 & COMP_LOOP_asn_itm_1;
  assign and_dcpl_247 = and_dcpl_246 & (~ (rem_12cyc_3_2[0]));
  assign and_dcpl_249 = and_dcpl_244 & (rem_12cyc_1_0[0]);
  assign and_dcpl_251 = (~ (rem_12cyc_3_2[1])) & (rem_12cyc_1_0[1]);
  assign and_dcpl_252 = and_dcpl_251 & (~ (rem_12cyc_1_0[0]));
  assign and_dcpl_254 = and_dcpl_251 & (rem_12cyc_1_0[0]);
  assign and_dcpl_256 = and_dcpl_246 & (rem_12cyc_3_2[0]);
  assign and_dcpl_261 = (rem_12cyc_3_2[1]) & (~ (rem_12cyc_1_0[1]));
  assign and_dcpl_266 = (rem_12cyc_3_2[1]) & (rem_12cyc_1_0[1]);
  assign and_dcpl_271 = ~((rem_12cyc_st_12_1_0!=2'b00));
  assign and_dcpl_272 = ~((rem_12cyc_st_12_3_2!=2'b00));
  assign and_dcpl_274 = (rem_12cyc_st_12_1_0==2'b01);
  assign and_dcpl_276 = (rem_12cyc_st_12_1_0==2'b10);
  assign and_dcpl_278 = (rem_12cyc_st_12_1_0==2'b11);
  assign and_dcpl_280 = (rem_12cyc_st_12_3_2==2'b01);
  assign and_dcpl_285 = (rem_12cyc_st_12_3_2==2'b10);
  assign and_dcpl_291 = ~((COMP_LOOP_acc_1_tmp[1:0]!=2'b00));
  assign and_dcpl_292 = ccs_ccore_start_rsci_idat & (~ (COMP_LOOP_acc_tmp[0]));
  assign and_dcpl_293 = and_dcpl_292 & (~ (COMP_LOOP_acc_tmp[1]));
  assign and_dcpl_294 = and_dcpl_293 & and_dcpl_291;
  assign and_dcpl_295 = ~((rem_12cyc_st_2_3_2!=2'b00));
  assign and_dcpl_296 = and_dcpl_295 & (~ (rem_12cyc_st_2_1_0[1]));
  assign and_dcpl_298 = (~ (rem_12cyc_st_2_1_0[0])) & main_stage_0_3 & COMP_LOOP_asn_itm_2;
  assign not_tmp_54 = ~(COMP_LOOP_asn_itm_1 & main_stage_0_2);
  assign or_tmp_2 = (rem_12cyc_1_0!=2'b00) | (rem_12cyc_3_2!=2'b00) | not_tmp_54;
  assign or_1_cse = (COMP_LOOP_acc_1_tmp[1:0]!=2'b00) | (COMP_LOOP_acc_tmp!=2'b00);
  assign nor_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_2));
  assign mux_12_nl = MUX_s_1_2_2(nor_nl, or_tmp_2, or_1_cse);
  assign and_dcpl_300 = mux_12_nl & and_dcpl_298 & and_dcpl_296;
  assign and_dcpl_301 = ~((rem_12cyc_st_3_3_2!=2'b00));
  assign and_dcpl_302 = and_dcpl_301 & (~ (rem_12cyc_st_3_1_0[1]));
  assign and_dcpl_304 = (~ (rem_12cyc_st_3_1_0[0])) & main_stage_0_4 & COMP_LOOP_asn_itm_3;
  assign or_6_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2!=2'b00) | (~ COMP_LOOP_asn_itm_2)
      | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp = or_6_cse & or_tmp_2;
  assign nor_516_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp));
  assign mux_13_nl = MUX_s_1_2_2(nor_516_nl, and_tmp, or_1_cse);
  assign and_dcpl_306 = mux_13_nl & and_dcpl_304 & and_dcpl_302;
  assign and_dcpl_307 = ~((rem_12cyc_st_4_3_2!=2'b00));
  assign and_dcpl_308 = and_dcpl_307 & (~ (rem_12cyc_st_4_1_0[1]));
  assign and_dcpl_310 = (~ (rem_12cyc_st_4_1_0[0])) & main_stage_0_5 & COMP_LOOP_asn_itm_4;
  assign or_10_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2!=2'b00) | (~ COMP_LOOP_asn_itm_3)
      | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_2 = or_6_cse & or_10_cse & or_tmp_2;
  assign nor_515_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_2));
  assign mux_14_nl = MUX_s_1_2_2(nor_515_nl, and_tmp_2, or_1_cse);
  assign and_dcpl_312 = mux_14_nl & and_dcpl_310 & and_dcpl_308;
  assign and_dcpl_313 = ~((rem_12cyc_st_5_3_2!=2'b00));
  assign and_dcpl_314 = and_dcpl_313 & (~ (rem_12cyc_st_5_1_0[1]));
  assign and_dcpl_316 = (~ (rem_12cyc_st_5_1_0[0])) & main_stage_0_6 & COMP_LOOP_asn_itm_5;
  assign or_15_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2!=2'b00) | (~ COMP_LOOP_asn_itm_4)
      | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_5 = or_6_cse & or_10_cse & or_15_cse & or_tmp_2;
  assign nor_514_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_5));
  assign mux_15_nl = MUX_s_1_2_2(nor_514_nl, and_tmp_5, or_1_cse);
  assign and_dcpl_318 = mux_15_nl & and_dcpl_316 & and_dcpl_314;
  assign or_21_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2!=2'b00) | (~ COMP_LOOP_asn_itm_5)
      | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_9 = or_6_cse & or_10_cse & or_15_cse & or_21_cse & or_tmp_2;
  assign nor_513_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_9));
  assign mux_16_nl = MUX_s_1_2_2(nor_513_nl, and_tmp_9, or_1_cse);
  assign and_dcpl_324 = mux_16_nl & and_dcpl_112 & and_dcpl_110;
  assign or_28_cse = (rem_12cyc_st_6_1_0!=2'b00) | (rem_12cyc_st_6_3_2!=2'b00);
  assign nor_511_nl = ~(and_dcpl_111 | (~ or_tmp_2));
  assign mux_17_nl = MUX_s_1_2_2(nor_511_nl, or_tmp_2, or_28_cse);
  assign and_tmp_13 = or_6_cse & or_10_cse & or_15_cse & or_21_cse & mux_17_nl;
  assign nor_512_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_13));
  assign mux_18_nl = MUX_s_1_2_2(nor_512_nl, and_tmp_13, or_1_cse);
  assign and_dcpl_330 = mux_18_nl & and_dcpl_85 & and_dcpl_83;
  assign or_37_cse = (rem_12cyc_st_7_1_0!=2'b00) | (rem_12cyc_st_7_3_2!=2'b00);
  assign nor_508_nl = ~(and_dcpl_84 | (~ or_tmp_2));
  assign mux_tmp_19 = MUX_s_1_2_2(nor_508_nl, or_tmp_2, or_37_cse);
  assign nor_509_nl = ~(and_dcpl_111 | (~ mux_tmp_19));
  assign mux_20_nl = MUX_s_1_2_2(nor_509_nl, mux_tmp_19, or_28_cse);
  assign and_tmp_17 = or_6_cse & or_10_cse & or_15_cse & or_21_cse & mux_20_nl;
  assign nor_510_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_17));
  assign mux_21_nl = MUX_s_1_2_2(nor_510_nl, and_tmp_17, or_1_cse);
  assign and_dcpl_336 = mux_21_nl & and_dcpl_58 & and_dcpl_56;
  assign or_48_cse = (rem_12cyc_st_8_1_0!=2'b00) | (rem_12cyc_st_8_3_2!=2'b00);
  assign nor_504_nl = ~(and_dcpl_57 | (~ or_tmp_2));
  assign mux_tmp_22 = MUX_s_1_2_2(nor_504_nl, or_tmp_2, or_48_cse);
  assign nor_505_nl = ~(and_dcpl_84 | (~ mux_tmp_22));
  assign mux_tmp_23 = MUX_s_1_2_2(nor_505_nl, mux_tmp_22, or_37_cse);
  assign nor_506_nl = ~(and_dcpl_111 | (~ mux_tmp_23));
  assign mux_24_nl = MUX_s_1_2_2(nor_506_nl, mux_tmp_23, or_28_cse);
  assign and_tmp_21 = or_6_cse & or_10_cse & or_15_cse & or_21_cse & mux_24_nl;
  assign nor_507_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_21));
  assign mux_25_nl = MUX_s_1_2_2(nor_507_nl, and_tmp_21, or_1_cse);
  assign and_dcpl_342 = mux_25_nl & and_dcpl_31 & and_dcpl_29;
  assign nor_499_nl = ~(and_dcpl_30 | (~ or_tmp_2));
  assign or_61_nl = (rem_12cyc_st_9_1_0!=2'b00) | (rem_12cyc_st_9_3_2!=2'b00);
  assign mux_tmp_26 = MUX_s_1_2_2(nor_499_nl, or_tmp_2, or_61_nl);
  assign nor_500_nl = ~(and_dcpl_57 | (~ mux_tmp_26));
  assign mux_tmp_27 = MUX_s_1_2_2(nor_500_nl, mux_tmp_26, or_48_cse);
  assign nor_501_nl = ~(and_dcpl_84 | (~ mux_tmp_27));
  assign mux_tmp_28 = MUX_s_1_2_2(nor_501_nl, mux_tmp_27, or_37_cse);
  assign nor_502_nl = ~(and_dcpl_111 | (~ mux_tmp_28));
  assign mux_29_nl = MUX_s_1_2_2(nor_502_nl, mux_tmp_28, or_28_cse);
  assign and_tmp_25 = or_6_cse & or_10_cse & or_15_cse & or_21_cse & mux_29_nl;
  assign nor_503_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_25));
  assign mux_30_nl = MUX_s_1_2_2(nor_503_nl, and_tmp_25, or_1_cse);
  assign and_dcpl_348 = mux_30_nl & and_dcpl_4 & and_dcpl_2;
  assign and_tmp_35 = ((~ main_stage_0_2) | (~ COMP_LOOP_asn_itm_1) | (rem_12cyc_3_2!=2'b00)
      | (rem_12cyc_1_0!=2'b00)) & ((~ main_stage_0_8) | (~ COMP_LOOP_asn_itm_7) |
      (rem_12cyc_st_7_1_0!=2'b00) | (rem_12cyc_st_7_3_2!=2'b00)) & ((~ main_stage_0_9)
      | (~ COMP_LOOP_asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b00) | (rem_12cyc_st_8_3_2!=2'b00))
      & ((~ main_stage_0_10) | (~ COMP_LOOP_asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b00)
      | (rem_12cyc_st_9_3_2!=2'b00)) & or_6_cse & or_10_cse & or_15_cse & or_21_cse
      & ((~ main_stage_0_7) | (~ COMP_LOOP_asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b00)
      | (rem_12cyc_st_6_3_2!=2'b00)) & ((~ main_stage_0_11) | (~ COMP_LOOP_asn_itm_10)
      | (rem_12cyc_st_10_1_0!=2'b00) | (rem_12cyc_st_10_3_2!=2'b00)) & ((COMP_LOOP_acc_tmp!=2'b00)
      | (COMP_LOOP_acc_1_tmp[1:0]!=2'b00) | (~ ccs_ccore_start_rsci_idat));
  assign and_dcpl_355 = (COMP_LOOP_acc_1_tmp[1:0]==2'b01);
  assign and_dcpl_356 = and_dcpl_293 & and_dcpl_355;
  assign and_dcpl_358 = (rem_12cyc_st_2_1_0[0]) & main_stage_0_3 & COMP_LOOP_asn_itm_2;
  assign or_tmp_80 = (rem_12cyc_1_0!=2'b01) | (rem_12cyc_3_2!=2'b00) | not_tmp_54;
  assign or_83_cse = (COMP_LOOP_acc_1_tmp[1:0]!=2'b01) | (COMP_LOOP_acc_tmp!=2'b00);
  assign nor_498_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_80));
  assign mux_31_nl = MUX_s_1_2_2(nor_498_nl, or_tmp_80, or_83_cse);
  assign and_dcpl_360 = mux_31_nl & and_dcpl_358 & and_dcpl_296;
  assign and_dcpl_362 = (rem_12cyc_st_3_1_0[0]) & main_stage_0_4 & COMP_LOOP_asn_itm_3;
  assign nand_276_cse = ~(COMP_LOOP_asn_itm_2 & main_stage_0_3 & (rem_12cyc_st_2_1_0[0]));
  assign or_88_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2!=2'b00);
  assign and_1168_nl = nand_276_cse & or_tmp_80;
  assign mux_tmp_32 = MUX_s_1_2_2(and_1168_nl, or_tmp_80, or_88_cse);
  assign nor_497_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_32));
  assign mux_33_nl = MUX_s_1_2_2(nor_497_nl, mux_tmp_32, or_83_cse);
  assign and_dcpl_364 = mux_33_nl & and_dcpl_362 & and_dcpl_302;
  assign and_dcpl_366 = (rem_12cyc_st_4_1_0[0]) & main_stage_0_5 & COMP_LOOP_asn_itm_4;
  assign nand_274_cse = ~(COMP_LOOP_asn_itm_3 & main_stage_0_4 & (rem_12cyc_st_3_1_0[0]));
  assign or_93_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2!=2'b00);
  assign and_1166_nl = nand_274_cse & or_tmp_80;
  assign mux_tmp_34 = MUX_s_1_2_2(and_1166_nl, or_tmp_80, or_93_cse);
  assign and_1167_nl = nand_276_cse & mux_tmp_34;
  assign mux_tmp_35 = MUX_s_1_2_2(and_1167_nl, mux_tmp_34, or_88_cse);
  assign nor_496_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_35));
  assign mux_36_nl = MUX_s_1_2_2(nor_496_nl, mux_tmp_35, or_83_cse);
  assign and_dcpl_368 = mux_36_nl & and_dcpl_366 & and_dcpl_308;
  assign and_dcpl_370 = (rem_12cyc_st_5_1_0[0]) & main_stage_0_6 & COMP_LOOP_asn_itm_5;
  assign nand_271_cse = ~(COMP_LOOP_asn_itm_4 & main_stage_0_5 & (rem_12cyc_st_4_1_0[0]));
  assign or_100_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2!=2'b00);
  assign and_1163_nl = nand_271_cse & or_tmp_80;
  assign mux_tmp_37 = MUX_s_1_2_2(and_1163_nl, or_tmp_80, or_100_cse);
  assign and_1164_nl = nand_274_cse & mux_tmp_37;
  assign mux_tmp_38 = MUX_s_1_2_2(and_1164_nl, mux_tmp_37, or_93_cse);
  assign and_1165_nl = nand_276_cse & mux_tmp_38;
  assign mux_tmp_39 = MUX_s_1_2_2(and_1165_nl, mux_tmp_38, or_88_cse);
  assign nor_495_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_39));
  assign mux_40_nl = MUX_s_1_2_2(nor_495_nl, mux_tmp_39, or_83_cse);
  assign and_dcpl_372 = mux_40_nl & and_dcpl_370 & and_dcpl_314;
  assign nand_267_cse = ~(COMP_LOOP_asn_itm_5 & main_stage_0_6 & (rem_12cyc_st_5_1_0[0]));
  assign or_109_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2!=2'b00);
  assign and_1159_nl = nand_267_cse & or_tmp_80;
  assign mux_tmp_41 = MUX_s_1_2_2(and_1159_nl, or_tmp_80, or_109_cse);
  assign and_1160_nl = nand_271_cse & mux_tmp_41;
  assign mux_tmp_42 = MUX_s_1_2_2(and_1160_nl, mux_tmp_41, or_100_cse);
  assign and_1161_nl = nand_274_cse & mux_tmp_42;
  assign mux_tmp_43 = MUX_s_1_2_2(and_1161_nl, mux_tmp_42, or_93_cse);
  assign and_1162_nl = nand_276_cse & mux_tmp_43;
  assign mux_tmp_44 = MUX_s_1_2_2(and_1162_nl, mux_tmp_43, or_88_cse);
  assign nor_494_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_44));
  assign mux_45_nl = MUX_s_1_2_2(nor_494_nl, mux_tmp_44, or_83_cse);
  assign and_dcpl_376 = mux_45_nl & and_dcpl_112 & and_dcpl_115;
  assign or_120_cse = (rem_12cyc_st_6_1_0!=2'b01) | (rem_12cyc_st_6_3_2!=2'b00);
  assign nor_492_nl = ~(and_dcpl_111 | (~ or_tmp_80));
  assign mux_tmp_46 = MUX_s_1_2_2(nor_492_nl, or_tmp_80, or_120_cse);
  assign and_1155_nl = nand_267_cse & mux_tmp_46;
  assign mux_tmp_47 = MUX_s_1_2_2(and_1155_nl, mux_tmp_46, or_109_cse);
  assign and_1156_nl = nand_271_cse & mux_tmp_47;
  assign mux_tmp_48 = MUX_s_1_2_2(and_1156_nl, mux_tmp_47, or_100_cse);
  assign and_1157_nl = nand_274_cse & mux_tmp_48;
  assign mux_tmp_49 = MUX_s_1_2_2(and_1157_nl, mux_tmp_48, or_93_cse);
  assign and_1158_nl = nand_276_cse & mux_tmp_49;
  assign mux_tmp_50 = MUX_s_1_2_2(and_1158_nl, mux_tmp_49, or_88_cse);
  assign nor_493_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_50));
  assign mux_51_nl = MUX_s_1_2_2(nor_493_nl, mux_tmp_50, or_83_cse);
  assign and_dcpl_379 = mux_51_nl & and_dcpl_85 & and_dcpl_87;
  assign or_133_cse = (rem_12cyc_st_7_1_0!=2'b01) | (rem_12cyc_st_7_3_2!=2'b00);
  assign nor_489_nl = ~(and_dcpl_84 | (~ or_tmp_80));
  assign mux_tmp_52 = MUX_s_1_2_2(nor_489_nl, or_tmp_80, or_133_cse);
  assign nor_490_nl = ~(and_dcpl_111 | (~ mux_tmp_52));
  assign mux_tmp_53 = MUX_s_1_2_2(nor_490_nl, mux_tmp_52, or_120_cse);
  assign and_1151_nl = nand_267_cse & mux_tmp_53;
  assign mux_tmp_54 = MUX_s_1_2_2(and_1151_nl, mux_tmp_53, or_109_cse);
  assign and_1152_nl = nand_271_cse & mux_tmp_54;
  assign mux_tmp_55 = MUX_s_1_2_2(and_1152_nl, mux_tmp_54, or_100_cse);
  assign and_1153_nl = nand_274_cse & mux_tmp_55;
  assign mux_tmp_56 = MUX_s_1_2_2(and_1153_nl, mux_tmp_55, or_93_cse);
  assign and_1154_nl = nand_276_cse & mux_tmp_56;
  assign mux_tmp_57 = MUX_s_1_2_2(and_1154_nl, mux_tmp_56, or_88_cse);
  assign nor_491_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_57));
  assign mux_58_nl = MUX_s_1_2_2(nor_491_nl, mux_tmp_57, or_83_cse);
  assign and_dcpl_382 = mux_58_nl & and_dcpl_58 & and_dcpl_60;
  assign or_148_cse = (rem_12cyc_st_8_1_0!=2'b01) | (rem_12cyc_st_8_3_2!=2'b00);
  assign nor_485_nl = ~(and_dcpl_57 | (~ or_tmp_80));
  assign mux_tmp_59 = MUX_s_1_2_2(nor_485_nl, or_tmp_80, or_148_cse);
  assign nor_486_nl = ~(and_dcpl_84 | (~ mux_tmp_59));
  assign mux_tmp_60 = MUX_s_1_2_2(nor_486_nl, mux_tmp_59, or_133_cse);
  assign nor_487_nl = ~(and_dcpl_111 | (~ mux_tmp_60));
  assign mux_tmp_61 = MUX_s_1_2_2(nor_487_nl, mux_tmp_60, or_120_cse);
  assign and_1147_nl = nand_267_cse & mux_tmp_61;
  assign mux_tmp_62 = MUX_s_1_2_2(and_1147_nl, mux_tmp_61, or_109_cse);
  assign and_1148_nl = nand_271_cse & mux_tmp_62;
  assign mux_tmp_63 = MUX_s_1_2_2(and_1148_nl, mux_tmp_62, or_100_cse);
  assign and_1149_nl = nand_274_cse & mux_tmp_63;
  assign mux_tmp_64 = MUX_s_1_2_2(and_1149_nl, mux_tmp_63, or_93_cse);
  assign and_1150_nl = nand_276_cse & mux_tmp_64;
  assign mux_tmp_65 = MUX_s_1_2_2(and_1150_nl, mux_tmp_64, or_88_cse);
  assign nor_488_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_65));
  assign mux_66_nl = MUX_s_1_2_2(nor_488_nl, mux_tmp_65, or_83_cse);
  assign and_dcpl_385 = mux_66_nl & and_dcpl_31 & and_dcpl_33;
  assign nor_480_nl = ~(and_dcpl_30 | (~ or_tmp_80));
  assign or_165_nl = (rem_12cyc_st_9_1_0!=2'b01) | (rem_12cyc_st_9_3_2!=2'b00);
  assign mux_tmp_67 = MUX_s_1_2_2(nor_480_nl, or_tmp_80, or_165_nl);
  assign nor_481_nl = ~(and_dcpl_57 | (~ mux_tmp_67));
  assign mux_tmp_68 = MUX_s_1_2_2(nor_481_nl, mux_tmp_67, or_148_cse);
  assign nor_482_nl = ~(and_dcpl_84 | (~ mux_tmp_68));
  assign mux_tmp_69 = MUX_s_1_2_2(nor_482_nl, mux_tmp_68, or_133_cse);
  assign nor_483_nl = ~(and_dcpl_111 | (~ mux_tmp_69));
  assign mux_tmp_70 = MUX_s_1_2_2(nor_483_nl, mux_tmp_69, or_120_cse);
  assign and_1143_nl = nand_267_cse & mux_tmp_70;
  assign mux_tmp_71 = MUX_s_1_2_2(and_1143_nl, mux_tmp_70, or_109_cse);
  assign and_1144_nl = nand_271_cse & mux_tmp_71;
  assign mux_tmp_72 = MUX_s_1_2_2(and_1144_nl, mux_tmp_71, or_100_cse);
  assign and_1145_nl = nand_274_cse & mux_tmp_72;
  assign mux_tmp_73 = MUX_s_1_2_2(and_1145_nl, mux_tmp_72, or_93_cse);
  assign and_1146_nl = nand_276_cse & mux_tmp_73;
  assign mux_tmp_74 = MUX_s_1_2_2(and_1146_nl, mux_tmp_73, or_88_cse);
  assign nor_484_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_74));
  assign mux_75_nl = MUX_s_1_2_2(nor_484_nl, mux_tmp_74, or_83_cse);
  assign and_dcpl_388 = mux_75_nl & and_dcpl_4 & and_dcpl_6;
  assign nand_250_cse = ~((COMP_LOOP_acc_1_tmp[0]) & ccs_ccore_start_rsci_idat);
  assign and_tmp_44 = ((~ main_stage_0_8) | (~ COMP_LOOP_asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b01)
      | (rem_12cyc_st_7_3_2!=2'b00)) & ((~ main_stage_0_9) | (~ COMP_LOOP_asn_itm_8)
      | (rem_12cyc_st_8_1_0!=2'b01) | (rem_12cyc_st_8_3_2!=2'b00)) & ((~ main_stage_0_10)
      | (~ COMP_LOOP_asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b01) | (rem_12cyc_st_9_3_2!=2'b00))
      & ((~ main_stage_0_3) | (~ COMP_LOOP_asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b01)
      | (rem_12cyc_st_2_3_2!=2'b00)) & ((~ main_stage_0_4) | (~ COMP_LOOP_asn_itm_3)
      | (rem_12cyc_st_3_1_0!=2'b01) | (rem_12cyc_st_3_3_2!=2'b00)) & ((~ main_stage_0_5)
      | (~ COMP_LOOP_asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b01) | (rem_12cyc_st_4_3_2!=2'b00))
      & ((~ main_stage_0_6) | (~ COMP_LOOP_asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b01)
      | (rem_12cyc_st_5_3_2!=2'b00)) & ((~ main_stage_0_7) | (~ COMP_LOOP_asn_itm_6)
      | (rem_12cyc_st_6_1_0!=2'b01) | (rem_12cyc_st_6_3_2!=2'b00)) & ((~ main_stage_0_11)
      | (~ COMP_LOOP_asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b01) | (rem_12cyc_st_10_3_2!=2'b00))
      & ((COMP_LOOP_acc_tmp!=2'b00) | (COMP_LOOP_acc_1_tmp[1]) | nand_250_cse);
  assign nor_479_nl = ~((rem_12cyc_1_0[0]) | (~ and_tmp_44));
  assign or_175_nl = (~ main_stage_0_2) | (~ COMP_LOOP_asn_itm_1) | (rem_12cyc_3_2!=2'b00)
      | (rem_12cyc_1_0[1]);
  assign mux_tmp_76 = MUX_s_1_2_2(nor_479_nl, and_tmp_44, or_175_nl);
  assign and_dcpl_393 = (COMP_LOOP_acc_1_tmp[1:0]==2'b10);
  assign and_dcpl_394 = and_dcpl_293 & and_dcpl_393;
  assign and_dcpl_395 = and_dcpl_295 & (rem_12cyc_st_2_1_0[1]);
  assign or_tmp_185 = (rem_12cyc_1_0!=2'b10) | (rem_12cyc_3_2!=2'b00) | not_tmp_54;
  assign or_190_cse = (COMP_LOOP_acc_1_tmp[1:0]!=2'b10) | (COMP_LOOP_acc_tmp!=2'b00);
  assign nor_478_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_185));
  assign mux_77_nl = MUX_s_1_2_2(nor_478_nl, or_tmp_185, or_190_cse);
  assign and_dcpl_397 = mux_77_nl & and_dcpl_298 & and_dcpl_395;
  assign and_dcpl_398 = and_dcpl_301 & (rem_12cyc_st_3_1_0[1]);
  assign or_195_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2!=2'b00) |
      (~ COMP_LOOP_asn_itm_2) | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp_45 = or_195_cse & or_tmp_185;
  assign nor_477_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_45));
  assign mux_78_nl = MUX_s_1_2_2(nor_477_nl, and_tmp_45, or_190_cse);
  assign and_dcpl_400 = mux_78_nl & and_dcpl_304 & and_dcpl_398;
  assign and_dcpl_401 = and_dcpl_307 & (rem_12cyc_st_4_1_0[1]);
  assign or_199_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2!=2'b00) |
      (~ COMP_LOOP_asn_itm_3) | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_47 = or_195_cse & or_199_cse & or_tmp_185;
  assign nor_476_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_47));
  assign mux_79_nl = MUX_s_1_2_2(nor_476_nl, and_tmp_47, or_190_cse);
  assign and_dcpl_403 = mux_79_nl & and_dcpl_310 & and_dcpl_401;
  assign and_dcpl_404 = and_dcpl_313 & (rem_12cyc_st_5_1_0[1]);
  assign or_204_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2!=2'b00) |
      (~ COMP_LOOP_asn_itm_4) | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_50 = or_195_cse & or_199_cse & or_204_cse & or_tmp_185;
  assign nor_475_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_50));
  assign mux_80_nl = MUX_s_1_2_2(nor_475_nl, and_tmp_50, or_190_cse);
  assign and_dcpl_406 = mux_80_nl & and_dcpl_316 & and_dcpl_404;
  assign or_210_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2!=2'b00) |
      (~ COMP_LOOP_asn_itm_5) | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_54 = or_195_cse & or_199_cse & or_204_cse & or_210_cse & or_tmp_185;
  assign nor_474_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_54));
  assign mux_81_nl = MUX_s_1_2_2(nor_474_nl, and_tmp_54, or_190_cse);
  assign and_dcpl_409 = mux_81_nl & and_dcpl_112 & and_dcpl_117;
  assign or_217_cse = (rem_12cyc_st_6_1_0!=2'b10) | (rem_12cyc_st_6_3_2!=2'b00);
  assign nor_472_nl = ~(and_dcpl_111 | (~ or_tmp_185));
  assign mux_82_nl = MUX_s_1_2_2(nor_472_nl, or_tmp_185, or_217_cse);
  assign and_tmp_58 = or_195_cse & or_199_cse & or_204_cse & or_210_cse & mux_82_nl;
  assign nor_473_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_58));
  assign mux_83_nl = MUX_s_1_2_2(nor_473_nl, and_tmp_58, or_190_cse);
  assign and_dcpl_413 = mux_83_nl & and_dcpl_85 & and_dcpl_90;
  assign or_226_cse = (rem_12cyc_st_7_1_0!=2'b10) | (rem_12cyc_st_7_3_2!=2'b00);
  assign nor_469_nl = ~(and_dcpl_84 | (~ or_tmp_185));
  assign mux_tmp_84 = MUX_s_1_2_2(nor_469_nl, or_tmp_185, or_226_cse);
  assign nor_470_nl = ~(and_dcpl_111 | (~ mux_tmp_84));
  assign mux_85_nl = MUX_s_1_2_2(nor_470_nl, mux_tmp_84, or_217_cse);
  assign and_tmp_62 = or_195_cse & or_199_cse & or_204_cse & or_210_cse & mux_85_nl;
  assign nor_471_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_62));
  assign mux_86_nl = MUX_s_1_2_2(nor_471_nl, and_tmp_62, or_190_cse);
  assign and_dcpl_417 = mux_86_nl & and_dcpl_58 & and_dcpl_63;
  assign or_237_cse = (rem_12cyc_st_8_1_0!=2'b10) | (rem_12cyc_st_8_3_2!=2'b00);
  assign nor_465_nl = ~(and_dcpl_57 | (~ or_tmp_185));
  assign mux_tmp_87 = MUX_s_1_2_2(nor_465_nl, or_tmp_185, or_237_cse);
  assign nor_466_nl = ~(and_dcpl_84 | (~ mux_tmp_87));
  assign mux_tmp_88 = MUX_s_1_2_2(nor_466_nl, mux_tmp_87, or_226_cse);
  assign nor_467_nl = ~(and_dcpl_111 | (~ mux_tmp_88));
  assign mux_89_nl = MUX_s_1_2_2(nor_467_nl, mux_tmp_88, or_217_cse);
  assign and_tmp_66 = or_195_cse & or_199_cse & or_204_cse & or_210_cse & mux_89_nl;
  assign nor_468_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_66));
  assign mux_90_nl = MUX_s_1_2_2(nor_468_nl, and_tmp_66, or_190_cse);
  assign and_dcpl_421 = mux_90_nl & and_dcpl_31 & and_dcpl_36;
  assign nor_460_nl = ~(and_dcpl_30 | (~ or_tmp_185));
  assign or_250_nl = (rem_12cyc_st_9_1_0!=2'b10) | (rem_12cyc_st_9_3_2!=2'b00);
  assign mux_tmp_91 = MUX_s_1_2_2(nor_460_nl, or_tmp_185, or_250_nl);
  assign nor_461_nl = ~(and_dcpl_57 | (~ mux_tmp_91));
  assign mux_tmp_92 = MUX_s_1_2_2(nor_461_nl, mux_tmp_91, or_237_cse);
  assign nor_462_nl = ~(and_dcpl_84 | (~ mux_tmp_92));
  assign mux_tmp_93 = MUX_s_1_2_2(nor_462_nl, mux_tmp_92, or_226_cse);
  assign nor_463_nl = ~(and_dcpl_111 | (~ mux_tmp_93));
  assign mux_94_nl = MUX_s_1_2_2(nor_463_nl, mux_tmp_93, or_217_cse);
  assign and_tmp_70 = or_195_cse & or_199_cse & or_204_cse & or_210_cse & mux_94_nl;
  assign nor_464_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_70));
  assign mux_95_nl = MUX_s_1_2_2(nor_464_nl, and_tmp_70, or_190_cse);
  assign and_dcpl_425 = mux_95_nl & and_dcpl_4 & and_dcpl_9;
  assign and_tmp_80 = ((~ main_stage_0_2) | (~ COMP_LOOP_asn_itm_1) | (rem_12cyc_3_2!=2'b00)
      | (rem_12cyc_1_0!=2'b10)) & ((~ main_stage_0_8) | (~ COMP_LOOP_asn_itm_7) |
      (rem_12cyc_st_7_1_0!=2'b10) | (rem_12cyc_st_7_3_2!=2'b00)) & ((~ main_stage_0_9)
      | (~ COMP_LOOP_asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b10) | (rem_12cyc_st_8_3_2!=2'b00))
      & ((~ main_stage_0_10) | (~ COMP_LOOP_asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b10)
      | (rem_12cyc_st_9_3_2!=2'b00)) & or_195_cse & or_199_cse & or_204_cse & or_210_cse
      & ((~ main_stage_0_7) | (~ COMP_LOOP_asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b10)
      | (rem_12cyc_st_6_3_2!=2'b00)) & ((~ main_stage_0_11) | (~ COMP_LOOP_asn_itm_10)
      | (rem_12cyc_st_10_1_0!=2'b10) | (rem_12cyc_st_10_3_2!=2'b00)) & ((COMP_LOOP_acc_tmp!=2'b00)
      | (COMP_LOOP_acc_1_tmp[1:0]!=2'b10) | (~ ccs_ccore_start_rsci_idat));
  assign and_dcpl_430 = (COMP_LOOP_acc_1_tmp[1:0]==2'b11);
  assign and_dcpl_431 = and_dcpl_293 & and_dcpl_430;
  assign or_tmp_263 = (rem_12cyc_1_0!=2'b11) | (rem_12cyc_3_2!=2'b00) | not_tmp_54;
  assign or_270_cse = (COMP_LOOP_acc_1_tmp[1:0]!=2'b11) | (COMP_LOOP_acc_tmp!=2'b00);
  assign nor_459_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_263));
  assign mux_96_nl = MUX_s_1_2_2(nor_459_nl, or_tmp_263, or_270_cse);
  assign and_dcpl_433 = mux_96_nl & and_dcpl_358 & and_dcpl_395;
  assign or_275_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2!=2'b00);
  assign and_1142_nl = nand_276_cse & or_tmp_263;
  assign mux_tmp_97 = MUX_s_1_2_2(and_1142_nl, or_tmp_263, or_275_cse);
  assign nor_458_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_97));
  assign mux_98_nl = MUX_s_1_2_2(nor_458_nl, mux_tmp_97, or_270_cse);
  assign and_dcpl_435 = mux_98_nl & and_dcpl_362 & and_dcpl_398;
  assign or_280_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2!=2'b00);
  assign and_1140_nl = nand_274_cse & or_tmp_263;
  assign mux_tmp_99 = MUX_s_1_2_2(and_1140_nl, or_tmp_263, or_280_cse);
  assign and_1141_nl = nand_276_cse & mux_tmp_99;
  assign mux_tmp_100 = MUX_s_1_2_2(and_1141_nl, mux_tmp_99, or_275_cse);
  assign nor_457_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_100));
  assign mux_101_nl = MUX_s_1_2_2(nor_457_nl, mux_tmp_100, or_270_cse);
  assign and_dcpl_437 = mux_101_nl & and_dcpl_366 & and_dcpl_401;
  assign or_287_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2!=2'b00);
  assign and_1137_nl = nand_271_cse & or_tmp_263;
  assign mux_tmp_102 = MUX_s_1_2_2(and_1137_nl, or_tmp_263, or_287_cse);
  assign and_1138_nl = nand_274_cse & mux_tmp_102;
  assign mux_tmp_103 = MUX_s_1_2_2(and_1138_nl, mux_tmp_102, or_280_cse);
  assign and_1139_nl = nand_276_cse & mux_tmp_103;
  assign mux_tmp_104 = MUX_s_1_2_2(and_1139_nl, mux_tmp_103, or_275_cse);
  assign nor_456_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_104));
  assign mux_105_nl = MUX_s_1_2_2(nor_456_nl, mux_tmp_104, or_270_cse);
  assign and_dcpl_439 = mux_105_nl & and_dcpl_370 & and_dcpl_404;
  assign or_296_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2!=2'b00);
  assign and_1133_nl = nand_267_cse & or_tmp_263;
  assign mux_tmp_106 = MUX_s_1_2_2(and_1133_nl, or_tmp_263, or_296_cse);
  assign and_1134_nl = nand_271_cse & mux_tmp_106;
  assign mux_tmp_107 = MUX_s_1_2_2(and_1134_nl, mux_tmp_106, or_287_cse);
  assign and_1135_nl = nand_274_cse & mux_tmp_107;
  assign mux_tmp_108 = MUX_s_1_2_2(and_1135_nl, mux_tmp_107, or_280_cse);
  assign and_1136_nl = nand_276_cse & mux_tmp_108;
  assign mux_tmp_109 = MUX_s_1_2_2(and_1136_nl, mux_tmp_108, or_275_cse);
  assign nor_455_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_109));
  assign mux_110_nl = MUX_s_1_2_2(nor_455_nl, mux_tmp_109, or_270_cse);
  assign and_dcpl_442 = mux_110_nl & and_dcpl_112 & and_dcpl_119;
  assign or_307_cse = (rem_12cyc_st_6_1_0!=2'b11) | (rem_12cyc_st_6_3_2!=2'b00);
  assign nor_453_nl = ~(and_dcpl_111 | (~ or_tmp_263));
  assign mux_tmp_111 = MUX_s_1_2_2(nor_453_nl, or_tmp_263, or_307_cse);
  assign and_1129_nl = nand_267_cse & mux_tmp_111;
  assign mux_tmp_112 = MUX_s_1_2_2(and_1129_nl, mux_tmp_111, or_296_cse);
  assign and_1130_nl = nand_271_cse & mux_tmp_112;
  assign mux_tmp_113 = MUX_s_1_2_2(and_1130_nl, mux_tmp_112, or_287_cse);
  assign and_1131_nl = nand_274_cse & mux_tmp_113;
  assign mux_tmp_114 = MUX_s_1_2_2(and_1131_nl, mux_tmp_113, or_280_cse);
  assign and_1132_nl = nand_276_cse & mux_tmp_114;
  assign mux_tmp_115 = MUX_s_1_2_2(and_1132_nl, mux_tmp_114, or_275_cse);
  assign nor_454_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_115));
  assign mux_116_nl = MUX_s_1_2_2(nor_454_nl, mux_tmp_115, or_270_cse);
  assign and_dcpl_445 = mux_116_nl & and_dcpl_85 & and_dcpl_92;
  assign or_320_cse = (rem_12cyc_st_7_1_0!=2'b11) | (rem_12cyc_st_7_3_2!=2'b00);
  assign nor_450_nl = ~(and_dcpl_84 | (~ or_tmp_263));
  assign mux_tmp_117 = MUX_s_1_2_2(nor_450_nl, or_tmp_263, or_320_cse);
  assign nor_451_nl = ~(and_dcpl_111 | (~ mux_tmp_117));
  assign mux_tmp_118 = MUX_s_1_2_2(nor_451_nl, mux_tmp_117, or_307_cse);
  assign and_1125_nl = nand_267_cse & mux_tmp_118;
  assign mux_tmp_119 = MUX_s_1_2_2(and_1125_nl, mux_tmp_118, or_296_cse);
  assign and_1126_nl = nand_271_cse & mux_tmp_119;
  assign mux_tmp_120 = MUX_s_1_2_2(and_1126_nl, mux_tmp_119, or_287_cse);
  assign and_1127_nl = nand_274_cse & mux_tmp_120;
  assign mux_tmp_121 = MUX_s_1_2_2(and_1127_nl, mux_tmp_120, or_280_cse);
  assign and_1128_nl = nand_276_cse & mux_tmp_121;
  assign mux_tmp_122 = MUX_s_1_2_2(and_1128_nl, mux_tmp_121, or_275_cse);
  assign nor_452_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_122));
  assign mux_123_nl = MUX_s_1_2_2(nor_452_nl, mux_tmp_122, or_270_cse);
  assign and_dcpl_448 = mux_123_nl & and_dcpl_58 & and_dcpl_65;
  assign or_335_cse = (rem_12cyc_st_8_1_0!=2'b11) | (rem_12cyc_st_8_3_2!=2'b00);
  assign nor_446_nl = ~(and_dcpl_57 | (~ or_tmp_263));
  assign mux_tmp_124 = MUX_s_1_2_2(nor_446_nl, or_tmp_263, or_335_cse);
  assign nor_447_nl = ~(and_dcpl_84 | (~ mux_tmp_124));
  assign mux_tmp_125 = MUX_s_1_2_2(nor_447_nl, mux_tmp_124, or_320_cse);
  assign nor_448_nl = ~(and_dcpl_111 | (~ mux_tmp_125));
  assign mux_tmp_126 = MUX_s_1_2_2(nor_448_nl, mux_tmp_125, or_307_cse);
  assign and_1121_nl = nand_267_cse & mux_tmp_126;
  assign mux_tmp_127 = MUX_s_1_2_2(and_1121_nl, mux_tmp_126, or_296_cse);
  assign and_1122_nl = nand_271_cse & mux_tmp_127;
  assign mux_tmp_128 = MUX_s_1_2_2(and_1122_nl, mux_tmp_127, or_287_cse);
  assign and_1123_nl = nand_274_cse & mux_tmp_128;
  assign mux_tmp_129 = MUX_s_1_2_2(and_1123_nl, mux_tmp_128, or_280_cse);
  assign and_1124_nl = nand_276_cse & mux_tmp_129;
  assign mux_tmp_130 = MUX_s_1_2_2(and_1124_nl, mux_tmp_129, or_275_cse);
  assign nor_449_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_130));
  assign mux_131_nl = MUX_s_1_2_2(nor_449_nl, mux_tmp_130, or_270_cse);
  assign and_dcpl_451 = mux_131_nl & and_dcpl_31 & and_dcpl_38;
  assign nor_441_nl = ~(and_dcpl_30 | (~ or_tmp_263));
  assign or_352_nl = (rem_12cyc_st_9_1_0!=2'b11) | (rem_12cyc_st_9_3_2!=2'b00);
  assign mux_tmp_132 = MUX_s_1_2_2(nor_441_nl, or_tmp_263, or_352_nl);
  assign nor_442_nl = ~(and_dcpl_57 | (~ mux_tmp_132));
  assign mux_tmp_133 = MUX_s_1_2_2(nor_442_nl, mux_tmp_132, or_335_cse);
  assign nor_443_nl = ~(and_dcpl_84 | (~ mux_tmp_133));
  assign mux_tmp_134 = MUX_s_1_2_2(nor_443_nl, mux_tmp_133, or_320_cse);
  assign nor_444_nl = ~(and_dcpl_111 | (~ mux_tmp_134));
  assign mux_tmp_135 = MUX_s_1_2_2(nor_444_nl, mux_tmp_134, or_307_cse);
  assign and_1117_nl = nand_267_cse & mux_tmp_135;
  assign mux_tmp_136 = MUX_s_1_2_2(and_1117_nl, mux_tmp_135, or_296_cse);
  assign and_1118_nl = nand_271_cse & mux_tmp_136;
  assign mux_tmp_137 = MUX_s_1_2_2(and_1118_nl, mux_tmp_136, or_287_cse);
  assign and_1119_nl = nand_274_cse & mux_tmp_137;
  assign mux_tmp_138 = MUX_s_1_2_2(and_1119_nl, mux_tmp_137, or_280_cse);
  assign and_1120_nl = nand_276_cse & mux_tmp_138;
  assign mux_tmp_139 = MUX_s_1_2_2(and_1120_nl, mux_tmp_138, or_275_cse);
  assign nor_445_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_139));
  assign mux_140_nl = MUX_s_1_2_2(nor_445_nl, mux_tmp_139, or_270_cse);
  assign and_dcpl_454 = mux_140_nl & and_dcpl_4 & and_dcpl_11;
  assign nand_222_cse = ~((COMP_LOOP_acc_1_tmp[1:0]==2'b11) & ccs_ccore_start_rsci_idat);
  assign and_tmp_89 = ((~ main_stage_0_8) | (~ COMP_LOOP_asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b11)
      | (rem_12cyc_st_7_3_2!=2'b00)) & ((~ main_stage_0_9) | (~ COMP_LOOP_asn_itm_8)
      | (rem_12cyc_st_8_1_0!=2'b11) | (rem_12cyc_st_8_3_2!=2'b00)) & ((~ main_stage_0_10)
      | (~ COMP_LOOP_asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b11) | (rem_12cyc_st_9_3_2!=2'b00))
      & ((~ main_stage_0_3) | (~ COMP_LOOP_asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b11)
      | (rem_12cyc_st_2_3_2!=2'b00)) & ((~ main_stage_0_4) | (~ COMP_LOOP_asn_itm_3)
      | (rem_12cyc_st_3_1_0!=2'b11) | (rem_12cyc_st_3_3_2!=2'b00)) & ((~ main_stage_0_5)
      | (~ COMP_LOOP_asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b11) | (rem_12cyc_st_4_3_2!=2'b00))
      & ((~ main_stage_0_6) | (~ COMP_LOOP_asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b11)
      | (rem_12cyc_st_5_3_2!=2'b00)) & ((~ main_stage_0_7) | (~ COMP_LOOP_asn_itm_6)
      | (rem_12cyc_st_6_1_0!=2'b11) | (rem_12cyc_st_6_3_2!=2'b00)) & ((~ main_stage_0_11)
      | (~ COMP_LOOP_asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b11) | (rem_12cyc_st_10_3_2!=2'b00))
      & ((COMP_LOOP_acc_tmp!=2'b00) | nand_222_cse);
  assign nand_223_cse = ~((rem_12cyc_1_0==2'b11));
  assign and_1116_nl = nand_223_cse & and_tmp_89;
  assign or_362_nl = (~ main_stage_0_2) | (~ COMP_LOOP_asn_itm_1) | (rem_12cyc_3_2!=2'b00);
  assign mux_tmp_141 = MUX_s_1_2_2(and_1116_nl, and_tmp_89, or_362_nl);
  assign and_dcpl_460 = ccs_ccore_start_rsci_idat & (COMP_LOOP_acc_tmp==2'b01);
  assign and_dcpl_461 = and_dcpl_460 & and_dcpl_291;
  assign and_dcpl_462 = (rem_12cyc_st_2_3_2==2'b01);
  assign and_dcpl_463 = and_dcpl_462 & (~ (rem_12cyc_st_2_1_0[1]));
  assign not_tmp_332 = ~((rem_12cyc_3_2[0]) & COMP_LOOP_asn_itm_1 & main_stage_0_2);
  assign or_tmp_368 = (rem_12cyc_1_0!=2'b00) | (rem_12cyc_3_2[1]) | not_tmp_332;
  assign nand_281_cse = ~((COMP_LOOP_acc_tmp[0]) & ccs_ccore_start_rsci_idat);
  assign or_377_cse = (COMP_LOOP_acc_1_tmp[1:0]!=2'b00) | (COMP_LOOP_acc_tmp[1]);
  assign and_1172_nl = nand_281_cse & or_tmp_368;
  assign mux_142_nl = MUX_s_1_2_2(and_1172_nl, or_tmp_368, or_377_cse);
  assign and_dcpl_465 = mux_142_nl & and_dcpl_298 & and_dcpl_463;
  assign and_dcpl_466 = (rem_12cyc_st_3_3_2==2'b01);
  assign and_dcpl_467 = and_dcpl_466 & (~ (rem_12cyc_st_3_1_0[1]));
  assign or_382_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2!=2'b01) | (~
      COMP_LOOP_asn_itm_2) | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp_90 = or_382_cse & or_tmp_368;
  assign and_1114_nl = nand_281_cse & and_tmp_90;
  assign mux_143_nl = MUX_s_1_2_2(and_1114_nl, and_tmp_90, or_377_cse);
  assign and_dcpl_469 = mux_143_nl & and_dcpl_304 & and_dcpl_467;
  assign and_dcpl_470 = (rem_12cyc_st_4_3_2==2'b01);
  assign and_dcpl_471 = and_dcpl_470 & (~ (rem_12cyc_st_4_1_0[1]));
  assign or_386_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2!=2'b01) | (~
      COMP_LOOP_asn_itm_3) | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_92 = or_382_cse & or_386_cse & or_tmp_368;
  assign and_1113_nl = nand_281_cse & and_tmp_92;
  assign mux_144_nl = MUX_s_1_2_2(and_1113_nl, and_tmp_92, or_377_cse);
  assign and_dcpl_473 = mux_144_nl & and_dcpl_310 & and_dcpl_471;
  assign and_dcpl_474 = (rem_12cyc_st_5_3_2==2'b01);
  assign and_dcpl_475 = and_dcpl_474 & (~ (rem_12cyc_st_5_1_0[1]));
  assign or_391_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2!=2'b01) | (~
      COMP_LOOP_asn_itm_4) | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_95 = or_382_cse & or_386_cse & or_391_cse & or_tmp_368;
  assign and_1112_nl = nand_281_cse & and_tmp_95;
  assign mux_145_nl = MUX_s_1_2_2(and_1112_nl, and_tmp_95, or_377_cse);
  assign and_dcpl_477 = mux_145_nl & and_dcpl_316 & and_dcpl_475;
  assign or_397_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2!=2'b01) | (~
      COMP_LOOP_asn_itm_5) | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_99 = or_382_cse & or_386_cse & or_391_cse & or_397_cse & or_tmp_368;
  assign and_1111_nl = nand_281_cse & and_tmp_99;
  assign mux_146_nl = MUX_s_1_2_2(and_1111_nl, and_tmp_99, or_377_cse);
  assign and_dcpl_480 = mux_146_nl & and_dcpl_121 & and_dcpl_110;
  assign nand_215_cse = ~((rem_12cyc_st_6_3_2[0]) & COMP_LOOP_asn_itm_6 & main_stage_0_7);
  assign or_404_cse = (rem_12cyc_st_6_1_0!=2'b00) | (rem_12cyc_st_6_3_2[1]);
  assign and_1109_nl = nand_215_cse & or_tmp_368;
  assign mux_147_nl = MUX_s_1_2_2(and_1109_nl, or_tmp_368, or_404_cse);
  assign and_tmp_103 = or_382_cse & or_386_cse & or_391_cse & or_397_cse & mux_147_nl;
  assign and_1110_nl = nand_281_cse & and_tmp_103;
  assign mux_148_nl = MUX_s_1_2_2(and_1110_nl, and_tmp_103, or_377_cse);
  assign and_dcpl_483 = mux_148_nl & and_dcpl_94 & and_dcpl_83;
  assign nand_212_cse = ~((rem_12cyc_st_7_3_2[0]) & COMP_LOOP_asn_itm_7 & main_stage_0_8);
  assign or_413_cse = (rem_12cyc_st_7_1_0!=2'b00) | (rem_12cyc_st_7_3_2[1]);
  assign and_1106_nl = nand_212_cse & or_tmp_368;
  assign mux_tmp_149 = MUX_s_1_2_2(and_1106_nl, or_tmp_368, or_413_cse);
  assign and_1107_nl = nand_215_cse & mux_tmp_149;
  assign mux_150_nl = MUX_s_1_2_2(and_1107_nl, mux_tmp_149, or_404_cse);
  assign and_tmp_107 = or_382_cse & or_386_cse & or_391_cse & or_397_cse & mux_150_nl;
  assign and_1108_nl = nand_281_cse & and_tmp_107;
  assign mux_151_nl = MUX_s_1_2_2(and_1108_nl, and_tmp_107, or_377_cse);
  assign and_dcpl_486 = mux_151_nl & and_dcpl_67 & and_dcpl_56;
  assign nand_208_cse = ~((rem_12cyc_st_8_3_2[0]) & COMP_LOOP_asn_itm_8 & main_stage_0_9);
  assign or_424_cse = (rem_12cyc_st_8_1_0!=2'b00) | (rem_12cyc_st_8_3_2[1]);
  assign and_1102_nl = nand_208_cse & or_tmp_368;
  assign mux_tmp_152 = MUX_s_1_2_2(and_1102_nl, or_tmp_368, or_424_cse);
  assign and_1103_nl = nand_212_cse & mux_tmp_152;
  assign mux_tmp_153 = MUX_s_1_2_2(and_1103_nl, mux_tmp_152, or_413_cse);
  assign and_1104_nl = nand_215_cse & mux_tmp_153;
  assign mux_154_nl = MUX_s_1_2_2(and_1104_nl, mux_tmp_153, or_404_cse);
  assign and_tmp_111 = or_382_cse & or_386_cse & or_391_cse & or_397_cse & mux_154_nl;
  assign and_1105_nl = nand_281_cse & and_tmp_111;
  assign mux_155_nl = MUX_s_1_2_2(and_1105_nl, and_tmp_111, or_377_cse);
  assign and_dcpl_489 = mux_155_nl & and_dcpl_40 & and_dcpl_29;
  assign nand_203_cse = ~((rem_12cyc_st_9_3_2[0]) & COMP_LOOP_asn_itm_9 & main_stage_0_10);
  assign and_1097_nl = nand_203_cse & or_tmp_368;
  assign or_437_nl = (rem_12cyc_st_9_1_0!=2'b00) | (rem_12cyc_st_9_3_2[1]);
  assign mux_tmp_156 = MUX_s_1_2_2(and_1097_nl, or_tmp_368, or_437_nl);
  assign and_1098_nl = nand_208_cse & mux_tmp_156;
  assign mux_tmp_157 = MUX_s_1_2_2(and_1098_nl, mux_tmp_156, or_424_cse);
  assign and_1099_nl = nand_212_cse & mux_tmp_157;
  assign mux_tmp_158 = MUX_s_1_2_2(and_1099_nl, mux_tmp_157, or_413_cse);
  assign and_1100_nl = nand_215_cse & mux_tmp_158;
  assign mux_159_nl = MUX_s_1_2_2(and_1100_nl, mux_tmp_158, or_404_cse);
  assign and_tmp_115 = or_382_cse & or_386_cse & or_391_cse & or_397_cse & mux_159_nl;
  assign and_1101_nl = nand_281_cse & and_tmp_115;
  assign mux_160_nl = MUX_s_1_2_2(and_1101_nl, and_tmp_115, or_377_cse);
  assign and_dcpl_492 = mux_160_nl & and_dcpl_13 & and_dcpl_2;
  assign and_tmp_125 = ((~ main_stage_0_2) | (~ COMP_LOOP_asn_itm_1) | (rem_12cyc_3_2!=2'b01)
      | (rem_12cyc_1_0!=2'b00)) & ((~ main_stage_0_8) | (~ COMP_LOOP_asn_itm_7) |
      (rem_12cyc_st_7_1_0!=2'b00) | (rem_12cyc_st_7_3_2!=2'b01)) & ((~ main_stage_0_9)
      | (~ COMP_LOOP_asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b00) | (rem_12cyc_st_8_3_2!=2'b01))
      & ((~ main_stage_0_10) | (~ COMP_LOOP_asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b00)
      | (rem_12cyc_st_9_3_2!=2'b01)) & or_382_cse & or_386_cse & or_391_cse & or_397_cse
      & ((~ main_stage_0_7) | (~ COMP_LOOP_asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b00)
      | (rem_12cyc_st_6_3_2!=2'b01)) & ((~ main_stage_0_11) | (~ COMP_LOOP_asn_itm_10)
      | (rem_12cyc_st_10_1_0!=2'b00) | (rem_12cyc_st_10_3_2!=2'b01)) & ((COMP_LOOP_acc_tmp!=2'b01)
      | (COMP_LOOP_acc_1_tmp[1:0]!=2'b00) | (~ ccs_ccore_start_rsci_idat));
  assign and_dcpl_498 = and_dcpl_460 & and_dcpl_355;
  assign or_tmp_446 = (rem_12cyc_1_0!=2'b01) | (rem_12cyc_3_2[1]) | not_tmp_332;
  assign or_458_cse = (COMP_LOOP_acc_1_tmp[1:0]!=2'b01) | (COMP_LOOP_acc_tmp[1]);
  assign and_1171_nl = nand_281_cse & or_tmp_446;
  assign mux_161_nl = MUX_s_1_2_2(and_1171_nl, or_tmp_446, or_458_cse);
  assign and_dcpl_500 = mux_161_nl & and_dcpl_358 & and_dcpl_463;
  assign or_463_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2!=2'b01);
  assign and_1094_nl = nand_276_cse & or_tmp_446;
  assign mux_tmp_162 = MUX_s_1_2_2(and_1094_nl, or_tmp_446, or_463_cse);
  assign and_1095_nl = nand_281_cse & mux_tmp_162;
  assign mux_163_nl = MUX_s_1_2_2(and_1095_nl, mux_tmp_162, or_458_cse);
  assign and_dcpl_502 = mux_163_nl & and_dcpl_362 & and_dcpl_467;
  assign nand_198_cse = ~((rem_12cyc_st_3_3_2[0]) & COMP_LOOP_asn_itm_3 & main_stage_0_4
      & (rem_12cyc_st_3_1_0[0]));
  assign or_468_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2[1]);
  assign and_1091_nl = nand_198_cse & or_tmp_446;
  assign mux_tmp_164 = MUX_s_1_2_2(and_1091_nl, or_tmp_446, or_468_cse);
  assign and_1092_nl = nand_276_cse & mux_tmp_164;
  assign mux_tmp_165 = MUX_s_1_2_2(and_1092_nl, mux_tmp_164, or_463_cse);
  assign and_1093_nl = nand_281_cse & mux_tmp_165;
  assign mux_166_nl = MUX_s_1_2_2(and_1093_nl, mux_tmp_165, or_458_cse);
  assign and_dcpl_504 = mux_166_nl & and_dcpl_366 & and_dcpl_471;
  assign or_475_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2!=2'b01);
  assign and_1087_nl = nand_271_cse & or_tmp_446;
  assign mux_tmp_167 = MUX_s_1_2_2(and_1087_nl, or_tmp_446, or_475_cse);
  assign and_1088_nl = nand_198_cse & mux_tmp_167;
  assign mux_tmp_168 = MUX_s_1_2_2(and_1088_nl, mux_tmp_167, or_468_cse);
  assign and_1089_nl = nand_276_cse & mux_tmp_168;
  assign mux_tmp_169 = MUX_s_1_2_2(and_1089_nl, mux_tmp_168, or_463_cse);
  assign and_1090_nl = nand_281_cse & mux_tmp_169;
  assign mux_170_nl = MUX_s_1_2_2(and_1090_nl, mux_tmp_169, or_458_cse);
  assign and_dcpl_506 = mux_170_nl & and_dcpl_370 & and_dcpl_475;
  assign nand_189_cse = ~((rem_12cyc_st_5_3_2[0]) & COMP_LOOP_asn_itm_5 & main_stage_0_6
      & (rem_12cyc_st_5_1_0[0]));
  assign or_484_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2[1]);
  assign and_1082_nl = nand_189_cse & or_tmp_446;
  assign mux_tmp_171 = MUX_s_1_2_2(and_1082_nl, or_tmp_446, or_484_cse);
  assign and_1083_nl = nand_271_cse & mux_tmp_171;
  assign mux_tmp_172 = MUX_s_1_2_2(and_1083_nl, mux_tmp_171, or_475_cse);
  assign and_1084_nl = nand_198_cse & mux_tmp_172;
  assign mux_tmp_173 = MUX_s_1_2_2(and_1084_nl, mux_tmp_172, or_468_cse);
  assign and_1085_nl = nand_276_cse & mux_tmp_173;
  assign mux_tmp_174 = MUX_s_1_2_2(and_1085_nl, mux_tmp_173, or_463_cse);
  assign and_1086_nl = nand_281_cse & mux_tmp_174;
  assign mux_175_nl = MUX_s_1_2_2(and_1086_nl, mux_tmp_174, or_458_cse);
  assign and_dcpl_508 = mux_175_nl & and_dcpl_121 & and_dcpl_115;
  assign or_495_cse = (rem_12cyc_st_6_1_0!=2'b01) | (rem_12cyc_st_6_3_2[1]);
  assign and_1076_nl = nand_215_cse & or_tmp_446;
  assign mux_tmp_176 = MUX_s_1_2_2(and_1076_nl, or_tmp_446, or_495_cse);
  assign and_1077_nl = nand_189_cse & mux_tmp_176;
  assign mux_tmp_177 = MUX_s_1_2_2(and_1077_nl, mux_tmp_176, or_484_cse);
  assign and_1078_nl = nand_271_cse & mux_tmp_177;
  assign mux_tmp_178 = MUX_s_1_2_2(and_1078_nl, mux_tmp_177, or_475_cse);
  assign and_1079_nl = nand_198_cse & mux_tmp_178;
  assign mux_tmp_179 = MUX_s_1_2_2(and_1079_nl, mux_tmp_178, or_468_cse);
  assign and_1080_nl = nand_276_cse & mux_tmp_179;
  assign mux_tmp_180 = MUX_s_1_2_2(and_1080_nl, mux_tmp_179, or_463_cse);
  assign and_1081_nl = nand_281_cse & mux_tmp_180;
  assign mux_181_nl = MUX_s_1_2_2(and_1081_nl, mux_tmp_180, or_458_cse);
  assign and_dcpl_510 = mux_181_nl & and_dcpl_94 & and_dcpl_87;
  assign or_508_cse = (rem_12cyc_st_7_1_0!=2'b01) | (rem_12cyc_st_7_3_2[1]);
  assign and_1069_nl = nand_212_cse & or_tmp_446;
  assign mux_tmp_182 = MUX_s_1_2_2(and_1069_nl, or_tmp_446, or_508_cse);
  assign and_1070_nl = nand_215_cse & mux_tmp_182;
  assign mux_tmp_183 = MUX_s_1_2_2(and_1070_nl, mux_tmp_182, or_495_cse);
  assign and_1071_nl = nand_189_cse & mux_tmp_183;
  assign mux_tmp_184 = MUX_s_1_2_2(and_1071_nl, mux_tmp_183, or_484_cse);
  assign and_1072_nl = nand_271_cse & mux_tmp_184;
  assign mux_tmp_185 = MUX_s_1_2_2(and_1072_nl, mux_tmp_184, or_475_cse);
  assign and_1073_nl = nand_198_cse & mux_tmp_185;
  assign mux_tmp_186 = MUX_s_1_2_2(and_1073_nl, mux_tmp_185, or_468_cse);
  assign and_1074_nl = nand_276_cse & mux_tmp_186;
  assign mux_tmp_187 = MUX_s_1_2_2(and_1074_nl, mux_tmp_186, or_463_cse);
  assign and_1075_nl = nand_281_cse & mux_tmp_187;
  assign mux_188_nl = MUX_s_1_2_2(and_1075_nl, mux_tmp_187, or_458_cse);
  assign and_dcpl_512 = mux_188_nl & and_dcpl_67 & and_dcpl_60;
  assign or_523_cse = (rem_12cyc_st_8_1_0!=2'b01) | (rem_12cyc_st_8_3_2[1]);
  assign and_1061_nl = nand_208_cse & or_tmp_446;
  assign mux_tmp_189 = MUX_s_1_2_2(and_1061_nl, or_tmp_446, or_523_cse);
  assign and_1062_nl = nand_212_cse & mux_tmp_189;
  assign mux_tmp_190 = MUX_s_1_2_2(and_1062_nl, mux_tmp_189, or_508_cse);
  assign and_1063_nl = nand_215_cse & mux_tmp_190;
  assign mux_tmp_191 = MUX_s_1_2_2(and_1063_nl, mux_tmp_190, or_495_cse);
  assign and_1064_nl = nand_189_cse & mux_tmp_191;
  assign mux_tmp_192 = MUX_s_1_2_2(and_1064_nl, mux_tmp_191, or_484_cse);
  assign and_1065_nl = nand_271_cse & mux_tmp_192;
  assign mux_tmp_193 = MUX_s_1_2_2(and_1065_nl, mux_tmp_192, or_475_cse);
  assign and_1066_nl = nand_198_cse & mux_tmp_193;
  assign mux_tmp_194 = MUX_s_1_2_2(and_1066_nl, mux_tmp_193, or_468_cse);
  assign and_1067_nl = nand_276_cse & mux_tmp_194;
  assign mux_tmp_195 = MUX_s_1_2_2(and_1067_nl, mux_tmp_194, or_463_cse);
  assign and_1068_nl = nand_281_cse & mux_tmp_195;
  assign mux_196_nl = MUX_s_1_2_2(and_1068_nl, mux_tmp_195, or_458_cse);
  assign and_dcpl_514 = mux_196_nl & and_dcpl_40 & and_dcpl_33;
  assign and_1052_nl = nand_203_cse & or_tmp_446;
  assign or_540_nl = (rem_12cyc_st_9_1_0!=2'b01) | (rem_12cyc_st_9_3_2[1]);
  assign mux_tmp_197 = MUX_s_1_2_2(and_1052_nl, or_tmp_446, or_540_nl);
  assign and_1053_nl = nand_208_cse & mux_tmp_197;
  assign mux_tmp_198 = MUX_s_1_2_2(and_1053_nl, mux_tmp_197, or_523_cse);
  assign and_1054_nl = nand_212_cse & mux_tmp_198;
  assign mux_tmp_199 = MUX_s_1_2_2(and_1054_nl, mux_tmp_198, or_508_cse);
  assign and_1055_nl = nand_215_cse & mux_tmp_199;
  assign mux_tmp_200 = MUX_s_1_2_2(and_1055_nl, mux_tmp_199, or_495_cse);
  assign and_1056_nl = nand_189_cse & mux_tmp_200;
  assign mux_tmp_201 = MUX_s_1_2_2(and_1056_nl, mux_tmp_200, or_484_cse);
  assign and_1057_nl = nand_271_cse & mux_tmp_201;
  assign mux_tmp_202 = MUX_s_1_2_2(and_1057_nl, mux_tmp_201, or_475_cse);
  assign and_1058_nl = nand_198_cse & mux_tmp_202;
  assign mux_tmp_203 = MUX_s_1_2_2(and_1058_nl, mux_tmp_202, or_468_cse);
  assign and_1059_nl = nand_276_cse & mux_tmp_203;
  assign mux_tmp_204 = MUX_s_1_2_2(and_1059_nl, mux_tmp_203, or_463_cse);
  assign and_1060_nl = nand_281_cse & mux_tmp_204;
  assign mux_205_nl = MUX_s_1_2_2(and_1060_nl, mux_tmp_204, or_458_cse);
  assign and_dcpl_516 = mux_205_nl & and_dcpl_13 & and_dcpl_6;
  assign and_tmp_134 = ((~ main_stage_0_8) | (~ COMP_LOOP_asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b01)
      | (rem_12cyc_st_7_3_2!=2'b01)) & ((~ main_stage_0_9) | (~ COMP_LOOP_asn_itm_8)
      | (rem_12cyc_st_8_1_0!=2'b01) | (rem_12cyc_st_8_3_2!=2'b01)) & ((~ main_stage_0_10)
      | (~ COMP_LOOP_asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b01) | (rem_12cyc_st_9_3_2!=2'b01))
      & ((~ main_stage_0_3) | (~ COMP_LOOP_asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b01)
      | (rem_12cyc_st_2_3_2!=2'b01)) & ((~ main_stage_0_4) | (~ COMP_LOOP_asn_itm_3)
      | (rem_12cyc_st_3_1_0!=2'b01) | (rem_12cyc_st_3_3_2!=2'b01)) & ((~ main_stage_0_5)
      | (~ COMP_LOOP_asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b01) | (rem_12cyc_st_4_3_2!=2'b01))
      & ((~ main_stage_0_6) | (~ COMP_LOOP_asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b01)
      | (rem_12cyc_st_5_3_2!=2'b01)) & ((~ main_stage_0_7) | (~ COMP_LOOP_asn_itm_6)
      | (rem_12cyc_st_6_1_0!=2'b01) | (rem_12cyc_st_6_3_2!=2'b01)) & ((~ main_stage_0_11)
      | (~ COMP_LOOP_asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b01) | (rem_12cyc_st_10_3_2!=2'b01))
      & ((COMP_LOOP_acc_tmp!=2'b01) | (COMP_LOOP_acc_1_tmp[1]) | nand_250_cse);
  assign nor_438_nl = ~((rem_12cyc_1_0[0]) | (~ and_tmp_134));
  assign or_550_nl = (~ main_stage_0_2) | (~ COMP_LOOP_asn_itm_1) | (rem_12cyc_3_2!=2'b01)
      | (rem_12cyc_1_0[1]);
  assign mux_tmp_206 = MUX_s_1_2_2(nor_438_nl, and_tmp_134, or_550_nl);
  assign and_dcpl_520 = and_dcpl_460 & and_dcpl_393;
  assign and_dcpl_521 = and_dcpl_462 & (rem_12cyc_st_2_1_0[1]);
  assign or_tmp_551 = (rem_12cyc_1_0!=2'b10) | (rem_12cyc_3_2[1]) | not_tmp_332;
  assign or_564_cse = (COMP_LOOP_acc_1_tmp[1:0]!=2'b10) | (COMP_LOOP_acc_tmp[1]);
  assign and_1170_nl = nand_281_cse & or_tmp_551;
  assign mux_207_nl = MUX_s_1_2_2(and_1170_nl, or_tmp_551, or_564_cse);
  assign and_dcpl_523 = mux_207_nl & and_dcpl_298 & and_dcpl_521;
  assign and_dcpl_524 = and_dcpl_466 & (rem_12cyc_st_3_1_0[1]);
  assign or_569_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2!=2'b01) |
      (~ COMP_LOOP_asn_itm_2) | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp_135 = or_569_cse & or_tmp_551;
  assign and_1050_nl = nand_281_cse & and_tmp_135;
  assign mux_208_nl = MUX_s_1_2_2(and_1050_nl, and_tmp_135, or_564_cse);
  assign and_dcpl_526 = mux_208_nl & and_dcpl_304 & and_dcpl_524;
  assign and_dcpl_527 = and_dcpl_470 & (rem_12cyc_st_4_1_0[1]);
  assign or_573_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2!=2'b01) |
      (~ COMP_LOOP_asn_itm_3) | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_137 = or_569_cse & or_573_cse & or_tmp_551;
  assign and_1049_nl = nand_281_cse & and_tmp_137;
  assign mux_209_nl = MUX_s_1_2_2(and_1049_nl, and_tmp_137, or_564_cse);
  assign and_dcpl_529 = mux_209_nl & and_dcpl_310 & and_dcpl_527;
  assign and_dcpl_530 = and_dcpl_474 & (rem_12cyc_st_5_1_0[1]);
  assign or_578_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2!=2'b01) |
      (~ COMP_LOOP_asn_itm_4) | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_140 = or_569_cse & or_573_cse & or_578_cse & or_tmp_551;
  assign and_1048_nl = nand_281_cse & and_tmp_140;
  assign mux_210_nl = MUX_s_1_2_2(and_1048_nl, and_tmp_140, or_564_cse);
  assign and_dcpl_532 = mux_210_nl & and_dcpl_316 & and_dcpl_530;
  assign or_584_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2!=2'b01) |
      (~ COMP_LOOP_asn_itm_5) | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_144 = or_569_cse & or_573_cse & or_578_cse & or_584_cse & or_tmp_551;
  assign and_1047_nl = nand_281_cse & and_tmp_144;
  assign mux_211_nl = MUX_s_1_2_2(and_1047_nl, and_tmp_144, or_564_cse);
  assign and_dcpl_534 = mux_211_nl & and_dcpl_121 & and_dcpl_117;
  assign or_591_cse = (rem_12cyc_st_6_1_0!=2'b10) | (rem_12cyc_st_6_3_2[1]);
  assign and_1045_nl = nand_215_cse & or_tmp_551;
  assign mux_212_nl = MUX_s_1_2_2(and_1045_nl, or_tmp_551, or_591_cse);
  assign and_tmp_148 = or_569_cse & or_573_cse & or_578_cse & or_584_cse & mux_212_nl;
  assign and_1046_nl = nand_281_cse & and_tmp_148;
  assign mux_213_nl = MUX_s_1_2_2(and_1046_nl, and_tmp_148, or_564_cse);
  assign and_dcpl_536 = mux_213_nl & and_dcpl_94 & and_dcpl_90;
  assign or_600_cse = (rem_12cyc_st_7_1_0!=2'b10) | (rem_12cyc_st_7_3_2[1]);
  assign and_1042_nl = nand_212_cse & or_tmp_551;
  assign mux_tmp_214 = MUX_s_1_2_2(and_1042_nl, or_tmp_551, or_600_cse);
  assign and_1043_nl = nand_215_cse & mux_tmp_214;
  assign mux_215_nl = MUX_s_1_2_2(and_1043_nl, mux_tmp_214, or_591_cse);
  assign and_tmp_152 = or_569_cse & or_573_cse & or_578_cse & or_584_cse & mux_215_nl;
  assign and_1044_nl = nand_281_cse & and_tmp_152;
  assign mux_216_nl = MUX_s_1_2_2(and_1044_nl, and_tmp_152, or_564_cse);
  assign and_dcpl_538 = mux_216_nl & and_dcpl_67 & and_dcpl_63;
  assign or_611_cse = (rem_12cyc_st_8_1_0!=2'b10) | (rem_12cyc_st_8_3_2[1]);
  assign and_1038_nl = nand_208_cse & or_tmp_551;
  assign mux_tmp_217 = MUX_s_1_2_2(and_1038_nl, or_tmp_551, or_611_cse);
  assign and_1039_nl = nand_212_cse & mux_tmp_217;
  assign mux_tmp_218 = MUX_s_1_2_2(and_1039_nl, mux_tmp_217, or_600_cse);
  assign and_1040_nl = nand_215_cse & mux_tmp_218;
  assign mux_219_nl = MUX_s_1_2_2(and_1040_nl, mux_tmp_218, or_591_cse);
  assign and_tmp_156 = or_569_cse & or_573_cse & or_578_cse & or_584_cse & mux_219_nl;
  assign and_1041_nl = nand_281_cse & and_tmp_156;
  assign mux_220_nl = MUX_s_1_2_2(and_1041_nl, and_tmp_156, or_564_cse);
  assign and_dcpl_540 = mux_220_nl & and_dcpl_40 & and_dcpl_36;
  assign and_1033_nl = nand_203_cse & or_tmp_551;
  assign or_624_nl = (rem_12cyc_st_9_1_0!=2'b10) | (rem_12cyc_st_9_3_2[1]);
  assign mux_tmp_221 = MUX_s_1_2_2(and_1033_nl, or_tmp_551, or_624_nl);
  assign and_1034_nl = nand_208_cse & mux_tmp_221;
  assign mux_tmp_222 = MUX_s_1_2_2(and_1034_nl, mux_tmp_221, or_611_cse);
  assign and_1035_nl = nand_212_cse & mux_tmp_222;
  assign mux_tmp_223 = MUX_s_1_2_2(and_1035_nl, mux_tmp_222, or_600_cse);
  assign and_1036_nl = nand_215_cse & mux_tmp_223;
  assign mux_224_nl = MUX_s_1_2_2(and_1036_nl, mux_tmp_223, or_591_cse);
  assign and_tmp_160 = or_569_cse & or_573_cse & or_578_cse & or_584_cse & mux_224_nl;
  assign and_1037_nl = nand_281_cse & and_tmp_160;
  assign mux_225_nl = MUX_s_1_2_2(and_1037_nl, and_tmp_160, or_564_cse);
  assign and_dcpl_542 = mux_225_nl & and_dcpl_13 & and_dcpl_9;
  assign and_tmp_170 = ((~ main_stage_0_2) | (~ COMP_LOOP_asn_itm_1) | (rem_12cyc_3_2!=2'b01)
      | (rem_12cyc_1_0!=2'b10)) & ((~ main_stage_0_8) | (~ COMP_LOOP_asn_itm_7) |
      (rem_12cyc_st_7_1_0!=2'b10) | (rem_12cyc_st_7_3_2!=2'b01)) & ((~ main_stage_0_9)
      | (~ COMP_LOOP_asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b10) | (rem_12cyc_st_8_3_2!=2'b01))
      & ((~ main_stage_0_10) | (~ COMP_LOOP_asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b10)
      | (rem_12cyc_st_9_3_2!=2'b01)) & or_569_cse & or_573_cse & or_578_cse & or_584_cse
      & ((~ main_stage_0_7) | (~ COMP_LOOP_asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b10)
      | (rem_12cyc_st_6_3_2!=2'b01)) & ((~ main_stage_0_11) | (~ COMP_LOOP_asn_itm_10)
      | (rem_12cyc_st_10_1_0!=2'b10) | (rem_12cyc_st_10_3_2!=2'b01)) & ((COMP_LOOP_acc_tmp!=2'b01)
      | (COMP_LOOP_acc_1_tmp[1:0]!=2'b10) | (~ ccs_ccore_start_rsci_idat));
  assign and_dcpl_546 = and_dcpl_460 & and_dcpl_430;
  assign or_tmp_629 = (rem_12cyc_1_0!=2'b11) | (rem_12cyc_3_2[1]) | not_tmp_332;
  assign or_643_cse = (COMP_LOOP_acc_1_tmp[1:0]!=2'b11) | (COMP_LOOP_acc_tmp[1]);
  assign and_1169_nl = nand_281_cse & or_tmp_629;
  assign mux_226_nl = MUX_s_1_2_2(and_1169_nl, or_tmp_629, or_643_cse);
  assign and_dcpl_548 = mux_226_nl & and_dcpl_358 & and_dcpl_521;
  assign or_648_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2!=2'b01);
  assign and_1030_nl = nand_276_cse & or_tmp_629;
  assign mux_tmp_227 = MUX_s_1_2_2(and_1030_nl, or_tmp_629, or_648_cse);
  assign and_1031_nl = nand_281_cse & mux_tmp_227;
  assign mux_228_nl = MUX_s_1_2_2(and_1031_nl, mux_tmp_227, or_643_cse);
  assign and_dcpl_550 = mux_228_nl & and_dcpl_362 & and_dcpl_524;
  assign or_653_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2[1]);
  assign and_1027_nl = nand_198_cse & or_tmp_629;
  assign mux_tmp_229 = MUX_s_1_2_2(and_1027_nl, or_tmp_629, or_653_cse);
  assign and_1028_nl = nand_276_cse & mux_tmp_229;
  assign mux_tmp_230 = MUX_s_1_2_2(and_1028_nl, mux_tmp_229, or_648_cse);
  assign and_1029_nl = nand_281_cse & mux_tmp_230;
  assign mux_231_nl = MUX_s_1_2_2(and_1029_nl, mux_tmp_230, or_643_cse);
  assign and_dcpl_552 = mux_231_nl & and_dcpl_366 & and_dcpl_527;
  assign or_660_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2!=2'b01);
  assign and_1023_nl = nand_271_cse & or_tmp_629;
  assign mux_tmp_232 = MUX_s_1_2_2(and_1023_nl, or_tmp_629, or_660_cse);
  assign and_1024_nl = nand_198_cse & mux_tmp_232;
  assign mux_tmp_233 = MUX_s_1_2_2(and_1024_nl, mux_tmp_232, or_653_cse);
  assign and_1025_nl = nand_276_cse & mux_tmp_233;
  assign mux_tmp_234 = MUX_s_1_2_2(and_1025_nl, mux_tmp_233, or_648_cse);
  assign and_1026_nl = nand_281_cse & mux_tmp_234;
  assign mux_235_nl = MUX_s_1_2_2(and_1026_nl, mux_tmp_234, or_643_cse);
  assign and_dcpl_554 = mux_235_nl & and_dcpl_370 & and_dcpl_530;
  assign or_669_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2[1]);
  assign and_1018_nl = nand_189_cse & or_tmp_629;
  assign mux_tmp_236 = MUX_s_1_2_2(and_1018_nl, or_tmp_629, or_669_cse);
  assign and_1019_nl = nand_271_cse & mux_tmp_236;
  assign mux_tmp_237 = MUX_s_1_2_2(and_1019_nl, mux_tmp_236, or_660_cse);
  assign and_1020_nl = nand_198_cse & mux_tmp_237;
  assign mux_tmp_238 = MUX_s_1_2_2(and_1020_nl, mux_tmp_237, or_653_cse);
  assign and_1021_nl = nand_276_cse & mux_tmp_238;
  assign mux_tmp_239 = MUX_s_1_2_2(and_1021_nl, mux_tmp_238, or_648_cse);
  assign and_1022_nl = nand_281_cse & mux_tmp_239;
  assign mux_240_nl = MUX_s_1_2_2(and_1022_nl, mux_tmp_239, or_643_cse);
  assign and_dcpl_556 = mux_240_nl & and_dcpl_121 & and_dcpl_119;
  assign or_680_cse = (rem_12cyc_st_6_1_0!=2'b11) | (rem_12cyc_st_6_3_2[1]);
  assign and_1012_nl = nand_215_cse & or_tmp_629;
  assign mux_tmp_241 = MUX_s_1_2_2(and_1012_nl, or_tmp_629, or_680_cse);
  assign and_1013_nl = nand_189_cse & mux_tmp_241;
  assign mux_tmp_242 = MUX_s_1_2_2(and_1013_nl, mux_tmp_241, or_669_cse);
  assign and_1014_nl = nand_271_cse & mux_tmp_242;
  assign mux_tmp_243 = MUX_s_1_2_2(and_1014_nl, mux_tmp_242, or_660_cse);
  assign and_1015_nl = nand_198_cse & mux_tmp_243;
  assign mux_tmp_244 = MUX_s_1_2_2(and_1015_nl, mux_tmp_243, or_653_cse);
  assign and_1016_nl = nand_276_cse & mux_tmp_244;
  assign mux_tmp_245 = MUX_s_1_2_2(and_1016_nl, mux_tmp_244, or_648_cse);
  assign and_1017_nl = nand_281_cse & mux_tmp_245;
  assign mux_246_nl = MUX_s_1_2_2(and_1017_nl, mux_tmp_245, or_643_cse);
  assign and_dcpl_558 = mux_246_nl & and_dcpl_94 & and_dcpl_92;
  assign or_693_cse = (rem_12cyc_st_7_1_0!=2'b11) | (rem_12cyc_st_7_3_2[1]);
  assign and_1005_nl = nand_212_cse & or_tmp_629;
  assign mux_tmp_247 = MUX_s_1_2_2(and_1005_nl, or_tmp_629, or_693_cse);
  assign and_1006_nl = nand_215_cse & mux_tmp_247;
  assign mux_tmp_248 = MUX_s_1_2_2(and_1006_nl, mux_tmp_247, or_680_cse);
  assign and_1007_nl = nand_189_cse & mux_tmp_248;
  assign mux_tmp_249 = MUX_s_1_2_2(and_1007_nl, mux_tmp_248, or_669_cse);
  assign and_1008_nl = nand_271_cse & mux_tmp_249;
  assign mux_tmp_250 = MUX_s_1_2_2(and_1008_nl, mux_tmp_249, or_660_cse);
  assign and_1009_nl = nand_198_cse & mux_tmp_250;
  assign mux_tmp_251 = MUX_s_1_2_2(and_1009_nl, mux_tmp_250, or_653_cse);
  assign and_1010_nl = nand_276_cse & mux_tmp_251;
  assign mux_tmp_252 = MUX_s_1_2_2(and_1010_nl, mux_tmp_251, or_648_cse);
  assign and_1011_nl = nand_281_cse & mux_tmp_252;
  assign mux_253_nl = MUX_s_1_2_2(and_1011_nl, mux_tmp_252, or_643_cse);
  assign and_dcpl_560 = mux_253_nl & and_dcpl_67 & and_dcpl_65;
  assign or_708_cse = (rem_12cyc_st_8_1_0!=2'b11) | (rem_12cyc_st_8_3_2[1]);
  assign and_997_nl = nand_208_cse & or_tmp_629;
  assign mux_tmp_254 = MUX_s_1_2_2(and_997_nl, or_tmp_629, or_708_cse);
  assign and_998_nl = nand_212_cse & mux_tmp_254;
  assign mux_tmp_255 = MUX_s_1_2_2(and_998_nl, mux_tmp_254, or_693_cse);
  assign and_999_nl = nand_215_cse & mux_tmp_255;
  assign mux_tmp_256 = MUX_s_1_2_2(and_999_nl, mux_tmp_255, or_680_cse);
  assign and_1000_nl = nand_189_cse & mux_tmp_256;
  assign mux_tmp_257 = MUX_s_1_2_2(and_1000_nl, mux_tmp_256, or_669_cse);
  assign and_1001_nl = nand_271_cse & mux_tmp_257;
  assign mux_tmp_258 = MUX_s_1_2_2(and_1001_nl, mux_tmp_257, or_660_cse);
  assign and_1002_nl = nand_198_cse & mux_tmp_258;
  assign mux_tmp_259 = MUX_s_1_2_2(and_1002_nl, mux_tmp_258, or_653_cse);
  assign and_1003_nl = nand_276_cse & mux_tmp_259;
  assign mux_tmp_260 = MUX_s_1_2_2(and_1003_nl, mux_tmp_259, or_648_cse);
  assign and_1004_nl = nand_281_cse & mux_tmp_260;
  assign mux_261_nl = MUX_s_1_2_2(and_1004_nl, mux_tmp_260, or_643_cse);
  assign and_dcpl_562 = mux_261_nl & and_dcpl_40 & and_dcpl_38;
  assign and_988_nl = nand_203_cse & or_tmp_629;
  assign or_725_nl = (rem_12cyc_st_9_1_0!=2'b11) | (rem_12cyc_st_9_3_2[1]);
  assign mux_tmp_262 = MUX_s_1_2_2(and_988_nl, or_tmp_629, or_725_nl);
  assign and_989_nl = nand_208_cse & mux_tmp_262;
  assign mux_tmp_263 = MUX_s_1_2_2(and_989_nl, mux_tmp_262, or_708_cse);
  assign and_990_nl = nand_212_cse & mux_tmp_263;
  assign mux_tmp_264 = MUX_s_1_2_2(and_990_nl, mux_tmp_263, or_693_cse);
  assign and_991_nl = nand_215_cse & mux_tmp_264;
  assign mux_tmp_265 = MUX_s_1_2_2(and_991_nl, mux_tmp_264, or_680_cse);
  assign and_992_nl = nand_189_cse & mux_tmp_265;
  assign mux_tmp_266 = MUX_s_1_2_2(and_992_nl, mux_tmp_265, or_669_cse);
  assign and_993_nl = nand_271_cse & mux_tmp_266;
  assign mux_tmp_267 = MUX_s_1_2_2(and_993_nl, mux_tmp_266, or_660_cse);
  assign and_994_nl = nand_198_cse & mux_tmp_267;
  assign mux_tmp_268 = MUX_s_1_2_2(and_994_nl, mux_tmp_267, or_653_cse);
  assign and_995_nl = nand_276_cse & mux_tmp_268;
  assign mux_tmp_269 = MUX_s_1_2_2(and_995_nl, mux_tmp_268, or_648_cse);
  assign and_996_nl = nand_281_cse & mux_tmp_269;
  assign mux_270_nl = MUX_s_1_2_2(and_996_nl, mux_tmp_269, or_643_cse);
  assign and_dcpl_564 = mux_270_nl & and_dcpl_13 & and_dcpl_11;
  assign and_tmp_179 = (~(main_stage_0_8 & COMP_LOOP_asn_itm_7 & (rem_12cyc_st_7_1_0==2'b11)
      & (rem_12cyc_st_7_3_2==2'b01))) & (~(main_stage_0_9 & COMP_LOOP_asn_itm_8 &
      (rem_12cyc_st_8_1_0==2'b11) & (rem_12cyc_st_8_3_2==2'b01))) & (~(main_stage_0_10
      & COMP_LOOP_asn_itm_9 & (rem_12cyc_st_9_1_0==2'b11) & (rem_12cyc_st_9_3_2==2'b01)))
      & (~(main_stage_0_3 & COMP_LOOP_asn_itm_2 & (rem_12cyc_st_2_1_0==2'b11) & (rem_12cyc_st_2_3_2==2'b01)))
      & (~(main_stage_0_4 & COMP_LOOP_asn_itm_3 & (rem_12cyc_st_3_1_0==2'b11) & (rem_12cyc_st_3_3_2==2'b01)))
      & (~(main_stage_0_5 & COMP_LOOP_asn_itm_4 & (rem_12cyc_st_4_1_0==2'b11) & (rem_12cyc_st_4_3_2==2'b01)))
      & (~(main_stage_0_6 & COMP_LOOP_asn_itm_5 & (rem_12cyc_st_5_1_0==2'b11) & (rem_12cyc_st_5_3_2==2'b01)))
      & (~(main_stage_0_7 & COMP_LOOP_asn_itm_6 & (rem_12cyc_st_6_1_0==2'b11) & (rem_12cyc_st_6_3_2==2'b01)))
      & (~(main_stage_0_11 & COMP_LOOP_asn_itm_10 & (rem_12cyc_st_10_1_0==2'b11)
      & (rem_12cyc_st_10_3_2==2'b01))) & ((COMP_LOOP_acc_tmp[1]) | (~((COMP_LOOP_acc_tmp[0])
      & (COMP_LOOP_acc_1_tmp[1:0]==2'b11) & ccs_ccore_start_rsci_idat)));
  assign and_987_nl = (~((rem_12cyc_3_2[0]) & (rem_12cyc_1_0==2'b11))) & and_tmp_179;
  assign or_735_nl = (~ main_stage_0_2) | (~ COMP_LOOP_asn_itm_1) | (rem_12cyc_3_2[1]);
  assign mux_tmp_271 = MUX_s_1_2_2(and_987_nl, and_tmp_179, or_735_nl);
  assign and_dcpl_568 = and_dcpl_292 & (COMP_LOOP_acc_tmp[1]);
  assign and_dcpl_569 = and_dcpl_568 & and_dcpl_291;
  assign and_dcpl_570 = (rem_12cyc_st_2_3_2==2'b10);
  assign and_dcpl_571 = and_dcpl_570 & (~ (rem_12cyc_st_2_1_0[1]));
  assign or_tmp_733 = (rem_12cyc_1_0!=2'b00) | (rem_12cyc_3_2!=2'b10) | not_tmp_54;
  assign or_748_cse = (COMP_LOOP_acc_1_tmp[1:0]!=2'b00) | (COMP_LOOP_acc_tmp!=2'b10);
  assign nor_435_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_733));
  assign mux_272_nl = MUX_s_1_2_2(nor_435_nl, or_tmp_733, or_748_cse);
  assign and_dcpl_573 = mux_272_nl & and_dcpl_298 & and_dcpl_571;
  assign and_dcpl_574 = (rem_12cyc_st_3_3_2==2'b10);
  assign and_dcpl_575 = and_dcpl_574 & (~ (rem_12cyc_st_3_1_0[1]));
  assign or_753_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2!=2'b10) | (~
      COMP_LOOP_asn_itm_2) | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp_180 = or_753_cse & or_tmp_733;
  assign nor_434_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_180));
  assign mux_273_nl = MUX_s_1_2_2(nor_434_nl, and_tmp_180, or_748_cse);
  assign and_dcpl_577 = mux_273_nl & and_dcpl_304 & and_dcpl_575;
  assign and_dcpl_578 = (rem_12cyc_st_4_3_2==2'b10);
  assign and_dcpl_579 = and_dcpl_578 & (~ (rem_12cyc_st_4_1_0[1]));
  assign or_757_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2!=2'b10) | (~
      COMP_LOOP_asn_itm_3) | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_182 = or_753_cse & or_757_cse & or_tmp_733;
  assign nor_433_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_182));
  assign mux_274_nl = MUX_s_1_2_2(nor_433_nl, and_tmp_182, or_748_cse);
  assign and_dcpl_581 = mux_274_nl & and_dcpl_310 & and_dcpl_579;
  assign and_dcpl_582 = (rem_12cyc_st_5_3_2==2'b10);
  assign and_dcpl_583 = and_dcpl_582 & (~ (rem_12cyc_st_5_1_0[1]));
  assign or_762_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2!=2'b10) | (~
      COMP_LOOP_asn_itm_4) | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_185 = or_753_cse & or_757_cse & or_762_cse & or_tmp_733;
  assign nor_432_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_185));
  assign mux_275_nl = MUX_s_1_2_2(nor_432_nl, and_tmp_185, or_748_cse);
  assign and_dcpl_585 = mux_275_nl & and_dcpl_316 & and_dcpl_583;
  assign or_768_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2!=2'b10) | (~
      COMP_LOOP_asn_itm_5) | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_189 = or_753_cse & or_757_cse & or_762_cse & or_768_cse & or_tmp_733;
  assign nor_431_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_189));
  assign mux_276_nl = MUX_s_1_2_2(nor_431_nl, and_tmp_189, or_748_cse);
  assign and_dcpl_589 = mux_276_nl & and_dcpl_112 & and_dcpl_126 & (~ (rem_12cyc_st_6_1_0[1]));
  assign or_775_cse = (rem_12cyc_st_6_1_0!=2'b00) | (rem_12cyc_st_6_3_2!=2'b10);
  assign nor_429_nl = ~(and_dcpl_111 | (~ or_tmp_733));
  assign mux_277_nl = MUX_s_1_2_2(nor_429_nl, or_tmp_733, or_775_cse);
  assign and_tmp_193 = or_753_cse & or_757_cse & or_762_cse & or_768_cse & mux_277_nl;
  assign nor_430_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_193));
  assign mux_278_nl = MUX_s_1_2_2(nor_430_nl, and_tmp_193, or_748_cse);
  assign and_dcpl_593 = mux_278_nl & and_dcpl_85 & and_dcpl_99 & (~ (rem_12cyc_st_7_1_0[0]));
  assign or_784_cse = (rem_12cyc_st_7_1_0!=2'b00) | (rem_12cyc_st_7_3_2!=2'b10);
  assign nor_426_nl = ~(and_dcpl_84 | (~ or_tmp_733));
  assign mux_tmp_279 = MUX_s_1_2_2(nor_426_nl, or_tmp_733, or_784_cse);
  assign nor_427_nl = ~(and_dcpl_111 | (~ mux_tmp_279));
  assign mux_280_nl = MUX_s_1_2_2(nor_427_nl, mux_tmp_279, or_775_cse);
  assign and_tmp_197 = or_753_cse & or_757_cse & or_762_cse & or_768_cse & mux_280_nl;
  assign nor_428_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_197));
  assign mux_281_nl = MUX_s_1_2_2(nor_428_nl, and_tmp_197, or_748_cse);
  assign and_dcpl_597 = mux_281_nl & and_dcpl_58 & and_dcpl_72 & (~ (rem_12cyc_st_8_1_0[0]));
  assign or_795_cse = (rem_12cyc_st_8_1_0!=2'b00) | (rem_12cyc_st_8_3_2!=2'b10);
  assign nor_422_nl = ~(and_dcpl_57 | (~ or_tmp_733));
  assign mux_tmp_282 = MUX_s_1_2_2(nor_422_nl, or_tmp_733, or_795_cse);
  assign nor_423_nl = ~(and_dcpl_84 | (~ mux_tmp_282));
  assign mux_tmp_283 = MUX_s_1_2_2(nor_423_nl, mux_tmp_282, or_784_cse);
  assign nor_424_nl = ~(and_dcpl_111 | (~ mux_tmp_283));
  assign mux_284_nl = MUX_s_1_2_2(nor_424_nl, mux_tmp_283, or_775_cse);
  assign and_tmp_201 = or_753_cse & or_757_cse & or_762_cse & or_768_cse & mux_284_nl;
  assign nor_425_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_201));
  assign mux_285_nl = MUX_s_1_2_2(nor_425_nl, and_tmp_201, or_748_cse);
  assign and_dcpl_601 = mux_285_nl & and_dcpl_31 & and_dcpl_45 & (~ (rem_12cyc_st_9_1_0[0]));
  assign nor_417_nl = ~(and_dcpl_30 | (~ or_tmp_733));
  assign or_808_nl = (rem_12cyc_st_9_1_0!=2'b00) | (rem_12cyc_st_9_3_2!=2'b10);
  assign mux_tmp_286 = MUX_s_1_2_2(nor_417_nl, or_tmp_733, or_808_nl);
  assign nor_418_nl = ~(and_dcpl_57 | (~ mux_tmp_286));
  assign mux_tmp_287 = MUX_s_1_2_2(nor_418_nl, mux_tmp_286, or_795_cse);
  assign nor_419_nl = ~(and_dcpl_84 | (~ mux_tmp_287));
  assign mux_tmp_288 = MUX_s_1_2_2(nor_419_nl, mux_tmp_287, or_784_cse);
  assign nor_420_nl = ~(and_dcpl_111 | (~ mux_tmp_288));
  assign mux_289_nl = MUX_s_1_2_2(nor_420_nl, mux_tmp_288, or_775_cse);
  assign and_tmp_205 = or_753_cse & or_757_cse & or_762_cse & or_768_cse & mux_289_nl;
  assign nor_421_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_205));
  assign mux_290_nl = MUX_s_1_2_2(nor_421_nl, and_tmp_205, or_748_cse);
  assign and_dcpl_605 = mux_290_nl & and_dcpl_4 & and_dcpl_18 & (~ (rem_12cyc_st_10_1_0[0]));
  assign or_tmp_808 = (COMP_LOOP_acc_tmp!=2'b10) | (COMP_LOOP_acc_1_tmp[1:0]!=2'b00)
      | (~ ccs_ccore_start_rsci_idat);
  assign nor_408_nl = ~((rem_12cyc_st_10_3_2[1]) | (~ or_tmp_808));
  assign or_823_nl = (~ main_stage_0_11) | (~ COMP_LOOP_asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b00)
      | (rem_12cyc_st_10_3_2[0]);
  assign mux_tmp_291 = MUX_s_1_2_2(nor_408_nl, or_tmp_808, or_823_nl);
  assign nor_409_nl = ~((rem_12cyc_st_6_3_2[1]) | (~ mux_tmp_291));
  assign or_822_nl = (~ main_stage_0_7) | (~ COMP_LOOP_asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b00)
      | (rem_12cyc_st_6_3_2[0]);
  assign mux_tmp_292 = MUX_s_1_2_2(nor_409_nl, mux_tmp_291, or_822_nl);
  assign nor_410_nl = ~((rem_12cyc_st_5_3_2[1]) | (~ mux_tmp_292));
  assign or_821_nl = (~ main_stage_0_6) | (~ COMP_LOOP_asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b00)
      | (rem_12cyc_st_5_3_2[0]);
  assign mux_tmp_293 = MUX_s_1_2_2(nor_410_nl, mux_tmp_292, or_821_nl);
  assign nor_411_nl = ~((rem_12cyc_st_4_3_2[1]) | (~ mux_tmp_293));
  assign or_820_nl = (~ main_stage_0_5) | (~ COMP_LOOP_asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b00)
      | (rem_12cyc_st_4_3_2[0]);
  assign mux_tmp_294 = MUX_s_1_2_2(nor_411_nl, mux_tmp_293, or_820_nl);
  assign nor_412_nl = ~((rem_12cyc_st_3_3_2[1]) | (~ mux_tmp_294));
  assign or_819_nl = (~ main_stage_0_4) | (~ COMP_LOOP_asn_itm_3) | (rem_12cyc_st_3_1_0!=2'b00)
      | (rem_12cyc_st_3_3_2[0]);
  assign mux_tmp_295 = MUX_s_1_2_2(nor_412_nl, mux_tmp_294, or_819_nl);
  assign nor_413_nl = ~((rem_12cyc_st_2_3_2[1]) | (~ mux_tmp_295));
  assign or_818_nl = (~ main_stage_0_3) | (~ COMP_LOOP_asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b00)
      | (rem_12cyc_st_2_3_2[0]);
  assign mux_tmp_296 = MUX_s_1_2_2(nor_413_nl, mux_tmp_295, or_818_nl);
  assign nor_414_nl = ~((rem_12cyc_st_9_3_2[1]) | (~ mux_tmp_296));
  assign or_817_nl = (~ main_stage_0_10) | (~ COMP_LOOP_asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b00)
      | (rem_12cyc_st_9_3_2[0]);
  assign mux_tmp_297 = MUX_s_1_2_2(nor_414_nl, mux_tmp_296, or_817_nl);
  assign nor_415_nl = ~((rem_12cyc_st_8_3_2[1]) | (~ mux_tmp_297));
  assign or_816_nl = (~ main_stage_0_9) | (~ COMP_LOOP_asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b00)
      | (rem_12cyc_st_8_3_2[0]);
  assign mux_tmp_298 = MUX_s_1_2_2(nor_415_nl, mux_tmp_297, or_816_nl);
  assign nor_416_nl = ~((rem_12cyc_st_7_3_2[1]) | (~ mux_tmp_298));
  assign or_815_nl = (~ main_stage_0_8) | (~ COMP_LOOP_asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b00)
      | (rem_12cyc_st_7_3_2[0]);
  assign mux_299_nl = MUX_s_1_2_2(nor_416_nl, mux_tmp_298, or_815_nl);
  assign and_tmp_206 = ((~ main_stage_0_2) | (~ COMP_LOOP_asn_itm_1) | (rem_12cyc_3_2!=2'b10)
      | (rem_12cyc_1_0!=2'b00)) & mux_299_nl;
  assign and_dcpl_610 = and_dcpl_568 & and_dcpl_355;
  assign or_tmp_820 = (rem_12cyc_1_0!=2'b01) | (rem_12cyc_3_2!=2'b10) | not_tmp_54;
  assign or_837_cse = (COMP_LOOP_acc_1_tmp[1:0]!=2'b01) | (COMP_LOOP_acc_tmp!=2'b10);
  assign nor_407_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_820));
  assign mux_300_nl = MUX_s_1_2_2(nor_407_nl, or_tmp_820, or_837_cse);
  assign and_dcpl_612 = mux_300_nl & and_dcpl_358 & and_dcpl_571;
  assign nand_84_cse = ~((rem_12cyc_st_2_3_2[1]) & COMP_LOOP_asn_itm_2 & main_stage_0_3
      & (rem_12cyc_st_2_1_0[0]));
  assign or_842_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2[0]);
  assign and_986_nl = nand_84_cse & or_tmp_820;
  assign mux_tmp_301 = MUX_s_1_2_2(and_986_nl, or_tmp_820, or_842_cse);
  assign nor_406_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_301));
  assign mux_302_nl = MUX_s_1_2_2(nor_406_nl, mux_tmp_301, or_837_cse);
  assign and_dcpl_614 = mux_302_nl & and_dcpl_362 & and_dcpl_575;
  assign or_847_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2!=2'b10);
  assign and_984_nl = nand_274_cse & or_tmp_820;
  assign mux_tmp_303 = MUX_s_1_2_2(and_984_nl, or_tmp_820, or_847_cse);
  assign and_985_nl = nand_84_cse & mux_tmp_303;
  assign mux_tmp_304 = MUX_s_1_2_2(and_985_nl, mux_tmp_303, or_842_cse);
  assign nor_405_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_304));
  assign mux_305_nl = MUX_s_1_2_2(nor_405_nl, mux_tmp_304, or_837_cse);
  assign and_dcpl_616 = mux_305_nl & and_dcpl_366 & and_dcpl_579;
  assign nand_79_cse = ~((rem_12cyc_st_4_3_2[1]) & COMP_LOOP_asn_itm_4 & main_stage_0_5
      & (rem_12cyc_st_4_1_0[0]));
  assign or_854_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2[0]);
  assign and_981_nl = nand_79_cse & or_tmp_820;
  assign mux_tmp_306 = MUX_s_1_2_2(and_981_nl, or_tmp_820, or_854_cse);
  assign and_982_nl = nand_274_cse & mux_tmp_306;
  assign mux_tmp_307 = MUX_s_1_2_2(and_982_nl, mux_tmp_306, or_847_cse);
  assign and_983_nl = nand_84_cse & mux_tmp_307;
  assign mux_tmp_308 = MUX_s_1_2_2(and_983_nl, mux_tmp_307, or_842_cse);
  assign nor_404_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_308));
  assign mux_309_nl = MUX_s_1_2_2(nor_404_nl, mux_tmp_308, or_837_cse);
  assign and_dcpl_618 = mux_309_nl & and_dcpl_370 & and_dcpl_583;
  assign or_863_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2!=2'b10);
  assign and_977_nl = nand_267_cse & or_tmp_820;
  assign mux_tmp_310 = MUX_s_1_2_2(and_977_nl, or_tmp_820, or_863_cse);
  assign and_978_nl = nand_79_cse & mux_tmp_310;
  assign mux_tmp_311 = MUX_s_1_2_2(and_978_nl, mux_tmp_310, or_854_cse);
  assign and_979_nl = nand_274_cse & mux_tmp_311;
  assign mux_tmp_312 = MUX_s_1_2_2(and_979_nl, mux_tmp_311, or_847_cse);
  assign and_980_nl = nand_84_cse & mux_tmp_312;
  assign mux_tmp_313 = MUX_s_1_2_2(and_980_nl, mux_tmp_312, or_842_cse);
  assign nor_403_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_313));
  assign mux_314_nl = MUX_s_1_2_2(nor_403_nl, mux_tmp_313, or_837_cse);
  assign and_dcpl_622 = mux_314_nl & and_dcpl_112 & and_dcpl_129 & (~ (rem_12cyc_st_6_1_0[1]));
  assign or_874_cse = (rem_12cyc_st_6_1_0!=2'b01) | (rem_12cyc_st_6_3_2!=2'b10);
  assign nor_401_nl = ~(and_dcpl_111 | (~ or_tmp_820));
  assign mux_tmp_315 = MUX_s_1_2_2(nor_401_nl, or_tmp_820, or_874_cse);
  assign and_973_nl = nand_267_cse & mux_tmp_315;
  assign mux_tmp_316 = MUX_s_1_2_2(and_973_nl, mux_tmp_315, or_863_cse);
  assign and_974_nl = nand_79_cse & mux_tmp_316;
  assign mux_tmp_317 = MUX_s_1_2_2(and_974_nl, mux_tmp_316, or_854_cse);
  assign and_975_nl = nand_274_cse & mux_tmp_317;
  assign mux_tmp_318 = MUX_s_1_2_2(and_975_nl, mux_tmp_317, or_847_cse);
  assign and_976_nl = nand_84_cse & mux_tmp_318;
  assign mux_tmp_319 = MUX_s_1_2_2(and_976_nl, mux_tmp_318, or_842_cse);
  assign nor_402_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_319));
  assign mux_320_nl = MUX_s_1_2_2(nor_402_nl, mux_tmp_319, or_837_cse);
  assign and_dcpl_625 = mux_320_nl & and_dcpl_85 & and_dcpl_99 & (rem_12cyc_st_7_1_0[0]);
  assign or_887_cse = (rem_12cyc_st_7_1_0!=2'b01) | (rem_12cyc_st_7_3_2!=2'b10);
  assign nor_398_nl = ~(and_dcpl_84 | (~ or_tmp_820));
  assign mux_tmp_321 = MUX_s_1_2_2(nor_398_nl, or_tmp_820, or_887_cse);
  assign nor_399_nl = ~(and_dcpl_111 | (~ mux_tmp_321));
  assign mux_tmp_322 = MUX_s_1_2_2(nor_399_nl, mux_tmp_321, or_874_cse);
  assign and_969_nl = nand_267_cse & mux_tmp_322;
  assign mux_tmp_323 = MUX_s_1_2_2(and_969_nl, mux_tmp_322, or_863_cse);
  assign and_970_nl = nand_79_cse & mux_tmp_323;
  assign mux_tmp_324 = MUX_s_1_2_2(and_970_nl, mux_tmp_323, or_854_cse);
  assign and_971_nl = nand_274_cse & mux_tmp_324;
  assign mux_tmp_325 = MUX_s_1_2_2(and_971_nl, mux_tmp_324, or_847_cse);
  assign and_972_nl = nand_84_cse & mux_tmp_325;
  assign mux_tmp_326 = MUX_s_1_2_2(and_972_nl, mux_tmp_325, or_842_cse);
  assign nor_400_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_326));
  assign mux_327_nl = MUX_s_1_2_2(nor_400_nl, mux_tmp_326, or_837_cse);
  assign and_dcpl_628 = mux_327_nl & and_dcpl_58 & and_dcpl_72 & (rem_12cyc_st_8_1_0[0]);
  assign or_902_cse = (rem_12cyc_st_8_1_0!=2'b01) | (rem_12cyc_st_8_3_2!=2'b10);
  assign nor_394_nl = ~(and_dcpl_57 | (~ or_tmp_820));
  assign mux_tmp_328 = MUX_s_1_2_2(nor_394_nl, or_tmp_820, or_902_cse);
  assign nor_395_nl = ~(and_dcpl_84 | (~ mux_tmp_328));
  assign mux_tmp_329 = MUX_s_1_2_2(nor_395_nl, mux_tmp_328, or_887_cse);
  assign nor_396_nl = ~(and_dcpl_111 | (~ mux_tmp_329));
  assign mux_tmp_330 = MUX_s_1_2_2(nor_396_nl, mux_tmp_329, or_874_cse);
  assign and_965_nl = nand_267_cse & mux_tmp_330;
  assign mux_tmp_331 = MUX_s_1_2_2(and_965_nl, mux_tmp_330, or_863_cse);
  assign and_966_nl = nand_79_cse & mux_tmp_331;
  assign mux_tmp_332 = MUX_s_1_2_2(and_966_nl, mux_tmp_331, or_854_cse);
  assign and_967_nl = nand_274_cse & mux_tmp_332;
  assign mux_tmp_333 = MUX_s_1_2_2(and_967_nl, mux_tmp_332, or_847_cse);
  assign and_968_nl = nand_84_cse & mux_tmp_333;
  assign mux_tmp_334 = MUX_s_1_2_2(and_968_nl, mux_tmp_333, or_842_cse);
  assign nor_397_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_334));
  assign mux_335_nl = MUX_s_1_2_2(nor_397_nl, mux_tmp_334, or_837_cse);
  assign and_dcpl_631 = mux_335_nl & and_dcpl_31 & and_dcpl_45 & (rem_12cyc_st_9_1_0[0]);
  assign nor_389_nl = ~(and_dcpl_30 | (~ or_tmp_820));
  assign or_919_nl = (rem_12cyc_st_9_1_0!=2'b01) | (rem_12cyc_st_9_3_2!=2'b10);
  assign mux_tmp_336 = MUX_s_1_2_2(nor_389_nl, or_tmp_820, or_919_nl);
  assign nor_390_nl = ~(and_dcpl_57 | (~ mux_tmp_336));
  assign mux_tmp_337 = MUX_s_1_2_2(nor_390_nl, mux_tmp_336, or_902_cse);
  assign nor_391_nl = ~(and_dcpl_84 | (~ mux_tmp_337));
  assign mux_tmp_338 = MUX_s_1_2_2(nor_391_nl, mux_tmp_337, or_887_cse);
  assign nor_392_nl = ~(and_dcpl_111 | (~ mux_tmp_338));
  assign mux_tmp_339 = MUX_s_1_2_2(nor_392_nl, mux_tmp_338, or_874_cse);
  assign and_961_nl = nand_267_cse & mux_tmp_339;
  assign mux_tmp_340 = MUX_s_1_2_2(and_961_nl, mux_tmp_339, or_863_cse);
  assign and_962_nl = nand_79_cse & mux_tmp_340;
  assign mux_tmp_341 = MUX_s_1_2_2(and_962_nl, mux_tmp_340, or_854_cse);
  assign and_963_nl = nand_274_cse & mux_tmp_341;
  assign mux_tmp_342 = MUX_s_1_2_2(and_963_nl, mux_tmp_341, or_847_cse);
  assign and_964_nl = nand_84_cse & mux_tmp_342;
  assign mux_tmp_343 = MUX_s_1_2_2(and_964_nl, mux_tmp_342, or_842_cse);
  assign nor_393_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_343));
  assign mux_344_nl = MUX_s_1_2_2(nor_393_nl, mux_tmp_343, or_837_cse);
  assign and_dcpl_634 = mux_344_nl & and_dcpl_4 & and_dcpl_18 & (rem_12cyc_st_10_1_0[0]);
  assign or_tmp_921 = (COMP_LOOP_acc_tmp!=2'b10) | (COMP_LOOP_acc_1_tmp[1]) | nand_250_cse;
  assign nor_379_nl = ~((rem_12cyc_st_10_3_2[1]) | (~ or_tmp_921));
  assign or_938_nl = (~ main_stage_0_11) | (~ COMP_LOOP_asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b01)
      | (rem_12cyc_st_10_3_2[0]);
  assign mux_tmp_345 = MUX_s_1_2_2(nor_379_nl, or_tmp_921, or_938_nl);
  assign nor_380_nl = ~((rem_12cyc_st_6_3_2[1]) | (~ mux_tmp_345));
  assign or_937_nl = (~ main_stage_0_7) | (~ COMP_LOOP_asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b01)
      | (rem_12cyc_st_6_3_2[0]);
  assign mux_tmp_346 = MUX_s_1_2_2(nor_380_nl, mux_tmp_345, or_937_nl);
  assign nor_381_nl = ~((rem_12cyc_st_5_3_2[1]) | (~ mux_tmp_346));
  assign or_936_nl = (~ main_stage_0_6) | (~ COMP_LOOP_asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b01)
      | (rem_12cyc_st_5_3_2[0]);
  assign mux_tmp_347 = MUX_s_1_2_2(nor_381_nl, mux_tmp_346, or_936_nl);
  assign nor_382_nl = ~((rem_12cyc_st_4_3_2[1]) | (~ mux_tmp_347));
  assign or_935_nl = (~ main_stage_0_5) | (~ COMP_LOOP_asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b01)
      | (rem_12cyc_st_4_3_2[0]);
  assign mux_tmp_348 = MUX_s_1_2_2(nor_382_nl, mux_tmp_347, or_935_nl);
  assign nor_383_nl = ~((rem_12cyc_st_3_3_2[1]) | (~ mux_tmp_348));
  assign or_934_nl = (~ main_stage_0_4) | (~ COMP_LOOP_asn_itm_3) | (rem_12cyc_st_3_1_0!=2'b01)
      | (rem_12cyc_st_3_3_2[0]);
  assign mux_tmp_349 = MUX_s_1_2_2(nor_383_nl, mux_tmp_348, or_934_nl);
  assign nor_384_nl = ~((rem_12cyc_st_2_3_2[1]) | (~ mux_tmp_349));
  assign or_933_nl = (~ main_stage_0_3) | (~ COMP_LOOP_asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b01)
      | (rem_12cyc_st_2_3_2[0]);
  assign mux_tmp_350 = MUX_s_1_2_2(nor_384_nl, mux_tmp_349, or_933_nl);
  assign nor_385_nl = ~((rem_12cyc_st_9_3_2[1]) | (~ mux_tmp_350));
  assign or_932_nl = (~ main_stage_0_10) | (~ COMP_LOOP_asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b01)
      | (rem_12cyc_st_9_3_2[0]);
  assign mux_tmp_351 = MUX_s_1_2_2(nor_385_nl, mux_tmp_350, or_932_nl);
  assign nor_386_nl = ~((rem_12cyc_st_8_3_2[1]) | (~ mux_tmp_351));
  assign or_931_nl = (~ main_stage_0_9) | (~ COMP_LOOP_asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b01)
      | (rem_12cyc_st_8_3_2[0]);
  assign mux_tmp_352 = MUX_s_1_2_2(nor_386_nl, mux_tmp_351, or_931_nl);
  assign nor_387_nl = ~((rem_12cyc_st_7_3_2[1]) | (~ mux_tmp_352));
  assign or_930_nl = (~ main_stage_0_8) | (~ COMP_LOOP_asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b01)
      | (rem_12cyc_st_7_3_2[0]);
  assign mux_tmp_353 = MUX_s_1_2_2(nor_387_nl, mux_tmp_352, or_930_nl);
  assign nor_388_nl = ~((rem_12cyc_1_0[0]) | (~ mux_tmp_353));
  assign or_929_nl = (~ main_stage_0_2) | (~ COMP_LOOP_asn_itm_1) | (rem_12cyc_3_2!=2'b10)
      | (rem_12cyc_1_0[1]);
  assign mux_tmp_354 = MUX_s_1_2_2(nor_388_nl, mux_tmp_353, or_929_nl);
  assign and_dcpl_638 = and_dcpl_568 & and_dcpl_393;
  assign and_dcpl_639 = and_dcpl_570 & (rem_12cyc_st_2_1_0[1]);
  assign or_tmp_934 = (rem_12cyc_1_0!=2'b10) | (rem_12cyc_3_2!=2'b10) | not_tmp_54;
  assign or_952_cse = (COMP_LOOP_acc_1_tmp[1:0]!=2'b10) | (COMP_LOOP_acc_tmp!=2'b10);
  assign nor_378_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_934));
  assign mux_355_nl = MUX_s_1_2_2(nor_378_nl, or_tmp_934, or_952_cse);
  assign and_dcpl_641 = mux_355_nl & and_dcpl_298 & and_dcpl_639;
  assign and_dcpl_642 = and_dcpl_574 & (rem_12cyc_st_3_1_0[1]);
  assign or_957_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2!=2'b10) |
      (~ COMP_LOOP_asn_itm_2) | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp_207 = or_957_cse & or_tmp_934;
  assign nor_377_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_207));
  assign mux_356_nl = MUX_s_1_2_2(nor_377_nl, and_tmp_207, or_952_cse);
  assign and_dcpl_644 = mux_356_nl & and_dcpl_304 & and_dcpl_642;
  assign and_dcpl_645 = and_dcpl_578 & (rem_12cyc_st_4_1_0[1]);
  assign or_961_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2!=2'b10) |
      (~ COMP_LOOP_asn_itm_3) | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_209 = or_957_cse & or_961_cse & or_tmp_934;
  assign nor_376_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_209));
  assign mux_357_nl = MUX_s_1_2_2(nor_376_nl, and_tmp_209, or_952_cse);
  assign and_dcpl_647 = mux_357_nl & and_dcpl_310 & and_dcpl_645;
  assign and_dcpl_648 = and_dcpl_582 & (rem_12cyc_st_5_1_0[1]);
  assign or_966_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2!=2'b10) |
      (~ COMP_LOOP_asn_itm_4) | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_212 = or_957_cse & or_961_cse & or_966_cse & or_tmp_934;
  assign nor_375_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_212));
  assign mux_358_nl = MUX_s_1_2_2(nor_375_nl, and_tmp_212, or_952_cse);
  assign and_dcpl_650 = mux_358_nl & and_dcpl_316 & and_dcpl_648;
  assign or_972_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2!=2'b10) |
      (~ COMP_LOOP_asn_itm_5) | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_216 = or_957_cse & or_961_cse & or_966_cse & or_972_cse & or_tmp_934;
  assign nor_374_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_216));
  assign mux_359_nl = MUX_s_1_2_2(nor_374_nl, and_tmp_216, or_952_cse);
  assign and_dcpl_653 = mux_359_nl & and_dcpl_112 & and_dcpl_126 & (rem_12cyc_st_6_1_0[1]);
  assign or_979_cse = (rem_12cyc_st_6_1_0!=2'b10) | (rem_12cyc_st_6_3_2!=2'b10);
  assign nor_372_nl = ~(and_dcpl_111 | (~ or_tmp_934));
  assign mux_360_nl = MUX_s_1_2_2(nor_372_nl, or_tmp_934, or_979_cse);
  assign and_tmp_220 = or_957_cse & or_961_cse & or_966_cse & or_972_cse & mux_360_nl;
  assign nor_373_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_220));
  assign mux_361_nl = MUX_s_1_2_2(nor_373_nl, and_tmp_220, or_952_cse);
  assign and_dcpl_657 = mux_361_nl & and_dcpl_85 & and_dcpl_104 & (~ (rem_12cyc_st_7_1_0[0]));
  assign or_988_cse = (rem_12cyc_st_7_1_0!=2'b10) | (rem_12cyc_st_7_3_2!=2'b10);
  assign nor_369_nl = ~(and_dcpl_84 | (~ or_tmp_934));
  assign mux_tmp_362 = MUX_s_1_2_2(nor_369_nl, or_tmp_934, or_988_cse);
  assign nor_370_nl = ~(and_dcpl_111 | (~ mux_tmp_362));
  assign mux_363_nl = MUX_s_1_2_2(nor_370_nl, mux_tmp_362, or_979_cse);
  assign and_tmp_224 = or_957_cse & or_961_cse & or_966_cse & or_972_cse & mux_363_nl;
  assign nor_371_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_224));
  assign mux_364_nl = MUX_s_1_2_2(nor_371_nl, and_tmp_224, or_952_cse);
  assign and_dcpl_661 = mux_364_nl & and_dcpl_58 & and_dcpl_77 & (~ (rem_12cyc_st_8_1_0[0]));
  assign or_999_cse = (rem_12cyc_st_8_1_0!=2'b10) | (rem_12cyc_st_8_3_2!=2'b10);
  assign nor_365_nl = ~(and_dcpl_57 | (~ or_tmp_934));
  assign mux_tmp_365 = MUX_s_1_2_2(nor_365_nl, or_tmp_934, or_999_cse);
  assign nor_366_nl = ~(and_dcpl_84 | (~ mux_tmp_365));
  assign mux_tmp_366 = MUX_s_1_2_2(nor_366_nl, mux_tmp_365, or_988_cse);
  assign nor_367_nl = ~(and_dcpl_111 | (~ mux_tmp_366));
  assign mux_367_nl = MUX_s_1_2_2(nor_367_nl, mux_tmp_366, or_979_cse);
  assign and_tmp_228 = or_957_cse & or_961_cse & or_966_cse & or_972_cse & mux_367_nl;
  assign nor_368_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_228));
  assign mux_368_nl = MUX_s_1_2_2(nor_368_nl, and_tmp_228, or_952_cse);
  assign and_dcpl_665 = mux_368_nl & and_dcpl_31 & and_dcpl_50 & (~ (rem_12cyc_st_9_1_0[0]));
  assign nor_360_nl = ~(and_dcpl_30 | (~ or_tmp_934));
  assign or_1012_nl = (rem_12cyc_st_9_1_0!=2'b10) | (rem_12cyc_st_9_3_2!=2'b10);
  assign mux_tmp_369 = MUX_s_1_2_2(nor_360_nl, or_tmp_934, or_1012_nl);
  assign nor_361_nl = ~(and_dcpl_57 | (~ mux_tmp_369));
  assign mux_tmp_370 = MUX_s_1_2_2(nor_361_nl, mux_tmp_369, or_999_cse);
  assign nor_362_nl = ~(and_dcpl_84 | (~ mux_tmp_370));
  assign mux_tmp_371 = MUX_s_1_2_2(nor_362_nl, mux_tmp_370, or_988_cse);
  assign nor_363_nl = ~(and_dcpl_111 | (~ mux_tmp_371));
  assign mux_372_nl = MUX_s_1_2_2(nor_363_nl, mux_tmp_371, or_979_cse);
  assign and_tmp_232 = or_957_cse & or_961_cse & or_966_cse & or_972_cse & mux_372_nl;
  assign nor_364_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_232));
  assign mux_373_nl = MUX_s_1_2_2(nor_364_nl, and_tmp_232, or_952_cse);
  assign and_dcpl_669 = mux_373_nl & and_dcpl_4 & and_dcpl_23 & (~ (rem_12cyc_st_10_1_0[0]));
  assign or_tmp_1009 = (COMP_LOOP_acc_tmp!=2'b10) | (COMP_LOOP_acc_1_tmp[1:0]!=2'b10)
      | (~ ccs_ccore_start_rsci_idat);
  assign nor_351_nl = ~((rem_12cyc_st_10_3_2[1]) | (~ or_tmp_1009));
  assign or_1027_nl = (~ main_stage_0_11) | (~ COMP_LOOP_asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b10)
      | (rem_12cyc_st_10_3_2[0]);
  assign mux_tmp_374 = MUX_s_1_2_2(nor_351_nl, or_tmp_1009, or_1027_nl);
  assign nor_352_nl = ~((rem_12cyc_st_6_3_2[1]) | (~ mux_tmp_374));
  assign or_1026_nl = (~ main_stage_0_7) | (~ COMP_LOOP_asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b10)
      | (rem_12cyc_st_6_3_2[0]);
  assign mux_tmp_375 = MUX_s_1_2_2(nor_352_nl, mux_tmp_374, or_1026_nl);
  assign nor_353_nl = ~((rem_12cyc_st_5_3_2[1]) | (~ mux_tmp_375));
  assign or_1025_nl = (~ main_stage_0_6) | (~ COMP_LOOP_asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b10)
      | (rem_12cyc_st_5_3_2[0]);
  assign mux_tmp_376 = MUX_s_1_2_2(nor_353_nl, mux_tmp_375, or_1025_nl);
  assign nor_354_nl = ~((rem_12cyc_st_4_3_2[1]) | (~ mux_tmp_376));
  assign or_1024_nl = (~ main_stage_0_5) | (~ COMP_LOOP_asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b10)
      | (rem_12cyc_st_4_3_2[0]);
  assign mux_tmp_377 = MUX_s_1_2_2(nor_354_nl, mux_tmp_376, or_1024_nl);
  assign nor_355_nl = ~((rem_12cyc_st_3_3_2[1]) | (~ mux_tmp_377));
  assign or_1023_nl = (~ main_stage_0_4) | (~ COMP_LOOP_asn_itm_3) | (rem_12cyc_st_3_1_0!=2'b10)
      | (rem_12cyc_st_3_3_2[0]);
  assign mux_tmp_378 = MUX_s_1_2_2(nor_355_nl, mux_tmp_377, or_1023_nl);
  assign nor_356_nl = ~((rem_12cyc_st_2_3_2[1]) | (~ mux_tmp_378));
  assign or_1022_nl = (~ main_stage_0_3) | (~ COMP_LOOP_asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b10)
      | (rem_12cyc_st_2_3_2[0]);
  assign mux_tmp_379 = MUX_s_1_2_2(nor_356_nl, mux_tmp_378, or_1022_nl);
  assign nor_357_nl = ~((rem_12cyc_st_9_3_2[1]) | (~ mux_tmp_379));
  assign or_1021_nl = (~ main_stage_0_10) | (~ COMP_LOOP_asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b10)
      | (rem_12cyc_st_9_3_2[0]);
  assign mux_tmp_380 = MUX_s_1_2_2(nor_357_nl, mux_tmp_379, or_1021_nl);
  assign nor_358_nl = ~((rem_12cyc_st_8_3_2[1]) | (~ mux_tmp_380));
  assign or_1020_nl = (~ main_stage_0_9) | (~ COMP_LOOP_asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b10)
      | (rem_12cyc_st_8_3_2[0]);
  assign mux_tmp_381 = MUX_s_1_2_2(nor_358_nl, mux_tmp_380, or_1020_nl);
  assign nor_359_nl = ~((rem_12cyc_st_7_3_2[1]) | (~ mux_tmp_381));
  assign or_1019_nl = (~ main_stage_0_8) | (~ COMP_LOOP_asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b10)
      | (rem_12cyc_st_7_3_2[0]);
  assign mux_382_nl = MUX_s_1_2_2(nor_359_nl, mux_tmp_381, or_1019_nl);
  assign and_tmp_233 = ((~ main_stage_0_2) | (~ COMP_LOOP_asn_itm_1) | (rem_12cyc_3_2!=2'b10)
      | (rem_12cyc_1_0!=2'b10)) & mux_382_nl;
  assign and_dcpl_673 = and_dcpl_568 & and_dcpl_430;
  assign or_tmp_1021 = (~((rem_12cyc_1_0==2'b11) & (rem_12cyc_3_2==2'b10))) | not_tmp_54;
  assign nand_57_cse = ~((COMP_LOOP_acc_1_tmp[1:0]==2'b11) & (COMP_LOOP_acc_tmp==2'b10));
  assign nor_350_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_1021));
  assign mux_383_nl = MUX_s_1_2_2(nor_350_nl, or_tmp_1021, nand_57_cse);
  assign and_dcpl_675 = mux_383_nl & and_dcpl_358 & and_dcpl_639;
  assign or_1045_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2[0]);
  assign and_960_nl = nand_84_cse & or_tmp_1021;
  assign mux_tmp_384 = MUX_s_1_2_2(and_960_nl, or_tmp_1021, or_1045_cse);
  assign nor_349_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_384));
  assign mux_385_nl = MUX_s_1_2_2(nor_349_nl, mux_tmp_384, nand_57_cse);
  assign and_dcpl_677 = mux_385_nl & and_dcpl_362 & and_dcpl_642;
  assign or_1050_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2!=2'b10);
  assign and_958_nl = nand_274_cse & or_tmp_1021;
  assign mux_tmp_386 = MUX_s_1_2_2(and_958_nl, or_tmp_1021, or_1050_cse);
  assign and_959_nl = nand_84_cse & mux_tmp_386;
  assign mux_tmp_387 = MUX_s_1_2_2(and_959_nl, mux_tmp_386, or_1045_cse);
  assign nor_348_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_387));
  assign mux_388_nl = MUX_s_1_2_2(nor_348_nl, mux_tmp_387, nand_57_cse);
  assign and_dcpl_679 = mux_388_nl & and_dcpl_366 & and_dcpl_645;
  assign or_1057_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2[0]);
  assign and_955_nl = nand_79_cse & or_tmp_1021;
  assign mux_tmp_389 = MUX_s_1_2_2(and_955_nl, or_tmp_1021, or_1057_cse);
  assign and_956_nl = nand_274_cse & mux_tmp_389;
  assign mux_tmp_390 = MUX_s_1_2_2(and_956_nl, mux_tmp_389, or_1050_cse);
  assign and_957_nl = nand_84_cse & mux_tmp_390;
  assign mux_tmp_391 = MUX_s_1_2_2(and_957_nl, mux_tmp_390, or_1045_cse);
  assign nor_347_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_391));
  assign mux_392_nl = MUX_s_1_2_2(nor_347_nl, mux_tmp_391, nand_57_cse);
  assign and_dcpl_681 = mux_392_nl & and_dcpl_370 & and_dcpl_648;
  assign or_1066_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2!=2'b10);
  assign and_951_nl = nand_267_cse & or_tmp_1021;
  assign mux_tmp_393 = MUX_s_1_2_2(and_951_nl, or_tmp_1021, or_1066_cse);
  assign and_952_nl = nand_79_cse & mux_tmp_393;
  assign mux_tmp_394 = MUX_s_1_2_2(and_952_nl, mux_tmp_393, or_1057_cse);
  assign and_953_nl = nand_274_cse & mux_tmp_394;
  assign mux_tmp_395 = MUX_s_1_2_2(and_953_nl, mux_tmp_394, or_1050_cse);
  assign and_954_nl = nand_84_cse & mux_tmp_395;
  assign mux_tmp_396 = MUX_s_1_2_2(and_954_nl, mux_tmp_395, or_1045_cse);
  assign nor_346_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_396));
  assign mux_397_nl = MUX_s_1_2_2(nor_346_nl, mux_tmp_396, nand_57_cse);
  assign and_dcpl_684 = mux_397_nl & and_dcpl_112 & and_dcpl_129 & (rem_12cyc_st_6_1_0[1]);
  assign nand_36_cse = ~((rem_12cyc_st_6_1_0==2'b11) & (rem_12cyc_st_6_3_2==2'b10));
  assign nor_344_nl = ~(and_dcpl_111 | (~ or_tmp_1021));
  assign mux_tmp_398 = MUX_s_1_2_2(nor_344_nl, or_tmp_1021, nand_36_cse);
  assign and_947_nl = nand_267_cse & mux_tmp_398;
  assign mux_tmp_399 = MUX_s_1_2_2(and_947_nl, mux_tmp_398, or_1066_cse);
  assign and_948_nl = nand_79_cse & mux_tmp_399;
  assign mux_tmp_400 = MUX_s_1_2_2(and_948_nl, mux_tmp_399, or_1057_cse);
  assign and_949_nl = nand_274_cse & mux_tmp_400;
  assign mux_tmp_401 = MUX_s_1_2_2(and_949_nl, mux_tmp_400, or_1050_cse);
  assign and_950_nl = nand_84_cse & mux_tmp_401;
  assign mux_tmp_402 = MUX_s_1_2_2(and_950_nl, mux_tmp_401, or_1045_cse);
  assign nor_345_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_402));
  assign mux_403_nl = MUX_s_1_2_2(nor_345_nl, mux_tmp_402, nand_57_cse);
  assign and_dcpl_687 = mux_403_nl & and_dcpl_85 & and_dcpl_104 & (rem_12cyc_st_7_1_0[0]);
  assign nand_29_cse = ~((rem_12cyc_st_7_1_0==2'b11) & (rem_12cyc_st_7_3_2==2'b10));
  assign nor_341_nl = ~(and_dcpl_84 | (~ or_tmp_1021));
  assign mux_tmp_404 = MUX_s_1_2_2(nor_341_nl, or_tmp_1021, nand_29_cse);
  assign nor_342_nl = ~(and_dcpl_111 | (~ mux_tmp_404));
  assign mux_tmp_405 = MUX_s_1_2_2(nor_342_nl, mux_tmp_404, nand_36_cse);
  assign and_943_nl = nand_267_cse & mux_tmp_405;
  assign mux_tmp_406 = MUX_s_1_2_2(and_943_nl, mux_tmp_405, or_1066_cse);
  assign and_944_nl = nand_79_cse & mux_tmp_406;
  assign mux_tmp_407 = MUX_s_1_2_2(and_944_nl, mux_tmp_406, or_1057_cse);
  assign and_945_nl = nand_274_cse & mux_tmp_407;
  assign mux_tmp_408 = MUX_s_1_2_2(and_945_nl, mux_tmp_407, or_1050_cse);
  assign and_946_nl = nand_84_cse & mux_tmp_408;
  assign mux_tmp_409 = MUX_s_1_2_2(and_946_nl, mux_tmp_408, or_1045_cse);
  assign nor_343_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_409));
  assign mux_410_nl = MUX_s_1_2_2(nor_343_nl, mux_tmp_409, nand_57_cse);
  assign and_dcpl_690 = mux_410_nl & and_dcpl_58 & and_dcpl_77 & (rem_12cyc_st_8_1_0[0]);
  assign nand_21_cse = ~((rem_12cyc_st_8_1_0==2'b11) & (rem_12cyc_st_8_3_2==2'b10));
  assign nor_337_nl = ~(and_dcpl_57 | (~ or_tmp_1021));
  assign mux_tmp_411 = MUX_s_1_2_2(nor_337_nl, or_tmp_1021, nand_21_cse);
  assign nor_338_nl = ~(and_dcpl_84 | (~ mux_tmp_411));
  assign mux_tmp_412 = MUX_s_1_2_2(nor_338_nl, mux_tmp_411, nand_29_cse);
  assign nor_339_nl = ~(and_dcpl_111 | (~ mux_tmp_412));
  assign mux_tmp_413 = MUX_s_1_2_2(nor_339_nl, mux_tmp_412, nand_36_cse);
  assign and_939_nl = nand_267_cse & mux_tmp_413;
  assign mux_tmp_414 = MUX_s_1_2_2(and_939_nl, mux_tmp_413, or_1066_cse);
  assign and_940_nl = nand_79_cse & mux_tmp_414;
  assign mux_tmp_415 = MUX_s_1_2_2(and_940_nl, mux_tmp_414, or_1057_cse);
  assign and_941_nl = nand_274_cse & mux_tmp_415;
  assign mux_tmp_416 = MUX_s_1_2_2(and_941_nl, mux_tmp_415, or_1050_cse);
  assign and_942_nl = nand_84_cse & mux_tmp_416;
  assign mux_tmp_417 = MUX_s_1_2_2(and_942_nl, mux_tmp_416, or_1045_cse);
  assign nor_340_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_417));
  assign mux_418_nl = MUX_s_1_2_2(nor_340_nl, mux_tmp_417, nand_57_cse);
  assign and_dcpl_693 = mux_418_nl & and_dcpl_31 & and_dcpl_50 & (rem_12cyc_st_9_1_0[0]);
  assign nor_332_nl = ~(and_dcpl_30 | (~ or_tmp_1021));
  assign nand_12_nl = ~((rem_12cyc_st_9_1_0==2'b11) & (rem_12cyc_st_9_3_2==2'b10));
  assign mux_tmp_419 = MUX_s_1_2_2(nor_332_nl, or_tmp_1021, nand_12_nl);
  assign nor_333_nl = ~(and_dcpl_57 | (~ mux_tmp_419));
  assign mux_tmp_420 = MUX_s_1_2_2(nor_333_nl, mux_tmp_419, nand_21_cse);
  assign nor_334_nl = ~(and_dcpl_84 | (~ mux_tmp_420));
  assign mux_tmp_421 = MUX_s_1_2_2(nor_334_nl, mux_tmp_420, nand_29_cse);
  assign nor_335_nl = ~(and_dcpl_111 | (~ mux_tmp_421));
  assign mux_tmp_422 = MUX_s_1_2_2(nor_335_nl, mux_tmp_421, nand_36_cse);
  assign and_935_nl = nand_267_cse & mux_tmp_422;
  assign mux_tmp_423 = MUX_s_1_2_2(and_935_nl, mux_tmp_422, or_1066_cse);
  assign and_936_nl = nand_79_cse & mux_tmp_423;
  assign mux_tmp_424 = MUX_s_1_2_2(and_936_nl, mux_tmp_423, or_1057_cse);
  assign and_937_nl = nand_274_cse & mux_tmp_424;
  assign mux_tmp_425 = MUX_s_1_2_2(and_937_nl, mux_tmp_424, or_1050_cse);
  assign and_938_nl = nand_84_cse & mux_tmp_425;
  assign mux_tmp_426 = MUX_s_1_2_2(and_938_nl, mux_tmp_425, or_1045_cse);
  assign nor_336_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_426));
  assign mux_427_nl = MUX_s_1_2_2(nor_336_nl, mux_tmp_426, nand_57_cse);
  assign and_dcpl_696 = mux_427_nl & and_dcpl_4 & and_dcpl_23 & (rem_12cyc_st_10_1_0[0]);
  assign or_tmp_1122 = (COMP_LOOP_acc_tmp!=2'b10) | nand_222_cse;
  assign nor_323_nl = ~((rem_12cyc_st_10_3_2[1]) | (~ or_tmp_1122));
  assign nand_1_nl = ~(main_stage_0_11 & COMP_LOOP_asn_itm_10 & (rem_12cyc_st_10_1_0==2'b11)
      & (~ (rem_12cyc_st_10_3_2[0])));
  assign mux_tmp_428 = MUX_s_1_2_2(nor_323_nl, or_tmp_1122, nand_1_nl);
  assign nor_324_nl = ~((rem_12cyc_st_6_3_2[1]) | (~ mux_tmp_428));
  assign nand_2_nl = ~(main_stage_0_7 & COMP_LOOP_asn_itm_6 & (rem_12cyc_st_6_1_0==2'b11)
      & (~ (rem_12cyc_st_6_3_2[0])));
  assign mux_tmp_429 = MUX_s_1_2_2(nor_324_nl, mux_tmp_428, nand_2_nl);
  assign nor_325_nl = ~((rem_12cyc_st_5_3_2[1]) | (~ mux_tmp_429));
  assign nand_3_nl = ~(main_stage_0_6 & COMP_LOOP_asn_itm_5 & (rem_12cyc_st_5_1_0==2'b11)
      & (~ (rem_12cyc_st_5_3_2[0])));
  assign mux_tmp_430 = MUX_s_1_2_2(nor_325_nl, mux_tmp_429, nand_3_nl);
  assign nor_326_nl = ~((rem_12cyc_st_4_3_2[1]) | (~ mux_tmp_430));
  assign nand_4_nl = ~(main_stage_0_5 & COMP_LOOP_asn_itm_4 & (rem_12cyc_st_4_1_0==2'b11)
      & (~ (rem_12cyc_st_4_3_2[0])));
  assign mux_tmp_431 = MUX_s_1_2_2(nor_326_nl, mux_tmp_430, nand_4_nl);
  assign nor_327_nl = ~((rem_12cyc_st_3_3_2[1]) | (~ mux_tmp_431));
  assign nand_5_nl = ~(main_stage_0_4 & COMP_LOOP_asn_itm_3 & (rem_12cyc_st_3_1_0==2'b11)
      & (~ (rem_12cyc_st_3_3_2[0])));
  assign mux_tmp_432 = MUX_s_1_2_2(nor_327_nl, mux_tmp_431, nand_5_nl);
  assign nor_328_nl = ~((rem_12cyc_st_2_3_2[1]) | (~ mux_tmp_432));
  assign nand_6_nl = ~(main_stage_0_3 & COMP_LOOP_asn_itm_2 & (rem_12cyc_st_2_1_0==2'b11)
      & (~ (rem_12cyc_st_2_3_2[0])));
  assign mux_tmp_433 = MUX_s_1_2_2(nor_328_nl, mux_tmp_432, nand_6_nl);
  assign nor_329_nl = ~((rem_12cyc_st_9_3_2[1]) | (~ mux_tmp_433));
  assign nand_7_nl = ~(main_stage_0_10 & COMP_LOOP_asn_itm_9 & (rem_12cyc_st_9_1_0==2'b11)
      & (~ (rem_12cyc_st_9_3_2[0])));
  assign mux_tmp_434 = MUX_s_1_2_2(nor_329_nl, mux_tmp_433, nand_7_nl);
  assign nor_330_nl = ~((rem_12cyc_st_8_3_2[1]) | (~ mux_tmp_434));
  assign nand_8_nl = ~(main_stage_0_9 & COMP_LOOP_asn_itm_8 & (rem_12cyc_st_8_1_0==2'b11)
      & (~ (rem_12cyc_st_8_3_2[0])));
  assign mux_tmp_435 = MUX_s_1_2_2(nor_330_nl, mux_tmp_434, nand_8_nl);
  assign nor_331_nl = ~((rem_12cyc_st_7_3_2[1]) | (~ mux_tmp_435));
  assign nand_9_nl = ~(main_stage_0_8 & COMP_LOOP_asn_itm_7 & (rem_12cyc_st_7_1_0==2'b11)
      & (~ (rem_12cyc_st_7_3_2[0])));
  assign mux_tmp_436 = MUX_s_1_2_2(nor_331_nl, mux_tmp_435, nand_9_nl);
  assign and_934_nl = nand_223_cse & mux_tmp_436;
  assign nand_11_nl = ~(main_stage_0_2 & COMP_LOOP_asn_itm_1 & (rem_12cyc_3_2==2'b10));
  assign mux_tmp_437 = MUX_s_1_2_2(and_934_nl, mux_tmp_436, nand_11_nl);
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_en ) begin
      return_rsci_d <= MUX_v_64_2_2(result_sva_duc_mx0, qelse_acc_nl, mux_11_nl);
      m_buf_sva_12 <= m_buf_sva_11;
      m_buf_sva_11 <= m_buf_sva_10;
      m_buf_sva_10 <= m_buf_sva_9;
      m_buf_sva_9 <= m_buf_sva_8;
      m_buf_sva_8 <= m_buf_sva_7;
      m_buf_sva_7 <= m_buf_sva_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      COMP_LOOP_asn_itm_12 <= 1'b0;
      COMP_LOOP_asn_itm_11 <= 1'b0;
      COMP_LOOP_asn_itm_10 <= 1'b0;
      COMP_LOOP_asn_itm_9 <= 1'b0;
      COMP_LOOP_asn_itm_8 <= 1'b0;
      COMP_LOOP_asn_itm_7 <= 1'b0;
      COMP_LOOP_asn_itm_6 <= 1'b0;
      COMP_LOOP_asn_itm_5 <= 1'b0;
      COMP_LOOP_asn_itm_4 <= 1'b0;
      COMP_LOOP_asn_itm_3 <= 1'b0;
      COMP_LOOP_asn_itm_2 <= 1'b0;
      COMP_LOOP_asn_itm_1 <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
      main_stage_0_5 <= 1'b0;
      main_stage_0_6 <= 1'b0;
      main_stage_0_7 <= 1'b0;
      main_stage_0_8 <= 1'b0;
      main_stage_0_9 <= 1'b0;
      main_stage_0_10 <= 1'b0;
      main_stage_0_11 <= 1'b0;
      main_stage_0_12 <= 1'b0;
      main_stage_0_13 <= 1'b0;
    end
    else if ( ccs_ccore_en ) begin
      COMP_LOOP_asn_itm_12 <= COMP_LOOP_asn_itm_11;
      COMP_LOOP_asn_itm_11 <= COMP_LOOP_asn_itm_10;
      COMP_LOOP_asn_itm_10 <= COMP_LOOP_asn_itm_9;
      COMP_LOOP_asn_itm_9 <= COMP_LOOP_asn_itm_8;
      COMP_LOOP_asn_itm_8 <= COMP_LOOP_asn_itm_7;
      COMP_LOOP_asn_itm_7 <= COMP_LOOP_asn_itm_6;
      COMP_LOOP_asn_itm_6 <= COMP_LOOP_asn_itm_5;
      COMP_LOOP_asn_itm_5 <= COMP_LOOP_asn_itm_4;
      COMP_LOOP_asn_itm_4 <= COMP_LOOP_asn_itm_3;
      COMP_LOOP_asn_itm_3 <= COMP_LOOP_asn_itm_2;
      COMP_LOOP_asn_itm_2 <= COMP_LOOP_asn_itm_1;
      COMP_LOOP_asn_itm_1 <= ccs_ccore_start_rsci_idat;
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
      main_stage_0_4 <= main_stage_0_3;
      main_stage_0_5 <= main_stage_0_4;
      main_stage_0_6 <= main_stage_0_5;
      main_stage_0_7 <= main_stage_0_6;
      main_stage_0_8 <= main_stage_0_7;
      main_stage_0_9 <= main_stage_0_8;
      main_stage_0_10 <= main_stage_0_9;
      main_stage_0_11 <= main_stage_0_10;
      main_stage_0_12 <= main_stage_0_11;
      main_stage_0_13 <= main_stage_0_12;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_sva_duc <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( COMP_LOOP_asn_itm_12 & main_stage_0_13 & ccs_ccore_en & (~((rem_12cyc_st_12_3_2==2'b11)))
        ) begin
      result_sva_duc <= result_sva_duc_mx0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_12_3_2 <= 2'b00;
      rem_12cyc_st_12_1_0 <= 2'b00;
    end
    else if ( COMP_LOOP_and_26_cse ) begin
      rem_12cyc_st_12_3_2 <= rem_12cyc_st_11_3_2;
      rem_12cyc_st_12_1_0 <= rem_12cyc_st_11_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_cse ) begin
      rem_12_cmp_1_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_3_2_63_0, mut_3_3_63_0,
          mut_3_4_63_0, mut_3_5_63_0, mut_3_6_63_0, mut_3_7_63_0, mut_3_8_63_0, mut_3_9_63_0,
          mut_3_10_63_0, mut_3_11_63_0, {and_dcpl_294 , and_dcpl_300 , and_dcpl_306
          , and_dcpl_312 , and_dcpl_318 , and_dcpl_324 , and_dcpl_330 , and_dcpl_336
          , and_dcpl_342 , and_dcpl_348 , and_tmp_35});
      rem_12_cmp_1_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_2_2_63_0, mut_2_3_63_0,
          mut_2_4_63_0, mut_2_5_63_0, mut_2_6_63_0, mut_2_7_63_0, mut_2_8_63_0, mut_2_9_63_0,
          mut_2_10_63_0, mut_2_11_63_0, {and_dcpl_294 , and_dcpl_300 , and_dcpl_306
          , and_dcpl_312 , and_dcpl_318 , and_dcpl_324 , and_dcpl_330 , and_dcpl_336
          , and_dcpl_342 , and_dcpl_348 , and_tmp_35});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_2_cse ) begin
      rem_12_cmp_2_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_5_2_63_0, mut_5_3_63_0,
          mut_5_4_63_0, mut_5_5_63_0, mut_5_6_63_0, mut_5_7_63_0, mut_5_8_63_0, mut_5_9_63_0,
          mut_5_10_63_0, mut_5_11_63_0, {and_dcpl_356 , and_dcpl_360 , and_dcpl_364
          , and_dcpl_368 , and_dcpl_372 , and_dcpl_376 , and_dcpl_379 , and_dcpl_382
          , and_dcpl_385 , and_dcpl_388 , mux_tmp_76});
      rem_12_cmp_2_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_4_2_63_0, mut_4_3_63_0,
          mut_4_4_63_0, mut_4_5_63_0, mut_4_6_63_0, mut_4_7_63_0, mut_4_8_63_0, mut_4_9_63_0,
          mut_4_10_63_0, mut_4_11_63_0, {and_dcpl_356 , and_dcpl_360 , and_dcpl_364
          , and_dcpl_368 , and_dcpl_372 , and_dcpl_376 , and_dcpl_379 , and_dcpl_382
          , and_dcpl_385 , and_dcpl_388 , mux_tmp_76});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_4_cse ) begin
      rem_12_cmp_3_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_7_2_63_0, mut_7_3_63_0,
          mut_7_4_63_0, mut_7_5_63_0, mut_7_6_63_0, mut_7_7_63_0, mut_7_8_63_0, mut_7_9_63_0,
          mut_7_10_63_0, mut_7_11_63_0, {and_dcpl_394 , and_dcpl_397 , and_dcpl_400
          , and_dcpl_403 , and_dcpl_406 , and_dcpl_409 , and_dcpl_413 , and_dcpl_417
          , and_dcpl_421 , and_dcpl_425 , and_tmp_80});
      rem_12_cmp_3_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_6_2_63_0, mut_6_3_63_0,
          mut_6_4_63_0, mut_6_5_63_0, mut_6_6_63_0, mut_6_7_63_0, mut_6_8_63_0, mut_6_9_63_0,
          mut_6_10_63_0, mut_6_11_63_0, {and_dcpl_394 , and_dcpl_397 , and_dcpl_400
          , and_dcpl_403 , and_dcpl_406 , and_dcpl_409 , and_dcpl_413 , and_dcpl_417
          , and_dcpl_421 , and_dcpl_425 , and_tmp_80});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_6_cse ) begin
      rem_12_cmp_4_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_9_2_63_0, mut_9_3_63_0,
          mut_9_4_63_0, mut_9_5_63_0, mut_9_6_63_0, mut_9_7_63_0, mut_9_8_63_0, mut_9_9_63_0,
          mut_9_10_63_0, mut_9_11_63_0, {and_dcpl_431 , and_dcpl_433 , and_dcpl_435
          , and_dcpl_437 , and_dcpl_439 , and_dcpl_442 , and_dcpl_445 , and_dcpl_448
          , and_dcpl_451 , and_dcpl_454 , mux_tmp_141});
      rem_12_cmp_4_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_8_2_63_0, mut_8_3_63_0,
          mut_8_4_63_0, mut_8_5_63_0, mut_8_6_63_0, mut_8_7_63_0, mut_8_8_63_0, mut_8_9_63_0,
          mut_8_10_63_0, mut_8_11_63_0, {and_dcpl_431 , and_dcpl_433 , and_dcpl_435
          , and_dcpl_437 , and_dcpl_439 , and_dcpl_442 , and_dcpl_445 , and_dcpl_448
          , and_dcpl_451 , and_dcpl_454 , mux_tmp_141});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_8_cse ) begin
      rem_12_cmp_5_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_11_2_63_0, mut_11_3_63_0,
          mut_11_4_63_0, mut_11_5_63_0, mut_11_6_63_0, mut_11_7_63_0, mut_11_8_63_0,
          mut_11_9_63_0, mut_11_10_63_0, mut_11_11_63_0, {and_dcpl_461 , and_dcpl_465
          , and_dcpl_469 , and_dcpl_473 , and_dcpl_477 , and_dcpl_480 , and_dcpl_483
          , and_dcpl_486 , and_dcpl_489 , and_dcpl_492 , and_tmp_125});
      rem_12_cmp_5_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_10_2_63_0, mut_10_3_63_0,
          mut_10_4_63_0, mut_10_5_63_0, mut_10_6_63_0, mut_10_7_63_0, mut_10_8_63_0,
          mut_10_9_63_0, mut_10_10_63_0, mut_10_11_63_0, {and_dcpl_461 , and_dcpl_465
          , and_dcpl_469 , and_dcpl_473 , and_dcpl_477 , and_dcpl_480 , and_dcpl_483
          , and_dcpl_486 , and_dcpl_489 , and_dcpl_492 , and_tmp_125});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_10_cse ) begin
      rem_12_cmp_6_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_13_2_63_0, mut_13_3_63_0,
          mut_13_4_63_0, mut_13_5_63_0, mut_13_6_63_0, mut_13_7_63_0, mut_13_8_63_0,
          mut_13_9_63_0, mut_13_10_63_0, mut_13_11_63_0, {and_dcpl_498 , and_dcpl_500
          , and_dcpl_502 , and_dcpl_504 , and_dcpl_506 , and_dcpl_508 , and_dcpl_510
          , and_dcpl_512 , and_dcpl_514 , and_dcpl_516 , mux_tmp_206});
      rem_12_cmp_6_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_12_2_63_0, mut_12_3_63_0,
          mut_12_4_63_0, mut_12_5_63_0, mut_12_6_63_0, mut_12_7_63_0, mut_12_8_63_0,
          mut_12_9_63_0, mut_12_10_63_0, mut_12_11_63_0, {and_dcpl_498 , and_dcpl_500
          , and_dcpl_502 , and_dcpl_504 , and_dcpl_506 , and_dcpl_508 , and_dcpl_510
          , and_dcpl_512 , and_dcpl_514 , and_dcpl_516 , mux_tmp_206});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_12_cse ) begin
      rem_12_cmp_7_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_15_2_63_0, mut_15_3_63_0,
          mut_15_4_63_0, mut_15_5_63_0, mut_15_6_63_0, mut_15_7_63_0, mut_15_8_63_0,
          mut_15_9_63_0, mut_15_10_63_0, mut_15_11_63_0, {and_dcpl_520 , and_dcpl_523
          , and_dcpl_526 , and_dcpl_529 , and_dcpl_532 , and_dcpl_534 , and_dcpl_536
          , and_dcpl_538 , and_dcpl_540 , and_dcpl_542 , and_tmp_170});
      rem_12_cmp_7_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_14_2_63_0, mut_14_3_63_0,
          mut_14_4_63_0, mut_14_5_63_0, mut_14_6_63_0, mut_14_7_63_0, mut_14_8_63_0,
          mut_14_9_63_0, mut_14_10_63_0, mut_14_11_63_0, {and_dcpl_520 , and_dcpl_523
          , and_dcpl_526 , and_dcpl_529 , and_dcpl_532 , and_dcpl_534 , and_dcpl_536
          , and_dcpl_538 , and_dcpl_540 , and_dcpl_542 , and_tmp_170});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_14_cse ) begin
      rem_12_cmp_8_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_17_2_63_0, mut_17_3_63_0,
          mut_17_4_63_0, mut_17_5_63_0, mut_17_6_63_0, mut_17_7_63_0, mut_17_8_63_0,
          mut_17_9_63_0, mut_17_10_63_0, mut_17_11_63_0, {and_dcpl_546 , and_dcpl_548
          , and_dcpl_550 , and_dcpl_552 , and_dcpl_554 , and_dcpl_556 , and_dcpl_558
          , and_dcpl_560 , and_dcpl_562 , and_dcpl_564 , mux_tmp_271});
      rem_12_cmp_8_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_16_2_63_0, mut_16_3_63_0,
          mut_16_4_63_0, mut_16_5_63_0, mut_16_6_63_0, mut_16_7_63_0, mut_16_8_63_0,
          mut_16_9_63_0, mut_16_10_63_0, mut_16_11_63_0, {and_dcpl_546 , and_dcpl_548
          , and_dcpl_550 , and_dcpl_552 , and_dcpl_554 , and_dcpl_556 , and_dcpl_558
          , and_dcpl_560 , and_dcpl_562 , and_dcpl_564 , mux_tmp_271});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_16_cse ) begin
      rem_12_cmp_9_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_19_2_63_0, mut_19_3_63_0,
          mut_19_4_63_0, mut_19_5_63_0, mut_19_6_63_0, mut_19_7_63_0, mut_19_8_63_0,
          mut_19_9_63_0, mut_19_10_63_0, mut_19_11_63_0, {and_dcpl_569 , and_dcpl_573
          , and_dcpl_577 , and_dcpl_581 , and_dcpl_585 , and_dcpl_589 , and_dcpl_593
          , and_dcpl_597 , and_dcpl_601 , and_dcpl_605 , and_tmp_206});
      rem_12_cmp_9_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_18_2_63_0, mut_18_3_63_0,
          mut_18_4_63_0, mut_18_5_63_0, mut_18_6_63_0, mut_18_7_63_0, mut_18_8_63_0,
          mut_18_9_63_0, mut_18_10_63_0, mut_18_11_63_0, {and_dcpl_569 , and_dcpl_573
          , and_dcpl_577 , and_dcpl_581 , and_dcpl_585 , and_dcpl_589 , and_dcpl_593
          , and_dcpl_597 , and_dcpl_601 , and_dcpl_605 , and_tmp_206});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_18_cse ) begin
      rem_12_cmp_10_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_21_2_63_0, mut_21_3_63_0,
          mut_21_4_63_0, mut_21_5_63_0, mut_21_6_63_0, mut_21_7_63_0, mut_21_8_63_0,
          mut_21_9_63_0, mut_21_10_63_0, mut_21_11_63_0, {and_dcpl_610 , and_dcpl_612
          , and_dcpl_614 , and_dcpl_616 , and_dcpl_618 , and_dcpl_622 , and_dcpl_625
          , and_dcpl_628 , and_dcpl_631 , and_dcpl_634 , mux_tmp_354});
      rem_12_cmp_10_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_20_2_63_0, mut_20_3_63_0,
          mut_20_4_63_0, mut_20_5_63_0, mut_20_6_63_0, mut_20_7_63_0, mut_20_8_63_0,
          mut_20_9_63_0, mut_20_10_63_0, mut_20_11_63_0, {and_dcpl_610 , and_dcpl_612
          , and_dcpl_614 , and_dcpl_616 , and_dcpl_618 , and_dcpl_622 , and_dcpl_625
          , and_dcpl_628 , and_dcpl_631 , and_dcpl_634 , mux_tmp_354});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_20_cse ) begin
      rem_12_cmp_11_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_23_2_63_0, mut_23_3_63_0,
          mut_23_4_63_0, mut_23_5_63_0, mut_23_6_63_0, mut_23_7_63_0, mut_23_8_63_0,
          mut_23_9_63_0, mut_23_10_63_0, mut_23_11_63_0, {and_dcpl_638 , and_dcpl_641
          , and_dcpl_644 , and_dcpl_647 , and_dcpl_650 , and_dcpl_653 , and_dcpl_657
          , and_dcpl_661 , and_dcpl_665 , and_dcpl_669 , and_tmp_233});
      rem_12_cmp_11_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_22_2_63_0, mut_22_3_63_0,
          mut_22_4_63_0, mut_22_5_63_0, mut_22_6_63_0, mut_22_7_63_0, mut_22_8_63_0,
          mut_22_9_63_0, mut_22_10_63_0, mut_22_11_63_0, {and_dcpl_638 , and_dcpl_641
          , and_dcpl_644 , and_dcpl_647 , and_dcpl_650 , and_dcpl_653 , and_dcpl_657
          , and_dcpl_661 , and_dcpl_665 , and_dcpl_669 , and_tmp_233});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_22_cse ) begin
      rem_12_cmp_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_1_2_63_0, mut_1_3_63_0,
          mut_1_4_63_0, mut_1_5_63_0, mut_1_6_63_0, mut_1_7_63_0, mut_1_8_63_0, mut_1_9_63_0,
          mut_1_10_63_0, mut_1_11_63_0, {and_dcpl_673 , and_dcpl_675 , and_dcpl_677
          , and_dcpl_679 , and_dcpl_681 , and_dcpl_684 , and_dcpl_687 , and_dcpl_690
          , and_dcpl_693 , and_dcpl_696 , mux_tmp_437});
      rem_12_cmp_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_2_63_0, mut_3_63_0,
          mut_4_63_0, mut_5_63_0, mut_6_63_0, mut_7_63_0, mut_8_63_0, mut_9_63_0,
          mut_10_63_0, mut_11_63_0, {and_dcpl_673 , and_dcpl_675 , and_dcpl_677 ,
          and_dcpl_679 , and_dcpl_681 , and_dcpl_684 , and_dcpl_687 , and_dcpl_690
          , and_dcpl_693 , and_dcpl_696 , mux_tmp_437});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_28_cse ) begin
      mut_3_11_63_0 <= mut_3_10_63_0;
      mut_2_11_63_0 <= mut_2_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_30_cse ) begin
      mut_5_11_63_0 <= mut_5_10_63_0;
      mut_4_11_63_0 <= mut_4_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_32_cse ) begin
      mut_7_11_63_0 <= mut_7_10_63_0;
      mut_6_11_63_0 <= mut_6_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_34_cse ) begin
      mut_9_11_63_0 <= mut_9_10_63_0;
      mut_8_11_63_0 <= mut_8_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_36_cse ) begin
      mut_11_11_63_0 <= mut_11_10_63_0;
      mut_10_11_63_0 <= mut_10_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_38_cse ) begin
      mut_13_11_63_0 <= mut_13_10_63_0;
      mut_12_11_63_0 <= mut_12_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_40_cse ) begin
      mut_15_11_63_0 <= mut_15_10_63_0;
      mut_14_11_63_0 <= mut_14_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_42_cse ) begin
      mut_17_11_63_0 <= mut_17_10_63_0;
      mut_16_11_63_0 <= mut_16_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_44_cse ) begin
      mut_19_11_63_0 <= mut_19_10_63_0;
      mut_18_11_63_0 <= mut_18_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_46_cse ) begin
      mut_21_11_63_0 <= mut_21_10_63_0;
      mut_20_11_63_0 <= mut_20_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_48_cse ) begin
      mut_23_11_63_0 <= mut_23_10_63_0;
      mut_22_11_63_0 <= mut_22_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_50_cse ) begin
      mut_1_11_63_0 <= mut_1_10_63_0;
      mut_11_63_0 <= mut_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_11_3_2 <= 2'b00;
      rem_12cyc_st_11_1_0 <= 2'b00;
    end
    else if ( COMP_LOOP_and_52_cse ) begin
      rem_12cyc_st_11_3_2 <= rem_12cyc_st_10_3_2;
      rem_12cyc_st_11_1_0 <= rem_12cyc_st_10_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_54_cse ) begin
      mut_3_10_63_0 <= mut_3_9_63_0;
      mut_2_10_63_0 <= mut_2_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_56_cse ) begin
      mut_5_10_63_0 <= mut_5_9_63_0;
      mut_4_10_63_0 <= mut_4_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_58_cse ) begin
      mut_7_10_63_0 <= mut_7_9_63_0;
      mut_6_10_63_0 <= mut_6_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_60_cse ) begin
      mut_9_10_63_0 <= mut_9_9_63_0;
      mut_8_10_63_0 <= mut_8_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_62_cse ) begin
      mut_11_10_63_0 <= mut_11_9_63_0;
      mut_10_10_63_0 <= mut_10_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_64_cse ) begin
      mut_13_10_63_0 <= mut_13_9_63_0;
      mut_12_10_63_0 <= mut_12_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_66_cse ) begin
      mut_15_10_63_0 <= mut_15_9_63_0;
      mut_14_10_63_0 <= mut_14_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_68_cse ) begin
      mut_17_10_63_0 <= mut_17_9_63_0;
      mut_16_10_63_0 <= mut_16_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_70_cse ) begin
      mut_19_10_63_0 <= mut_19_9_63_0;
      mut_18_10_63_0 <= mut_18_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_72_cse ) begin
      mut_21_10_63_0 <= mut_21_9_63_0;
      mut_20_10_63_0 <= mut_20_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_74_cse ) begin
      mut_23_10_63_0 <= mut_23_9_63_0;
      mut_22_10_63_0 <= mut_22_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_76_cse ) begin
      mut_1_10_63_0 <= mut_1_9_63_0;
      mut_10_63_0 <= mut_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_10_3_2 <= 2'b00;
      rem_12cyc_st_10_1_0 <= 2'b00;
    end
    else if ( COMP_LOOP_and_78_cse ) begin
      rem_12cyc_st_10_3_2 <= rem_12cyc_st_9_3_2;
      rem_12cyc_st_10_1_0 <= rem_12cyc_st_9_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_80_cse ) begin
      mut_3_9_63_0 <= mut_3_8_63_0;
      mut_2_9_63_0 <= mut_2_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_82_cse ) begin
      mut_5_9_63_0 <= mut_5_8_63_0;
      mut_4_9_63_0 <= mut_4_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_84_cse ) begin
      mut_7_9_63_0 <= mut_7_8_63_0;
      mut_6_9_63_0 <= mut_6_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_86_cse ) begin
      mut_9_9_63_0 <= mut_9_8_63_0;
      mut_8_9_63_0 <= mut_8_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_88_cse ) begin
      mut_11_9_63_0 <= mut_11_8_63_0;
      mut_10_9_63_0 <= mut_10_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_90_cse ) begin
      mut_13_9_63_0 <= mut_13_8_63_0;
      mut_12_9_63_0 <= mut_12_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_92_cse ) begin
      mut_15_9_63_0 <= mut_15_8_63_0;
      mut_14_9_63_0 <= mut_14_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_94_cse ) begin
      mut_17_9_63_0 <= mut_17_8_63_0;
      mut_16_9_63_0 <= mut_16_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_96_cse ) begin
      mut_19_9_63_0 <= mut_19_8_63_0;
      mut_18_9_63_0 <= mut_18_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_98_cse ) begin
      mut_21_9_63_0 <= mut_21_8_63_0;
      mut_20_9_63_0 <= mut_20_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_100_cse ) begin
      mut_23_9_63_0 <= mut_23_8_63_0;
      mut_22_9_63_0 <= mut_22_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_102_cse ) begin
      mut_1_9_63_0 <= mut_1_8_63_0;
      mut_9_63_0 <= mut_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_9_3_2 <= 2'b00;
      rem_12cyc_st_9_1_0 <= 2'b00;
    end
    else if ( COMP_LOOP_and_104_cse ) begin
      rem_12cyc_st_9_3_2 <= rem_12cyc_st_8_3_2;
      rem_12cyc_st_9_1_0 <= rem_12cyc_st_8_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_106_cse ) begin
      mut_3_8_63_0 <= mut_3_7_63_0;
      mut_2_8_63_0 <= mut_2_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_108_cse ) begin
      mut_5_8_63_0 <= mut_5_7_63_0;
      mut_4_8_63_0 <= mut_4_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_110_cse ) begin
      mut_7_8_63_0 <= mut_7_7_63_0;
      mut_6_8_63_0 <= mut_6_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_112_cse ) begin
      mut_9_8_63_0 <= mut_9_7_63_0;
      mut_8_8_63_0 <= mut_8_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_114_cse ) begin
      mut_11_8_63_0 <= mut_11_7_63_0;
      mut_10_8_63_0 <= mut_10_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_116_cse ) begin
      mut_13_8_63_0 <= mut_13_7_63_0;
      mut_12_8_63_0 <= mut_12_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_118_cse ) begin
      mut_15_8_63_0 <= mut_15_7_63_0;
      mut_14_8_63_0 <= mut_14_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_120_cse ) begin
      mut_17_8_63_0 <= mut_17_7_63_0;
      mut_16_8_63_0 <= mut_16_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_122_cse ) begin
      mut_19_8_63_0 <= mut_19_7_63_0;
      mut_18_8_63_0 <= mut_18_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_124_cse ) begin
      mut_21_8_63_0 <= mut_21_7_63_0;
      mut_20_8_63_0 <= mut_20_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_126_cse ) begin
      mut_23_8_63_0 <= mut_23_7_63_0;
      mut_22_8_63_0 <= mut_22_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_128_cse ) begin
      mut_1_8_63_0 <= mut_1_7_63_0;
      mut_8_63_0 <= mut_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_8_3_2 <= 2'b00;
      rem_12cyc_st_8_1_0 <= 2'b00;
    end
    else if ( COMP_LOOP_and_130_cse ) begin
      rem_12cyc_st_8_3_2 <= rem_12cyc_st_7_3_2;
      rem_12cyc_st_8_1_0 <= rem_12cyc_st_7_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_132_cse ) begin
      mut_3_7_63_0 <= mut_3_6_63_0;
      mut_2_7_63_0 <= mut_2_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_134_cse ) begin
      mut_5_7_63_0 <= mut_5_6_63_0;
      mut_4_7_63_0 <= mut_4_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_136_cse ) begin
      mut_7_7_63_0 <= mut_7_6_63_0;
      mut_6_7_63_0 <= mut_6_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_138_cse ) begin
      mut_9_7_63_0 <= mut_9_6_63_0;
      mut_8_7_63_0 <= mut_8_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_140_cse ) begin
      mut_11_7_63_0 <= mut_11_6_63_0;
      mut_10_7_63_0 <= mut_10_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_142_cse ) begin
      mut_13_7_63_0 <= mut_13_6_63_0;
      mut_12_7_63_0 <= mut_12_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_144_cse ) begin
      mut_15_7_63_0 <= mut_15_6_63_0;
      mut_14_7_63_0 <= mut_14_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_146_cse ) begin
      mut_17_7_63_0 <= mut_17_6_63_0;
      mut_16_7_63_0 <= mut_16_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_148_cse ) begin
      mut_19_7_63_0 <= mut_19_6_63_0;
      mut_18_7_63_0 <= mut_18_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_150_cse ) begin
      mut_21_7_63_0 <= mut_21_6_63_0;
      mut_20_7_63_0 <= mut_20_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_152_cse ) begin
      mut_23_7_63_0 <= mut_23_6_63_0;
      mut_22_7_63_0 <= mut_22_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_154_cse ) begin
      mut_1_7_63_0 <= mut_1_6_63_0;
      mut_7_63_0 <= mut_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_7_3_2 <= 2'b00;
      rem_12cyc_st_7_1_0 <= 2'b00;
    end
    else if ( COMP_LOOP_and_156_cse ) begin
      rem_12cyc_st_7_3_2 <= rem_12cyc_st_6_3_2;
      rem_12cyc_st_7_1_0 <= rem_12cyc_st_6_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_158_cse ) begin
      mut_3_6_63_0 <= mut_3_5_63_0;
      mut_2_6_63_0 <= mut_2_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_160_cse ) begin
      mut_5_6_63_0 <= mut_5_5_63_0;
      mut_4_6_63_0 <= mut_4_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_162_cse ) begin
      mut_7_6_63_0 <= mut_7_5_63_0;
      mut_6_6_63_0 <= mut_6_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_164_cse ) begin
      mut_9_6_63_0 <= mut_9_5_63_0;
      mut_8_6_63_0 <= mut_8_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_166_cse ) begin
      mut_11_6_63_0 <= mut_11_5_63_0;
      mut_10_6_63_0 <= mut_10_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_168_cse ) begin
      mut_13_6_63_0 <= mut_13_5_63_0;
      mut_12_6_63_0 <= mut_12_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_170_cse ) begin
      mut_15_6_63_0 <= mut_15_5_63_0;
      mut_14_6_63_0 <= mut_14_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_172_cse ) begin
      mut_17_6_63_0 <= mut_17_5_63_0;
      mut_16_6_63_0 <= mut_16_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_174_cse ) begin
      mut_19_6_63_0 <= mut_19_5_63_0;
      mut_18_6_63_0 <= mut_18_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_176_cse ) begin
      mut_21_6_63_0 <= mut_21_5_63_0;
      mut_20_6_63_0 <= mut_20_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_178_cse ) begin
      mut_23_6_63_0 <= mut_23_5_63_0;
      mut_22_6_63_0 <= mut_22_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_180_cse ) begin
      mut_1_6_63_0 <= mut_1_5_63_0;
      mut_6_63_0 <= mut_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_182_cse ) begin
      m_buf_sva_6 <= m_buf_sva_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_6_3_2 <= 2'b00;
      rem_12cyc_st_6_1_0 <= 2'b00;
    end
    else if ( COMP_LOOP_and_182_cse ) begin
      rem_12cyc_st_6_3_2 <= rem_12cyc_st_5_3_2;
      rem_12cyc_st_6_1_0 <= rem_12cyc_st_5_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_184_cse ) begin
      mut_3_5_63_0 <= mut_3_4_63_0;
      mut_2_5_63_0 <= mut_2_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_186_cse ) begin
      mut_5_5_63_0 <= mut_5_4_63_0;
      mut_4_5_63_0 <= mut_4_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_188_cse ) begin
      mut_7_5_63_0 <= mut_7_4_63_0;
      mut_6_5_63_0 <= mut_6_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_190_cse ) begin
      mut_9_5_63_0 <= mut_9_4_63_0;
      mut_8_5_63_0 <= mut_8_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_192_cse ) begin
      mut_11_5_63_0 <= mut_11_4_63_0;
      mut_10_5_63_0 <= mut_10_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_194_cse ) begin
      mut_13_5_63_0 <= mut_13_4_63_0;
      mut_12_5_63_0 <= mut_12_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_196_cse ) begin
      mut_15_5_63_0 <= mut_15_4_63_0;
      mut_14_5_63_0 <= mut_14_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_198_cse ) begin
      mut_17_5_63_0 <= mut_17_4_63_0;
      mut_16_5_63_0 <= mut_16_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_200_cse ) begin
      mut_19_5_63_0 <= mut_19_4_63_0;
      mut_18_5_63_0 <= mut_18_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_202_cse ) begin
      mut_21_5_63_0 <= mut_21_4_63_0;
      mut_20_5_63_0 <= mut_20_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_204_cse ) begin
      mut_23_5_63_0 <= mut_23_4_63_0;
      mut_22_5_63_0 <= mut_22_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_206_cse ) begin
      mut_1_5_63_0 <= mut_1_4_63_0;
      mut_5_63_0 <= mut_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_208_cse ) begin
      m_buf_sva_5 <= m_buf_sva_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_5_3_2 <= 2'b00;
      rem_12cyc_st_5_1_0 <= 2'b00;
    end
    else if ( COMP_LOOP_and_208_cse ) begin
      rem_12cyc_st_5_3_2 <= rem_12cyc_st_4_3_2;
      rem_12cyc_st_5_1_0 <= rem_12cyc_st_4_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_210_cse ) begin
      mut_3_4_63_0 <= mut_3_3_63_0;
      mut_2_4_63_0 <= mut_2_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_212_cse ) begin
      mut_5_4_63_0 <= mut_5_3_63_0;
      mut_4_4_63_0 <= mut_4_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_214_cse ) begin
      mut_7_4_63_0 <= mut_7_3_63_0;
      mut_6_4_63_0 <= mut_6_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_216_cse ) begin
      mut_9_4_63_0 <= mut_9_3_63_0;
      mut_8_4_63_0 <= mut_8_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_218_cse ) begin
      mut_11_4_63_0 <= mut_11_3_63_0;
      mut_10_4_63_0 <= mut_10_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_220_cse ) begin
      mut_13_4_63_0 <= mut_13_3_63_0;
      mut_12_4_63_0 <= mut_12_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_222_cse ) begin
      mut_15_4_63_0 <= mut_15_3_63_0;
      mut_14_4_63_0 <= mut_14_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_224_cse ) begin
      mut_17_4_63_0 <= mut_17_3_63_0;
      mut_16_4_63_0 <= mut_16_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_226_cse ) begin
      mut_19_4_63_0 <= mut_19_3_63_0;
      mut_18_4_63_0 <= mut_18_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_228_cse ) begin
      mut_21_4_63_0 <= mut_21_3_63_0;
      mut_20_4_63_0 <= mut_20_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_230_cse ) begin
      mut_23_4_63_0 <= mut_23_3_63_0;
      mut_22_4_63_0 <= mut_22_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_232_cse ) begin
      mut_1_4_63_0 <= mut_1_3_63_0;
      mut_4_63_0 <= mut_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_234_cse ) begin
      m_buf_sva_4 <= m_buf_sva_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_4_3_2 <= 2'b00;
      rem_12cyc_st_4_1_0 <= 2'b00;
    end
    else if ( COMP_LOOP_and_234_cse ) begin
      rem_12cyc_st_4_3_2 <= rem_12cyc_st_3_3_2;
      rem_12cyc_st_4_1_0 <= rem_12cyc_st_3_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_236_cse ) begin
      mut_3_3_63_0 <= mut_3_2_63_0;
      mut_2_3_63_0 <= mut_2_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_238_cse ) begin
      mut_5_3_63_0 <= mut_5_2_63_0;
      mut_4_3_63_0 <= mut_4_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_240_cse ) begin
      mut_7_3_63_0 <= mut_7_2_63_0;
      mut_6_3_63_0 <= mut_6_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_242_cse ) begin
      mut_9_3_63_0 <= mut_9_2_63_0;
      mut_8_3_63_0 <= mut_8_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_244_cse ) begin
      mut_11_3_63_0 <= mut_11_2_63_0;
      mut_10_3_63_0 <= mut_10_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_246_cse ) begin
      mut_13_3_63_0 <= mut_13_2_63_0;
      mut_12_3_63_0 <= mut_12_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_248_cse ) begin
      mut_15_3_63_0 <= mut_15_2_63_0;
      mut_14_3_63_0 <= mut_14_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_250_cse ) begin
      mut_17_3_63_0 <= mut_17_2_63_0;
      mut_16_3_63_0 <= mut_16_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_252_cse ) begin
      mut_19_3_63_0 <= mut_19_2_63_0;
      mut_18_3_63_0 <= mut_18_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_254_cse ) begin
      mut_21_3_63_0 <= mut_21_2_63_0;
      mut_20_3_63_0 <= mut_20_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_256_cse ) begin
      mut_23_3_63_0 <= mut_23_2_63_0;
      mut_22_3_63_0 <= mut_22_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_258_cse ) begin
      mut_1_3_63_0 <= mut_1_2_63_0;
      mut_3_63_0 <= mut_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_260_cse ) begin
      m_buf_sva_3 <= m_buf_sva_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_3_3_2 <= 2'b00;
      rem_12cyc_st_3_1_0 <= 2'b00;
    end
    else if ( COMP_LOOP_and_260_cse ) begin
      rem_12cyc_st_3_3_2 <= rem_12cyc_st_2_3_2;
      rem_12cyc_st_3_1_0 <= rem_12cyc_st_2_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_262_cse ) begin
      mut_3_2_63_0 <= rem_12_cmp_1_b_63_0;
      mut_2_2_63_0 <= rem_12_cmp_1_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_264_cse ) begin
      mut_5_2_63_0 <= rem_12_cmp_2_b_63_0;
      mut_4_2_63_0 <= rem_12_cmp_2_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_266_cse ) begin
      mut_7_2_63_0 <= rem_12_cmp_3_b_63_0;
      mut_6_2_63_0 <= rem_12_cmp_3_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_268_cse ) begin
      mut_9_2_63_0 <= rem_12_cmp_4_b_63_0;
      mut_8_2_63_0 <= rem_12_cmp_4_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_270_cse ) begin
      mut_11_2_63_0 <= rem_12_cmp_5_b_63_0;
      mut_10_2_63_0 <= rem_12_cmp_5_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_272_cse ) begin
      mut_13_2_63_0 <= rem_12_cmp_6_b_63_0;
      mut_12_2_63_0 <= rem_12_cmp_6_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_274_cse ) begin
      mut_15_2_63_0 <= rem_12_cmp_7_b_63_0;
      mut_14_2_63_0 <= rem_12_cmp_7_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_276_cse ) begin
      mut_17_2_63_0 <= rem_12_cmp_8_b_63_0;
      mut_16_2_63_0 <= rem_12_cmp_8_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_278_cse ) begin
      mut_19_2_63_0 <= rem_12_cmp_9_b_63_0;
      mut_18_2_63_0 <= rem_12_cmp_9_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_280_cse ) begin
      mut_21_2_63_0 <= rem_12_cmp_10_b_63_0;
      mut_20_2_63_0 <= rem_12_cmp_10_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_282_cse ) begin
      mut_23_2_63_0 <= rem_12_cmp_11_b_63_0;
      mut_22_2_63_0 <= rem_12_cmp_11_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_284_cse ) begin
      mut_1_2_63_0 <= rem_12_cmp_b_63_0;
      mut_2_63_0 <= rem_12_cmp_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_286_cse ) begin
      m_buf_sva_2 <= m_buf_sva_1;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_2_3_2 <= 2'b00;
      rem_12cyc_st_2_1_0 <= 2'b00;
    end
    else if ( COMP_LOOP_and_286_cse ) begin
      rem_12cyc_st_2_3_2 <= rem_12cyc_3_2;
      rem_12cyc_st_2_1_0 <= rem_12cyc_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( COMP_LOOP_and_24_cse ) begin
      m_buf_sva_1 <= m_rsci_idat;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_3_2 <= 2'b00;
      rem_12cyc_1_0 <= 2'b00;
    end
    else if ( COMP_LOOP_and_24_cse ) begin
      rem_12cyc_3_2 <= COMP_LOOP_acc_tmp;
      rem_12cyc_1_0 <= COMP_LOOP_acc_1_tmp[1:0];
    end
  end
  assign nl_qelse_acc_nl = result_sva_duc_mx0 + m_buf_sva_12;
  assign qelse_acc_nl = nl_qelse_acc_nl[63:0];
  assign mux_8_nl = MUX_s_1_2_2((rem_12_cmp_1_z[63]), (rem_12_cmp_3_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_7_nl = MUX_s_1_2_2((rem_12_cmp_2_z[63]), (rem_12_cmp_4_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_9_nl = MUX_s_1_2_2(mux_8_nl, mux_7_nl, rem_12cyc_st_12_1_0[0]);
  assign mux_5_nl = MUX_s_1_2_2((rem_12_cmp_9_z[63]), (rem_12_cmp_11_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_4_nl = MUX_s_1_2_2((rem_12_cmp_10_z[63]), (rem_12_cmp_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_6_nl = MUX_s_1_2_2(mux_5_nl, mux_4_nl, rem_12cyc_st_12_1_0[0]);
  assign mux_10_nl = MUX_s_1_2_2(mux_9_nl, mux_6_nl, rem_12cyc_st_12_3_2[1]);
  assign mux_1_nl = MUX_s_1_2_2((rem_12_cmp_5_z[63]), (rem_12_cmp_7_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_nl = MUX_s_1_2_2((rem_12_cmp_6_z[63]), (rem_12_cmp_8_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_2_nl = MUX_s_1_2_2(mux_1_nl, mux_nl, rem_12cyc_st_12_1_0[0]);
  assign mux_3_nl = MUX_s_1_2_2(mux_2_nl, (result_sva_duc[63]), rem_12cyc_st_12_3_2[1]);
  assign mux_11_nl = MUX_s_1_2_2(mux_10_nl, mux_3_nl, rem_12cyc_st_12_3_2[0]);

  function automatic [63:0] MUX1HOT_v_64_11_2;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [10:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    MUX1HOT_v_64_11_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_13_2;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [12:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    MUX1HOT_v_64_13_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    modulo
// ------------------------------------------------------------------


module modulo (
  base_rsc_dat, m_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [63:0] base_rsc_dat;
  input [63:0] m_rsc_dat;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  modulo_core modulo_core_inst (
      .base_rsc_dat(base_rsc_dat),
      .m_rsc_dat(m_rsc_dat),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Mon Aug  2 20:58:11 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_40_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_40_6_64_64_64_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output [63:0] q_d;
  input [5:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_39_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_39_6_64_64_64_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output [63:0] q_d;
  input [5:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_38_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_38_6_64_64_64_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output [63:0] q_d;
  input [5:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_37_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_37_6_64_64_64_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output [63:0] q_d;
  input [5:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_36_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_36_6_64_64_64_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output [63:0] q_d;
  input [5:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_35_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_35_6_64_64_64_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output [63:0] q_d;
  input [5:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_34_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_34_6_64_64_64_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output [63:0] q_d;
  input [5:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_33_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_33_6_64_64_64_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output [63:0] q_d;
  input [5:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_32_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_32_6_64_64_64_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output [63:0] q_d;
  input [5:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_31_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_31_6_64_64_64_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output [63:0] q_d;
  input [5:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_30_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_30_6_64_64_64_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output [63:0] q_d;
  input [5:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_29_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_29_6_64_64_64_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output [63:0] q_d;
  input [5:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_28_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_28_6_64_64_64_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output [63:0] q_d;
  input [5:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_27_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_27_6_64_64_64_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output [63:0] q_d;
  input [5:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_26_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_26_6_64_64_64_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output [63:0] q_d;
  input [5:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_25_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_25_6_64_64_64_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output [63:0] q_d;
  input [5:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module inPlaceNTT_DIF_core_core_fsm (
  clk, rst, fsm_output, COMP_LOOP_C_31_tr0, COMP_LOOP_C_62_tr0, COMP_LOOP_C_93_tr0,
      COMP_LOOP_C_124_tr0, COMP_LOOP_C_155_tr0, COMP_LOOP_C_186_tr0, COMP_LOOP_C_217_tr0,
      COMP_LOOP_C_248_tr0, COMP_LOOP_C_279_tr0, COMP_LOOP_C_310_tr0, COMP_LOOP_C_341_tr0,
      COMP_LOOP_C_372_tr0, COMP_LOOP_C_403_tr0, COMP_LOOP_C_434_tr0, COMP_LOOP_C_465_tr0,
      COMP_LOOP_C_496_tr0, VEC_LOOP_C_0_tr0, STAGE_LOOP_C_1_tr0
);
  input clk;
  input rst;
  output [8:0] fsm_output;
  reg [8:0] fsm_output;
  input COMP_LOOP_C_31_tr0;
  input COMP_LOOP_C_62_tr0;
  input COMP_LOOP_C_93_tr0;
  input COMP_LOOP_C_124_tr0;
  input COMP_LOOP_C_155_tr0;
  input COMP_LOOP_C_186_tr0;
  input COMP_LOOP_C_217_tr0;
  input COMP_LOOP_C_248_tr0;
  input COMP_LOOP_C_279_tr0;
  input COMP_LOOP_C_310_tr0;
  input COMP_LOOP_C_341_tr0;
  input COMP_LOOP_C_372_tr0;
  input COMP_LOOP_C_403_tr0;
  input COMP_LOOP_C_434_tr0;
  input COMP_LOOP_C_465_tr0;
  input COMP_LOOP_C_496_tr0;
  input VEC_LOOP_C_0_tr0;
  input STAGE_LOOP_C_1_tr0;


  // FSM State Type Declaration for inPlaceNTT_DIF_core_core_fsm_1
  parameter
    main_C_0 = 9'd0,
    STAGE_LOOP_C_0 = 9'd1,
    COMP_LOOP_C_0 = 9'd2,
    COMP_LOOP_C_1 = 9'd3,
    COMP_LOOP_C_2 = 9'd4,
    COMP_LOOP_C_3 = 9'd5,
    COMP_LOOP_C_4 = 9'd6,
    COMP_LOOP_C_5 = 9'd7,
    COMP_LOOP_C_6 = 9'd8,
    COMP_LOOP_C_7 = 9'd9,
    COMP_LOOP_C_8 = 9'd10,
    COMP_LOOP_C_9 = 9'd11,
    COMP_LOOP_C_10 = 9'd12,
    COMP_LOOP_C_11 = 9'd13,
    COMP_LOOP_C_12 = 9'd14,
    COMP_LOOP_C_13 = 9'd15,
    COMP_LOOP_C_14 = 9'd16,
    COMP_LOOP_C_15 = 9'd17,
    COMP_LOOP_C_16 = 9'd18,
    COMP_LOOP_C_17 = 9'd19,
    COMP_LOOP_C_18 = 9'd20,
    COMP_LOOP_C_19 = 9'd21,
    COMP_LOOP_C_20 = 9'd22,
    COMP_LOOP_C_21 = 9'd23,
    COMP_LOOP_C_22 = 9'd24,
    COMP_LOOP_C_23 = 9'd25,
    COMP_LOOP_C_24 = 9'd26,
    COMP_LOOP_C_25 = 9'd27,
    COMP_LOOP_C_26 = 9'd28,
    COMP_LOOP_C_27 = 9'd29,
    COMP_LOOP_C_28 = 9'd30,
    COMP_LOOP_C_29 = 9'd31,
    COMP_LOOP_C_30 = 9'd32,
    COMP_LOOP_C_31 = 9'd33,
    COMP_LOOP_C_32 = 9'd34,
    COMP_LOOP_C_33 = 9'd35,
    COMP_LOOP_C_34 = 9'd36,
    COMP_LOOP_C_35 = 9'd37,
    COMP_LOOP_C_36 = 9'd38,
    COMP_LOOP_C_37 = 9'd39,
    COMP_LOOP_C_38 = 9'd40,
    COMP_LOOP_C_39 = 9'd41,
    COMP_LOOP_C_40 = 9'd42,
    COMP_LOOP_C_41 = 9'd43,
    COMP_LOOP_C_42 = 9'd44,
    COMP_LOOP_C_43 = 9'd45,
    COMP_LOOP_C_44 = 9'd46,
    COMP_LOOP_C_45 = 9'd47,
    COMP_LOOP_C_46 = 9'd48,
    COMP_LOOP_C_47 = 9'd49,
    COMP_LOOP_C_48 = 9'd50,
    COMP_LOOP_C_49 = 9'd51,
    COMP_LOOP_C_50 = 9'd52,
    COMP_LOOP_C_51 = 9'd53,
    COMP_LOOP_C_52 = 9'd54,
    COMP_LOOP_C_53 = 9'd55,
    COMP_LOOP_C_54 = 9'd56,
    COMP_LOOP_C_55 = 9'd57,
    COMP_LOOP_C_56 = 9'd58,
    COMP_LOOP_C_57 = 9'd59,
    COMP_LOOP_C_58 = 9'd60,
    COMP_LOOP_C_59 = 9'd61,
    COMP_LOOP_C_60 = 9'd62,
    COMP_LOOP_C_61 = 9'd63,
    COMP_LOOP_C_62 = 9'd64,
    COMP_LOOP_C_63 = 9'd65,
    COMP_LOOP_C_64 = 9'd66,
    COMP_LOOP_C_65 = 9'd67,
    COMP_LOOP_C_66 = 9'd68,
    COMP_LOOP_C_67 = 9'd69,
    COMP_LOOP_C_68 = 9'd70,
    COMP_LOOP_C_69 = 9'd71,
    COMP_LOOP_C_70 = 9'd72,
    COMP_LOOP_C_71 = 9'd73,
    COMP_LOOP_C_72 = 9'd74,
    COMP_LOOP_C_73 = 9'd75,
    COMP_LOOP_C_74 = 9'd76,
    COMP_LOOP_C_75 = 9'd77,
    COMP_LOOP_C_76 = 9'd78,
    COMP_LOOP_C_77 = 9'd79,
    COMP_LOOP_C_78 = 9'd80,
    COMP_LOOP_C_79 = 9'd81,
    COMP_LOOP_C_80 = 9'd82,
    COMP_LOOP_C_81 = 9'd83,
    COMP_LOOP_C_82 = 9'd84,
    COMP_LOOP_C_83 = 9'd85,
    COMP_LOOP_C_84 = 9'd86,
    COMP_LOOP_C_85 = 9'd87,
    COMP_LOOP_C_86 = 9'd88,
    COMP_LOOP_C_87 = 9'd89,
    COMP_LOOP_C_88 = 9'd90,
    COMP_LOOP_C_89 = 9'd91,
    COMP_LOOP_C_90 = 9'd92,
    COMP_LOOP_C_91 = 9'd93,
    COMP_LOOP_C_92 = 9'd94,
    COMP_LOOP_C_93 = 9'd95,
    COMP_LOOP_C_94 = 9'd96,
    COMP_LOOP_C_95 = 9'd97,
    COMP_LOOP_C_96 = 9'd98,
    COMP_LOOP_C_97 = 9'd99,
    COMP_LOOP_C_98 = 9'd100,
    COMP_LOOP_C_99 = 9'd101,
    COMP_LOOP_C_100 = 9'd102,
    COMP_LOOP_C_101 = 9'd103,
    COMP_LOOP_C_102 = 9'd104,
    COMP_LOOP_C_103 = 9'd105,
    COMP_LOOP_C_104 = 9'd106,
    COMP_LOOP_C_105 = 9'd107,
    COMP_LOOP_C_106 = 9'd108,
    COMP_LOOP_C_107 = 9'd109,
    COMP_LOOP_C_108 = 9'd110,
    COMP_LOOP_C_109 = 9'd111,
    COMP_LOOP_C_110 = 9'd112,
    COMP_LOOP_C_111 = 9'd113,
    COMP_LOOP_C_112 = 9'd114,
    COMP_LOOP_C_113 = 9'd115,
    COMP_LOOP_C_114 = 9'd116,
    COMP_LOOP_C_115 = 9'd117,
    COMP_LOOP_C_116 = 9'd118,
    COMP_LOOP_C_117 = 9'd119,
    COMP_LOOP_C_118 = 9'd120,
    COMP_LOOP_C_119 = 9'd121,
    COMP_LOOP_C_120 = 9'd122,
    COMP_LOOP_C_121 = 9'd123,
    COMP_LOOP_C_122 = 9'd124,
    COMP_LOOP_C_123 = 9'd125,
    COMP_LOOP_C_124 = 9'd126,
    COMP_LOOP_C_125 = 9'd127,
    COMP_LOOP_C_126 = 9'd128,
    COMP_LOOP_C_127 = 9'd129,
    COMP_LOOP_C_128 = 9'd130,
    COMP_LOOP_C_129 = 9'd131,
    COMP_LOOP_C_130 = 9'd132,
    COMP_LOOP_C_131 = 9'd133,
    COMP_LOOP_C_132 = 9'd134,
    COMP_LOOP_C_133 = 9'd135,
    COMP_LOOP_C_134 = 9'd136,
    COMP_LOOP_C_135 = 9'd137,
    COMP_LOOP_C_136 = 9'd138,
    COMP_LOOP_C_137 = 9'd139,
    COMP_LOOP_C_138 = 9'd140,
    COMP_LOOP_C_139 = 9'd141,
    COMP_LOOP_C_140 = 9'd142,
    COMP_LOOP_C_141 = 9'd143,
    COMP_LOOP_C_142 = 9'd144,
    COMP_LOOP_C_143 = 9'd145,
    COMP_LOOP_C_144 = 9'd146,
    COMP_LOOP_C_145 = 9'd147,
    COMP_LOOP_C_146 = 9'd148,
    COMP_LOOP_C_147 = 9'd149,
    COMP_LOOP_C_148 = 9'd150,
    COMP_LOOP_C_149 = 9'd151,
    COMP_LOOP_C_150 = 9'd152,
    COMP_LOOP_C_151 = 9'd153,
    COMP_LOOP_C_152 = 9'd154,
    COMP_LOOP_C_153 = 9'd155,
    COMP_LOOP_C_154 = 9'd156,
    COMP_LOOP_C_155 = 9'd157,
    COMP_LOOP_C_156 = 9'd158,
    COMP_LOOP_C_157 = 9'd159,
    COMP_LOOP_C_158 = 9'd160,
    COMP_LOOP_C_159 = 9'd161,
    COMP_LOOP_C_160 = 9'd162,
    COMP_LOOP_C_161 = 9'd163,
    COMP_LOOP_C_162 = 9'd164,
    COMP_LOOP_C_163 = 9'd165,
    COMP_LOOP_C_164 = 9'd166,
    COMP_LOOP_C_165 = 9'd167,
    COMP_LOOP_C_166 = 9'd168,
    COMP_LOOP_C_167 = 9'd169,
    COMP_LOOP_C_168 = 9'd170,
    COMP_LOOP_C_169 = 9'd171,
    COMP_LOOP_C_170 = 9'd172,
    COMP_LOOP_C_171 = 9'd173,
    COMP_LOOP_C_172 = 9'd174,
    COMP_LOOP_C_173 = 9'd175,
    COMP_LOOP_C_174 = 9'd176,
    COMP_LOOP_C_175 = 9'd177,
    COMP_LOOP_C_176 = 9'd178,
    COMP_LOOP_C_177 = 9'd179,
    COMP_LOOP_C_178 = 9'd180,
    COMP_LOOP_C_179 = 9'd181,
    COMP_LOOP_C_180 = 9'd182,
    COMP_LOOP_C_181 = 9'd183,
    COMP_LOOP_C_182 = 9'd184,
    COMP_LOOP_C_183 = 9'd185,
    COMP_LOOP_C_184 = 9'd186,
    COMP_LOOP_C_185 = 9'd187,
    COMP_LOOP_C_186 = 9'd188,
    COMP_LOOP_C_187 = 9'd189,
    COMP_LOOP_C_188 = 9'd190,
    COMP_LOOP_C_189 = 9'd191,
    COMP_LOOP_C_190 = 9'd192,
    COMP_LOOP_C_191 = 9'd193,
    COMP_LOOP_C_192 = 9'd194,
    COMP_LOOP_C_193 = 9'd195,
    COMP_LOOP_C_194 = 9'd196,
    COMP_LOOP_C_195 = 9'd197,
    COMP_LOOP_C_196 = 9'd198,
    COMP_LOOP_C_197 = 9'd199,
    COMP_LOOP_C_198 = 9'd200,
    COMP_LOOP_C_199 = 9'd201,
    COMP_LOOP_C_200 = 9'd202,
    COMP_LOOP_C_201 = 9'd203,
    COMP_LOOP_C_202 = 9'd204,
    COMP_LOOP_C_203 = 9'd205,
    COMP_LOOP_C_204 = 9'd206,
    COMP_LOOP_C_205 = 9'd207,
    COMP_LOOP_C_206 = 9'd208,
    COMP_LOOP_C_207 = 9'd209,
    COMP_LOOP_C_208 = 9'd210,
    COMP_LOOP_C_209 = 9'd211,
    COMP_LOOP_C_210 = 9'd212,
    COMP_LOOP_C_211 = 9'd213,
    COMP_LOOP_C_212 = 9'd214,
    COMP_LOOP_C_213 = 9'd215,
    COMP_LOOP_C_214 = 9'd216,
    COMP_LOOP_C_215 = 9'd217,
    COMP_LOOP_C_216 = 9'd218,
    COMP_LOOP_C_217 = 9'd219,
    COMP_LOOP_C_218 = 9'd220,
    COMP_LOOP_C_219 = 9'd221,
    COMP_LOOP_C_220 = 9'd222,
    COMP_LOOP_C_221 = 9'd223,
    COMP_LOOP_C_222 = 9'd224,
    COMP_LOOP_C_223 = 9'd225,
    COMP_LOOP_C_224 = 9'd226,
    COMP_LOOP_C_225 = 9'd227,
    COMP_LOOP_C_226 = 9'd228,
    COMP_LOOP_C_227 = 9'd229,
    COMP_LOOP_C_228 = 9'd230,
    COMP_LOOP_C_229 = 9'd231,
    COMP_LOOP_C_230 = 9'd232,
    COMP_LOOP_C_231 = 9'd233,
    COMP_LOOP_C_232 = 9'd234,
    COMP_LOOP_C_233 = 9'd235,
    COMP_LOOP_C_234 = 9'd236,
    COMP_LOOP_C_235 = 9'd237,
    COMP_LOOP_C_236 = 9'd238,
    COMP_LOOP_C_237 = 9'd239,
    COMP_LOOP_C_238 = 9'd240,
    COMP_LOOP_C_239 = 9'd241,
    COMP_LOOP_C_240 = 9'd242,
    COMP_LOOP_C_241 = 9'd243,
    COMP_LOOP_C_242 = 9'd244,
    COMP_LOOP_C_243 = 9'd245,
    COMP_LOOP_C_244 = 9'd246,
    COMP_LOOP_C_245 = 9'd247,
    COMP_LOOP_C_246 = 9'd248,
    COMP_LOOP_C_247 = 9'd249,
    COMP_LOOP_C_248 = 9'd250,
    COMP_LOOP_C_249 = 9'd251,
    COMP_LOOP_C_250 = 9'd252,
    COMP_LOOP_C_251 = 9'd253,
    COMP_LOOP_C_252 = 9'd254,
    COMP_LOOP_C_253 = 9'd255,
    COMP_LOOP_C_254 = 9'd256,
    COMP_LOOP_C_255 = 9'd257,
    COMP_LOOP_C_256 = 9'd258,
    COMP_LOOP_C_257 = 9'd259,
    COMP_LOOP_C_258 = 9'd260,
    COMP_LOOP_C_259 = 9'd261,
    COMP_LOOP_C_260 = 9'd262,
    COMP_LOOP_C_261 = 9'd263,
    COMP_LOOP_C_262 = 9'd264,
    COMP_LOOP_C_263 = 9'd265,
    COMP_LOOP_C_264 = 9'd266,
    COMP_LOOP_C_265 = 9'd267,
    COMP_LOOP_C_266 = 9'd268,
    COMP_LOOP_C_267 = 9'd269,
    COMP_LOOP_C_268 = 9'd270,
    COMP_LOOP_C_269 = 9'd271,
    COMP_LOOP_C_270 = 9'd272,
    COMP_LOOP_C_271 = 9'd273,
    COMP_LOOP_C_272 = 9'd274,
    COMP_LOOP_C_273 = 9'd275,
    COMP_LOOP_C_274 = 9'd276,
    COMP_LOOP_C_275 = 9'd277,
    COMP_LOOP_C_276 = 9'd278,
    COMP_LOOP_C_277 = 9'd279,
    COMP_LOOP_C_278 = 9'd280,
    COMP_LOOP_C_279 = 9'd281,
    COMP_LOOP_C_280 = 9'd282,
    COMP_LOOP_C_281 = 9'd283,
    COMP_LOOP_C_282 = 9'd284,
    COMP_LOOP_C_283 = 9'd285,
    COMP_LOOP_C_284 = 9'd286,
    COMP_LOOP_C_285 = 9'd287,
    COMP_LOOP_C_286 = 9'd288,
    COMP_LOOP_C_287 = 9'd289,
    COMP_LOOP_C_288 = 9'd290,
    COMP_LOOP_C_289 = 9'd291,
    COMP_LOOP_C_290 = 9'd292,
    COMP_LOOP_C_291 = 9'd293,
    COMP_LOOP_C_292 = 9'd294,
    COMP_LOOP_C_293 = 9'd295,
    COMP_LOOP_C_294 = 9'd296,
    COMP_LOOP_C_295 = 9'd297,
    COMP_LOOP_C_296 = 9'd298,
    COMP_LOOP_C_297 = 9'd299,
    COMP_LOOP_C_298 = 9'd300,
    COMP_LOOP_C_299 = 9'd301,
    COMP_LOOP_C_300 = 9'd302,
    COMP_LOOP_C_301 = 9'd303,
    COMP_LOOP_C_302 = 9'd304,
    COMP_LOOP_C_303 = 9'd305,
    COMP_LOOP_C_304 = 9'd306,
    COMP_LOOP_C_305 = 9'd307,
    COMP_LOOP_C_306 = 9'd308,
    COMP_LOOP_C_307 = 9'd309,
    COMP_LOOP_C_308 = 9'd310,
    COMP_LOOP_C_309 = 9'd311,
    COMP_LOOP_C_310 = 9'd312,
    COMP_LOOP_C_311 = 9'd313,
    COMP_LOOP_C_312 = 9'd314,
    COMP_LOOP_C_313 = 9'd315,
    COMP_LOOP_C_314 = 9'd316,
    COMP_LOOP_C_315 = 9'd317,
    COMP_LOOP_C_316 = 9'd318,
    COMP_LOOP_C_317 = 9'd319,
    COMP_LOOP_C_318 = 9'd320,
    COMP_LOOP_C_319 = 9'd321,
    COMP_LOOP_C_320 = 9'd322,
    COMP_LOOP_C_321 = 9'd323,
    COMP_LOOP_C_322 = 9'd324,
    COMP_LOOP_C_323 = 9'd325,
    COMP_LOOP_C_324 = 9'd326,
    COMP_LOOP_C_325 = 9'd327,
    COMP_LOOP_C_326 = 9'd328,
    COMP_LOOP_C_327 = 9'd329,
    COMP_LOOP_C_328 = 9'd330,
    COMP_LOOP_C_329 = 9'd331,
    COMP_LOOP_C_330 = 9'd332,
    COMP_LOOP_C_331 = 9'd333,
    COMP_LOOP_C_332 = 9'd334,
    COMP_LOOP_C_333 = 9'd335,
    COMP_LOOP_C_334 = 9'd336,
    COMP_LOOP_C_335 = 9'd337,
    COMP_LOOP_C_336 = 9'd338,
    COMP_LOOP_C_337 = 9'd339,
    COMP_LOOP_C_338 = 9'd340,
    COMP_LOOP_C_339 = 9'd341,
    COMP_LOOP_C_340 = 9'd342,
    COMP_LOOP_C_341 = 9'd343,
    COMP_LOOP_C_342 = 9'd344,
    COMP_LOOP_C_343 = 9'd345,
    COMP_LOOP_C_344 = 9'd346,
    COMP_LOOP_C_345 = 9'd347,
    COMP_LOOP_C_346 = 9'd348,
    COMP_LOOP_C_347 = 9'd349,
    COMP_LOOP_C_348 = 9'd350,
    COMP_LOOP_C_349 = 9'd351,
    COMP_LOOP_C_350 = 9'd352,
    COMP_LOOP_C_351 = 9'd353,
    COMP_LOOP_C_352 = 9'd354,
    COMP_LOOP_C_353 = 9'd355,
    COMP_LOOP_C_354 = 9'd356,
    COMP_LOOP_C_355 = 9'd357,
    COMP_LOOP_C_356 = 9'd358,
    COMP_LOOP_C_357 = 9'd359,
    COMP_LOOP_C_358 = 9'd360,
    COMP_LOOP_C_359 = 9'd361,
    COMP_LOOP_C_360 = 9'd362,
    COMP_LOOP_C_361 = 9'd363,
    COMP_LOOP_C_362 = 9'd364,
    COMP_LOOP_C_363 = 9'd365,
    COMP_LOOP_C_364 = 9'd366,
    COMP_LOOP_C_365 = 9'd367,
    COMP_LOOP_C_366 = 9'd368,
    COMP_LOOP_C_367 = 9'd369,
    COMP_LOOP_C_368 = 9'd370,
    COMP_LOOP_C_369 = 9'd371,
    COMP_LOOP_C_370 = 9'd372,
    COMP_LOOP_C_371 = 9'd373,
    COMP_LOOP_C_372 = 9'd374,
    COMP_LOOP_C_373 = 9'd375,
    COMP_LOOP_C_374 = 9'd376,
    COMP_LOOP_C_375 = 9'd377,
    COMP_LOOP_C_376 = 9'd378,
    COMP_LOOP_C_377 = 9'd379,
    COMP_LOOP_C_378 = 9'd380,
    COMP_LOOP_C_379 = 9'd381,
    COMP_LOOP_C_380 = 9'd382,
    COMP_LOOP_C_381 = 9'd383,
    COMP_LOOP_C_382 = 9'd384,
    COMP_LOOP_C_383 = 9'd385,
    COMP_LOOP_C_384 = 9'd386,
    COMP_LOOP_C_385 = 9'd387,
    COMP_LOOP_C_386 = 9'd388,
    COMP_LOOP_C_387 = 9'd389,
    COMP_LOOP_C_388 = 9'd390,
    COMP_LOOP_C_389 = 9'd391,
    COMP_LOOP_C_390 = 9'd392,
    COMP_LOOP_C_391 = 9'd393,
    COMP_LOOP_C_392 = 9'd394,
    COMP_LOOP_C_393 = 9'd395,
    COMP_LOOP_C_394 = 9'd396,
    COMP_LOOP_C_395 = 9'd397,
    COMP_LOOP_C_396 = 9'd398,
    COMP_LOOP_C_397 = 9'd399,
    COMP_LOOP_C_398 = 9'd400,
    COMP_LOOP_C_399 = 9'd401,
    COMP_LOOP_C_400 = 9'd402,
    COMP_LOOP_C_401 = 9'd403,
    COMP_LOOP_C_402 = 9'd404,
    COMP_LOOP_C_403 = 9'd405,
    COMP_LOOP_C_404 = 9'd406,
    COMP_LOOP_C_405 = 9'd407,
    COMP_LOOP_C_406 = 9'd408,
    COMP_LOOP_C_407 = 9'd409,
    COMP_LOOP_C_408 = 9'd410,
    COMP_LOOP_C_409 = 9'd411,
    COMP_LOOP_C_410 = 9'd412,
    COMP_LOOP_C_411 = 9'd413,
    COMP_LOOP_C_412 = 9'd414,
    COMP_LOOP_C_413 = 9'd415,
    COMP_LOOP_C_414 = 9'd416,
    COMP_LOOP_C_415 = 9'd417,
    COMP_LOOP_C_416 = 9'd418,
    COMP_LOOP_C_417 = 9'd419,
    COMP_LOOP_C_418 = 9'd420,
    COMP_LOOP_C_419 = 9'd421,
    COMP_LOOP_C_420 = 9'd422,
    COMP_LOOP_C_421 = 9'd423,
    COMP_LOOP_C_422 = 9'd424,
    COMP_LOOP_C_423 = 9'd425,
    COMP_LOOP_C_424 = 9'd426,
    COMP_LOOP_C_425 = 9'd427,
    COMP_LOOP_C_426 = 9'd428,
    COMP_LOOP_C_427 = 9'd429,
    COMP_LOOP_C_428 = 9'd430,
    COMP_LOOP_C_429 = 9'd431,
    COMP_LOOP_C_430 = 9'd432,
    COMP_LOOP_C_431 = 9'd433,
    COMP_LOOP_C_432 = 9'd434,
    COMP_LOOP_C_433 = 9'd435,
    COMP_LOOP_C_434 = 9'd436,
    COMP_LOOP_C_435 = 9'd437,
    COMP_LOOP_C_436 = 9'd438,
    COMP_LOOP_C_437 = 9'd439,
    COMP_LOOP_C_438 = 9'd440,
    COMP_LOOP_C_439 = 9'd441,
    COMP_LOOP_C_440 = 9'd442,
    COMP_LOOP_C_441 = 9'd443,
    COMP_LOOP_C_442 = 9'd444,
    COMP_LOOP_C_443 = 9'd445,
    COMP_LOOP_C_444 = 9'd446,
    COMP_LOOP_C_445 = 9'd447,
    COMP_LOOP_C_446 = 9'd448,
    COMP_LOOP_C_447 = 9'd449,
    COMP_LOOP_C_448 = 9'd450,
    COMP_LOOP_C_449 = 9'd451,
    COMP_LOOP_C_450 = 9'd452,
    COMP_LOOP_C_451 = 9'd453,
    COMP_LOOP_C_452 = 9'd454,
    COMP_LOOP_C_453 = 9'd455,
    COMP_LOOP_C_454 = 9'd456,
    COMP_LOOP_C_455 = 9'd457,
    COMP_LOOP_C_456 = 9'd458,
    COMP_LOOP_C_457 = 9'd459,
    COMP_LOOP_C_458 = 9'd460,
    COMP_LOOP_C_459 = 9'd461,
    COMP_LOOP_C_460 = 9'd462,
    COMP_LOOP_C_461 = 9'd463,
    COMP_LOOP_C_462 = 9'd464,
    COMP_LOOP_C_463 = 9'd465,
    COMP_LOOP_C_464 = 9'd466,
    COMP_LOOP_C_465 = 9'd467,
    COMP_LOOP_C_466 = 9'd468,
    COMP_LOOP_C_467 = 9'd469,
    COMP_LOOP_C_468 = 9'd470,
    COMP_LOOP_C_469 = 9'd471,
    COMP_LOOP_C_470 = 9'd472,
    COMP_LOOP_C_471 = 9'd473,
    COMP_LOOP_C_472 = 9'd474,
    COMP_LOOP_C_473 = 9'd475,
    COMP_LOOP_C_474 = 9'd476,
    COMP_LOOP_C_475 = 9'd477,
    COMP_LOOP_C_476 = 9'd478,
    COMP_LOOP_C_477 = 9'd479,
    COMP_LOOP_C_478 = 9'd480,
    COMP_LOOP_C_479 = 9'd481,
    COMP_LOOP_C_480 = 9'd482,
    COMP_LOOP_C_481 = 9'd483,
    COMP_LOOP_C_482 = 9'd484,
    COMP_LOOP_C_483 = 9'd485,
    COMP_LOOP_C_484 = 9'd486,
    COMP_LOOP_C_485 = 9'd487,
    COMP_LOOP_C_486 = 9'd488,
    COMP_LOOP_C_487 = 9'd489,
    COMP_LOOP_C_488 = 9'd490,
    COMP_LOOP_C_489 = 9'd491,
    COMP_LOOP_C_490 = 9'd492,
    COMP_LOOP_C_491 = 9'd493,
    COMP_LOOP_C_492 = 9'd494,
    COMP_LOOP_C_493 = 9'd495,
    COMP_LOOP_C_494 = 9'd496,
    COMP_LOOP_C_495 = 9'd497,
    COMP_LOOP_C_496 = 9'd498,
    VEC_LOOP_C_0 = 9'd499,
    STAGE_LOOP_C_1 = 9'd500,
    main_C_1 = 9'd501;

  reg [8:0] state_var;
  reg [8:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : inPlaceNTT_DIF_core_core_fsm_1
    case (state_var)
      STAGE_LOOP_C_0 : begin
        fsm_output = 9'b000000001;
        state_var_NS = COMP_LOOP_C_0;
      end
      COMP_LOOP_C_0 : begin
        fsm_output = 9'b000000010;
        state_var_NS = COMP_LOOP_C_1;
      end
      COMP_LOOP_C_1 : begin
        fsm_output = 9'b000000011;
        state_var_NS = COMP_LOOP_C_2;
      end
      COMP_LOOP_C_2 : begin
        fsm_output = 9'b000000100;
        state_var_NS = COMP_LOOP_C_3;
      end
      COMP_LOOP_C_3 : begin
        fsm_output = 9'b000000101;
        state_var_NS = COMP_LOOP_C_4;
      end
      COMP_LOOP_C_4 : begin
        fsm_output = 9'b000000110;
        state_var_NS = COMP_LOOP_C_5;
      end
      COMP_LOOP_C_5 : begin
        fsm_output = 9'b000000111;
        state_var_NS = COMP_LOOP_C_6;
      end
      COMP_LOOP_C_6 : begin
        fsm_output = 9'b000001000;
        state_var_NS = COMP_LOOP_C_7;
      end
      COMP_LOOP_C_7 : begin
        fsm_output = 9'b000001001;
        state_var_NS = COMP_LOOP_C_8;
      end
      COMP_LOOP_C_8 : begin
        fsm_output = 9'b000001010;
        state_var_NS = COMP_LOOP_C_9;
      end
      COMP_LOOP_C_9 : begin
        fsm_output = 9'b000001011;
        state_var_NS = COMP_LOOP_C_10;
      end
      COMP_LOOP_C_10 : begin
        fsm_output = 9'b000001100;
        state_var_NS = COMP_LOOP_C_11;
      end
      COMP_LOOP_C_11 : begin
        fsm_output = 9'b000001101;
        state_var_NS = COMP_LOOP_C_12;
      end
      COMP_LOOP_C_12 : begin
        fsm_output = 9'b000001110;
        state_var_NS = COMP_LOOP_C_13;
      end
      COMP_LOOP_C_13 : begin
        fsm_output = 9'b000001111;
        state_var_NS = COMP_LOOP_C_14;
      end
      COMP_LOOP_C_14 : begin
        fsm_output = 9'b000010000;
        state_var_NS = COMP_LOOP_C_15;
      end
      COMP_LOOP_C_15 : begin
        fsm_output = 9'b000010001;
        state_var_NS = COMP_LOOP_C_16;
      end
      COMP_LOOP_C_16 : begin
        fsm_output = 9'b000010010;
        state_var_NS = COMP_LOOP_C_17;
      end
      COMP_LOOP_C_17 : begin
        fsm_output = 9'b000010011;
        state_var_NS = COMP_LOOP_C_18;
      end
      COMP_LOOP_C_18 : begin
        fsm_output = 9'b000010100;
        state_var_NS = COMP_LOOP_C_19;
      end
      COMP_LOOP_C_19 : begin
        fsm_output = 9'b000010101;
        state_var_NS = COMP_LOOP_C_20;
      end
      COMP_LOOP_C_20 : begin
        fsm_output = 9'b000010110;
        state_var_NS = COMP_LOOP_C_21;
      end
      COMP_LOOP_C_21 : begin
        fsm_output = 9'b000010111;
        state_var_NS = COMP_LOOP_C_22;
      end
      COMP_LOOP_C_22 : begin
        fsm_output = 9'b000011000;
        state_var_NS = COMP_LOOP_C_23;
      end
      COMP_LOOP_C_23 : begin
        fsm_output = 9'b000011001;
        state_var_NS = COMP_LOOP_C_24;
      end
      COMP_LOOP_C_24 : begin
        fsm_output = 9'b000011010;
        state_var_NS = COMP_LOOP_C_25;
      end
      COMP_LOOP_C_25 : begin
        fsm_output = 9'b000011011;
        state_var_NS = COMP_LOOP_C_26;
      end
      COMP_LOOP_C_26 : begin
        fsm_output = 9'b000011100;
        state_var_NS = COMP_LOOP_C_27;
      end
      COMP_LOOP_C_27 : begin
        fsm_output = 9'b000011101;
        state_var_NS = COMP_LOOP_C_28;
      end
      COMP_LOOP_C_28 : begin
        fsm_output = 9'b000011110;
        state_var_NS = COMP_LOOP_C_29;
      end
      COMP_LOOP_C_29 : begin
        fsm_output = 9'b000011111;
        state_var_NS = COMP_LOOP_C_30;
      end
      COMP_LOOP_C_30 : begin
        fsm_output = 9'b000100000;
        state_var_NS = COMP_LOOP_C_31;
      end
      COMP_LOOP_C_31 : begin
        fsm_output = 9'b000100001;
        if ( COMP_LOOP_C_31_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_32;
        end
      end
      COMP_LOOP_C_32 : begin
        fsm_output = 9'b000100010;
        state_var_NS = COMP_LOOP_C_33;
      end
      COMP_LOOP_C_33 : begin
        fsm_output = 9'b000100011;
        state_var_NS = COMP_LOOP_C_34;
      end
      COMP_LOOP_C_34 : begin
        fsm_output = 9'b000100100;
        state_var_NS = COMP_LOOP_C_35;
      end
      COMP_LOOP_C_35 : begin
        fsm_output = 9'b000100101;
        state_var_NS = COMP_LOOP_C_36;
      end
      COMP_LOOP_C_36 : begin
        fsm_output = 9'b000100110;
        state_var_NS = COMP_LOOP_C_37;
      end
      COMP_LOOP_C_37 : begin
        fsm_output = 9'b000100111;
        state_var_NS = COMP_LOOP_C_38;
      end
      COMP_LOOP_C_38 : begin
        fsm_output = 9'b000101000;
        state_var_NS = COMP_LOOP_C_39;
      end
      COMP_LOOP_C_39 : begin
        fsm_output = 9'b000101001;
        state_var_NS = COMP_LOOP_C_40;
      end
      COMP_LOOP_C_40 : begin
        fsm_output = 9'b000101010;
        state_var_NS = COMP_LOOP_C_41;
      end
      COMP_LOOP_C_41 : begin
        fsm_output = 9'b000101011;
        state_var_NS = COMP_LOOP_C_42;
      end
      COMP_LOOP_C_42 : begin
        fsm_output = 9'b000101100;
        state_var_NS = COMP_LOOP_C_43;
      end
      COMP_LOOP_C_43 : begin
        fsm_output = 9'b000101101;
        state_var_NS = COMP_LOOP_C_44;
      end
      COMP_LOOP_C_44 : begin
        fsm_output = 9'b000101110;
        state_var_NS = COMP_LOOP_C_45;
      end
      COMP_LOOP_C_45 : begin
        fsm_output = 9'b000101111;
        state_var_NS = COMP_LOOP_C_46;
      end
      COMP_LOOP_C_46 : begin
        fsm_output = 9'b000110000;
        state_var_NS = COMP_LOOP_C_47;
      end
      COMP_LOOP_C_47 : begin
        fsm_output = 9'b000110001;
        state_var_NS = COMP_LOOP_C_48;
      end
      COMP_LOOP_C_48 : begin
        fsm_output = 9'b000110010;
        state_var_NS = COMP_LOOP_C_49;
      end
      COMP_LOOP_C_49 : begin
        fsm_output = 9'b000110011;
        state_var_NS = COMP_LOOP_C_50;
      end
      COMP_LOOP_C_50 : begin
        fsm_output = 9'b000110100;
        state_var_NS = COMP_LOOP_C_51;
      end
      COMP_LOOP_C_51 : begin
        fsm_output = 9'b000110101;
        state_var_NS = COMP_LOOP_C_52;
      end
      COMP_LOOP_C_52 : begin
        fsm_output = 9'b000110110;
        state_var_NS = COMP_LOOP_C_53;
      end
      COMP_LOOP_C_53 : begin
        fsm_output = 9'b000110111;
        state_var_NS = COMP_LOOP_C_54;
      end
      COMP_LOOP_C_54 : begin
        fsm_output = 9'b000111000;
        state_var_NS = COMP_LOOP_C_55;
      end
      COMP_LOOP_C_55 : begin
        fsm_output = 9'b000111001;
        state_var_NS = COMP_LOOP_C_56;
      end
      COMP_LOOP_C_56 : begin
        fsm_output = 9'b000111010;
        state_var_NS = COMP_LOOP_C_57;
      end
      COMP_LOOP_C_57 : begin
        fsm_output = 9'b000111011;
        state_var_NS = COMP_LOOP_C_58;
      end
      COMP_LOOP_C_58 : begin
        fsm_output = 9'b000111100;
        state_var_NS = COMP_LOOP_C_59;
      end
      COMP_LOOP_C_59 : begin
        fsm_output = 9'b000111101;
        state_var_NS = COMP_LOOP_C_60;
      end
      COMP_LOOP_C_60 : begin
        fsm_output = 9'b000111110;
        state_var_NS = COMP_LOOP_C_61;
      end
      COMP_LOOP_C_61 : begin
        fsm_output = 9'b000111111;
        state_var_NS = COMP_LOOP_C_62;
      end
      COMP_LOOP_C_62 : begin
        fsm_output = 9'b001000000;
        if ( COMP_LOOP_C_62_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_63;
        end
      end
      COMP_LOOP_C_63 : begin
        fsm_output = 9'b001000001;
        state_var_NS = COMP_LOOP_C_64;
      end
      COMP_LOOP_C_64 : begin
        fsm_output = 9'b001000010;
        state_var_NS = COMP_LOOP_C_65;
      end
      COMP_LOOP_C_65 : begin
        fsm_output = 9'b001000011;
        state_var_NS = COMP_LOOP_C_66;
      end
      COMP_LOOP_C_66 : begin
        fsm_output = 9'b001000100;
        state_var_NS = COMP_LOOP_C_67;
      end
      COMP_LOOP_C_67 : begin
        fsm_output = 9'b001000101;
        state_var_NS = COMP_LOOP_C_68;
      end
      COMP_LOOP_C_68 : begin
        fsm_output = 9'b001000110;
        state_var_NS = COMP_LOOP_C_69;
      end
      COMP_LOOP_C_69 : begin
        fsm_output = 9'b001000111;
        state_var_NS = COMP_LOOP_C_70;
      end
      COMP_LOOP_C_70 : begin
        fsm_output = 9'b001001000;
        state_var_NS = COMP_LOOP_C_71;
      end
      COMP_LOOP_C_71 : begin
        fsm_output = 9'b001001001;
        state_var_NS = COMP_LOOP_C_72;
      end
      COMP_LOOP_C_72 : begin
        fsm_output = 9'b001001010;
        state_var_NS = COMP_LOOP_C_73;
      end
      COMP_LOOP_C_73 : begin
        fsm_output = 9'b001001011;
        state_var_NS = COMP_LOOP_C_74;
      end
      COMP_LOOP_C_74 : begin
        fsm_output = 9'b001001100;
        state_var_NS = COMP_LOOP_C_75;
      end
      COMP_LOOP_C_75 : begin
        fsm_output = 9'b001001101;
        state_var_NS = COMP_LOOP_C_76;
      end
      COMP_LOOP_C_76 : begin
        fsm_output = 9'b001001110;
        state_var_NS = COMP_LOOP_C_77;
      end
      COMP_LOOP_C_77 : begin
        fsm_output = 9'b001001111;
        state_var_NS = COMP_LOOP_C_78;
      end
      COMP_LOOP_C_78 : begin
        fsm_output = 9'b001010000;
        state_var_NS = COMP_LOOP_C_79;
      end
      COMP_LOOP_C_79 : begin
        fsm_output = 9'b001010001;
        state_var_NS = COMP_LOOP_C_80;
      end
      COMP_LOOP_C_80 : begin
        fsm_output = 9'b001010010;
        state_var_NS = COMP_LOOP_C_81;
      end
      COMP_LOOP_C_81 : begin
        fsm_output = 9'b001010011;
        state_var_NS = COMP_LOOP_C_82;
      end
      COMP_LOOP_C_82 : begin
        fsm_output = 9'b001010100;
        state_var_NS = COMP_LOOP_C_83;
      end
      COMP_LOOP_C_83 : begin
        fsm_output = 9'b001010101;
        state_var_NS = COMP_LOOP_C_84;
      end
      COMP_LOOP_C_84 : begin
        fsm_output = 9'b001010110;
        state_var_NS = COMP_LOOP_C_85;
      end
      COMP_LOOP_C_85 : begin
        fsm_output = 9'b001010111;
        state_var_NS = COMP_LOOP_C_86;
      end
      COMP_LOOP_C_86 : begin
        fsm_output = 9'b001011000;
        state_var_NS = COMP_LOOP_C_87;
      end
      COMP_LOOP_C_87 : begin
        fsm_output = 9'b001011001;
        state_var_NS = COMP_LOOP_C_88;
      end
      COMP_LOOP_C_88 : begin
        fsm_output = 9'b001011010;
        state_var_NS = COMP_LOOP_C_89;
      end
      COMP_LOOP_C_89 : begin
        fsm_output = 9'b001011011;
        state_var_NS = COMP_LOOP_C_90;
      end
      COMP_LOOP_C_90 : begin
        fsm_output = 9'b001011100;
        state_var_NS = COMP_LOOP_C_91;
      end
      COMP_LOOP_C_91 : begin
        fsm_output = 9'b001011101;
        state_var_NS = COMP_LOOP_C_92;
      end
      COMP_LOOP_C_92 : begin
        fsm_output = 9'b001011110;
        state_var_NS = COMP_LOOP_C_93;
      end
      COMP_LOOP_C_93 : begin
        fsm_output = 9'b001011111;
        if ( COMP_LOOP_C_93_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_94;
        end
      end
      COMP_LOOP_C_94 : begin
        fsm_output = 9'b001100000;
        state_var_NS = COMP_LOOP_C_95;
      end
      COMP_LOOP_C_95 : begin
        fsm_output = 9'b001100001;
        state_var_NS = COMP_LOOP_C_96;
      end
      COMP_LOOP_C_96 : begin
        fsm_output = 9'b001100010;
        state_var_NS = COMP_LOOP_C_97;
      end
      COMP_LOOP_C_97 : begin
        fsm_output = 9'b001100011;
        state_var_NS = COMP_LOOP_C_98;
      end
      COMP_LOOP_C_98 : begin
        fsm_output = 9'b001100100;
        state_var_NS = COMP_LOOP_C_99;
      end
      COMP_LOOP_C_99 : begin
        fsm_output = 9'b001100101;
        state_var_NS = COMP_LOOP_C_100;
      end
      COMP_LOOP_C_100 : begin
        fsm_output = 9'b001100110;
        state_var_NS = COMP_LOOP_C_101;
      end
      COMP_LOOP_C_101 : begin
        fsm_output = 9'b001100111;
        state_var_NS = COMP_LOOP_C_102;
      end
      COMP_LOOP_C_102 : begin
        fsm_output = 9'b001101000;
        state_var_NS = COMP_LOOP_C_103;
      end
      COMP_LOOP_C_103 : begin
        fsm_output = 9'b001101001;
        state_var_NS = COMP_LOOP_C_104;
      end
      COMP_LOOP_C_104 : begin
        fsm_output = 9'b001101010;
        state_var_NS = COMP_LOOP_C_105;
      end
      COMP_LOOP_C_105 : begin
        fsm_output = 9'b001101011;
        state_var_NS = COMP_LOOP_C_106;
      end
      COMP_LOOP_C_106 : begin
        fsm_output = 9'b001101100;
        state_var_NS = COMP_LOOP_C_107;
      end
      COMP_LOOP_C_107 : begin
        fsm_output = 9'b001101101;
        state_var_NS = COMP_LOOP_C_108;
      end
      COMP_LOOP_C_108 : begin
        fsm_output = 9'b001101110;
        state_var_NS = COMP_LOOP_C_109;
      end
      COMP_LOOP_C_109 : begin
        fsm_output = 9'b001101111;
        state_var_NS = COMP_LOOP_C_110;
      end
      COMP_LOOP_C_110 : begin
        fsm_output = 9'b001110000;
        state_var_NS = COMP_LOOP_C_111;
      end
      COMP_LOOP_C_111 : begin
        fsm_output = 9'b001110001;
        state_var_NS = COMP_LOOP_C_112;
      end
      COMP_LOOP_C_112 : begin
        fsm_output = 9'b001110010;
        state_var_NS = COMP_LOOP_C_113;
      end
      COMP_LOOP_C_113 : begin
        fsm_output = 9'b001110011;
        state_var_NS = COMP_LOOP_C_114;
      end
      COMP_LOOP_C_114 : begin
        fsm_output = 9'b001110100;
        state_var_NS = COMP_LOOP_C_115;
      end
      COMP_LOOP_C_115 : begin
        fsm_output = 9'b001110101;
        state_var_NS = COMP_LOOP_C_116;
      end
      COMP_LOOP_C_116 : begin
        fsm_output = 9'b001110110;
        state_var_NS = COMP_LOOP_C_117;
      end
      COMP_LOOP_C_117 : begin
        fsm_output = 9'b001110111;
        state_var_NS = COMP_LOOP_C_118;
      end
      COMP_LOOP_C_118 : begin
        fsm_output = 9'b001111000;
        state_var_NS = COMP_LOOP_C_119;
      end
      COMP_LOOP_C_119 : begin
        fsm_output = 9'b001111001;
        state_var_NS = COMP_LOOP_C_120;
      end
      COMP_LOOP_C_120 : begin
        fsm_output = 9'b001111010;
        state_var_NS = COMP_LOOP_C_121;
      end
      COMP_LOOP_C_121 : begin
        fsm_output = 9'b001111011;
        state_var_NS = COMP_LOOP_C_122;
      end
      COMP_LOOP_C_122 : begin
        fsm_output = 9'b001111100;
        state_var_NS = COMP_LOOP_C_123;
      end
      COMP_LOOP_C_123 : begin
        fsm_output = 9'b001111101;
        state_var_NS = COMP_LOOP_C_124;
      end
      COMP_LOOP_C_124 : begin
        fsm_output = 9'b001111110;
        if ( COMP_LOOP_C_124_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_125;
        end
      end
      COMP_LOOP_C_125 : begin
        fsm_output = 9'b001111111;
        state_var_NS = COMP_LOOP_C_126;
      end
      COMP_LOOP_C_126 : begin
        fsm_output = 9'b010000000;
        state_var_NS = COMP_LOOP_C_127;
      end
      COMP_LOOP_C_127 : begin
        fsm_output = 9'b010000001;
        state_var_NS = COMP_LOOP_C_128;
      end
      COMP_LOOP_C_128 : begin
        fsm_output = 9'b010000010;
        state_var_NS = COMP_LOOP_C_129;
      end
      COMP_LOOP_C_129 : begin
        fsm_output = 9'b010000011;
        state_var_NS = COMP_LOOP_C_130;
      end
      COMP_LOOP_C_130 : begin
        fsm_output = 9'b010000100;
        state_var_NS = COMP_LOOP_C_131;
      end
      COMP_LOOP_C_131 : begin
        fsm_output = 9'b010000101;
        state_var_NS = COMP_LOOP_C_132;
      end
      COMP_LOOP_C_132 : begin
        fsm_output = 9'b010000110;
        state_var_NS = COMP_LOOP_C_133;
      end
      COMP_LOOP_C_133 : begin
        fsm_output = 9'b010000111;
        state_var_NS = COMP_LOOP_C_134;
      end
      COMP_LOOP_C_134 : begin
        fsm_output = 9'b010001000;
        state_var_NS = COMP_LOOP_C_135;
      end
      COMP_LOOP_C_135 : begin
        fsm_output = 9'b010001001;
        state_var_NS = COMP_LOOP_C_136;
      end
      COMP_LOOP_C_136 : begin
        fsm_output = 9'b010001010;
        state_var_NS = COMP_LOOP_C_137;
      end
      COMP_LOOP_C_137 : begin
        fsm_output = 9'b010001011;
        state_var_NS = COMP_LOOP_C_138;
      end
      COMP_LOOP_C_138 : begin
        fsm_output = 9'b010001100;
        state_var_NS = COMP_LOOP_C_139;
      end
      COMP_LOOP_C_139 : begin
        fsm_output = 9'b010001101;
        state_var_NS = COMP_LOOP_C_140;
      end
      COMP_LOOP_C_140 : begin
        fsm_output = 9'b010001110;
        state_var_NS = COMP_LOOP_C_141;
      end
      COMP_LOOP_C_141 : begin
        fsm_output = 9'b010001111;
        state_var_NS = COMP_LOOP_C_142;
      end
      COMP_LOOP_C_142 : begin
        fsm_output = 9'b010010000;
        state_var_NS = COMP_LOOP_C_143;
      end
      COMP_LOOP_C_143 : begin
        fsm_output = 9'b010010001;
        state_var_NS = COMP_LOOP_C_144;
      end
      COMP_LOOP_C_144 : begin
        fsm_output = 9'b010010010;
        state_var_NS = COMP_LOOP_C_145;
      end
      COMP_LOOP_C_145 : begin
        fsm_output = 9'b010010011;
        state_var_NS = COMP_LOOP_C_146;
      end
      COMP_LOOP_C_146 : begin
        fsm_output = 9'b010010100;
        state_var_NS = COMP_LOOP_C_147;
      end
      COMP_LOOP_C_147 : begin
        fsm_output = 9'b010010101;
        state_var_NS = COMP_LOOP_C_148;
      end
      COMP_LOOP_C_148 : begin
        fsm_output = 9'b010010110;
        state_var_NS = COMP_LOOP_C_149;
      end
      COMP_LOOP_C_149 : begin
        fsm_output = 9'b010010111;
        state_var_NS = COMP_LOOP_C_150;
      end
      COMP_LOOP_C_150 : begin
        fsm_output = 9'b010011000;
        state_var_NS = COMP_LOOP_C_151;
      end
      COMP_LOOP_C_151 : begin
        fsm_output = 9'b010011001;
        state_var_NS = COMP_LOOP_C_152;
      end
      COMP_LOOP_C_152 : begin
        fsm_output = 9'b010011010;
        state_var_NS = COMP_LOOP_C_153;
      end
      COMP_LOOP_C_153 : begin
        fsm_output = 9'b010011011;
        state_var_NS = COMP_LOOP_C_154;
      end
      COMP_LOOP_C_154 : begin
        fsm_output = 9'b010011100;
        state_var_NS = COMP_LOOP_C_155;
      end
      COMP_LOOP_C_155 : begin
        fsm_output = 9'b010011101;
        if ( COMP_LOOP_C_155_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_156;
        end
      end
      COMP_LOOP_C_156 : begin
        fsm_output = 9'b010011110;
        state_var_NS = COMP_LOOP_C_157;
      end
      COMP_LOOP_C_157 : begin
        fsm_output = 9'b010011111;
        state_var_NS = COMP_LOOP_C_158;
      end
      COMP_LOOP_C_158 : begin
        fsm_output = 9'b010100000;
        state_var_NS = COMP_LOOP_C_159;
      end
      COMP_LOOP_C_159 : begin
        fsm_output = 9'b010100001;
        state_var_NS = COMP_LOOP_C_160;
      end
      COMP_LOOP_C_160 : begin
        fsm_output = 9'b010100010;
        state_var_NS = COMP_LOOP_C_161;
      end
      COMP_LOOP_C_161 : begin
        fsm_output = 9'b010100011;
        state_var_NS = COMP_LOOP_C_162;
      end
      COMP_LOOP_C_162 : begin
        fsm_output = 9'b010100100;
        state_var_NS = COMP_LOOP_C_163;
      end
      COMP_LOOP_C_163 : begin
        fsm_output = 9'b010100101;
        state_var_NS = COMP_LOOP_C_164;
      end
      COMP_LOOP_C_164 : begin
        fsm_output = 9'b010100110;
        state_var_NS = COMP_LOOP_C_165;
      end
      COMP_LOOP_C_165 : begin
        fsm_output = 9'b010100111;
        state_var_NS = COMP_LOOP_C_166;
      end
      COMP_LOOP_C_166 : begin
        fsm_output = 9'b010101000;
        state_var_NS = COMP_LOOP_C_167;
      end
      COMP_LOOP_C_167 : begin
        fsm_output = 9'b010101001;
        state_var_NS = COMP_LOOP_C_168;
      end
      COMP_LOOP_C_168 : begin
        fsm_output = 9'b010101010;
        state_var_NS = COMP_LOOP_C_169;
      end
      COMP_LOOP_C_169 : begin
        fsm_output = 9'b010101011;
        state_var_NS = COMP_LOOP_C_170;
      end
      COMP_LOOP_C_170 : begin
        fsm_output = 9'b010101100;
        state_var_NS = COMP_LOOP_C_171;
      end
      COMP_LOOP_C_171 : begin
        fsm_output = 9'b010101101;
        state_var_NS = COMP_LOOP_C_172;
      end
      COMP_LOOP_C_172 : begin
        fsm_output = 9'b010101110;
        state_var_NS = COMP_LOOP_C_173;
      end
      COMP_LOOP_C_173 : begin
        fsm_output = 9'b010101111;
        state_var_NS = COMP_LOOP_C_174;
      end
      COMP_LOOP_C_174 : begin
        fsm_output = 9'b010110000;
        state_var_NS = COMP_LOOP_C_175;
      end
      COMP_LOOP_C_175 : begin
        fsm_output = 9'b010110001;
        state_var_NS = COMP_LOOP_C_176;
      end
      COMP_LOOP_C_176 : begin
        fsm_output = 9'b010110010;
        state_var_NS = COMP_LOOP_C_177;
      end
      COMP_LOOP_C_177 : begin
        fsm_output = 9'b010110011;
        state_var_NS = COMP_LOOP_C_178;
      end
      COMP_LOOP_C_178 : begin
        fsm_output = 9'b010110100;
        state_var_NS = COMP_LOOP_C_179;
      end
      COMP_LOOP_C_179 : begin
        fsm_output = 9'b010110101;
        state_var_NS = COMP_LOOP_C_180;
      end
      COMP_LOOP_C_180 : begin
        fsm_output = 9'b010110110;
        state_var_NS = COMP_LOOP_C_181;
      end
      COMP_LOOP_C_181 : begin
        fsm_output = 9'b010110111;
        state_var_NS = COMP_LOOP_C_182;
      end
      COMP_LOOP_C_182 : begin
        fsm_output = 9'b010111000;
        state_var_NS = COMP_LOOP_C_183;
      end
      COMP_LOOP_C_183 : begin
        fsm_output = 9'b010111001;
        state_var_NS = COMP_LOOP_C_184;
      end
      COMP_LOOP_C_184 : begin
        fsm_output = 9'b010111010;
        state_var_NS = COMP_LOOP_C_185;
      end
      COMP_LOOP_C_185 : begin
        fsm_output = 9'b010111011;
        state_var_NS = COMP_LOOP_C_186;
      end
      COMP_LOOP_C_186 : begin
        fsm_output = 9'b010111100;
        if ( COMP_LOOP_C_186_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_187;
        end
      end
      COMP_LOOP_C_187 : begin
        fsm_output = 9'b010111101;
        state_var_NS = COMP_LOOP_C_188;
      end
      COMP_LOOP_C_188 : begin
        fsm_output = 9'b010111110;
        state_var_NS = COMP_LOOP_C_189;
      end
      COMP_LOOP_C_189 : begin
        fsm_output = 9'b010111111;
        state_var_NS = COMP_LOOP_C_190;
      end
      COMP_LOOP_C_190 : begin
        fsm_output = 9'b011000000;
        state_var_NS = COMP_LOOP_C_191;
      end
      COMP_LOOP_C_191 : begin
        fsm_output = 9'b011000001;
        state_var_NS = COMP_LOOP_C_192;
      end
      COMP_LOOP_C_192 : begin
        fsm_output = 9'b011000010;
        state_var_NS = COMP_LOOP_C_193;
      end
      COMP_LOOP_C_193 : begin
        fsm_output = 9'b011000011;
        state_var_NS = COMP_LOOP_C_194;
      end
      COMP_LOOP_C_194 : begin
        fsm_output = 9'b011000100;
        state_var_NS = COMP_LOOP_C_195;
      end
      COMP_LOOP_C_195 : begin
        fsm_output = 9'b011000101;
        state_var_NS = COMP_LOOP_C_196;
      end
      COMP_LOOP_C_196 : begin
        fsm_output = 9'b011000110;
        state_var_NS = COMP_LOOP_C_197;
      end
      COMP_LOOP_C_197 : begin
        fsm_output = 9'b011000111;
        state_var_NS = COMP_LOOP_C_198;
      end
      COMP_LOOP_C_198 : begin
        fsm_output = 9'b011001000;
        state_var_NS = COMP_LOOP_C_199;
      end
      COMP_LOOP_C_199 : begin
        fsm_output = 9'b011001001;
        state_var_NS = COMP_LOOP_C_200;
      end
      COMP_LOOP_C_200 : begin
        fsm_output = 9'b011001010;
        state_var_NS = COMP_LOOP_C_201;
      end
      COMP_LOOP_C_201 : begin
        fsm_output = 9'b011001011;
        state_var_NS = COMP_LOOP_C_202;
      end
      COMP_LOOP_C_202 : begin
        fsm_output = 9'b011001100;
        state_var_NS = COMP_LOOP_C_203;
      end
      COMP_LOOP_C_203 : begin
        fsm_output = 9'b011001101;
        state_var_NS = COMP_LOOP_C_204;
      end
      COMP_LOOP_C_204 : begin
        fsm_output = 9'b011001110;
        state_var_NS = COMP_LOOP_C_205;
      end
      COMP_LOOP_C_205 : begin
        fsm_output = 9'b011001111;
        state_var_NS = COMP_LOOP_C_206;
      end
      COMP_LOOP_C_206 : begin
        fsm_output = 9'b011010000;
        state_var_NS = COMP_LOOP_C_207;
      end
      COMP_LOOP_C_207 : begin
        fsm_output = 9'b011010001;
        state_var_NS = COMP_LOOP_C_208;
      end
      COMP_LOOP_C_208 : begin
        fsm_output = 9'b011010010;
        state_var_NS = COMP_LOOP_C_209;
      end
      COMP_LOOP_C_209 : begin
        fsm_output = 9'b011010011;
        state_var_NS = COMP_LOOP_C_210;
      end
      COMP_LOOP_C_210 : begin
        fsm_output = 9'b011010100;
        state_var_NS = COMP_LOOP_C_211;
      end
      COMP_LOOP_C_211 : begin
        fsm_output = 9'b011010101;
        state_var_NS = COMP_LOOP_C_212;
      end
      COMP_LOOP_C_212 : begin
        fsm_output = 9'b011010110;
        state_var_NS = COMP_LOOP_C_213;
      end
      COMP_LOOP_C_213 : begin
        fsm_output = 9'b011010111;
        state_var_NS = COMP_LOOP_C_214;
      end
      COMP_LOOP_C_214 : begin
        fsm_output = 9'b011011000;
        state_var_NS = COMP_LOOP_C_215;
      end
      COMP_LOOP_C_215 : begin
        fsm_output = 9'b011011001;
        state_var_NS = COMP_LOOP_C_216;
      end
      COMP_LOOP_C_216 : begin
        fsm_output = 9'b011011010;
        state_var_NS = COMP_LOOP_C_217;
      end
      COMP_LOOP_C_217 : begin
        fsm_output = 9'b011011011;
        if ( COMP_LOOP_C_217_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_218;
        end
      end
      COMP_LOOP_C_218 : begin
        fsm_output = 9'b011011100;
        state_var_NS = COMP_LOOP_C_219;
      end
      COMP_LOOP_C_219 : begin
        fsm_output = 9'b011011101;
        state_var_NS = COMP_LOOP_C_220;
      end
      COMP_LOOP_C_220 : begin
        fsm_output = 9'b011011110;
        state_var_NS = COMP_LOOP_C_221;
      end
      COMP_LOOP_C_221 : begin
        fsm_output = 9'b011011111;
        state_var_NS = COMP_LOOP_C_222;
      end
      COMP_LOOP_C_222 : begin
        fsm_output = 9'b011100000;
        state_var_NS = COMP_LOOP_C_223;
      end
      COMP_LOOP_C_223 : begin
        fsm_output = 9'b011100001;
        state_var_NS = COMP_LOOP_C_224;
      end
      COMP_LOOP_C_224 : begin
        fsm_output = 9'b011100010;
        state_var_NS = COMP_LOOP_C_225;
      end
      COMP_LOOP_C_225 : begin
        fsm_output = 9'b011100011;
        state_var_NS = COMP_LOOP_C_226;
      end
      COMP_LOOP_C_226 : begin
        fsm_output = 9'b011100100;
        state_var_NS = COMP_LOOP_C_227;
      end
      COMP_LOOP_C_227 : begin
        fsm_output = 9'b011100101;
        state_var_NS = COMP_LOOP_C_228;
      end
      COMP_LOOP_C_228 : begin
        fsm_output = 9'b011100110;
        state_var_NS = COMP_LOOP_C_229;
      end
      COMP_LOOP_C_229 : begin
        fsm_output = 9'b011100111;
        state_var_NS = COMP_LOOP_C_230;
      end
      COMP_LOOP_C_230 : begin
        fsm_output = 9'b011101000;
        state_var_NS = COMP_LOOP_C_231;
      end
      COMP_LOOP_C_231 : begin
        fsm_output = 9'b011101001;
        state_var_NS = COMP_LOOP_C_232;
      end
      COMP_LOOP_C_232 : begin
        fsm_output = 9'b011101010;
        state_var_NS = COMP_LOOP_C_233;
      end
      COMP_LOOP_C_233 : begin
        fsm_output = 9'b011101011;
        state_var_NS = COMP_LOOP_C_234;
      end
      COMP_LOOP_C_234 : begin
        fsm_output = 9'b011101100;
        state_var_NS = COMP_LOOP_C_235;
      end
      COMP_LOOP_C_235 : begin
        fsm_output = 9'b011101101;
        state_var_NS = COMP_LOOP_C_236;
      end
      COMP_LOOP_C_236 : begin
        fsm_output = 9'b011101110;
        state_var_NS = COMP_LOOP_C_237;
      end
      COMP_LOOP_C_237 : begin
        fsm_output = 9'b011101111;
        state_var_NS = COMP_LOOP_C_238;
      end
      COMP_LOOP_C_238 : begin
        fsm_output = 9'b011110000;
        state_var_NS = COMP_LOOP_C_239;
      end
      COMP_LOOP_C_239 : begin
        fsm_output = 9'b011110001;
        state_var_NS = COMP_LOOP_C_240;
      end
      COMP_LOOP_C_240 : begin
        fsm_output = 9'b011110010;
        state_var_NS = COMP_LOOP_C_241;
      end
      COMP_LOOP_C_241 : begin
        fsm_output = 9'b011110011;
        state_var_NS = COMP_LOOP_C_242;
      end
      COMP_LOOP_C_242 : begin
        fsm_output = 9'b011110100;
        state_var_NS = COMP_LOOP_C_243;
      end
      COMP_LOOP_C_243 : begin
        fsm_output = 9'b011110101;
        state_var_NS = COMP_LOOP_C_244;
      end
      COMP_LOOP_C_244 : begin
        fsm_output = 9'b011110110;
        state_var_NS = COMP_LOOP_C_245;
      end
      COMP_LOOP_C_245 : begin
        fsm_output = 9'b011110111;
        state_var_NS = COMP_LOOP_C_246;
      end
      COMP_LOOP_C_246 : begin
        fsm_output = 9'b011111000;
        state_var_NS = COMP_LOOP_C_247;
      end
      COMP_LOOP_C_247 : begin
        fsm_output = 9'b011111001;
        state_var_NS = COMP_LOOP_C_248;
      end
      COMP_LOOP_C_248 : begin
        fsm_output = 9'b011111010;
        if ( COMP_LOOP_C_248_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_249;
        end
      end
      COMP_LOOP_C_249 : begin
        fsm_output = 9'b011111011;
        state_var_NS = COMP_LOOP_C_250;
      end
      COMP_LOOP_C_250 : begin
        fsm_output = 9'b011111100;
        state_var_NS = COMP_LOOP_C_251;
      end
      COMP_LOOP_C_251 : begin
        fsm_output = 9'b011111101;
        state_var_NS = COMP_LOOP_C_252;
      end
      COMP_LOOP_C_252 : begin
        fsm_output = 9'b011111110;
        state_var_NS = COMP_LOOP_C_253;
      end
      COMP_LOOP_C_253 : begin
        fsm_output = 9'b011111111;
        state_var_NS = COMP_LOOP_C_254;
      end
      COMP_LOOP_C_254 : begin
        fsm_output = 9'b100000000;
        state_var_NS = COMP_LOOP_C_255;
      end
      COMP_LOOP_C_255 : begin
        fsm_output = 9'b100000001;
        state_var_NS = COMP_LOOP_C_256;
      end
      COMP_LOOP_C_256 : begin
        fsm_output = 9'b100000010;
        state_var_NS = COMP_LOOP_C_257;
      end
      COMP_LOOP_C_257 : begin
        fsm_output = 9'b100000011;
        state_var_NS = COMP_LOOP_C_258;
      end
      COMP_LOOP_C_258 : begin
        fsm_output = 9'b100000100;
        state_var_NS = COMP_LOOP_C_259;
      end
      COMP_LOOP_C_259 : begin
        fsm_output = 9'b100000101;
        state_var_NS = COMP_LOOP_C_260;
      end
      COMP_LOOP_C_260 : begin
        fsm_output = 9'b100000110;
        state_var_NS = COMP_LOOP_C_261;
      end
      COMP_LOOP_C_261 : begin
        fsm_output = 9'b100000111;
        state_var_NS = COMP_LOOP_C_262;
      end
      COMP_LOOP_C_262 : begin
        fsm_output = 9'b100001000;
        state_var_NS = COMP_LOOP_C_263;
      end
      COMP_LOOP_C_263 : begin
        fsm_output = 9'b100001001;
        state_var_NS = COMP_LOOP_C_264;
      end
      COMP_LOOP_C_264 : begin
        fsm_output = 9'b100001010;
        state_var_NS = COMP_LOOP_C_265;
      end
      COMP_LOOP_C_265 : begin
        fsm_output = 9'b100001011;
        state_var_NS = COMP_LOOP_C_266;
      end
      COMP_LOOP_C_266 : begin
        fsm_output = 9'b100001100;
        state_var_NS = COMP_LOOP_C_267;
      end
      COMP_LOOP_C_267 : begin
        fsm_output = 9'b100001101;
        state_var_NS = COMP_LOOP_C_268;
      end
      COMP_LOOP_C_268 : begin
        fsm_output = 9'b100001110;
        state_var_NS = COMP_LOOP_C_269;
      end
      COMP_LOOP_C_269 : begin
        fsm_output = 9'b100001111;
        state_var_NS = COMP_LOOP_C_270;
      end
      COMP_LOOP_C_270 : begin
        fsm_output = 9'b100010000;
        state_var_NS = COMP_LOOP_C_271;
      end
      COMP_LOOP_C_271 : begin
        fsm_output = 9'b100010001;
        state_var_NS = COMP_LOOP_C_272;
      end
      COMP_LOOP_C_272 : begin
        fsm_output = 9'b100010010;
        state_var_NS = COMP_LOOP_C_273;
      end
      COMP_LOOP_C_273 : begin
        fsm_output = 9'b100010011;
        state_var_NS = COMP_LOOP_C_274;
      end
      COMP_LOOP_C_274 : begin
        fsm_output = 9'b100010100;
        state_var_NS = COMP_LOOP_C_275;
      end
      COMP_LOOP_C_275 : begin
        fsm_output = 9'b100010101;
        state_var_NS = COMP_LOOP_C_276;
      end
      COMP_LOOP_C_276 : begin
        fsm_output = 9'b100010110;
        state_var_NS = COMP_LOOP_C_277;
      end
      COMP_LOOP_C_277 : begin
        fsm_output = 9'b100010111;
        state_var_NS = COMP_LOOP_C_278;
      end
      COMP_LOOP_C_278 : begin
        fsm_output = 9'b100011000;
        state_var_NS = COMP_LOOP_C_279;
      end
      COMP_LOOP_C_279 : begin
        fsm_output = 9'b100011001;
        if ( COMP_LOOP_C_279_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_280;
        end
      end
      COMP_LOOP_C_280 : begin
        fsm_output = 9'b100011010;
        state_var_NS = COMP_LOOP_C_281;
      end
      COMP_LOOP_C_281 : begin
        fsm_output = 9'b100011011;
        state_var_NS = COMP_LOOP_C_282;
      end
      COMP_LOOP_C_282 : begin
        fsm_output = 9'b100011100;
        state_var_NS = COMP_LOOP_C_283;
      end
      COMP_LOOP_C_283 : begin
        fsm_output = 9'b100011101;
        state_var_NS = COMP_LOOP_C_284;
      end
      COMP_LOOP_C_284 : begin
        fsm_output = 9'b100011110;
        state_var_NS = COMP_LOOP_C_285;
      end
      COMP_LOOP_C_285 : begin
        fsm_output = 9'b100011111;
        state_var_NS = COMP_LOOP_C_286;
      end
      COMP_LOOP_C_286 : begin
        fsm_output = 9'b100100000;
        state_var_NS = COMP_LOOP_C_287;
      end
      COMP_LOOP_C_287 : begin
        fsm_output = 9'b100100001;
        state_var_NS = COMP_LOOP_C_288;
      end
      COMP_LOOP_C_288 : begin
        fsm_output = 9'b100100010;
        state_var_NS = COMP_LOOP_C_289;
      end
      COMP_LOOP_C_289 : begin
        fsm_output = 9'b100100011;
        state_var_NS = COMP_LOOP_C_290;
      end
      COMP_LOOP_C_290 : begin
        fsm_output = 9'b100100100;
        state_var_NS = COMP_LOOP_C_291;
      end
      COMP_LOOP_C_291 : begin
        fsm_output = 9'b100100101;
        state_var_NS = COMP_LOOP_C_292;
      end
      COMP_LOOP_C_292 : begin
        fsm_output = 9'b100100110;
        state_var_NS = COMP_LOOP_C_293;
      end
      COMP_LOOP_C_293 : begin
        fsm_output = 9'b100100111;
        state_var_NS = COMP_LOOP_C_294;
      end
      COMP_LOOP_C_294 : begin
        fsm_output = 9'b100101000;
        state_var_NS = COMP_LOOP_C_295;
      end
      COMP_LOOP_C_295 : begin
        fsm_output = 9'b100101001;
        state_var_NS = COMP_LOOP_C_296;
      end
      COMP_LOOP_C_296 : begin
        fsm_output = 9'b100101010;
        state_var_NS = COMP_LOOP_C_297;
      end
      COMP_LOOP_C_297 : begin
        fsm_output = 9'b100101011;
        state_var_NS = COMP_LOOP_C_298;
      end
      COMP_LOOP_C_298 : begin
        fsm_output = 9'b100101100;
        state_var_NS = COMP_LOOP_C_299;
      end
      COMP_LOOP_C_299 : begin
        fsm_output = 9'b100101101;
        state_var_NS = COMP_LOOP_C_300;
      end
      COMP_LOOP_C_300 : begin
        fsm_output = 9'b100101110;
        state_var_NS = COMP_LOOP_C_301;
      end
      COMP_LOOP_C_301 : begin
        fsm_output = 9'b100101111;
        state_var_NS = COMP_LOOP_C_302;
      end
      COMP_LOOP_C_302 : begin
        fsm_output = 9'b100110000;
        state_var_NS = COMP_LOOP_C_303;
      end
      COMP_LOOP_C_303 : begin
        fsm_output = 9'b100110001;
        state_var_NS = COMP_LOOP_C_304;
      end
      COMP_LOOP_C_304 : begin
        fsm_output = 9'b100110010;
        state_var_NS = COMP_LOOP_C_305;
      end
      COMP_LOOP_C_305 : begin
        fsm_output = 9'b100110011;
        state_var_NS = COMP_LOOP_C_306;
      end
      COMP_LOOP_C_306 : begin
        fsm_output = 9'b100110100;
        state_var_NS = COMP_LOOP_C_307;
      end
      COMP_LOOP_C_307 : begin
        fsm_output = 9'b100110101;
        state_var_NS = COMP_LOOP_C_308;
      end
      COMP_LOOP_C_308 : begin
        fsm_output = 9'b100110110;
        state_var_NS = COMP_LOOP_C_309;
      end
      COMP_LOOP_C_309 : begin
        fsm_output = 9'b100110111;
        state_var_NS = COMP_LOOP_C_310;
      end
      COMP_LOOP_C_310 : begin
        fsm_output = 9'b100111000;
        if ( COMP_LOOP_C_310_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_311;
        end
      end
      COMP_LOOP_C_311 : begin
        fsm_output = 9'b100111001;
        state_var_NS = COMP_LOOP_C_312;
      end
      COMP_LOOP_C_312 : begin
        fsm_output = 9'b100111010;
        state_var_NS = COMP_LOOP_C_313;
      end
      COMP_LOOP_C_313 : begin
        fsm_output = 9'b100111011;
        state_var_NS = COMP_LOOP_C_314;
      end
      COMP_LOOP_C_314 : begin
        fsm_output = 9'b100111100;
        state_var_NS = COMP_LOOP_C_315;
      end
      COMP_LOOP_C_315 : begin
        fsm_output = 9'b100111101;
        state_var_NS = COMP_LOOP_C_316;
      end
      COMP_LOOP_C_316 : begin
        fsm_output = 9'b100111110;
        state_var_NS = COMP_LOOP_C_317;
      end
      COMP_LOOP_C_317 : begin
        fsm_output = 9'b100111111;
        state_var_NS = COMP_LOOP_C_318;
      end
      COMP_LOOP_C_318 : begin
        fsm_output = 9'b101000000;
        state_var_NS = COMP_LOOP_C_319;
      end
      COMP_LOOP_C_319 : begin
        fsm_output = 9'b101000001;
        state_var_NS = COMP_LOOP_C_320;
      end
      COMP_LOOP_C_320 : begin
        fsm_output = 9'b101000010;
        state_var_NS = COMP_LOOP_C_321;
      end
      COMP_LOOP_C_321 : begin
        fsm_output = 9'b101000011;
        state_var_NS = COMP_LOOP_C_322;
      end
      COMP_LOOP_C_322 : begin
        fsm_output = 9'b101000100;
        state_var_NS = COMP_LOOP_C_323;
      end
      COMP_LOOP_C_323 : begin
        fsm_output = 9'b101000101;
        state_var_NS = COMP_LOOP_C_324;
      end
      COMP_LOOP_C_324 : begin
        fsm_output = 9'b101000110;
        state_var_NS = COMP_LOOP_C_325;
      end
      COMP_LOOP_C_325 : begin
        fsm_output = 9'b101000111;
        state_var_NS = COMP_LOOP_C_326;
      end
      COMP_LOOP_C_326 : begin
        fsm_output = 9'b101001000;
        state_var_NS = COMP_LOOP_C_327;
      end
      COMP_LOOP_C_327 : begin
        fsm_output = 9'b101001001;
        state_var_NS = COMP_LOOP_C_328;
      end
      COMP_LOOP_C_328 : begin
        fsm_output = 9'b101001010;
        state_var_NS = COMP_LOOP_C_329;
      end
      COMP_LOOP_C_329 : begin
        fsm_output = 9'b101001011;
        state_var_NS = COMP_LOOP_C_330;
      end
      COMP_LOOP_C_330 : begin
        fsm_output = 9'b101001100;
        state_var_NS = COMP_LOOP_C_331;
      end
      COMP_LOOP_C_331 : begin
        fsm_output = 9'b101001101;
        state_var_NS = COMP_LOOP_C_332;
      end
      COMP_LOOP_C_332 : begin
        fsm_output = 9'b101001110;
        state_var_NS = COMP_LOOP_C_333;
      end
      COMP_LOOP_C_333 : begin
        fsm_output = 9'b101001111;
        state_var_NS = COMP_LOOP_C_334;
      end
      COMP_LOOP_C_334 : begin
        fsm_output = 9'b101010000;
        state_var_NS = COMP_LOOP_C_335;
      end
      COMP_LOOP_C_335 : begin
        fsm_output = 9'b101010001;
        state_var_NS = COMP_LOOP_C_336;
      end
      COMP_LOOP_C_336 : begin
        fsm_output = 9'b101010010;
        state_var_NS = COMP_LOOP_C_337;
      end
      COMP_LOOP_C_337 : begin
        fsm_output = 9'b101010011;
        state_var_NS = COMP_LOOP_C_338;
      end
      COMP_LOOP_C_338 : begin
        fsm_output = 9'b101010100;
        state_var_NS = COMP_LOOP_C_339;
      end
      COMP_LOOP_C_339 : begin
        fsm_output = 9'b101010101;
        state_var_NS = COMP_LOOP_C_340;
      end
      COMP_LOOP_C_340 : begin
        fsm_output = 9'b101010110;
        state_var_NS = COMP_LOOP_C_341;
      end
      COMP_LOOP_C_341 : begin
        fsm_output = 9'b101010111;
        if ( COMP_LOOP_C_341_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_342;
        end
      end
      COMP_LOOP_C_342 : begin
        fsm_output = 9'b101011000;
        state_var_NS = COMP_LOOP_C_343;
      end
      COMP_LOOP_C_343 : begin
        fsm_output = 9'b101011001;
        state_var_NS = COMP_LOOP_C_344;
      end
      COMP_LOOP_C_344 : begin
        fsm_output = 9'b101011010;
        state_var_NS = COMP_LOOP_C_345;
      end
      COMP_LOOP_C_345 : begin
        fsm_output = 9'b101011011;
        state_var_NS = COMP_LOOP_C_346;
      end
      COMP_LOOP_C_346 : begin
        fsm_output = 9'b101011100;
        state_var_NS = COMP_LOOP_C_347;
      end
      COMP_LOOP_C_347 : begin
        fsm_output = 9'b101011101;
        state_var_NS = COMP_LOOP_C_348;
      end
      COMP_LOOP_C_348 : begin
        fsm_output = 9'b101011110;
        state_var_NS = COMP_LOOP_C_349;
      end
      COMP_LOOP_C_349 : begin
        fsm_output = 9'b101011111;
        state_var_NS = COMP_LOOP_C_350;
      end
      COMP_LOOP_C_350 : begin
        fsm_output = 9'b101100000;
        state_var_NS = COMP_LOOP_C_351;
      end
      COMP_LOOP_C_351 : begin
        fsm_output = 9'b101100001;
        state_var_NS = COMP_LOOP_C_352;
      end
      COMP_LOOP_C_352 : begin
        fsm_output = 9'b101100010;
        state_var_NS = COMP_LOOP_C_353;
      end
      COMP_LOOP_C_353 : begin
        fsm_output = 9'b101100011;
        state_var_NS = COMP_LOOP_C_354;
      end
      COMP_LOOP_C_354 : begin
        fsm_output = 9'b101100100;
        state_var_NS = COMP_LOOP_C_355;
      end
      COMP_LOOP_C_355 : begin
        fsm_output = 9'b101100101;
        state_var_NS = COMP_LOOP_C_356;
      end
      COMP_LOOP_C_356 : begin
        fsm_output = 9'b101100110;
        state_var_NS = COMP_LOOP_C_357;
      end
      COMP_LOOP_C_357 : begin
        fsm_output = 9'b101100111;
        state_var_NS = COMP_LOOP_C_358;
      end
      COMP_LOOP_C_358 : begin
        fsm_output = 9'b101101000;
        state_var_NS = COMP_LOOP_C_359;
      end
      COMP_LOOP_C_359 : begin
        fsm_output = 9'b101101001;
        state_var_NS = COMP_LOOP_C_360;
      end
      COMP_LOOP_C_360 : begin
        fsm_output = 9'b101101010;
        state_var_NS = COMP_LOOP_C_361;
      end
      COMP_LOOP_C_361 : begin
        fsm_output = 9'b101101011;
        state_var_NS = COMP_LOOP_C_362;
      end
      COMP_LOOP_C_362 : begin
        fsm_output = 9'b101101100;
        state_var_NS = COMP_LOOP_C_363;
      end
      COMP_LOOP_C_363 : begin
        fsm_output = 9'b101101101;
        state_var_NS = COMP_LOOP_C_364;
      end
      COMP_LOOP_C_364 : begin
        fsm_output = 9'b101101110;
        state_var_NS = COMP_LOOP_C_365;
      end
      COMP_LOOP_C_365 : begin
        fsm_output = 9'b101101111;
        state_var_NS = COMP_LOOP_C_366;
      end
      COMP_LOOP_C_366 : begin
        fsm_output = 9'b101110000;
        state_var_NS = COMP_LOOP_C_367;
      end
      COMP_LOOP_C_367 : begin
        fsm_output = 9'b101110001;
        state_var_NS = COMP_LOOP_C_368;
      end
      COMP_LOOP_C_368 : begin
        fsm_output = 9'b101110010;
        state_var_NS = COMP_LOOP_C_369;
      end
      COMP_LOOP_C_369 : begin
        fsm_output = 9'b101110011;
        state_var_NS = COMP_LOOP_C_370;
      end
      COMP_LOOP_C_370 : begin
        fsm_output = 9'b101110100;
        state_var_NS = COMP_LOOP_C_371;
      end
      COMP_LOOP_C_371 : begin
        fsm_output = 9'b101110101;
        state_var_NS = COMP_LOOP_C_372;
      end
      COMP_LOOP_C_372 : begin
        fsm_output = 9'b101110110;
        if ( COMP_LOOP_C_372_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_373;
        end
      end
      COMP_LOOP_C_373 : begin
        fsm_output = 9'b101110111;
        state_var_NS = COMP_LOOP_C_374;
      end
      COMP_LOOP_C_374 : begin
        fsm_output = 9'b101111000;
        state_var_NS = COMP_LOOP_C_375;
      end
      COMP_LOOP_C_375 : begin
        fsm_output = 9'b101111001;
        state_var_NS = COMP_LOOP_C_376;
      end
      COMP_LOOP_C_376 : begin
        fsm_output = 9'b101111010;
        state_var_NS = COMP_LOOP_C_377;
      end
      COMP_LOOP_C_377 : begin
        fsm_output = 9'b101111011;
        state_var_NS = COMP_LOOP_C_378;
      end
      COMP_LOOP_C_378 : begin
        fsm_output = 9'b101111100;
        state_var_NS = COMP_LOOP_C_379;
      end
      COMP_LOOP_C_379 : begin
        fsm_output = 9'b101111101;
        state_var_NS = COMP_LOOP_C_380;
      end
      COMP_LOOP_C_380 : begin
        fsm_output = 9'b101111110;
        state_var_NS = COMP_LOOP_C_381;
      end
      COMP_LOOP_C_381 : begin
        fsm_output = 9'b101111111;
        state_var_NS = COMP_LOOP_C_382;
      end
      COMP_LOOP_C_382 : begin
        fsm_output = 9'b110000000;
        state_var_NS = COMP_LOOP_C_383;
      end
      COMP_LOOP_C_383 : begin
        fsm_output = 9'b110000001;
        state_var_NS = COMP_LOOP_C_384;
      end
      COMP_LOOP_C_384 : begin
        fsm_output = 9'b110000010;
        state_var_NS = COMP_LOOP_C_385;
      end
      COMP_LOOP_C_385 : begin
        fsm_output = 9'b110000011;
        state_var_NS = COMP_LOOP_C_386;
      end
      COMP_LOOP_C_386 : begin
        fsm_output = 9'b110000100;
        state_var_NS = COMP_LOOP_C_387;
      end
      COMP_LOOP_C_387 : begin
        fsm_output = 9'b110000101;
        state_var_NS = COMP_LOOP_C_388;
      end
      COMP_LOOP_C_388 : begin
        fsm_output = 9'b110000110;
        state_var_NS = COMP_LOOP_C_389;
      end
      COMP_LOOP_C_389 : begin
        fsm_output = 9'b110000111;
        state_var_NS = COMP_LOOP_C_390;
      end
      COMP_LOOP_C_390 : begin
        fsm_output = 9'b110001000;
        state_var_NS = COMP_LOOP_C_391;
      end
      COMP_LOOP_C_391 : begin
        fsm_output = 9'b110001001;
        state_var_NS = COMP_LOOP_C_392;
      end
      COMP_LOOP_C_392 : begin
        fsm_output = 9'b110001010;
        state_var_NS = COMP_LOOP_C_393;
      end
      COMP_LOOP_C_393 : begin
        fsm_output = 9'b110001011;
        state_var_NS = COMP_LOOP_C_394;
      end
      COMP_LOOP_C_394 : begin
        fsm_output = 9'b110001100;
        state_var_NS = COMP_LOOP_C_395;
      end
      COMP_LOOP_C_395 : begin
        fsm_output = 9'b110001101;
        state_var_NS = COMP_LOOP_C_396;
      end
      COMP_LOOP_C_396 : begin
        fsm_output = 9'b110001110;
        state_var_NS = COMP_LOOP_C_397;
      end
      COMP_LOOP_C_397 : begin
        fsm_output = 9'b110001111;
        state_var_NS = COMP_LOOP_C_398;
      end
      COMP_LOOP_C_398 : begin
        fsm_output = 9'b110010000;
        state_var_NS = COMP_LOOP_C_399;
      end
      COMP_LOOP_C_399 : begin
        fsm_output = 9'b110010001;
        state_var_NS = COMP_LOOP_C_400;
      end
      COMP_LOOP_C_400 : begin
        fsm_output = 9'b110010010;
        state_var_NS = COMP_LOOP_C_401;
      end
      COMP_LOOP_C_401 : begin
        fsm_output = 9'b110010011;
        state_var_NS = COMP_LOOP_C_402;
      end
      COMP_LOOP_C_402 : begin
        fsm_output = 9'b110010100;
        state_var_NS = COMP_LOOP_C_403;
      end
      COMP_LOOP_C_403 : begin
        fsm_output = 9'b110010101;
        if ( COMP_LOOP_C_403_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_404;
        end
      end
      COMP_LOOP_C_404 : begin
        fsm_output = 9'b110010110;
        state_var_NS = COMP_LOOP_C_405;
      end
      COMP_LOOP_C_405 : begin
        fsm_output = 9'b110010111;
        state_var_NS = COMP_LOOP_C_406;
      end
      COMP_LOOP_C_406 : begin
        fsm_output = 9'b110011000;
        state_var_NS = COMP_LOOP_C_407;
      end
      COMP_LOOP_C_407 : begin
        fsm_output = 9'b110011001;
        state_var_NS = COMP_LOOP_C_408;
      end
      COMP_LOOP_C_408 : begin
        fsm_output = 9'b110011010;
        state_var_NS = COMP_LOOP_C_409;
      end
      COMP_LOOP_C_409 : begin
        fsm_output = 9'b110011011;
        state_var_NS = COMP_LOOP_C_410;
      end
      COMP_LOOP_C_410 : begin
        fsm_output = 9'b110011100;
        state_var_NS = COMP_LOOP_C_411;
      end
      COMP_LOOP_C_411 : begin
        fsm_output = 9'b110011101;
        state_var_NS = COMP_LOOP_C_412;
      end
      COMP_LOOP_C_412 : begin
        fsm_output = 9'b110011110;
        state_var_NS = COMP_LOOP_C_413;
      end
      COMP_LOOP_C_413 : begin
        fsm_output = 9'b110011111;
        state_var_NS = COMP_LOOP_C_414;
      end
      COMP_LOOP_C_414 : begin
        fsm_output = 9'b110100000;
        state_var_NS = COMP_LOOP_C_415;
      end
      COMP_LOOP_C_415 : begin
        fsm_output = 9'b110100001;
        state_var_NS = COMP_LOOP_C_416;
      end
      COMP_LOOP_C_416 : begin
        fsm_output = 9'b110100010;
        state_var_NS = COMP_LOOP_C_417;
      end
      COMP_LOOP_C_417 : begin
        fsm_output = 9'b110100011;
        state_var_NS = COMP_LOOP_C_418;
      end
      COMP_LOOP_C_418 : begin
        fsm_output = 9'b110100100;
        state_var_NS = COMP_LOOP_C_419;
      end
      COMP_LOOP_C_419 : begin
        fsm_output = 9'b110100101;
        state_var_NS = COMP_LOOP_C_420;
      end
      COMP_LOOP_C_420 : begin
        fsm_output = 9'b110100110;
        state_var_NS = COMP_LOOP_C_421;
      end
      COMP_LOOP_C_421 : begin
        fsm_output = 9'b110100111;
        state_var_NS = COMP_LOOP_C_422;
      end
      COMP_LOOP_C_422 : begin
        fsm_output = 9'b110101000;
        state_var_NS = COMP_LOOP_C_423;
      end
      COMP_LOOP_C_423 : begin
        fsm_output = 9'b110101001;
        state_var_NS = COMP_LOOP_C_424;
      end
      COMP_LOOP_C_424 : begin
        fsm_output = 9'b110101010;
        state_var_NS = COMP_LOOP_C_425;
      end
      COMP_LOOP_C_425 : begin
        fsm_output = 9'b110101011;
        state_var_NS = COMP_LOOP_C_426;
      end
      COMP_LOOP_C_426 : begin
        fsm_output = 9'b110101100;
        state_var_NS = COMP_LOOP_C_427;
      end
      COMP_LOOP_C_427 : begin
        fsm_output = 9'b110101101;
        state_var_NS = COMP_LOOP_C_428;
      end
      COMP_LOOP_C_428 : begin
        fsm_output = 9'b110101110;
        state_var_NS = COMP_LOOP_C_429;
      end
      COMP_LOOP_C_429 : begin
        fsm_output = 9'b110101111;
        state_var_NS = COMP_LOOP_C_430;
      end
      COMP_LOOP_C_430 : begin
        fsm_output = 9'b110110000;
        state_var_NS = COMP_LOOP_C_431;
      end
      COMP_LOOP_C_431 : begin
        fsm_output = 9'b110110001;
        state_var_NS = COMP_LOOP_C_432;
      end
      COMP_LOOP_C_432 : begin
        fsm_output = 9'b110110010;
        state_var_NS = COMP_LOOP_C_433;
      end
      COMP_LOOP_C_433 : begin
        fsm_output = 9'b110110011;
        state_var_NS = COMP_LOOP_C_434;
      end
      COMP_LOOP_C_434 : begin
        fsm_output = 9'b110110100;
        if ( COMP_LOOP_C_434_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_435;
        end
      end
      COMP_LOOP_C_435 : begin
        fsm_output = 9'b110110101;
        state_var_NS = COMP_LOOP_C_436;
      end
      COMP_LOOP_C_436 : begin
        fsm_output = 9'b110110110;
        state_var_NS = COMP_LOOP_C_437;
      end
      COMP_LOOP_C_437 : begin
        fsm_output = 9'b110110111;
        state_var_NS = COMP_LOOP_C_438;
      end
      COMP_LOOP_C_438 : begin
        fsm_output = 9'b110111000;
        state_var_NS = COMP_LOOP_C_439;
      end
      COMP_LOOP_C_439 : begin
        fsm_output = 9'b110111001;
        state_var_NS = COMP_LOOP_C_440;
      end
      COMP_LOOP_C_440 : begin
        fsm_output = 9'b110111010;
        state_var_NS = COMP_LOOP_C_441;
      end
      COMP_LOOP_C_441 : begin
        fsm_output = 9'b110111011;
        state_var_NS = COMP_LOOP_C_442;
      end
      COMP_LOOP_C_442 : begin
        fsm_output = 9'b110111100;
        state_var_NS = COMP_LOOP_C_443;
      end
      COMP_LOOP_C_443 : begin
        fsm_output = 9'b110111101;
        state_var_NS = COMP_LOOP_C_444;
      end
      COMP_LOOP_C_444 : begin
        fsm_output = 9'b110111110;
        state_var_NS = COMP_LOOP_C_445;
      end
      COMP_LOOP_C_445 : begin
        fsm_output = 9'b110111111;
        state_var_NS = COMP_LOOP_C_446;
      end
      COMP_LOOP_C_446 : begin
        fsm_output = 9'b111000000;
        state_var_NS = COMP_LOOP_C_447;
      end
      COMP_LOOP_C_447 : begin
        fsm_output = 9'b111000001;
        state_var_NS = COMP_LOOP_C_448;
      end
      COMP_LOOP_C_448 : begin
        fsm_output = 9'b111000010;
        state_var_NS = COMP_LOOP_C_449;
      end
      COMP_LOOP_C_449 : begin
        fsm_output = 9'b111000011;
        state_var_NS = COMP_LOOP_C_450;
      end
      COMP_LOOP_C_450 : begin
        fsm_output = 9'b111000100;
        state_var_NS = COMP_LOOP_C_451;
      end
      COMP_LOOP_C_451 : begin
        fsm_output = 9'b111000101;
        state_var_NS = COMP_LOOP_C_452;
      end
      COMP_LOOP_C_452 : begin
        fsm_output = 9'b111000110;
        state_var_NS = COMP_LOOP_C_453;
      end
      COMP_LOOP_C_453 : begin
        fsm_output = 9'b111000111;
        state_var_NS = COMP_LOOP_C_454;
      end
      COMP_LOOP_C_454 : begin
        fsm_output = 9'b111001000;
        state_var_NS = COMP_LOOP_C_455;
      end
      COMP_LOOP_C_455 : begin
        fsm_output = 9'b111001001;
        state_var_NS = COMP_LOOP_C_456;
      end
      COMP_LOOP_C_456 : begin
        fsm_output = 9'b111001010;
        state_var_NS = COMP_LOOP_C_457;
      end
      COMP_LOOP_C_457 : begin
        fsm_output = 9'b111001011;
        state_var_NS = COMP_LOOP_C_458;
      end
      COMP_LOOP_C_458 : begin
        fsm_output = 9'b111001100;
        state_var_NS = COMP_LOOP_C_459;
      end
      COMP_LOOP_C_459 : begin
        fsm_output = 9'b111001101;
        state_var_NS = COMP_LOOP_C_460;
      end
      COMP_LOOP_C_460 : begin
        fsm_output = 9'b111001110;
        state_var_NS = COMP_LOOP_C_461;
      end
      COMP_LOOP_C_461 : begin
        fsm_output = 9'b111001111;
        state_var_NS = COMP_LOOP_C_462;
      end
      COMP_LOOP_C_462 : begin
        fsm_output = 9'b111010000;
        state_var_NS = COMP_LOOP_C_463;
      end
      COMP_LOOP_C_463 : begin
        fsm_output = 9'b111010001;
        state_var_NS = COMP_LOOP_C_464;
      end
      COMP_LOOP_C_464 : begin
        fsm_output = 9'b111010010;
        state_var_NS = COMP_LOOP_C_465;
      end
      COMP_LOOP_C_465 : begin
        fsm_output = 9'b111010011;
        if ( COMP_LOOP_C_465_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_466;
        end
      end
      COMP_LOOP_C_466 : begin
        fsm_output = 9'b111010100;
        state_var_NS = COMP_LOOP_C_467;
      end
      COMP_LOOP_C_467 : begin
        fsm_output = 9'b111010101;
        state_var_NS = COMP_LOOP_C_468;
      end
      COMP_LOOP_C_468 : begin
        fsm_output = 9'b111010110;
        state_var_NS = COMP_LOOP_C_469;
      end
      COMP_LOOP_C_469 : begin
        fsm_output = 9'b111010111;
        state_var_NS = COMP_LOOP_C_470;
      end
      COMP_LOOP_C_470 : begin
        fsm_output = 9'b111011000;
        state_var_NS = COMP_LOOP_C_471;
      end
      COMP_LOOP_C_471 : begin
        fsm_output = 9'b111011001;
        state_var_NS = COMP_LOOP_C_472;
      end
      COMP_LOOP_C_472 : begin
        fsm_output = 9'b111011010;
        state_var_NS = COMP_LOOP_C_473;
      end
      COMP_LOOP_C_473 : begin
        fsm_output = 9'b111011011;
        state_var_NS = COMP_LOOP_C_474;
      end
      COMP_LOOP_C_474 : begin
        fsm_output = 9'b111011100;
        state_var_NS = COMP_LOOP_C_475;
      end
      COMP_LOOP_C_475 : begin
        fsm_output = 9'b111011101;
        state_var_NS = COMP_LOOP_C_476;
      end
      COMP_LOOP_C_476 : begin
        fsm_output = 9'b111011110;
        state_var_NS = COMP_LOOP_C_477;
      end
      COMP_LOOP_C_477 : begin
        fsm_output = 9'b111011111;
        state_var_NS = COMP_LOOP_C_478;
      end
      COMP_LOOP_C_478 : begin
        fsm_output = 9'b111100000;
        state_var_NS = COMP_LOOP_C_479;
      end
      COMP_LOOP_C_479 : begin
        fsm_output = 9'b111100001;
        state_var_NS = COMP_LOOP_C_480;
      end
      COMP_LOOP_C_480 : begin
        fsm_output = 9'b111100010;
        state_var_NS = COMP_LOOP_C_481;
      end
      COMP_LOOP_C_481 : begin
        fsm_output = 9'b111100011;
        state_var_NS = COMP_LOOP_C_482;
      end
      COMP_LOOP_C_482 : begin
        fsm_output = 9'b111100100;
        state_var_NS = COMP_LOOP_C_483;
      end
      COMP_LOOP_C_483 : begin
        fsm_output = 9'b111100101;
        state_var_NS = COMP_LOOP_C_484;
      end
      COMP_LOOP_C_484 : begin
        fsm_output = 9'b111100110;
        state_var_NS = COMP_LOOP_C_485;
      end
      COMP_LOOP_C_485 : begin
        fsm_output = 9'b111100111;
        state_var_NS = COMP_LOOP_C_486;
      end
      COMP_LOOP_C_486 : begin
        fsm_output = 9'b111101000;
        state_var_NS = COMP_LOOP_C_487;
      end
      COMP_LOOP_C_487 : begin
        fsm_output = 9'b111101001;
        state_var_NS = COMP_LOOP_C_488;
      end
      COMP_LOOP_C_488 : begin
        fsm_output = 9'b111101010;
        state_var_NS = COMP_LOOP_C_489;
      end
      COMP_LOOP_C_489 : begin
        fsm_output = 9'b111101011;
        state_var_NS = COMP_LOOP_C_490;
      end
      COMP_LOOP_C_490 : begin
        fsm_output = 9'b111101100;
        state_var_NS = COMP_LOOP_C_491;
      end
      COMP_LOOP_C_491 : begin
        fsm_output = 9'b111101101;
        state_var_NS = COMP_LOOP_C_492;
      end
      COMP_LOOP_C_492 : begin
        fsm_output = 9'b111101110;
        state_var_NS = COMP_LOOP_C_493;
      end
      COMP_LOOP_C_493 : begin
        fsm_output = 9'b111101111;
        state_var_NS = COMP_LOOP_C_494;
      end
      COMP_LOOP_C_494 : begin
        fsm_output = 9'b111110000;
        state_var_NS = COMP_LOOP_C_495;
      end
      COMP_LOOP_C_495 : begin
        fsm_output = 9'b111110001;
        state_var_NS = COMP_LOOP_C_496;
      end
      COMP_LOOP_C_496 : begin
        fsm_output = 9'b111110010;
        if ( COMP_LOOP_C_496_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_C_0 : begin
        fsm_output = 9'b111110011;
        if ( VEC_LOOP_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      STAGE_LOOP_C_1 : begin
        fsm_output = 9'b111110100;
        if ( STAGE_LOOP_C_1_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = STAGE_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 9'b111110101;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 9'b000000000;
        state_var_NS = STAGE_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_core_wait_dp
// ------------------------------------------------------------------


module inPlaceNTT_DIF_core_wait_dp (
  ensig_cgo_iro, ensig_cgo, COMP_LOOP_1_modulo_cmp_ccs_ccore_en
);
  input ensig_cgo_iro;
  input ensig_cgo;
  output COMP_LOOP_1_modulo_cmp_ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  assign COMP_LOOP_1_modulo_cmp_ccs_ccore_en = ensig_cgo | ensig_cgo_iro;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_core
// ------------------------------------------------------------------


module inPlaceNTT_DIF_core (
  clk, rst, vec_rsc_triosy_0_0_lz, vec_rsc_triosy_0_1_lz, vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz, vec_rsc_triosy_0_4_lz, vec_rsc_triosy_0_5_lz, vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz, vec_rsc_triosy_0_8_lz, vec_rsc_triosy_0_9_lz, vec_rsc_triosy_0_10_lz,
      vec_rsc_triosy_0_11_lz, vec_rsc_triosy_0_12_lz, vec_rsc_triosy_0_13_lz, vec_rsc_triosy_0_14_lz,
      vec_rsc_triosy_0_15_lz, p_rsc_dat, p_rsc_triosy_lz, r_rsc_triosy_lz, twiddle_rsc_triosy_0_0_lz,
      twiddle_rsc_triosy_0_1_lz, twiddle_rsc_triosy_0_2_lz, twiddle_rsc_triosy_0_3_lz,
      twiddle_rsc_triosy_0_4_lz, twiddle_rsc_triosy_0_5_lz, twiddle_rsc_triosy_0_6_lz,
      twiddle_rsc_triosy_0_7_lz, twiddle_rsc_triosy_0_8_lz, twiddle_rsc_triosy_0_9_lz,
      twiddle_rsc_triosy_0_10_lz, twiddle_rsc_triosy_0_11_lz, twiddle_rsc_triosy_0_12_lz,
      twiddle_rsc_triosy_0_13_lz, twiddle_rsc_triosy_0_14_lz, twiddle_rsc_triosy_0_15_lz,
      vec_rsc_0_0_i_q_d, vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_1_i_q_d,
      vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_2_i_q_d, vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_q_d, vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_4_i_q_d,
      vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_5_i_q_d, vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_q_d, vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_7_i_q_d,
      vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_8_i_q_d, vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_9_i_q_d, vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_10_i_q_d,
      vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_11_i_q_d, vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_12_i_q_d, vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_13_i_q_d,
      vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_14_i_q_d, vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_15_i_q_d, vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_0_i_q_d,
      twiddle_rsc_0_0_i_radr_d, twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_1_i_q_d, twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_3_i_q_d, twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_4_i_q_d, twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_5_i_q_d, twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_6_i_q_d, twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_7_i_q_d, twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_8_i_q_d, twiddle_rsc_0_8_i_radr_d, twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_9_i_q_d, twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_10_i_q_d, twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_11_i_q_d, twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_12_i_q_d, twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_13_i_q_d, twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_14_i_q_d, twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_15_i_q_d, twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_0_i_d_d_pff, vec_rsc_0_0_i_radr_d_pff, vec_rsc_0_0_i_wadr_d_pff,
      vec_rsc_0_0_i_we_d_pff, vec_rsc_0_1_i_we_d_pff, vec_rsc_0_2_i_we_d_pff, vec_rsc_0_3_i_we_d_pff,
      vec_rsc_0_4_i_we_d_pff, vec_rsc_0_5_i_we_d_pff, vec_rsc_0_6_i_we_d_pff, vec_rsc_0_7_i_we_d_pff,
      vec_rsc_0_8_i_we_d_pff, vec_rsc_0_9_i_we_d_pff, vec_rsc_0_10_i_we_d_pff, vec_rsc_0_11_i_we_d_pff,
      vec_rsc_0_12_i_we_d_pff, vec_rsc_0_13_i_we_d_pff, vec_rsc_0_14_i_we_d_pff,
      vec_rsc_0_15_i_we_d_pff, twiddle_rsc_0_1_i_radr_d_pff, twiddle_rsc_0_2_i_radr_d_pff,
      twiddle_rsc_0_4_i_radr_d_pff
);
  input clk;
  input rst;
  output vec_rsc_triosy_0_0_lz;
  output vec_rsc_triosy_0_1_lz;
  output vec_rsc_triosy_0_2_lz;
  output vec_rsc_triosy_0_3_lz;
  output vec_rsc_triosy_0_4_lz;
  output vec_rsc_triosy_0_5_lz;
  output vec_rsc_triosy_0_6_lz;
  output vec_rsc_triosy_0_7_lz;
  output vec_rsc_triosy_0_8_lz;
  output vec_rsc_triosy_0_9_lz;
  output vec_rsc_triosy_0_10_lz;
  output vec_rsc_triosy_0_11_lz;
  output vec_rsc_triosy_0_12_lz;
  output vec_rsc_triosy_0_13_lz;
  output vec_rsc_triosy_0_14_lz;
  output vec_rsc_triosy_0_15_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  output r_rsc_triosy_lz;
  output twiddle_rsc_triosy_0_0_lz;
  output twiddle_rsc_triosy_0_1_lz;
  output twiddle_rsc_triosy_0_2_lz;
  output twiddle_rsc_triosy_0_3_lz;
  output twiddle_rsc_triosy_0_4_lz;
  output twiddle_rsc_triosy_0_5_lz;
  output twiddle_rsc_triosy_0_6_lz;
  output twiddle_rsc_triosy_0_7_lz;
  output twiddle_rsc_triosy_0_8_lz;
  output twiddle_rsc_triosy_0_9_lz;
  output twiddle_rsc_triosy_0_10_lz;
  output twiddle_rsc_triosy_0_11_lz;
  output twiddle_rsc_triosy_0_12_lz;
  output twiddle_rsc_triosy_0_13_lz;
  output twiddle_rsc_triosy_0_14_lz;
  output twiddle_rsc_triosy_0_15_lz;
  input [63:0] vec_rsc_0_0_i_q_d;
  output vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_1_i_q_d;
  output vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_2_i_q_d;
  output vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_3_i_q_d;
  output vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_4_i_q_d;
  output vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_5_i_q_d;
  output vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_6_i_q_d;
  output vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_7_i_q_d;
  output vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_8_i_q_d;
  output vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_9_i_q_d;
  output vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_10_i_q_d;
  output vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_11_i_q_d;
  output vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_12_i_q_d;
  output vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_13_i_q_d;
  output vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_14_i_q_d;
  output vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_15_i_q_d;
  output vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_0_i_q_d;
  output [5:0] twiddle_rsc_0_0_i_radr_d;
  output twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_1_i_q_d;
  output twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_2_i_q_d;
  output twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_3_i_q_d;
  output twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_4_i_q_d;
  output twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_5_i_q_d;
  output twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_6_i_q_d;
  output twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_7_i_q_d;
  output twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_8_i_q_d;
  output [5:0] twiddle_rsc_0_8_i_radr_d;
  output twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_9_i_q_d;
  output twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_10_i_q_d;
  output twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_11_i_q_d;
  output twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_12_i_q_d;
  output twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_13_i_q_d;
  output twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_14_i_q_d;
  output twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_15_i_q_d;
  output twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d;
  output [63:0] vec_rsc_0_0_i_d_d_pff;
  output [5:0] vec_rsc_0_0_i_radr_d_pff;
  output [5:0] vec_rsc_0_0_i_wadr_d_pff;
  output vec_rsc_0_0_i_we_d_pff;
  output vec_rsc_0_1_i_we_d_pff;
  output vec_rsc_0_2_i_we_d_pff;
  output vec_rsc_0_3_i_we_d_pff;
  output vec_rsc_0_4_i_we_d_pff;
  output vec_rsc_0_5_i_we_d_pff;
  output vec_rsc_0_6_i_we_d_pff;
  output vec_rsc_0_7_i_we_d_pff;
  output vec_rsc_0_8_i_we_d_pff;
  output vec_rsc_0_9_i_we_d_pff;
  output vec_rsc_0_10_i_we_d_pff;
  output vec_rsc_0_11_i_we_d_pff;
  output vec_rsc_0_12_i_we_d_pff;
  output vec_rsc_0_13_i_we_d_pff;
  output vec_rsc_0_14_i_we_d_pff;
  output vec_rsc_0_15_i_we_d_pff;
  output [5:0] twiddle_rsc_0_1_i_radr_d_pff;
  output [5:0] twiddle_rsc_0_2_i_radr_d_pff;
  output [5:0] twiddle_rsc_0_4_i_radr_d_pff;


  // Interconnect Declarations
  wire [63:0] p_rsci_idat;
  wire [63:0] COMP_LOOP_1_modulo_cmp_return_rsc_z;
  wire COMP_LOOP_1_modulo_cmp_ccs_ccore_en;
  wire [8:0] fsm_output;
  wire or_dcpl_5;
  wire and_dcpl_5;
  wire nor_tmp_10;
  wire or_tmp_29;
  wire nor_tmp_47;
  wire nor_tmp_115;
  wire mux_tmp_439;
  wire mux_tmp_538;
  wire mux_tmp_929;
  wire nand_tmp_13;
  wire and_dcpl_45;
  wire and_dcpl_46;
  wire and_dcpl_47;
  wire and_dcpl_48;
  wire and_dcpl_51;
  wire and_dcpl_53;
  wire and_dcpl_54;
  wire and_dcpl_55;
  wire and_dcpl_57;
  wire and_dcpl_58;
  wire nor_tmp_339;
  wire mux_tmp_1062;
  wire mux_tmp_1065;
  wire mux_tmp_1067;
  wire and_dcpl_60;
  wire and_dcpl_61;
  wire and_dcpl_62;
  wire and_dcpl_63;
  wire and_dcpl_64;
  wire and_dcpl_65;
  wire and_dcpl_66;
  wire and_dcpl_67;
  wire and_dcpl_69;
  wire and_dcpl_70;
  wire and_dcpl_71;
  wire and_dcpl_72;
  wire and_dcpl_74;
  wire and_dcpl_75;
  wire and_dcpl_77;
  wire and_dcpl_79;
  wire and_dcpl_81;
  wire and_dcpl_82;
  wire and_dcpl_83;
  wire and_dcpl_85;
  wire and_dcpl_86;
  wire and_dcpl_87;
  wire and_dcpl_88;
  wire and_dcpl_89;
  wire and_dcpl_91;
  wire and_dcpl_92;
  wire and_dcpl_93;
  wire and_dcpl_95;
  wire and_dcpl_96;
  wire and_dcpl_97;
  wire and_dcpl_99;
  wire and_dcpl_100;
  wire and_dcpl_102;
  wire and_dcpl_103;
  wire and_dcpl_104;
  wire and_dcpl_105;
  wire and_dcpl_107;
  wire and_dcpl_108;
  wire and_dcpl_110;
  wire and_dcpl_111;
  wire and_dcpl_112;
  wire and_dcpl_113;
  wire and_dcpl_115;
  wire and_dcpl_116;
  wire and_dcpl_118;
  wire and_dcpl_119;
  wire and_dcpl_120;
  wire and_dcpl_121;
  wire and_dcpl_123;
  wire and_dcpl_124;
  wire and_dcpl_125;
  wire and_dcpl_127;
  wire and_dcpl_128;
  wire and_dcpl_130;
  wire and_dcpl_131;
  wire and_dcpl_136;
  wire and_dcpl_141;
  wire and_dcpl_146;
  wire and_dcpl_151;
  wire and_dcpl_156;
  wire and_dcpl_161;
  wire and_dcpl_166;
  wire not_tmp_395;
  wire not_tmp_399;
  wire and_dcpl_171;
  wire and_dcpl_175;
  wire and_dcpl_180;
  wire and_dcpl_181;
  wire and_dcpl_182;
  wire and_dcpl_183;
  wire and_dcpl_184;
  wire and_dcpl_186;
  wire or_tmp_2077;
  wire and_dcpl_188;
  wire and_dcpl_189;
  wire and_dcpl_190;
  wire and_dcpl_191;
  wire and_dcpl_192;
  wire and_dcpl_193;
  wire and_dcpl_195;
  wire and_dcpl_196;
  wire and_dcpl_197;
  wire and_dcpl_198;
  wire and_dcpl_202;
  wire and_dcpl_207;
  wire mux_tmp_2224;
  wire mux_tmp_2225;
  wire mux_tmp_2229;
  wire or_tmp_2258;
  wire mux_tmp_2237;
  wire not_tmp_676;
  wire nor_tmp_480;
  wire mux_tmp_2238;
  wire or_tmp_2266;
  wire mux_tmp_2245;
  wire mux_tmp_2246;
  wire mux_tmp_2249;
  wire and_dcpl_220;
  wire and_dcpl_222;
  wire and_dcpl_223;
  wire and_dcpl_225;
  wire and_dcpl_226;
  wire and_dcpl_227;
  wire and_dcpl_228;
  wire and_dcpl_229;
  wire and_dcpl_230;
  wire and_dcpl_231;
  wire and_dcpl_232;
  wire and_dcpl_233;
  wire and_dcpl_234;
  wire and_dcpl_235;
  wire and_dcpl_236;
  wire or_tmp_2274;
  wire mux_tmp_2256;
  wire mux_tmp_2257;
  wire mux_tmp_2258;
  wire mux_tmp_2259;
  wire or_tmp_2277;
  wire or_tmp_2279;
  wire mux_tmp_2264;
  wire or_dcpl_182;
  wire or_dcpl_183;
  wire or_dcpl_184;
  wire mux_tmp_2282;
  wire nor_tmp_489;
  wire mux_tmp_2288;
  wire mux_tmp_2291;
  wire mux_tmp_2292;
  wire not_tmp_703;
  wire or_tmp_2300;
  wire or_dcpl_190;
  wire and_dcpl_248;
  wire and_dcpl_252;
  wire and_dcpl_255;
  wire nor_tmp_499;
  wire mux_tmp_2311;
  wire and_dcpl_258;
  wire mux_tmp_2318;
  wire and_dcpl_262;
  wire nor_tmp_507;
  wire and_tmp_28;
  wire mux_tmp_2325;
  wire mux_tmp_2328;
  wire nor_tmp_509;
  wire and_dcpl_266;
  wire not_tmp_727;
  wire and_dcpl_270;
  wire nor_tmp_515;
  wire mux_tmp_2344;
  wire mux_tmp_2347;
  wire mux_tmp_2348;
  wire mux_tmp_2351;
  wire and_dcpl_271;
  wire mux_tmp_2357;
  wire mux_tmp_2365;
  wire mux_tmp_2369;
  wire nor_tmp_528;
  wire nor_tmp_530;
  wire mux_tmp_2384;
  wire nor_tmp_537;
  wire mux_tmp_2392;
  wire mux_tmp_2395;
  wire nor_tmp_538;
  wire mux_tmp_2401;
  wire nor_tmp_544;
  wire mux_tmp_2410;
  wire nor_tmp_547;
  wire nor_tmp_548;
  wire not_tmp_762;
  wire or_dcpl_207;
  wire and_dcpl_277;
  wire or_tmp_2358;
  wire mux_tmp_2447;
  wire nand_tmp_100;
  wire mux_tmp_2450;
  wire or_tmp_2362;
  wire and_dcpl_286;
  wire or_tmp_2384;
  reg COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm;
  wire [7:0] COMP_LOOP_acc_13_psp_sva_1;
  wire [8:0] nl_COMP_LOOP_acc_13_psp_sva_1;
  wire [9:0] COMP_LOOP_acc_1_cse_4_sva_1;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_4_sva_1;
  reg [9:0] VEC_LOOP_j_10_0_sva_9_0;
  reg COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm;
  reg COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm;
  reg COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm;
  reg COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm;
  reg COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm;
  reg [9:0] COMP_LOOP_10_tmp_mul_idiv_sva;
  reg COMP_LOOP_tmp_nor_itm;
  reg COMP_LOOP_tmp_nor_13_itm;
  reg COMP_LOOP_tmp_nor_1_itm;
  reg COMP_LOOP_tmp_nor_14_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm;
  reg COMP_LOOP_tmp_nor_3_itm;
  reg COMP_LOOP_tmp_nor_16_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm;
  reg [6:0] COMP_LOOP_9_tmp_lshift_itm;
  reg COMP_LOOP_tmp_nor_6_itm;
  reg COMP_LOOP_tmp_nor_19_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_itm;
  reg [8:0] COMP_LOOP_11_tmp_mul_idiv_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_2_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_6_sva;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_6_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_10_sva;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_10_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_14_sva;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_14_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_4_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_8_sva;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_8_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_12_sva;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_12_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_sva;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_2_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_6_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_10_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_14_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_4_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_8_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_12_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_1_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_5_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_9_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_13_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_3_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_7_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_11_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_15_sva;
  reg [8:0] COMP_LOOP_acc_11_psp_sva;
  wire [9:0] nl_COMP_LOOP_acc_11_psp_sva;
  reg [8:0] COMP_LOOP_acc_14_psp_sva;
  wire [9:0] nl_COMP_LOOP_acc_14_psp_sva;
  reg [8:0] COMP_LOOP_acc_17_psp_sva;
  wire [9:0] nl_COMP_LOOP_acc_17_psp_sva;
  reg [8:0] COMP_LOOP_acc_20_psp_sva;
  wire [9:0] nl_COMP_LOOP_acc_20_psp_sva;
  reg [7:0] COMP_LOOP_acc_13_psp_sva;
  reg [6:0] COMP_LOOP_acc_16_psp_sva;
  wire [7:0] nl_COMP_LOOP_acc_16_psp_sva;
  reg [7:0] COMP_LOOP_acc_19_psp_sva;
  wire [8:0] nl_COMP_LOOP_acc_19_psp_sva;
  reg [7:0] COMP_LOOP_13_tmp_mul_idiv_sva;
  reg [7:0] COMP_LOOP_5_tmp_mul_idiv_sva;
  reg [10:0] STAGE_LOOP_lshift_psp_sva;
  reg [5:0] COMP_LOOP_k_10_4_sva_5_0;
  wire [9:0] COMP_LOOP_acc_1_cse_2_sva_1;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_2_sva_1;
  wire nor_1796_tmp;
  wire nor_1798_tmp;
  wire and_342_tmp;
  wire and_341_tmp;
  wire and_332_tmp;
  wire and_314_m1c;
  reg [5:0] reg_COMP_LOOP_k_10_4_ftd;
  wire mux_1128_cse;
  wire nand_271_cse;
  wire nand_272_cse;
  wire mux_1191_cse;
  wire nor_346_cse;
  wire nor_351_cse;
  wire nor_1528_cse;
  wire nand_265_cse;
  wire mux_1378_cse;
  wire nand_219_cse;
  wire mux_1628_cse;
  wire nand_211_cse;
  wire nand_212_cse;
  wire mux_1691_cse;
  wire and_523_cse;
  wire mux_1878_cse;
  wire nand_122_cse;
  wire nand_121_cse;
  reg reg_vec_rsc_triosy_0_15_obj_ld_cse;
  reg reg_ensig_cgo_cse;
  wire and_421_cse;
  wire and_831_cse;
  wire and_407_cse;
  wire and_733_cse;
  wire or_432_cse;
  wire and_674_cse;
  wire and_675_cse;
  wire nand_301_cse;
  wire COMP_LOOP_tmp_or_2_cse;
  wire COMP_LOOP_tmp_or_1_cse;
  wire COMP_LOOP_tmp_or_21_cse;
  wire COMP_LOOP_tmp_or_29_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_nor_14_cse;
  wire and_570_cse;
  wire or_2729_cse;
  wire and_712_cse;
  wire nor_1792_cse;
  wire nor_1630_cse;
  wire nor_1624_cse;
  wire or_36_cse;
  wire mux_228_cse;
  wire nor_572_cse;
  wire or_2732_cse;
  wire or_455_cse;
  wire or_454_cse;
  wire mux_464_cse;
  wire or_610_cse;
  wire mux_1116_cse;
  wire nor_1523_cse;
  wire nor_1526_cse;
  wire nor_1527_cse;
  wire mux_1241_cse;
  wire nor_1402_cse;
  wire nor_1405_cse;
  wire nor_1406_cse;
  wire mux_1366_cse;
  wire nor_1286_cse;
  wire nor_1289_cse;
  wire nor_1290_cse;
  wire nand_268_cse;
  wire mux_1491_cse;
  wire nand_261_cse;
  wire nand_226_cse;
  wire and_529_cse;
  wire nor_1173_cse;
  wire nor_1174_cse;
  wire mux_1616_cse;
  wire nand_222_cse;
  wire nand_223_cse;
  wire nor_1056_cse;
  wire nor_1059_cse;
  wire nor_1060_cse;
  wire mux_1741_cse;
  wire and_506_cse;
  wire nor_944_cse;
  wire nor_945_cse;
  wire mux_1866_cse;
  wire nand_184_cse;
  wire nand_185_cse;
  wire and_490_cse;
  wire nor_837_cse;
  wire nor_838_cse;
  wire nand_170_cse;
  wire mux_1991_cse;
  wire nand_157_cse;
  wire and_450_cse;
  wire and_836_cse;
  wire and_453_cse;
  wire nor_1767_cse;
  wire or_2589_cse;
  wire or_2697_cse;
  wire or_2487_cse;
  wire or_2486_cse;
  wire or_2612_cse;
  wire or_2635_cse;
  wire nor_1554_cse;
  wire nor_1435_cse;
  wire nor_1317_cse;
  wire nor_1200_cse;
  wire mux_1441_cse;
  wire nor_1086_cse;
  wire nor_970_cse;
  wire nor_860_cse;
  wire nor_761_cse;
  wire mux_1941_cse;
  wire mux_955_cse;
  wire and_728_cse;
  wire mux_559_cse;
  wire or_2626_cse;
  wire or_2621_cse;
  wire and_655_cse;
  wire or_611_cse;
  wire mux_952_cse;
  wire mux_949_cse;
  wire mux_965_cse;
  wire mux_2255_rmff;
  reg [63:0] COMP_LOOP_10_acc_8_itm;
  reg [63:0] p_sva;
  reg [5:0] COMP_LOOP_acc_psp_sva;
  wire [6:0] nl_COMP_LOOP_acc_psp_sva;
  wire mux_2303_itm;
  wire mux_2383_itm;
  wire mux_2398_itm;
  wire mux_2410_itm;
  wire mux_2424_itm;
  wire mux_2435_itm;
  wire mux_2442_itm;
  wire mux_2444_itm;
  wire mux_2449_itm;
  wire [5:0] COMP_LOOP_1_tmp_lshift_itm;
  wire [10:0] z_out;
  wire [9:0] z_out_1;
  wire and_dcpl_356;
  wire [10:0] z_out_2;
  wire and_dcpl_360;
  wire and_dcpl_362;
  wire and_dcpl_366;
  wire and_dcpl_367;
  wire and_dcpl_370;
  wire and_dcpl_373;
  wire and_dcpl_374;
  wire and_dcpl_376;
  wire and_dcpl_377;
  wire and_dcpl_378;
  wire and_dcpl_380;
  wire and_dcpl_383;
  wire and_dcpl_384;
  wire and_dcpl_385;
  wire and_dcpl_386;
  wire and_dcpl_387;
  wire and_dcpl_389;
  wire and_dcpl_390;
  wire and_dcpl_391;
  wire and_dcpl_394;
  wire and_dcpl_395;
  wire and_dcpl_396;
  wire and_dcpl_397;
  wire and_dcpl_399;
  wire and_dcpl_400;
  wire and_dcpl_401;
  wire and_dcpl_404;
  wire and_dcpl_405;
  wire and_dcpl_406;
  wire and_dcpl_409;
  wire and_dcpl_410;
  wire and_dcpl_411;
  wire and_dcpl_412;
  wire and_dcpl_413;
  wire and_dcpl_414;
  wire and_dcpl_415;
  wire and_dcpl_416;
  wire and_dcpl_417;
  wire and_dcpl_418;
  wire and_dcpl_419;
  wire and_dcpl_420;
  wire and_dcpl_421;
  wire and_dcpl_422;
  wire and_dcpl_425;
  wire and_dcpl_426;
  wire and_dcpl_427;
  wire and_dcpl_428;
  wire and_dcpl_429;
  wire and_dcpl_430;
  wire and_dcpl_431;
  wire [63:0] z_out_3;
  wire [127:0] nl_z_out_3;
  wire and_dcpl_447;
  wire [3:0] z_out_4;
  wire [4:0] nl_z_out_4;
  wire and_dcpl_465;
  wire and_dcpl_467;
  wire and_dcpl_475;
  wire and_dcpl_477;
  wire and_dcpl_480;
  wire and_dcpl_482;
  wire and_dcpl_484;
  wire and_dcpl_486;
  wire and_dcpl_495;
  wire and_dcpl_571;
  wire and_dcpl_577;
  wire and_dcpl_589;
  wire [63:0] z_out_7;
  reg [3:0] STAGE_LOOP_i_3_0_sva;
  reg [3:0] COMP_LOOP_1_tmp_acc_cse_sva;
  reg [9:0] COMP_LOOP_2_tmp_lshift_ncse_sva;
  reg [63:0] tmp_33_sva_1;
  reg [63:0] tmp_33_sva_2;
  reg [63:0] tmp_33_sva_3;
  reg [63:0] tmp_33_sva_4;
  reg [63:0] tmp_33_sva_5;
  reg [63:0] tmp_33_sva_6;
  reg [63:0] tmp_33_sva_7;
  reg [63:0] tmp_33_sva_8;
  reg [63:0] tmp_33_sva_9;
  reg [63:0] tmp_33_sva_10;
  reg [63:0] tmp_33_sva_11;
  reg [63:0] tmp_33_sva_12;
  reg [63:0] tmp_33_sva_13;
  reg [63:0] tmp_33_sva_14;
  reg [63:0] tmp_33_sva_15;
  reg [8:0] COMP_LOOP_3_tmp_lshift_ncse_sva;
  reg [63:0] tmp_36_sva_1;
  reg [63:0] tmp_36_sva_2;
  reg COMP_LOOP_COMP_LOOP_nor_itm;
  reg COMP_LOOP_COMP_LOOP_and_6_itm;
  reg COMP_LOOP_COMP_LOOP_and_10_itm;
  reg COMP_LOOP_COMP_LOOP_and_12_itm;
  reg COMP_LOOP_COMP_LOOP_and_13_itm;
  reg COMP_LOOP_COMP_LOOP_and_14_itm;
  reg COMP_LOOP_COMP_LOOP_and_62_itm;
  reg COMP_LOOP_COMP_LOOP_and_64_itm;
  reg COMP_LOOP_COMP_LOOP_and_65_itm;
  reg COMP_LOOP_COMP_LOOP_and_66_itm;
  reg COMP_LOOP_COMP_LOOP_and_68_itm;
  reg COMP_LOOP_COMP_LOOP_and_69_itm;
  reg COMP_LOOP_COMP_LOOP_and_70_itm;
  reg COMP_LOOP_COMP_LOOP_and_72_itm;
  reg COMP_LOOP_COMP_LOOP_nor_5_itm;
  reg COMP_LOOP_nor_51_itm;
  reg COMP_LOOP_nor_52_itm;
  reg COMP_LOOP_COMP_LOOP_and_77_itm;
  reg COMP_LOOP_nor_54_itm;
  reg COMP_LOOP_COMP_LOOP_and_79_itm;
  reg COMP_LOOP_COMP_LOOP_and_80_itm;
  reg COMP_LOOP_COMP_LOOP_and_81_itm;
  reg COMP_LOOP_nor_57_itm;
  reg COMP_LOOP_COMP_LOOP_and_83_itm;
  reg COMP_LOOP_COMP_LOOP_and_84_itm;
  reg COMP_LOOP_COMP_LOOP_and_85_itm;
  reg COMP_LOOP_COMP_LOOP_and_86_itm;
  reg COMP_LOOP_COMP_LOOP_and_87_itm;
  reg COMP_LOOP_COMP_LOOP_and_88_itm;
  reg COMP_LOOP_COMP_LOOP_and_89_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_nor_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_itm;
  reg COMP_LOOP_COMP_LOOP_nor_9_itm;
  reg COMP_LOOP_nor_91_itm;
  reg COMP_LOOP_nor_92_itm;
  reg COMP_LOOP_COMP_LOOP_and_137_itm;
  reg COMP_LOOP_nor_94_itm;
  reg COMP_LOOP_COMP_LOOP_and_139_itm;
  reg COMP_LOOP_COMP_LOOP_and_140_itm;
  reg COMP_LOOP_COMP_LOOP_and_141_itm;
  reg COMP_LOOP_nor_97_itm;
  reg COMP_LOOP_COMP_LOOP_and_143_itm;
  reg COMP_LOOP_COMP_LOOP_and_144_itm;
  reg COMP_LOOP_COMP_LOOP_and_145_itm;
  reg COMP_LOOP_COMP_LOOP_and_146_itm;
  reg COMP_LOOP_COMP_LOOP_and_147_itm;
  reg COMP_LOOP_COMP_LOOP_and_148_itm;
  reg COMP_LOOP_COMP_LOOP_and_149_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_1_itm;
  reg COMP_LOOP_COMP_LOOP_and_185_itm;
  reg COMP_LOOP_COMP_LOOP_nor_13_itm;
  reg COMP_LOOP_nor_131_itm;
  reg COMP_LOOP_nor_132_itm;
  reg COMP_LOOP_COMP_LOOP_and_197_itm;
  reg COMP_LOOP_nor_134_itm;
  reg COMP_LOOP_COMP_LOOP_and_199_itm;
  reg COMP_LOOP_COMP_LOOP_and_200_itm;
  reg COMP_LOOP_COMP_LOOP_and_201_itm;
  reg COMP_LOOP_nor_137_itm;
  reg COMP_LOOP_COMP_LOOP_and_203_itm;
  reg COMP_LOOP_COMP_LOOP_and_204_itm;
  reg COMP_LOOP_COMP_LOOP_and_205_itm;
  reg COMP_LOOP_COMP_LOOP_and_206_itm;
  reg COMP_LOOP_COMP_LOOP_and_207_itm;
  reg COMP_LOOP_COMP_LOOP_and_208_itm;
  reg COMP_LOOP_COMP_LOOP_and_209_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_2_itm;
  reg COMP_LOOP_COMP_LOOP_and_244_itm;
  reg COMP_LOOP_COMP_LOOP_nor_17_itm;
  reg COMP_LOOP_nor_171_itm;
  reg COMP_LOOP_nor_172_itm;
  reg COMP_LOOP_COMP_LOOP_and_257_itm;
  reg COMP_LOOP_nor_174_itm;
  reg COMP_LOOP_COMP_LOOP_and_259_itm;
  reg COMP_LOOP_COMP_LOOP_and_260_itm;
  reg COMP_LOOP_COMP_LOOP_and_261_itm;
  reg COMP_LOOP_nor_177_itm;
  reg COMP_LOOP_COMP_LOOP_and_263_itm;
  reg COMP_LOOP_COMP_LOOP_and_264_itm;
  reg COMP_LOOP_COMP_LOOP_and_265_itm;
  reg COMP_LOOP_COMP_LOOP_and_266_itm;
  reg COMP_LOOP_COMP_LOOP_and_267_itm;
  reg COMP_LOOP_COMP_LOOP_and_268_itm;
  reg COMP_LOOP_COMP_LOOP_and_269_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_3_itm;
  reg COMP_LOOP_COMP_LOOP_nor_21_itm;
  reg COMP_LOOP_nor_211_itm;
  reg COMP_LOOP_nor_212_itm;
  reg COMP_LOOP_COMP_LOOP_and_317_itm;
  reg COMP_LOOP_nor_214_itm;
  reg COMP_LOOP_COMP_LOOP_and_319_itm;
  reg COMP_LOOP_COMP_LOOP_and_320_itm;
  reg COMP_LOOP_COMP_LOOP_and_321_itm;
  reg COMP_LOOP_nor_217_itm;
  reg COMP_LOOP_COMP_LOOP_and_323_itm;
  reg COMP_LOOP_COMP_LOOP_and_324_itm;
  reg COMP_LOOP_COMP_LOOP_and_325_itm;
  reg COMP_LOOP_COMP_LOOP_and_326_itm;
  reg COMP_LOOP_COMP_LOOP_and_327_itm;
  reg COMP_LOOP_COMP_LOOP_and_328_itm;
  reg COMP_LOOP_COMP_LOOP_and_329_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_4_itm;
  reg COMP_LOOP_COMP_LOOP_nor_25_itm;
  reg COMP_LOOP_nor_251_itm;
  reg COMP_LOOP_nor_252_itm;
  reg COMP_LOOP_COMP_LOOP_and_377_itm;
  reg COMP_LOOP_nor_254_itm;
  reg COMP_LOOP_COMP_LOOP_and_379_itm;
  reg COMP_LOOP_COMP_LOOP_and_380_itm;
  reg COMP_LOOP_COMP_LOOP_and_381_itm;
  reg COMP_LOOP_nor_257_itm;
  reg COMP_LOOP_COMP_LOOP_and_383_itm;
  reg COMP_LOOP_COMP_LOOP_and_384_itm;
  reg COMP_LOOP_COMP_LOOP_and_385_itm;
  reg COMP_LOOP_COMP_LOOP_and_386_itm;
  reg COMP_LOOP_COMP_LOOP_and_387_itm;
  reg COMP_LOOP_COMP_LOOP_and_388_itm;
  reg COMP_LOOP_COMP_LOOP_and_389_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_5_itm;
  reg COMP_LOOP_COMP_LOOP_nor_29_itm;
  reg COMP_LOOP_nor_291_itm;
  reg COMP_LOOP_nor_292_itm;
  reg COMP_LOOP_COMP_LOOP_and_437_itm;
  reg COMP_LOOP_nor_294_itm;
  reg COMP_LOOP_COMP_LOOP_and_439_itm;
  reg COMP_LOOP_COMP_LOOP_and_440_itm;
  reg COMP_LOOP_COMP_LOOP_and_441_itm;
  reg COMP_LOOP_nor_297_itm;
  reg COMP_LOOP_COMP_LOOP_and_443_itm;
  reg COMP_LOOP_COMP_LOOP_and_444_itm;
  reg COMP_LOOP_COMP_LOOP_and_445_itm;
  reg COMP_LOOP_COMP_LOOP_and_446_itm;
  reg COMP_LOOP_COMP_LOOP_and_447_itm;
  reg COMP_LOOP_COMP_LOOP_and_448_itm;
  reg COMP_LOOP_COMP_LOOP_and_449_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_6_itm;
  reg COMP_LOOP_COMP_LOOP_nor_33_itm;
  reg COMP_LOOP_nor_331_itm;
  reg COMP_LOOP_nor_332_itm;
  reg COMP_LOOP_COMP_LOOP_and_497_itm;
  reg COMP_LOOP_nor_334_itm;
  reg COMP_LOOP_COMP_LOOP_and_499_itm;
  reg COMP_LOOP_COMP_LOOP_and_500_itm;
  reg COMP_LOOP_COMP_LOOP_and_501_itm;
  reg COMP_LOOP_nor_337_itm;
  reg COMP_LOOP_COMP_LOOP_and_503_itm;
  reg COMP_LOOP_COMP_LOOP_and_504_itm;
  reg COMP_LOOP_COMP_LOOP_and_505_itm;
  reg COMP_LOOP_COMP_LOOP_and_506_itm;
  reg COMP_LOOP_COMP_LOOP_and_507_itm;
  reg COMP_LOOP_COMP_LOOP_and_508_itm;
  reg COMP_LOOP_COMP_LOOP_and_509_itm;
  reg [63:0] COMP_LOOP_tmp_mux_itm;
  reg COMP_LOOP_COMP_LOOP_nor_37_itm;
  reg COMP_LOOP_nor_371_itm;
  reg COMP_LOOP_nor_372_itm;
  reg COMP_LOOP_COMP_LOOP_and_557_itm;
  reg COMP_LOOP_nor_374_itm;
  reg COMP_LOOP_COMP_LOOP_and_559_itm;
  reg COMP_LOOP_COMP_LOOP_and_560_itm;
  reg COMP_LOOP_COMP_LOOP_and_561_itm;
  reg COMP_LOOP_nor_377_itm;
  reg COMP_LOOP_COMP_LOOP_and_563_itm;
  reg COMP_LOOP_COMP_LOOP_and_564_itm;
  reg COMP_LOOP_COMP_LOOP_and_565_itm;
  reg COMP_LOOP_COMP_LOOP_and_566_itm;
  reg COMP_LOOP_COMP_LOOP_and_567_itm;
  reg COMP_LOOP_COMP_LOOP_and_568_itm;
  reg COMP_LOOP_COMP_LOOP_and_569_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_7_itm;
  reg COMP_LOOP_COMP_LOOP_nor_41_itm;
  reg COMP_LOOP_nor_411_itm;
  reg COMP_LOOP_nor_412_itm;
  reg COMP_LOOP_COMP_LOOP_and_617_itm;
  reg COMP_LOOP_nor_414_itm;
  reg COMP_LOOP_COMP_LOOP_and_619_itm;
  reg COMP_LOOP_COMP_LOOP_and_620_itm;
  reg COMP_LOOP_COMP_LOOP_and_621_itm;
  reg COMP_LOOP_nor_417_itm;
  reg COMP_LOOP_COMP_LOOP_and_623_itm;
  reg COMP_LOOP_COMP_LOOP_and_624_itm;
  reg COMP_LOOP_COMP_LOOP_and_625_itm;
  reg COMP_LOOP_COMP_LOOP_and_626_itm;
  reg COMP_LOOP_COMP_LOOP_and_627_itm;
  reg COMP_LOOP_COMP_LOOP_and_628_itm;
  reg COMP_LOOP_COMP_LOOP_and_629_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_8_itm;
  reg COMP_LOOP_COMP_LOOP_nor_45_itm;
  reg COMP_LOOP_nor_451_itm;
  reg COMP_LOOP_nor_452_itm;
  reg COMP_LOOP_COMP_LOOP_and_677_itm;
  reg COMP_LOOP_nor_454_itm;
  reg COMP_LOOP_COMP_LOOP_and_679_itm;
  reg COMP_LOOP_COMP_LOOP_and_680_itm;
  reg COMP_LOOP_COMP_LOOP_and_681_itm;
  reg COMP_LOOP_nor_457_itm;
  reg COMP_LOOP_COMP_LOOP_and_683_itm;
  reg COMP_LOOP_COMP_LOOP_and_684_itm;
  reg COMP_LOOP_COMP_LOOP_and_685_itm;
  reg COMP_LOOP_COMP_LOOP_and_686_itm;
  reg COMP_LOOP_COMP_LOOP_and_687_itm;
  reg COMP_LOOP_COMP_LOOP_and_688_itm;
  reg COMP_LOOP_COMP_LOOP_and_689_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_9_itm;
  reg COMP_LOOP_COMP_LOOP_nor_49_itm;
  reg COMP_LOOP_nor_491_itm;
  reg COMP_LOOP_nor_492_itm;
  reg COMP_LOOP_COMP_LOOP_and_737_itm;
  reg COMP_LOOP_nor_494_itm;
  reg COMP_LOOP_COMP_LOOP_and_739_itm;
  reg COMP_LOOP_COMP_LOOP_and_740_itm;
  reg COMP_LOOP_COMP_LOOP_and_741_itm;
  reg COMP_LOOP_nor_497_itm;
  reg COMP_LOOP_COMP_LOOP_and_743_itm;
  reg COMP_LOOP_COMP_LOOP_and_744_itm;
  reg COMP_LOOP_COMP_LOOP_and_745_itm;
  reg COMP_LOOP_COMP_LOOP_and_746_itm;
  reg COMP_LOOP_COMP_LOOP_and_747_itm;
  reg COMP_LOOP_COMP_LOOP_and_748_itm;
  reg COMP_LOOP_COMP_LOOP_and_749_itm;
  reg COMP_LOOP_COMP_LOOP_nor_53_itm;
  reg COMP_LOOP_nor_531_itm;
  reg COMP_LOOP_nor_532_itm;
  reg COMP_LOOP_COMP_LOOP_and_797_itm;
  reg COMP_LOOP_nor_534_itm;
  reg COMP_LOOP_COMP_LOOP_and_799_itm;
  reg COMP_LOOP_COMP_LOOP_and_800_itm;
  reg COMP_LOOP_COMP_LOOP_and_801_itm;
  reg COMP_LOOP_nor_537_itm;
  reg COMP_LOOP_COMP_LOOP_and_803_itm;
  reg COMP_LOOP_COMP_LOOP_and_804_itm;
  reg COMP_LOOP_COMP_LOOP_and_805_itm;
  reg COMP_LOOP_COMP_LOOP_and_806_itm;
  reg COMP_LOOP_COMP_LOOP_and_807_itm;
  reg COMP_LOOP_COMP_LOOP_and_808_itm;
  reg COMP_LOOP_COMP_LOOP_and_809_itm;
  reg COMP_LOOP_COMP_LOOP_nor_57_itm;
  reg COMP_LOOP_nor_571_itm;
  reg COMP_LOOP_nor_572_itm;
  reg COMP_LOOP_COMP_LOOP_and_857_itm;
  reg COMP_LOOP_nor_574_itm;
  reg COMP_LOOP_COMP_LOOP_and_859_itm;
  reg COMP_LOOP_COMP_LOOP_and_860_itm;
  reg COMP_LOOP_COMP_LOOP_and_861_itm;
  reg COMP_LOOP_nor_577_itm;
  reg COMP_LOOP_COMP_LOOP_and_863_itm;
  reg COMP_LOOP_COMP_LOOP_and_864_itm;
  reg COMP_LOOP_COMP_LOOP_and_865_itm;
  reg COMP_LOOP_COMP_LOOP_and_866_itm;
  reg COMP_LOOP_COMP_LOOP_and_867_itm;
  reg COMP_LOOP_COMP_LOOP_and_868_itm;
  reg COMP_LOOP_COMP_LOOP_and_869_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_nor_12_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_12_itm;
  reg COMP_LOOP_COMP_LOOP_nor_61_itm;
  reg COMP_LOOP_nor_611_itm;
  reg COMP_LOOP_nor_612_itm;
  reg COMP_LOOP_COMP_LOOP_and_917_itm;
  reg COMP_LOOP_nor_614_itm;
  reg COMP_LOOP_COMP_LOOP_and_919_itm;
  reg COMP_LOOP_COMP_LOOP_and_920_itm;
  reg COMP_LOOP_COMP_LOOP_and_921_itm;
  reg COMP_LOOP_nor_617_itm;
  reg COMP_LOOP_COMP_LOOP_and_923_itm;
  reg COMP_LOOP_COMP_LOOP_and_924_itm;
  reg COMP_LOOP_COMP_LOOP_and_925_itm;
  reg COMP_LOOP_COMP_LOOP_and_926_itm;
  reg COMP_LOOP_COMP_LOOP_and_927_itm;
  reg COMP_LOOP_COMP_LOOP_and_928_itm;
  reg COMP_LOOP_COMP_LOOP_and_929_itm;
  wire STAGE_LOOP_i_3_0_sva_mx0c1;
  wire VEC_LOOP_j_10_0_sva_9_0_mx0c0;
  wire [6:0] COMP_LOOP_k_10_4_sva_2;
  wire [7:0] nl_COMP_LOOP_k_10_4_sva_2;
  wire [63:0] COMP_LOOP_tmp_mux1h_4_itm_mx0w3;
  wire [63:0] tmp_33_sva_13_mx0w1;
  wire COMP_LOOP_10_acc_8_itm_mx0c2;
  wire COMP_LOOP_10_acc_8_itm_mx0c3;
  wire COMP_LOOP_10_acc_8_itm_mx0c6;
  wire COMP_LOOP_10_acc_8_itm_mx0c9;
  wire COMP_LOOP_10_acc_8_itm_mx0c12;
  wire COMP_LOOP_10_acc_8_itm_mx0c15;
  wire COMP_LOOP_10_acc_8_itm_mx0c18;
  wire COMP_LOOP_10_acc_8_itm_mx0c21;
  wire COMP_LOOP_10_acc_8_itm_mx0c24;
  wire COMP_LOOP_10_acc_8_itm_mx0c27;
  wire COMP_LOOP_10_acc_8_itm_mx0c30;
  wire COMP_LOOP_10_acc_8_itm_mx0c33;
  wire COMP_LOOP_10_acc_8_itm_mx0c36;
  wire COMP_LOOP_10_acc_8_itm_mx0c39;
  wire COMP_LOOP_10_acc_8_itm_mx0c42;
  wire COMP_LOOP_10_acc_8_itm_mx0c47;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_155;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_157;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_159;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_161;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_167;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_nor_16_rgt;
  wire COMP_LOOP_tmp_and_14_rgt;
  wire COMP_LOOP_tmp_and_15_rgt;
  wire COMP_LOOP_tmp_and_16_rgt;
  wire COMP_LOOP_or_17_ssc;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_cse;
  wire COMP_LOOP_or_27_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_17_cse;
  wire COMP_LOOP_tmp_nor_cse;
  wire COMP_LOOP_tmp_nor_1_cse;
  wire COMP_LOOP_or_23_cse;
  wire COMP_LOOP_tmp_nor_3_cse;
  wire COMP_LOOP_tmp_nor_6_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_nor_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_19_cse;
  wire COMP_LOOP_or_31_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_20_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_21_cse;
  wire nor_724_cse;
  wire COMP_LOOP_tmp_or_19_cse;
  wire nor_712_cse;
  wire nor_704_cse;
  wire mux_2131_cse;
  wire nor_691_cse;
  wire nor_682_cse;
  wire nor_670_cse;
  wire nor_662_cse;
  wire COMP_LOOP_tmp_or_46_cse;
  wire nor_647_cse;
  wire nor_639_cse;
  wire nor_627_cse;
  wire nor_619_cse;
  wire mux_2208_cse;
  wire nor_606_cse;
  wire nor_597_cse;
  wire nor_589_cse;
  wire and_427_cse;
  wire mux_2465_cse;
  wire mux_2169_cse;
  wire and_1025_cse;
  wire and_1028_cse;
  wire and_1044_cse;
  wire and_1046_cse;
  wire and_1051_cse;
  wire and_1052_cse;
  wire and_1055_cse;
  wire and_1056_cse;
  wire and_1060_cse;
  wire and_1061_cse;
  wire and_1064_cse;
  wire and_1037_cse;
  wire and_1040_cse;
  wire or_tmp_2410;
  wire or_2259_cse_1;
  wire and_1189_cse;
  wire and_1191_cse;
  wire and_1190_cse;
  wire nand_324_cse;
  wire COMP_LOOP_nor_itm;
  wire COMP_LOOP_or_40_itm;
  wire COMP_LOOP_nor_621_itm;
  wire COMP_LOOP_or_41_itm;
  wire COMP_LOOP_or_43_itm;
  wire COMP_LOOP_nor_622_itm;
  wire COMP_LOOP_or_47_itm;
  wire COMP_LOOP_or_52_itm;
  wire COMP_LOOP_or_54_itm;
  wire COMP_LOOP_or_18_itm;
  wire [9:0] COMP_LOOP_1_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_2_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_3_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_4_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_5_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_6_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_7_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_8_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_9_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_10_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_11_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_12_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_13_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_14_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_15_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_16_acc_10_itm_10_1_1;
  wire STAGE_LOOP_acc_itm_4_1;
  wire [63:0] COMP_LOOP_mux_361_cse;

  wire[0:0] nor_1871_nl;
  wire[0:0] and_1183_nl;
  wire[0:0] nor_1589_nl;
  wire[0:0] nor_1590_nl;
  wire[0:0] mux_1190_nl;
  wire[0:0] nor_1529_nl;
  wire[0:0] nor_1530_nl;
  wire[0:0] nor_1352_nl;
  wire[0:0] nor_1353_nl;
  wire[0:0] nor_1291_nl;
  wire[0:0] mux_1440_nl;
  wire[0:0] nor_1293_nl;
  wire[0:0] nor_1121_nl;
  wire[0:0] nor_1122_nl;
  wire[0:0] mux_1690_nl;
  wire[0:0] nor_1061_nl;
  wire[0:0] nor_1062_nl;
  wire[0:0] and_503_nl;
  wire[0:0] nor_893_nl;
  wire[0:0] and_493_nl;
  wire[0:0] mux_1940_nl;
  wire[0:0] nor_839_nl;
  wire[0:0] mux_2254_nl;
  wire[0:0] mux_2253_nl;
  wire[0:0] mux_2252_nl;
  wire[0:0] mux_2251_nl;
  wire[0:0] mux_2250_nl;
  wire[0:0] mux_2249_nl;
  wire[0:0] mux_2245_nl;
  wire[0:0] mux_2242_nl;
  wire[0:0] VEC_LOOP_j_not_1_nl;
  wire[0:0] nor_1870_nl;
  wire[0:0] and_nl;
  wire[0:0] nand_nl;
  wire[0:0] mux_1074_nl;
  wire[0:0] nor_1622_nl;
  wire[0:0] and_568_nl;
  wire[0:0] mux_2558_nl;
  wire[0:0] or_nl;
  wire[0:0] mux_nl;
  wire[0:0] nand_325_nl;
  wire[0:0] nand_323_nl;
  wire[0:0] mux_2309_nl;
  wire[0:0] mux_2308_nl;
  wire[0:0] mux_2312_nl;
  wire[0:0] and_270_nl;
  wire[0:0] mux_2314_nl;
  wire[0:0] nand_320_nl;
  wire[0:0] mux_2315_nl;
  wire[0:0] nand_111_nl;
  wire[10:0] COMP_LOOP_3_acc_nl;
  wire[11:0] nl_COMP_LOOP_3_acc_nl;
  wire[0:0] mux_2317_nl;
  wire[0:0] mux_2316_nl;
  wire[0:0] mux_2319_nl;
  wire[0:0] mux_2318_nl;
  wire[8:0] COMP_LOOP_acc_12_nl;
  wire[9:0] nl_COMP_LOOP_acc_12_nl;
  wire[0:0] mux_2321_nl;
  wire[0:0] mux_2320_nl;
  wire[0:0] nand_110_nl;
  wire[0:0] mux_2326_nl;
  wire[0:0] and_823_nl;
  wire[10:0] COMP_LOOP_5_acc_nl;
  wire[11:0] nl_COMP_LOOP_5_acc_nl;
  wire[0:0] mux_2327_nl;
  wire[0:0] and_412_nl;
  wire[0:0] mux_2332_nl;
  wire[0:0] mux_2331_nl;
  wire[10:0] COMP_LOOP_6_acc_nl;
  wire[11:0] nl_COMP_LOOP_6_acc_nl;
  wire[0:0] mux_2335_nl;
  wire[0:0] mux_2334_nl;
  wire[0:0] mux_2333_nl;
  wire[0:0] and_408_nl;
  wire[0:0] mux_2338_nl;
  wire[0:0] mux_2336_nl;
  wire[0:0] mux_2340_nl;
  wire[0:0] mux_2339_nl;
  wire[10:0] COMP_LOOP_7_acc_nl;
  wire[11:0] nl_COMP_LOOP_7_acc_nl;
  wire[0:0] mux_2341_nl;
  wire[0:0] and_405_nl;
  wire[0:0] mux_2346_nl;
  wire[0:0] mux_2345_nl;
  wire[0:0] mux_2349_nl;
  wire[0:0] mux_2348_nl;
  wire[7:0] COMP_LOOP_acc_15_nl;
  wire[8:0] nl_COMP_LOOP_acc_15_nl;
  wire[0:0] mux_2352_nl;
  wire[0:0] mux_2351_nl;
  wire[0:0] mux_2350_nl;
  wire[0:0] mux_2354_nl;
  wire[0:0] and_296_nl;
  wire[0:0] mux_2355_nl;
  wire[0:0] and_397_nl;
  wire[10:0] COMP_LOOP_9_acc_nl;
  wire[11:0] nl_COMP_LOOP_9_acc_nl;
  wire[0:0] mux_2356_nl;
  wire[0:0] and_299_nl;
  wire[0:0] mux_2364_nl;
  wire[0:0] mux_2368_nl;
  wire[10:0] COMP_LOOP_10_acc_nl;
  wire[11:0] nl_COMP_LOOP_10_acc_nl;
  wire[0:0] mux_2372_nl;
  wire[0:0] mux_2371_nl;
  wire[0:0] mux_2375_nl;
  wire[0:0] mux_2378_nl;
  wire[10:0] COMP_LOOP_11_acc_nl;
  wire[11:0] nl_COMP_LOOP_11_acc_nl;
  wire[0:0] and_390_nl;
  wire[0:0] mux_2389_nl;
  wire[0:0] mux_2392_nl;
  wire[0:0] mux_2391_nl;
  wire[8:0] COMP_LOOP_acc_18_nl;
  wire[9:0] nl_COMP_LOOP_acc_18_nl;
  wire[0:0] mux_2395_nl;
  wire[0:0] mux_2394_nl;
  wire[0:0] mux_2400_nl;
  wire[0:0] mux_2399_nl;
  wire[0:0] nor_581_nl;
  wire[0:0] and_379_nl;
  wire[0:0] and_380_nl;
  wire[0:0] mux_2402_nl;
  wire[10:0] COMP_LOOP_13_acc_nl;
  wire[11:0] nl_COMP_LOOP_13_acc_nl;
  wire[0:0] mux_2405_nl;
  wire[0:0] mux_2415_nl;
  wire[0:0] mux_2418_nl;
  wire[0:0] mux_2417_nl;
  wire[10:0] COMP_LOOP_14_acc_nl;
  wire[11:0] nl_COMP_LOOP_14_acc_nl;
  wire[0:0] mux_2422_nl;
  wire[0:0] mux_2421_nl;
  wire[0:0] mux_2426_nl;
  wire[0:0] mux_2425_nl;
  wire[0:0] nor_580_nl;
  wire[0:0] mux_2428_nl;
  wire[10:0] COMP_LOOP_15_acc_nl;
  wire[11:0] nl_COMP_LOOP_15_acc_nl;
  wire[0:0] mux_2431_nl;
  wire[0:0] mux_2436_nl;
  wire[0:0] mux_2438_nl;
  wire[6:0] COMP_LOOP_acc_21_nl;
  wire[7:0] nl_COMP_LOOP_acc_21_nl;
  wire[0:0] nor_298_nl;
  wire[0:0] or_614_nl;
  wire[0:0] mux_951_nl;
  wire[0:0] nor_1642_nl;
  wire[0:0] and_303_nl;
  wire[0:0] and_363_nl;
  wire[10:0] COMP_LOOP_1_acc_nl;
  wire[11:0] nl_COMP_LOOP_1_acc_nl;
  wire[0:0] and_304_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_17_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_19_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_20_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_21_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_23_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_24_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_25_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_26_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_27_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_28_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_29_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_nor_1_nl;
  wire[0:0] COMP_LOOP_nor_11_nl;
  wire[0:0] COMP_LOOP_nor_12_nl;
  wire[0:0] COMP_LOOP_nor_14_nl;
  wire[0:0] COMP_LOOP_nor_17_nl;
  wire[0:0] and_311_nl;
  wire[0:0] mux_2565_nl;
  wire[0:0] mux_2564_nl;
  wire[0:0] or_2758_nl;
  wire[0:0] mux_2563_nl;
  wire[0:0] mux_2562_nl;
  wire[0:0] mux_2561_nl;
  wire[0:0] mux_2560_nl;
  wire[0:0] or_2756_nl;
  wire[0:0] or_2754_nl;
  wire[0:0] COMP_LOOP_tmp_or_33_nl;
  wire[0:0] COMP_LOOP_tmp_and_55_nl;
  wire[0:0] COMP_LOOP_tmp_and_56_nl;
  wire[0:0] COMP_LOOP_tmp_and_57_nl;
  wire[0:0] COMP_LOOP_tmp_and_58_nl;
  wire[0:0] COMP_LOOP_tmp_and_59_nl;
  wire[0:0] mux_2463_nl;
  wire[0:0] mux_2462_nl;
  wire[0:0] mux_2461_nl;
  wire[0:0] mux_2460_nl;
  wire[0:0] mux_2459_nl;
  wire[0:0] mux_2458_nl;
  wire[0:0] or_2563_nl;
  wire[63:0] COMP_LOOP_acc_23_nl;
  wire[64:0] nl_COMP_LOOP_acc_23_nl;
  wire[63:0] COMP_LOOP_COMP_LOOP_mux_9_nl;
  wire[0:0] COMP_LOOP_or_nl;
  wire[0:0] COMP_LOOP_or_1_nl;
  wire[0:0] COMP_LOOP_or_2_nl;
  wire[0:0] COMP_LOOP_or_3_nl;
  wire[0:0] COMP_LOOP_or_4_nl;
  wire[0:0] COMP_LOOP_or_5_nl;
  wire[0:0] COMP_LOOP_or_6_nl;
  wire[0:0] COMP_LOOP_or_7_nl;
  wire[0:0] COMP_LOOP_or_8_nl;
  wire[0:0] COMP_LOOP_or_9_nl;
  wire[0:0] COMP_LOOP_or_10_nl;
  wire[0:0] COMP_LOOP_or_11_nl;
  wire[0:0] COMP_LOOP_or_12_nl;
  wire[0:0] COMP_LOOP_or_13_nl;
  wire[0:0] COMP_LOOP_or_14_nl;
  wire[0:0] COMP_LOOP_or_15_nl;
  wire[0:0] COMP_LOOP_or_21_nl;
  wire[0:0] COMP_LOOP_or_22_nl;
  wire[0:0] COMP_LOOP_tmp_and_42_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_1_nl;
  wire[0:0] COMP_LOOP_tmp_and_43_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl;
  wire[0:0] COMP_LOOP_tmp_and_44_nl;
  wire[0:0] COMP_LOOP_tmp_and_45_nl;
  wire[0:0] COMP_LOOP_tmp_and_46_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_7_nl;
  wire[0:0] COMP_LOOP_tmp_and_47_nl;
  wire[0:0] COMP_LOOP_tmp_and_48_nl;
  wire[0:0] COMP_LOOP_tmp_and_49_nl;
  wire[0:0] COMP_LOOP_tmp_and_50_nl;
  wire[0:0] COMP_LOOP_tmp_and_51_nl;
  wire[0:0] COMP_LOOP_tmp_and_52_nl;
  wire[0:0] COMP_LOOP_tmp_and_53_nl;
  wire[0:0] and_336_nl;
  wire[0:0] and_340_nl;
  wire[0:0] mux_2504_nl;
  wire[0:0] mux_2503_nl;
  wire[0:0] mux_2502_nl;
  wire[0:0] mux_2501_nl;
  wire[0:0] or_2595_nl;
  wire[0:0] mux_2500_nl;
  wire[0:0] mux_2499_nl;
  wire[0:0] or_2593_nl;
  wire[0:0] or_2591_nl;
  wire[0:0] COMP_LOOP_tmp_and_36_nl;
  wire[0:0] COMP_LOOP_tmp_and_37_nl;
  wire[0:0] COMP_LOOP_tmp_and_38_nl;
  wire[0:0] COMP_LOOP_tmp_and_39_nl;
  wire[0:0] COMP_LOOP_tmp_and_40_nl;
  wire[0:0] COMP_LOOP_tmp_and_41_nl;
  wire[0:0] COMP_LOOP_tmp_and_20_nl;
  wire[0:0] COMP_LOOP_tmp_and_21_nl;
  wire[0:0] COMP_LOOP_tmp_and_22_nl;
  wire[0:0] COMP_LOOP_tmp_and_23_nl;
  wire[0:0] COMP_LOOP_tmp_and_24_nl;
  wire[0:0] COMP_LOOP_tmp_and_25_nl;
  wire[0:0] COMP_LOOP_tmp_and_26_nl;
  wire[0:0] COMP_LOOP_tmp_and_27_nl;
  wire[0:0] COMP_LOOP_tmp_and_28_nl;
  wire[0:0] COMP_LOOP_tmp_and_29_nl;
  wire[0:0] COMP_LOOP_tmp_and_30_nl;
  wire[0:0] COMP_LOOP_tmp_and_31_nl;
  wire[0:0] COMP_LOOP_tmp_and_32_nl;
  wire[0:0] COMP_LOOP_tmp_and_33_nl;
  wire[0:0] COMP_LOOP_tmp_and_34_nl;
  wire[0:0] COMP_LOOP_tmp_and_35_nl;
  wire[0:0] COMP_LOOP_tmp_and_nl;
  wire[0:0] COMP_LOOP_tmp_and_17_nl;
  wire[0:0] COMP_LOOP_tmp_and_18_nl;
  wire[0:0] mux_2518_nl;
  wire[0:0] mux_2517_nl;
  wire[0:0] mux_2516_nl;
  wire[0:0] mux_2515_nl;
  wire[0:0] mux_2514_nl;
  wire[0:0] mux_2520_nl;
  wire[0:0] mux_2519_nl;
  wire[0:0] and_357_nl;
  wire[0:0] mux_2532_nl;
  wire[0:0] mux_2531_nl;
  wire[0:0] mux_2530_nl;
  wire[0:0] mux_2529_nl;
  wire[0:0] mux_2528_nl;
  wire[0:0] mux_2527_nl;
  wire[0:0] mux_2526_nl;
  wire[0:0] COMP_LOOP_tmp_and_7_nl;
  wire[0:0] COMP_LOOP_tmp_and_8_nl;
  wire[0:0] COMP_LOOP_tmp_and_9_nl;
  wire[0:0] COMP_LOOP_tmp_and_10_nl;
  wire[0:0] COMP_LOOP_tmp_and_11_nl;
  wire[0:0] COMP_LOOP_tmp_and_12_nl;
  wire[0:0] mux_2542_nl;
  wire[0:0] nor_568_nl;
  wire[0:0] mux_2541_nl;
  wire[0:0] mux_2540_nl;
  wire[0:0] mux_2539_nl;
  wire[0:0] mux_2546_nl;
  wire[0:0] mux_2545_nl;
  wire[0:0] mux_2544_nl;
  wire[0:0] mux_2543_nl;
  wire[0:0] and_352_nl;
  wire[0:0] COMP_LOOP_tmp_and_2_nl;
  wire[0:0] COMP_LOOP_tmp_and_3_nl;
  wire[0:0] COMP_LOOP_tmp_and_4_nl;
  wire[0:0] COMP_LOOP_tmp_and_5_nl;
  wire[0:0] COMP_LOOP_tmp_and_6_nl;
  wire[0:0] mux_2553_nl;
  wire[0:0] mux_2552_nl;
  wire[0:0] mux_2551_nl;
  wire[0:0] mux_561_nl;
  wire[0:0] mux_560_nl;
  wire[0:0] mux_2556_nl;
  wire[0:0] mux_2555_nl;
  wire[0:0] mux_2554_nl;
  wire[0:0] or_2625_nl;
  wire[10:0] COMP_LOOP_1_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_1_acc_10_nl;
  wire[10:0] COMP_LOOP_2_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_2_acc_10_nl;
  wire[10:0] COMP_LOOP_3_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_3_acc_10_nl;
  wire[10:0] COMP_LOOP_4_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_4_acc_10_nl;
  wire[10:0] COMP_LOOP_5_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_5_acc_10_nl;
  wire[10:0] COMP_LOOP_6_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_6_acc_10_nl;
  wire[10:0] COMP_LOOP_7_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_7_acc_10_nl;
  wire[10:0] COMP_LOOP_8_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_8_acc_10_nl;
  wire[10:0] COMP_LOOP_9_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_9_acc_10_nl;
  wire[10:0] COMP_LOOP_10_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_10_acc_10_nl;
  wire[10:0] COMP_LOOP_11_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_11_acc_10_nl;
  wire[10:0] COMP_LOOP_12_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_12_acc_10_nl;
  wire[10:0] COMP_LOOP_13_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_13_acc_10_nl;
  wire[10:0] COMP_LOOP_14_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_14_acc_10_nl;
  wire[10:0] COMP_LOOP_15_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_15_acc_10_nl;
  wire[10:0] COMP_LOOP_16_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_16_acc_10_nl;
  wire[0:0] and_313_nl;
  wire[0:0] mux_1080_nl;
  wire[0:0] and_565_nl;
  wire[0:0] or_714_nl;
  wire[0:0] nand_22_nl;
  wire[0:0] mux_1083_nl;
  wire[0:0] nand_23_nl;
  wire[0:0] mux_1085_nl;
  wire[0:0] or_712_nl;
  wire[0:0] or_762_nl;
  wire[0:0] mux_1115_nl;
  wire[0:0] or_760_nl;
  wire[0:0] or_758_nl;
  wire[0:0] nor_1479_nl;
  wire[0:0] mux_1240_nl;
  wire[0:0] nor_1480_nl;
  wire[0:0] nor_1481_nl;
  wire[0:0] or_1150_nl;
  wire[0:0] mux_1365_nl;
  wire[0:0] or_1148_nl;
  wire[0:0] or_1146_nl;
  wire[0:0] nor_1242_nl;
  wire[0:0] mux_1490_nl;
  wire[0:0] nor_1243_nl;
  wire[0:0] nor_1244_nl;
  wire[0:0] or_1538_nl;
  wire[0:0] mux_1615_nl;
  wire[0:0] or_1536_nl;
  wire[0:0] or_1534_nl;
  wire[0:0] nor_1012_nl;
  wire[0:0] mux_1740_nl;
  wire[0:0] nor_1013_nl;
  wire[0:0] nor_1014_nl;
  wire[0:0] nand_322_nl;
  wire[0:0] mux_1865_nl;
  wire[0:0] or_1922_nl;
  wire[0:0] or_1920_nl;
  wire[0:0] and_835_nl;
  wire[0:0] mux_1990_nl;
  wire[0:0] nor_795_nl;
  wire[0:0] nor_796_nl;
  wire[0:0] or_2430_nl;
  wire[0:0] or_2434_nl;
  wire[0:0] or_2435_nl;
  wire[0:0] or_2443_nl;
  wire[0:0] mux_2263_nl;
  wire[0:0] or_2444_nl;
  wire[0:0] or_2440_nl;
  wire[0:0] mux_2267_nl;
  wire[0:0] nand_114_nl;
  wire[0:0] nand_113_nl;
  wire[0:0] or_2455_nl;
  wire[0:0] or_2482_nl;
  wire[0:0] or_2481_nl;
  wire[0:0] mux_2302_nl;
  wire[0:0] mux_2306_nl;
  wire[0:0] mux_2305_nl;
  wire[0:0] and_416_nl;
  wire[0:0] mux_22_nl;
  wire[0:0] mux_2325_nl;
  wire[0:0] mux_2324_nl;
  wire[0:0] mux_2323_nl;
  wire[0:0] or_2497_nl;
  wire[0:0] mux_61_nl;
  wire[0:0] mux_2328_nl;
  wire[0:0] and_411_nl;
  wire[0:0] mux_2329_nl;
  wire[0:0] mux_2343_nl;
  wire[0:0] mux_2342_nl;
  wire[0:0] and_403_nl;
  wire[0:0] or_2507_nl;
  wire[0:0] or_2506_nl;
  wire[0:0] and_401_nl;
  wire[0:0] mux_2353_nl;
  wire[0:0] and_398_nl;
  wire[0:0] mux_2359_nl;
  wire[0:0] mux_2358_nl;
  wire[0:0] mux_2357_nl;
  wire[0:0] and_396_nl;
  wire[0:0] mux_2362_nl;
  wire[0:0] mux_2361_nl;
  wire[0:0] and_566_nl;
  wire[0:0] mux_2374_nl;
  wire[0:0] and_392_nl;
  wire[0:0] mux_2382_nl;
  wire[0:0] mux_2381_nl;
  wire[0:0] and_388_nl;
  wire[0:0] mux_2387_nl;
  wire[0:0] mux_2386_nl;
  wire[0:0] mux_2397_nl;
  wire[0:0] mux_2409_nl;
  wire[0:0] mux_2408_nl;
  wire[0:0] mux_2407_nl;
  wire[0:0] and_376_nl;
  wire[0:0] mux_2413_nl;
  wire[0:0] mux_2412_nl;
  wire[0:0] and_372_nl;
  wire[0:0] and_370_nl;
  wire[0:0] mux_2434_nl;
  wire[0:0] mux_2433_nl;
  wire[0:0] and_366_nl;
  wire[0:0] mux_2441_nl;
  wire[0:0] mux_2440_nl;
  wire[0:0] mux_2443_nl;
  wire[0:0] mux_2448_nl;
  wire[0:0] or_427_nl;
  wire[0:0] or_2571_nl;
  wire[0:0] mux_2468_nl;
  wire[0:0] and_361_nl;
  wire[0:0] nor_577_nl;
  wire[0:0] nor_576_nl;
  wire[0:0] mux_2471_nl;
  wire[0:0] nand_103_nl;
  wire[0:0] and_360_nl;
  wire[0:0] mux_2470_nl;
  wire[0:0] nand_101_nl;
  wire[0:0] mux_2467_nl;
  wire[0:0] or_2569_nl;
  wire[4:0] STAGE_LOOP_acc_nl;
  wire[5:0] nl_STAGE_LOOP_acc_nl;
  wire[0:0] mux_2498_nl;
  wire[0:0] nor_575_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] or_44_nl;
  wire[0:0] mux_2509_nl;
  wire[0:0] mux_2508_nl;
  wire[0:0] mux_2507_nl;
  wire[0:0] nand_107_nl;
  wire[0:0] mux_2512_nl;
  wire[0:0] nor_570_nl;
  wire[0:0] mux_2511_nl;
  wire[0:0] mux_2510_nl;
  wire[0:0] mux_2525_nl;
  wire[0:0] mux_2524_nl;
  wire[0:0] mux_2523_nl;
  wire[0:0] and_354_nl;
  wire[0:0] mux_2522_nl;
  wire[0:0] and_356_nl;
  wire[0:0] mux_2538_nl;
  wire[0:0] mux_2537_nl;
  wire[0:0] mux_2536_nl;
  wire[0:0] mux_234_nl;
  wire[0:0] nor_1750_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] mux_232_nl;
  wire[0:0] mux_1089_nl;
  wire[0:0] mux_1088_nl;
  wire[0:0] or_715_nl;
  wire[0:0] mux_1087_nl;
  wire[0:0] or_711_nl;
  wire[0:0] and_94_nl;
  wire[0:0] and_99_nl;
  wire[0:0] and_106_nl;
  wire[0:0] and_110_nl;
  wire[0:0] and_116_nl;
  wire[0:0] and_120_nl;
  wire[0:0] and_124_nl;
  wire[0:0] and_127_nl;
  wire[0:0] and_132_nl;
  wire[0:0] and_135_nl;
  wire[0:0] and_140_nl;
  wire[0:0] and_143_nl;
  wire[0:0] and_148_nl;
  wire[0:0] and_152_nl;
  wire[0:0] and_155_nl;
  wire[0:0] and_158_nl;
  wire[0:0] and_159_nl;
  wire[0:0] and_160_nl;
  wire[0:0] and_161_nl;
  wire[0:0] and_163_nl;
  wire[0:0] and_164_nl;
  wire[0:0] and_165_nl;
  wire[0:0] and_166_nl;
  wire[0:0] and_168_nl;
  wire[0:0] and_169_nl;
  wire[0:0] and_170_nl;
  wire[0:0] and_171_nl;
  wire[0:0] and_173_nl;
  wire[0:0] and_174_nl;
  wire[0:0] and_175_nl;
  wire[0:0] and_176_nl;
  wire[0:0] and_178_nl;
  wire[0:0] and_179_nl;
  wire[0:0] and_180_nl;
  wire[0:0] and_181_nl;
  wire[0:0] and_183_nl;
  wire[0:0] and_184_nl;
  wire[0:0] and_185_nl;
  wire[0:0] and_186_nl;
  wire[0:0] and_188_nl;
  wire[0:0] and_189_nl;
  wire[0:0] and_190_nl;
  wire[0:0] and_191_nl;
  wire[0:0] and_193_nl;
  wire[0:0] and_194_nl;
  wire[0:0] and_195_nl;
  wire[0:0] and_196_nl;
  wire[0:0] nor_1596_nl;
  wire[0:0] mux_1119_nl;
  wire[0:0] mux_1118_nl;
  wire[0:0] nor_1597_nl;
  wire[0:0] mux_1117_nl;
  wire[0:0] or_763_nl;
  wire[0:0] mux_1114_nl;
  wire[0:0] mux_1113_nl;
  wire[0:0] or_757_nl;
  wire[0:0] or_755_nl;
  wire[0:0] mux_1112_nl;
  wire[0:0] or_753_nl;
  wire[0:0] or_752_nl;
  wire[0:0] mux_1111_nl;
  wire[0:0] mux_1110_nl;
  wire[0:0] mux_1109_nl;
  wire[0:0] nor_1598_nl;
  wire[0:0] nor_1599_nl;
  wire[0:0] mux_1108_nl;
  wire[0:0] nor_1600_nl;
  wire[0:0] nor_1601_nl;
  wire[0:0] mux_1107_nl;
  wire[0:0] mux_1106_nl;
  wire[0:0] nor_1602_nl;
  wire[0:0] nor_1603_nl;
  wire[0:0] mux_1105_nl;
  wire[0:0] nor_1604_nl;
  wire[0:0] nor_1605_nl;
  wire[0:0] mux_1104_nl;
  wire[0:0] mux_1103_nl;
  wire[0:0] mux_1102_nl;
  wire[0:0] mux_1101_nl;
  wire[0:0] nor_1606_nl;
  wire[0:0] nor_1607_nl;
  wire[0:0] mux_1100_nl;
  wire[0:0] nor_1608_nl;
  wire[0:0] nor_1609_nl;
  wire[0:0] mux_1099_nl;
  wire[0:0] mux_1098_nl;
  wire[0:0] nor_1610_nl;
  wire[0:0] nor_1611_nl;
  wire[0:0] mux_1097_nl;
  wire[0:0] nor_1612_nl;
  wire[0:0] nor_1613_nl;
  wire[0:0] mux_1096_nl;
  wire[0:0] mux_1095_nl;
  wire[0:0] mux_1094_nl;
  wire[0:0] nor_1614_nl;
  wire[0:0] nor_1615_nl;
  wire[0:0] mux_1093_nl;
  wire[0:0] nor_1616_nl;
  wire[0:0] nor_1617_nl;
  wire[0:0] mux_1092_nl;
  wire[0:0] mux_1091_nl;
  wire[0:0] nor_1618_nl;
  wire[0:0] nor_1619_nl;
  wire[0:0] mux_1090_nl;
  wire[0:0] nor_1620_nl;
  wire[0:0] nor_1621_nl;
  wire[0:0] mux_1150_nl;
  wire[0:0] mux_1149_nl;
  wire[0:0] mux_1148_nl;
  wire[0:0] nor_1569_nl;
  wire[0:0] mux_1147_nl;
  wire[0:0] mux_1146_nl;
  wire[0:0] nor_1570_nl;
  wire[0:0] nor_1571_nl;
  wire[0:0] nor_1572_nl;
  wire[0:0] mux_1145_nl;
  wire[0:0] mux_1144_nl;
  wire[0:0] mux_1143_nl;
  wire[0:0] nor_1573_nl;
  wire[0:0] nor_1574_nl;
  wire[0:0] nor_1575_nl;
  wire[0:0] nor_1576_nl;
  wire[0:0] mux_1142_nl;
  wire[0:0] mux_1141_nl;
  wire[0:0] mux_1140_nl;
  wire[0:0] nor_1577_nl;
  wire[0:0] mux_1139_nl;
  wire[0:0] nor_1578_nl;
  wire[0:0] nor_1579_nl;
  wire[0:0] nor_1580_nl;
  wire[0:0] mux_1138_nl;
  wire[0:0] nor_1581_nl;
  wire[0:0] mux_1137_nl;
  wire[0:0] mux_1136_nl;
  wire[0:0] nor_1582_nl;
  wire[0:0] nor_1583_nl;
  wire[0:0] nor_1584_nl;
  wire[0:0] mux_1135_nl;
  wire[0:0] mux_1134_nl;
  wire[0:0] mux_1133_nl;
  wire[0:0] and_561_nl;
  wire[0:0] mux_1132_nl;
  wire[0:0] nor_1585_nl;
  wire[0:0] nor_1586_nl;
  wire[0:0] nor_1587_nl;
  wire[0:0] mux_1131_nl;
  wire[0:0] or_785_nl;
  wire[0:0] or_783_nl;
  wire[0:0] mux_1130_nl;
  wire[0:0] nor_1588_nl;
  wire[0:0] mux_1129_nl;
  wire[0:0] or_781_nl;
  wire[0:0] or_779_nl;
  wire[0:0] and_562_nl;
  wire[0:0] mux_1127_nl;
  wire[0:0] nor_1591_nl;
  wire[0:0] mux_1126_nl;
  wire[0:0] mux_1125_nl;
  wire[0:0] or_775_nl;
  wire[0:0] or_773_nl;
  wire[0:0] mux_1124_nl;
  wire[0:0] or_772_nl;
  wire[0:0] or_770_nl;
  wire[0:0] and_563_nl;
  wire[0:0] mux_1123_nl;
  wire[0:0] mux_1122_nl;
  wire[0:0] nor_1592_nl;
  wire[0:0] nor_1593_nl;
  wire[0:0] mux_1121_nl;
  wire[0:0] nor_1594_nl;
  wire[0:0] nor_1595_nl;
  wire[0:0] nor_1539_nl;
  wire[0:0] mux_1181_nl;
  wire[0:0] mux_1180_nl;
  wire[0:0] and_560_nl;
  wire[0:0] mux_1179_nl;
  wire[0:0] nor_1540_nl;
  wire[0:0] mux_1176_nl;
  wire[0:0] mux_1175_nl;
  wire[0:0] nor_1541_nl;
  wire[0:0] nor_1542_nl;
  wire[0:0] mux_1174_nl;
  wire[0:0] nor_1543_nl;
  wire[0:0] nor_1544_nl;
  wire[0:0] mux_1173_nl;
  wire[0:0] mux_1172_nl;
  wire[0:0] mux_1171_nl;
  wire[0:0] nor_1545_nl;
  wire[0:0] nor_1546_nl;
  wire[0:0] mux_1170_nl;
  wire[0:0] nor_1547_nl;
  wire[0:0] nor_1548_nl;
  wire[0:0] mux_1169_nl;
  wire[0:0] mux_1168_nl;
  wire[0:0] nor_1549_nl;
  wire[0:0] nor_1550_nl;
  wire[0:0] mux_1167_nl;
  wire[0:0] nor_1551_nl;
  wire[0:0] nor_1552_nl;
  wire[0:0] mux_1166_nl;
  wire[0:0] mux_1165_nl;
  wire[0:0] mux_1164_nl;
  wire[0:0] mux_1163_nl;
  wire[0:0] nor_1553_nl;
  wire[0:0] mux_1162_nl;
  wire[0:0] nor_1556_nl;
  wire[0:0] mux_1161_nl;
  wire[0:0] mux_1160_nl;
  wire[0:0] nor_1557_nl;
  wire[0:0] mux_1159_nl;
  wire[0:0] nor_1560_nl;
  wire[0:0] mux_1158_nl;
  wire[0:0] mux_1157_nl;
  wire[0:0] mux_1156_nl;
  wire[0:0] nor_1561_nl;
  wire[0:0] nor_1562_nl;
  wire[0:0] mux_1155_nl;
  wire[0:0] nor_1563_nl;
  wire[0:0] nor_1564_nl;
  wire[0:0] mux_1154_nl;
  wire[0:0] mux_1153_nl;
  wire[0:0] nor_1565_nl;
  wire[0:0] nor_1566_nl;
  wire[0:0] mux_1152_nl;
  wire[0:0] nor_1567_nl;
  wire[0:0] nor_1568_nl;
  wire[0:0] mux_1213_nl;
  wire[0:0] mux_1212_nl;
  wire[0:0] mux_1211_nl;
  wire[0:0] mux_1210_nl;
  wire[0:0] nor_1506_nl;
  wire[0:0] nor_1507_nl;
  wire[0:0] mux_1209_nl;
  wire[0:0] nor_1508_nl;
  wire[0:0] nor_1509_nl;
  wire[0:0] mux_1208_nl;
  wire[0:0] mux_1207_nl;
  wire[0:0] nor_1510_nl;
  wire[0:0] nor_1511_nl;
  wire[0:0] nor_1512_nl;
  wire[0:0] mux_1206_nl;
  wire[0:0] mux_1205_nl;
  wire[0:0] mux_1204_nl;
  wire[0:0] nor_1513_nl;
  wire[0:0] nor_1514_nl;
  wire[0:0] mux_1203_nl;
  wire[0:0] nor_1515_nl;
  wire[0:0] nor_1516_nl;
  wire[0:0] mux_1202_nl;
  wire[0:0] mux_1201_nl;
  wire[0:0] nor_1517_nl;
  wire[0:0] nor_1518_nl;
  wire[0:0] mux_1200_nl;
  wire[0:0] mux_1199_nl;
  wire[0:0] nor_1519_nl;
  wire[0:0] nor_1520_nl;
  wire[0:0] nor_1521_nl;
  wire[0:0] and_557_nl;
  wire[0:0] mux_1198_nl;
  wire[0:0] mux_1197_nl;
  wire[0:0] mux_1196_nl;
  wire[0:0] mux_1195_nl;
  wire[0:0] and_558_nl;
  wire[0:0] mux_1194_nl;
  wire[0:0] nor_1524_nl;
  wire[0:0] nor_1525_nl;
  wire[0:0] mux_1193_nl;
  wire[0:0] mux_1192_nl;
  wire[0:0] and_559_nl;
  wire[0:0] mux_1189_nl;
  wire[0:0] mux_1188_nl;
  wire[0:0] mux_1187_nl;
  wire[0:0] nor_1531_nl;
  wire[0:0] nor_1532_nl;
  wire[0:0] mux_1186_nl;
  wire[0:0] nor_1533_nl;
  wire[0:0] nor_1534_nl;
  wire[0:0] mux_1185_nl;
  wire[0:0] mux_1184_nl;
  wire[0:0] nor_1535_nl;
  wire[0:0] nor_1536_nl;
  wire[0:0] mux_1183_nl;
  wire[0:0] nor_1537_nl;
  wire[0:0] nor_1538_nl;
  wire[0:0] nor_1477_nl;
  wire[0:0] mux_1244_nl;
  wire[0:0] mux_1243_nl;
  wire[0:0] nor_1478_nl;
  wire[0:0] mux_1242_nl;
  wire[0:0] nand_31_nl;
  wire[0:0] mux_1239_nl;
  wire[0:0] mux_1238_nl;
  wire[0:0] or_952_nl;
  wire[0:0] or_950_nl;
  wire[0:0] mux_1237_nl;
  wire[0:0] or_948_nl;
  wire[0:0] or_947_nl;
  wire[0:0] mux_1236_nl;
  wire[0:0] mux_1235_nl;
  wire[0:0] mux_1234_nl;
  wire[0:0] nor_1482_nl;
  wire[0:0] nor_1483_nl;
  wire[0:0] mux_1233_nl;
  wire[0:0] nor_1484_nl;
  wire[0:0] nor_1485_nl;
  wire[0:0] mux_1232_nl;
  wire[0:0] mux_1231_nl;
  wire[0:0] nor_1486_nl;
  wire[0:0] nor_1487_nl;
  wire[0:0] mux_1230_nl;
  wire[0:0] nor_1488_nl;
  wire[0:0] nor_1489_nl;
  wire[0:0] mux_1229_nl;
  wire[0:0] mux_1228_nl;
  wire[0:0] mux_1227_nl;
  wire[0:0] mux_1226_nl;
  wire[0:0] nor_1490_nl;
  wire[0:0] nor_1491_nl;
  wire[0:0] mux_1225_nl;
  wire[0:0] nor_1492_nl;
  wire[0:0] nor_1493_nl;
  wire[0:0] mux_1224_nl;
  wire[0:0] mux_1223_nl;
  wire[0:0] nor_1494_nl;
  wire[0:0] nor_1495_nl;
  wire[0:0] mux_1222_nl;
  wire[0:0] nor_1496_nl;
  wire[0:0] nor_1497_nl;
  wire[0:0] mux_1221_nl;
  wire[0:0] mux_1220_nl;
  wire[0:0] mux_1219_nl;
  wire[0:0] nor_1498_nl;
  wire[0:0] nor_1499_nl;
  wire[0:0] mux_1218_nl;
  wire[0:0] nor_1500_nl;
  wire[0:0] nor_1501_nl;
  wire[0:0] mux_1217_nl;
  wire[0:0] mux_1216_nl;
  wire[0:0] nor_1502_nl;
  wire[0:0] nor_1503_nl;
  wire[0:0] mux_1215_nl;
  wire[0:0] nor_1504_nl;
  wire[0:0] nor_1505_nl;
  wire[0:0] mux_1275_nl;
  wire[0:0] mux_1274_nl;
  wire[0:0] mux_1273_nl;
  wire[0:0] nor_1450_nl;
  wire[0:0] mux_1272_nl;
  wire[0:0] mux_1271_nl;
  wire[0:0] nor_1451_nl;
  wire[0:0] nor_1452_nl;
  wire[0:0] nor_1453_nl;
  wire[0:0] mux_1270_nl;
  wire[0:0] mux_1269_nl;
  wire[0:0] mux_1268_nl;
  wire[0:0] nor_1454_nl;
  wire[0:0] nor_1455_nl;
  wire[0:0] nor_1456_nl;
  wire[0:0] nor_1457_nl;
  wire[0:0] mux_1267_nl;
  wire[0:0] mux_1266_nl;
  wire[0:0] mux_1265_nl;
  wire[0:0] nor_1458_nl;
  wire[0:0] mux_1264_nl;
  wire[0:0] nor_1459_nl;
  wire[0:0] nor_1460_nl;
  wire[0:0] nor_1461_nl;
  wire[0:0] mux_1263_nl;
  wire[0:0] nor_1462_nl;
  wire[0:0] mux_1262_nl;
  wire[0:0] mux_1261_nl;
  wire[0:0] nor_1463_nl;
  wire[0:0] nor_1464_nl;
  wire[0:0] nor_1465_nl;
  wire[0:0] mux_1260_nl;
  wire[0:0] mux_1259_nl;
  wire[0:0] mux_1258_nl;
  wire[0:0] and_554_nl;
  wire[0:0] mux_1257_nl;
  wire[0:0] nor_1466_nl;
  wire[0:0] nor_1467_nl;
  wire[0:0] nor_1468_nl;
  wire[0:0] mux_1256_nl;
  wire[0:0] or_979_nl;
  wire[0:0] or_977_nl;
  wire[0:0] mux_1255_nl;
  wire[0:0] nor_1469_nl;
  wire[0:0] mux_1254_nl;
  wire[0:0] or_975_nl;
  wire[0:0] or_973_nl;
  wire[0:0] and_555_nl;
  wire[0:0] mux_1252_nl;
  wire[0:0] nor_1472_nl;
  wire[0:0] mux_1251_nl;
  wire[0:0] mux_1250_nl;
  wire[0:0] or_969_nl;
  wire[0:0] or_967_nl;
  wire[0:0] mux_1249_nl;
  wire[0:0] or_966_nl;
  wire[0:0] or_964_nl;
  wire[0:0] and_556_nl;
  wire[0:0] mux_1248_nl;
  wire[0:0] mux_1247_nl;
  wire[0:0] nor_1473_nl;
  wire[0:0] nor_1474_nl;
  wire[0:0] mux_1246_nl;
  wire[0:0] nor_1475_nl;
  wire[0:0] nor_1476_nl;
  wire[0:0] nor_1418_nl;
  wire[0:0] mux_1306_nl;
  wire[0:0] mux_1305_nl;
  wire[0:0] and_552_nl;
  wire[0:0] mux_1304_nl;
  wire[0:0] and_553_nl;
  wire[0:0] mux_1301_nl;
  wire[0:0] mux_1300_nl;
  wire[0:0] nor_1422_nl;
  wire[0:0] nor_1423_nl;
  wire[0:0] mux_1299_nl;
  wire[0:0] nor_1424_nl;
  wire[0:0] nor_1425_nl;
  wire[0:0] mux_1298_nl;
  wire[0:0] mux_1297_nl;
  wire[0:0] mux_1296_nl;
  wire[0:0] nor_1426_nl;
  wire[0:0] nor_1427_nl;
  wire[0:0] mux_1295_nl;
  wire[0:0] nor_1428_nl;
  wire[0:0] nor_1429_nl;
  wire[0:0] mux_1294_nl;
  wire[0:0] mux_1293_nl;
  wire[0:0] nor_1430_nl;
  wire[0:0] nor_1431_nl;
  wire[0:0] mux_1292_nl;
  wire[0:0] nor_1432_nl;
  wire[0:0] nor_1433_nl;
  wire[0:0] mux_1291_nl;
  wire[0:0] mux_1290_nl;
  wire[0:0] mux_1289_nl;
  wire[0:0] mux_1288_nl;
  wire[0:0] nor_1434_nl;
  wire[0:0] mux_1287_nl;
  wire[0:0] nor_1437_nl;
  wire[0:0] mux_1286_nl;
  wire[0:0] mux_1285_nl;
  wire[0:0] nor_1438_nl;
  wire[0:0] mux_1284_nl;
  wire[0:0] nor_1441_nl;
  wire[0:0] mux_1283_nl;
  wire[0:0] mux_1282_nl;
  wire[0:0] mux_1281_nl;
  wire[0:0] nor_1442_nl;
  wire[0:0] nor_1443_nl;
  wire[0:0] mux_1280_nl;
  wire[0:0] nor_1444_nl;
  wire[0:0] nor_1445_nl;
  wire[0:0] mux_1279_nl;
  wire[0:0] mux_1278_nl;
  wire[0:0] nor_1446_nl;
  wire[0:0] nor_1447_nl;
  wire[0:0] mux_1277_nl;
  wire[0:0] nor_1448_nl;
  wire[0:0] nor_1449_nl;
  wire[0:0] mux_1338_nl;
  wire[0:0] mux_1337_nl;
  wire[0:0] mux_1336_nl;
  wire[0:0] mux_1335_nl;
  wire[0:0] nor_1385_nl;
  wire[0:0] nor_1386_nl;
  wire[0:0] mux_1334_nl;
  wire[0:0] nor_1387_nl;
  wire[0:0] nor_1388_nl;
  wire[0:0] mux_1333_nl;
  wire[0:0] mux_1332_nl;
  wire[0:0] nor_1389_nl;
  wire[0:0] nor_1390_nl;
  wire[0:0] nor_1391_nl;
  wire[0:0] mux_1331_nl;
  wire[0:0] mux_1330_nl;
  wire[0:0] mux_1329_nl;
  wire[0:0] nor_1392_nl;
  wire[0:0] nor_1393_nl;
  wire[0:0] mux_1328_nl;
  wire[0:0] nor_1394_nl;
  wire[0:0] nor_1395_nl;
  wire[0:0] mux_1327_nl;
  wire[0:0] mux_1326_nl;
  wire[0:0] nor_1396_nl;
  wire[0:0] nor_1397_nl;
  wire[0:0] mux_1325_nl;
  wire[0:0] mux_1324_nl;
  wire[0:0] nor_1398_nl;
  wire[0:0] nor_1399_nl;
  wire[0:0] nor_1400_nl;
  wire[0:0] and_549_nl;
  wire[0:0] mux_1323_nl;
  wire[0:0] mux_1322_nl;
  wire[0:0] mux_1321_nl;
  wire[0:0] mux_1320_nl;
  wire[0:0] and_550_nl;
  wire[0:0] mux_1319_nl;
  wire[0:0] nor_1403_nl;
  wire[0:0] nor_1404_nl;
  wire[0:0] mux_1318_nl;
  wire[0:0] mux_1317_nl;
  wire[0:0] and_551_nl;
  wire[0:0] mux_1314_nl;
  wire[0:0] mux_1313_nl;
  wire[0:0] mux_1312_nl;
  wire[0:0] nor_1410_nl;
  wire[0:0] nor_1411_nl;
  wire[0:0] mux_1311_nl;
  wire[0:0] nor_1412_nl;
  wire[0:0] nor_1413_nl;
  wire[0:0] mux_1310_nl;
  wire[0:0] mux_1309_nl;
  wire[0:0] nor_1414_nl;
  wire[0:0] nor_1415_nl;
  wire[0:0] mux_1308_nl;
  wire[0:0] nor_1416_nl;
  wire[0:0] nor_1417_nl;
  wire[0:0] nor_1359_nl;
  wire[0:0] mux_1369_nl;
  wire[0:0] mux_1368_nl;
  wire[0:0] nor_1360_nl;
  wire[0:0] mux_1367_nl;
  wire[0:0] or_1151_nl;
  wire[0:0] mux_1364_nl;
  wire[0:0] mux_1363_nl;
  wire[0:0] or_1145_nl;
  wire[0:0] or_1143_nl;
  wire[0:0] mux_1362_nl;
  wire[0:0] or_1141_nl;
  wire[0:0] or_1140_nl;
  wire[0:0] mux_1361_nl;
  wire[0:0] mux_1360_nl;
  wire[0:0] mux_1359_nl;
  wire[0:0] nor_1361_nl;
  wire[0:0] nor_1362_nl;
  wire[0:0] mux_1358_nl;
  wire[0:0] nor_1363_nl;
  wire[0:0] nor_1364_nl;
  wire[0:0] mux_1357_nl;
  wire[0:0] mux_1356_nl;
  wire[0:0] nor_1365_nl;
  wire[0:0] nor_1366_nl;
  wire[0:0] mux_1355_nl;
  wire[0:0] nor_1367_nl;
  wire[0:0] nor_1368_nl;
  wire[0:0] mux_1354_nl;
  wire[0:0] mux_1353_nl;
  wire[0:0] mux_1352_nl;
  wire[0:0] mux_1351_nl;
  wire[0:0] nor_1369_nl;
  wire[0:0] nor_1370_nl;
  wire[0:0] mux_1350_nl;
  wire[0:0] nor_1371_nl;
  wire[0:0] nor_1372_nl;
  wire[0:0] mux_1349_nl;
  wire[0:0] mux_1348_nl;
  wire[0:0] nor_1373_nl;
  wire[0:0] nor_1374_nl;
  wire[0:0] mux_1347_nl;
  wire[0:0] nor_1375_nl;
  wire[0:0] nor_1376_nl;
  wire[0:0] mux_1346_nl;
  wire[0:0] mux_1345_nl;
  wire[0:0] mux_1344_nl;
  wire[0:0] nor_1377_nl;
  wire[0:0] nor_1378_nl;
  wire[0:0] mux_1343_nl;
  wire[0:0] nor_1379_nl;
  wire[0:0] nor_1380_nl;
  wire[0:0] mux_1342_nl;
  wire[0:0] mux_1341_nl;
  wire[0:0] nor_1381_nl;
  wire[0:0] nor_1382_nl;
  wire[0:0] mux_1340_nl;
  wire[0:0] nor_1383_nl;
  wire[0:0] nor_1384_nl;
  wire[0:0] mux_1400_nl;
  wire[0:0] mux_1399_nl;
  wire[0:0] mux_1398_nl;
  wire[0:0] nor_1332_nl;
  wire[0:0] mux_1397_nl;
  wire[0:0] mux_1396_nl;
  wire[0:0] nor_1333_nl;
  wire[0:0] nor_1334_nl;
  wire[0:0] nor_1335_nl;
  wire[0:0] mux_1395_nl;
  wire[0:0] mux_1394_nl;
  wire[0:0] mux_1393_nl;
  wire[0:0] nor_1336_nl;
  wire[0:0] nor_1337_nl;
  wire[0:0] nor_1338_nl;
  wire[0:0] nor_1339_nl;
  wire[0:0] mux_1392_nl;
  wire[0:0] mux_1391_nl;
  wire[0:0] mux_1390_nl;
  wire[0:0] nor_1340_nl;
  wire[0:0] mux_1389_nl;
  wire[0:0] nor_1341_nl;
  wire[0:0] nor_1342_nl;
  wire[0:0] nor_1343_nl;
  wire[0:0] mux_1388_nl;
  wire[0:0] nor_1344_nl;
  wire[0:0] mux_1387_nl;
  wire[0:0] mux_1386_nl;
  wire[0:0] nor_1345_nl;
  wire[0:0] nor_1346_nl;
  wire[0:0] nor_1347_nl;
  wire[0:0] mux_1385_nl;
  wire[0:0] mux_1384_nl;
  wire[0:0] mux_1383_nl;
  wire[0:0] and_546_nl;
  wire[0:0] mux_1382_nl;
  wire[0:0] nor_1348_nl;
  wire[0:0] nor_1349_nl;
  wire[0:0] nor_1350_nl;
  wire[0:0] mux_1381_nl;
  wire[0:0] or_1173_nl;
  wire[0:0] or_1171_nl;
  wire[0:0] mux_1380_nl;
  wire[0:0] nor_1351_nl;
  wire[0:0] mux_1379_nl;
  wire[0:0] or_1169_nl;
  wire[0:0] or_1167_nl;
  wire[0:0] and_547_nl;
  wire[0:0] mux_1377_nl;
  wire[0:0] nor_1354_nl;
  wire[0:0] mux_1376_nl;
  wire[0:0] mux_1375_nl;
  wire[0:0] or_1163_nl;
  wire[0:0] or_1161_nl;
  wire[0:0] mux_1374_nl;
  wire[0:0] or_1160_nl;
  wire[0:0] or_1158_nl;
  wire[0:0] and_548_nl;
  wire[0:0] mux_1373_nl;
  wire[0:0] mux_1372_nl;
  wire[0:0] nor_1355_nl;
  wire[0:0] nor_1356_nl;
  wire[0:0] mux_1371_nl;
  wire[0:0] nor_1357_nl;
  wire[0:0] nor_1358_nl;
  wire[0:0] nor_1302_nl;
  wire[0:0] mux_1431_nl;
  wire[0:0] mux_1430_nl;
  wire[0:0] and_545_nl;
  wire[0:0] mux_1429_nl;
  wire[0:0] nor_1303_nl;
  wire[0:0] mux_1426_nl;
  wire[0:0] mux_1425_nl;
  wire[0:0] nor_1304_nl;
  wire[0:0] nor_1305_nl;
  wire[0:0] mux_1424_nl;
  wire[0:0] nor_1306_nl;
  wire[0:0] nor_1307_nl;
  wire[0:0] mux_1423_nl;
  wire[0:0] mux_1422_nl;
  wire[0:0] mux_1421_nl;
  wire[0:0] nor_1308_nl;
  wire[0:0] nor_1309_nl;
  wire[0:0] mux_1420_nl;
  wire[0:0] nor_1310_nl;
  wire[0:0] nor_1311_nl;
  wire[0:0] mux_1419_nl;
  wire[0:0] mux_1418_nl;
  wire[0:0] nor_1312_nl;
  wire[0:0] nor_1313_nl;
  wire[0:0] mux_1417_nl;
  wire[0:0] nor_1314_nl;
  wire[0:0] nor_1315_nl;
  wire[0:0] mux_1416_nl;
  wire[0:0] mux_1415_nl;
  wire[0:0] mux_1414_nl;
  wire[0:0] mux_1413_nl;
  wire[0:0] nor_1316_nl;
  wire[0:0] mux_1412_nl;
  wire[0:0] nor_1319_nl;
  wire[0:0] mux_1411_nl;
  wire[0:0] mux_1410_nl;
  wire[0:0] nor_1320_nl;
  wire[0:0] mux_1409_nl;
  wire[0:0] nor_1323_nl;
  wire[0:0] mux_1408_nl;
  wire[0:0] mux_1407_nl;
  wire[0:0] mux_1406_nl;
  wire[0:0] nor_1324_nl;
  wire[0:0] nor_1325_nl;
  wire[0:0] mux_1405_nl;
  wire[0:0] nor_1326_nl;
  wire[0:0] nor_1327_nl;
  wire[0:0] mux_1404_nl;
  wire[0:0] mux_1403_nl;
  wire[0:0] nor_1328_nl;
  wire[0:0] nor_1329_nl;
  wire[0:0] mux_1402_nl;
  wire[0:0] nor_1330_nl;
  wire[0:0] nor_1331_nl;
  wire[0:0] mux_1463_nl;
  wire[0:0] mux_1462_nl;
  wire[0:0] mux_1461_nl;
  wire[0:0] mux_1460_nl;
  wire[0:0] nor_1269_nl;
  wire[0:0] nor_1270_nl;
  wire[0:0] mux_1459_nl;
  wire[0:0] nor_1271_nl;
  wire[0:0] nor_1272_nl;
  wire[0:0] mux_1458_nl;
  wire[0:0] mux_1457_nl;
  wire[0:0] nor_1273_nl;
  wire[0:0] nor_1274_nl;
  wire[0:0] nor_1275_nl;
  wire[0:0] mux_1456_nl;
  wire[0:0] mux_1455_nl;
  wire[0:0] mux_1454_nl;
  wire[0:0] nor_1276_nl;
  wire[0:0] nor_1277_nl;
  wire[0:0] mux_1453_nl;
  wire[0:0] nor_1278_nl;
  wire[0:0] nor_1279_nl;
  wire[0:0] mux_1452_nl;
  wire[0:0] mux_1451_nl;
  wire[0:0] nor_1280_nl;
  wire[0:0] nor_1281_nl;
  wire[0:0] mux_1450_nl;
  wire[0:0] mux_1449_nl;
  wire[0:0] nor_1282_nl;
  wire[0:0] nor_1283_nl;
  wire[0:0] nor_1284_nl;
  wire[0:0] and_542_nl;
  wire[0:0] mux_1448_nl;
  wire[0:0] mux_1447_nl;
  wire[0:0] mux_1446_nl;
  wire[0:0] mux_1445_nl;
  wire[0:0] and_543_nl;
  wire[0:0] mux_1444_nl;
  wire[0:0] nor_1287_nl;
  wire[0:0] nor_1288_nl;
  wire[0:0] mux_1443_nl;
  wire[0:0] mux_1442_nl;
  wire[0:0] and_544_nl;
  wire[0:0] mux_1439_nl;
  wire[0:0] mux_1438_nl;
  wire[0:0] mux_1437_nl;
  wire[0:0] nor_1294_nl;
  wire[0:0] nor_1295_nl;
  wire[0:0] mux_1436_nl;
  wire[0:0] nor_1296_nl;
  wire[0:0] nor_1297_nl;
  wire[0:0] mux_1435_nl;
  wire[0:0] mux_1434_nl;
  wire[0:0] nor_1298_nl;
  wire[0:0] nor_1299_nl;
  wire[0:0] mux_1433_nl;
  wire[0:0] nor_1300_nl;
  wire[0:0] nor_1301_nl;
  wire[0:0] nor_1240_nl;
  wire[0:0] mux_1494_nl;
  wire[0:0] mux_1493_nl;
  wire[0:0] nor_1241_nl;
  wire[0:0] mux_1492_nl;
  wire[0:0] nand_47_nl;
  wire[0:0] mux_1489_nl;
  wire[0:0] mux_1488_nl;
  wire[0:0] or_1340_nl;
  wire[0:0] or_1338_nl;
  wire[0:0] mux_1487_nl;
  wire[0:0] or_1336_nl;
  wire[0:0] or_1335_nl;
  wire[0:0] mux_1486_nl;
  wire[0:0] mux_1485_nl;
  wire[0:0] mux_1484_nl;
  wire[0:0] nor_1245_nl;
  wire[0:0] nor_1246_nl;
  wire[0:0] mux_1483_nl;
  wire[0:0] nor_1247_nl;
  wire[0:0] nor_1248_nl;
  wire[0:0] mux_1482_nl;
  wire[0:0] mux_1481_nl;
  wire[0:0] nor_1249_nl;
  wire[0:0] nor_1250_nl;
  wire[0:0] mux_1480_nl;
  wire[0:0] nor_1251_nl;
  wire[0:0] nor_1252_nl;
  wire[0:0] mux_1479_nl;
  wire[0:0] mux_1478_nl;
  wire[0:0] mux_1477_nl;
  wire[0:0] mux_1476_nl;
  wire[0:0] nor_1253_nl;
  wire[0:0] nor_1254_nl;
  wire[0:0] mux_1475_nl;
  wire[0:0] nor_1255_nl;
  wire[0:0] nor_1256_nl;
  wire[0:0] mux_1474_nl;
  wire[0:0] mux_1473_nl;
  wire[0:0] nor_1257_nl;
  wire[0:0] nor_1258_nl;
  wire[0:0] mux_1472_nl;
  wire[0:0] nor_1259_nl;
  wire[0:0] nor_1260_nl;
  wire[0:0] mux_1471_nl;
  wire[0:0] mux_1470_nl;
  wire[0:0] mux_1469_nl;
  wire[0:0] nor_1261_nl;
  wire[0:0] nor_1262_nl;
  wire[0:0] mux_1468_nl;
  wire[0:0] nor_1263_nl;
  wire[0:0] nor_1264_nl;
  wire[0:0] mux_1467_nl;
  wire[0:0] mux_1466_nl;
  wire[0:0] nor_1265_nl;
  wire[0:0] nor_1266_nl;
  wire[0:0] mux_1465_nl;
  wire[0:0] nor_1267_nl;
  wire[0:0] nor_1268_nl;
  wire[0:0] mux_1525_nl;
  wire[0:0] mux_1524_nl;
  wire[0:0] mux_1523_nl;
  wire[0:0] nor_1213_nl;
  wire[0:0] mux_1522_nl;
  wire[0:0] mux_1521_nl;
  wire[0:0] nor_1214_nl;
  wire[0:0] nor_1215_nl;
  wire[0:0] nor_1216_nl;
  wire[0:0] mux_1520_nl;
  wire[0:0] mux_1519_nl;
  wire[0:0] mux_1518_nl;
  wire[0:0] nor_1217_nl;
  wire[0:0] nor_1218_nl;
  wire[0:0] nor_1219_nl;
  wire[0:0] nor_1220_nl;
  wire[0:0] mux_1517_nl;
  wire[0:0] mux_1516_nl;
  wire[0:0] mux_1515_nl;
  wire[0:0] nor_1221_nl;
  wire[0:0] mux_1514_nl;
  wire[0:0] nor_1222_nl;
  wire[0:0] nor_1223_nl;
  wire[0:0] nor_1224_nl;
  wire[0:0] mux_1513_nl;
  wire[0:0] nor_1225_nl;
  wire[0:0] mux_1512_nl;
  wire[0:0] mux_1511_nl;
  wire[0:0] nor_1226_nl;
  wire[0:0] nor_1227_nl;
  wire[0:0] nor_1228_nl;
  wire[0:0] mux_1510_nl;
  wire[0:0] mux_1509_nl;
  wire[0:0] mux_1508_nl;
  wire[0:0] and_539_nl;
  wire[0:0] mux_1507_nl;
  wire[0:0] nor_1229_nl;
  wire[0:0] nor_1230_nl;
  wire[0:0] nor_1231_nl;
  wire[0:0] mux_1506_nl;
  wire[0:0] or_1367_nl;
  wire[0:0] or_1365_nl;
  wire[0:0] mux_1505_nl;
  wire[0:0] nor_1232_nl;
  wire[0:0] mux_1504_nl;
  wire[0:0] or_1363_nl;
  wire[0:0] or_1361_nl;
  wire[0:0] and_540_nl;
  wire[0:0] mux_1502_nl;
  wire[0:0] nor_1235_nl;
  wire[0:0] mux_1501_nl;
  wire[0:0] mux_1500_nl;
  wire[0:0] or_1357_nl;
  wire[0:0] or_1355_nl;
  wire[0:0] mux_1499_nl;
  wire[0:0] or_1354_nl;
  wire[0:0] or_1352_nl;
  wire[0:0] and_541_nl;
  wire[0:0] mux_1498_nl;
  wire[0:0] mux_1497_nl;
  wire[0:0] nor_1236_nl;
  wire[0:0] nor_1237_nl;
  wire[0:0] mux_1496_nl;
  wire[0:0] nor_1238_nl;
  wire[0:0] nor_1239_nl;
  wire[0:0] nor_1184_nl;
  wire[0:0] mux_1556_nl;
  wire[0:0] mux_1555_nl;
  wire[0:0] and_534_nl;
  wire[0:0] mux_1554_nl;
  wire[0:0] and_535_nl;
  wire[0:0] mux_1551_nl;
  wire[0:0] mux_1550_nl;
  wire[0:0] nor_1188_nl;
  wire[0:0] nor_1189_nl;
  wire[0:0] mux_1549_nl;
  wire[0:0] nor_1190_nl;
  wire[0:0] nor_1191_nl;
  wire[0:0] mux_1548_nl;
  wire[0:0] mux_1547_nl;
  wire[0:0] mux_1546_nl;
  wire[0:0] nor_1192_nl;
  wire[0:0] nor_1193_nl;
  wire[0:0] mux_1545_nl;
  wire[0:0] and_536_nl;
  wire[0:0] nor_1194_nl;
  wire[0:0] mux_1544_nl;
  wire[0:0] mux_1543_nl;
  wire[0:0] and_842_nl;
  wire[0:0] nor_1196_nl;
  wire[0:0] mux_1542_nl;
  wire[0:0] nor_1197_nl;
  wire[0:0] nor_1198_nl;
  wire[0:0] mux_1541_nl;
  wire[0:0] mux_1540_nl;
  wire[0:0] mux_1539_nl;
  wire[0:0] mux_1538_nl;
  wire[0:0] nor_1199_nl;
  wire[0:0] mux_1537_nl;
  wire[0:0] nor_1201_nl;
  wire[0:0] mux_1536_nl;
  wire[0:0] mux_1535_nl;
  wire[0:0] and_853_nl;
  wire[0:0] mux_1534_nl;
  wire[0:0] nor_1205_nl;
  wire[0:0] mux_1533_nl;
  wire[0:0] mux_1532_nl;
  wire[0:0] mux_1531_nl;
  wire[0:0] nor_1206_nl;
  wire[0:0] nor_1207_nl;
  wire[0:0] mux_1530_nl;
  wire[0:0] and_538_nl;
  wire[0:0] nor_1208_nl;
  wire[0:0] mux_1529_nl;
  wire[0:0] mux_1528_nl;
  wire[0:0] and_872_nl;
  wire[0:0] nor_1210_nl;
  wire[0:0] mux_1527_nl;
  wire[0:0] nor_1211_nl;
  wire[0:0] nor_1212_nl;
  wire[0:0] mux_1588_nl;
  wire[0:0] mux_1587_nl;
  wire[0:0] mux_1586_nl;
  wire[0:0] mux_1585_nl;
  wire[0:0] nor_1154_nl;
  wire[0:0] nor_1155_nl;
  wire[0:0] mux_1584_nl;
  wire[0:0] nor_1156_nl;
  wire[0:0] nor_1157_nl;
  wire[0:0] mux_1583_nl;
  wire[0:0] mux_1582_nl;
  wire[0:0] nor_1158_nl;
  wire[0:0] nor_1159_nl;
  wire[0:0] nor_1160_nl;
  wire[0:0] mux_1581_nl;
  wire[0:0] mux_1580_nl;
  wire[0:0] mux_1579_nl;
  wire[0:0] nor_1161_nl;
  wire[0:0] and_852_nl;
  wire[0:0] mux_1578_nl;
  wire[0:0] and_858_nl;
  wire[0:0] nor_1164_nl;
  wire[0:0] mux_1577_nl;
  wire[0:0] mux_1576_nl;
  wire[0:0] and_870_nl;
  wire[0:0] and_871_nl;
  wire[0:0] mux_1575_nl;
  wire[0:0] mux_1574_nl;
  wire[0:0] nor_1167_nl;
  wire[0:0] nor_1168_nl;
  wire[0:0] nor_1169_nl;
  wire[0:0] and_528_nl;
  wire[0:0] mux_1573_nl;
  wire[0:0] mux_1572_nl;
  wire[0:0] mux_1571_nl;
  wire[0:0] mux_1570_nl;
  wire[0:0] and_530_nl;
  wire[0:0] mux_1569_nl;
  wire[0:0] nor_1171_nl;
  wire[0:0] nor_1172_nl;
  wire[0:0] mux_1568_nl;
  wire[0:0] mux_1567_nl;
  wire[0:0] and_531_nl;
  wire[0:0] mux_1564_nl;
  wire[0:0] mux_1563_nl;
  wire[0:0] mux_1562_nl;
  wire[0:0] nor_1178_nl;
  wire[0:0] nor_1179_nl;
  wire[0:0] mux_1561_nl;
  wire[0:0] nor_1180_nl;
  wire[0:0] nor_1181_nl;
  wire[0:0] mux_1560_nl;
  wire[0:0] mux_1559_nl;
  wire[0:0] and_532_nl;
  wire[0:0] nor_1182_nl;
  wire[0:0] mux_1558_nl;
  wire[0:0] and_533_nl;
  wire[0:0] nor_1183_nl;
  wire[0:0] nor_1128_nl;
  wire[0:0] mux_1619_nl;
  wire[0:0] mux_1618_nl;
  wire[0:0] nor_1129_nl;
  wire[0:0] mux_1617_nl;
  wire[0:0] or_1539_nl;
  wire[0:0] mux_1614_nl;
  wire[0:0] mux_1613_nl;
  wire[0:0] or_1533_nl;
  wire[0:0] or_1531_nl;
  wire[0:0] mux_1612_nl;
  wire[0:0] or_1529_nl;
  wire[0:0] or_1528_nl;
  wire[0:0] mux_1611_nl;
  wire[0:0] mux_1610_nl;
  wire[0:0] mux_1609_nl;
  wire[0:0] nor_1130_nl;
  wire[0:0] nor_1131_nl;
  wire[0:0] mux_1608_nl;
  wire[0:0] nor_1132_nl;
  wire[0:0] nor_1133_nl;
  wire[0:0] mux_1607_nl;
  wire[0:0] mux_1606_nl;
  wire[0:0] nor_1134_nl;
  wire[0:0] nor_1135_nl;
  wire[0:0] mux_1605_nl;
  wire[0:0] nor_1136_nl;
  wire[0:0] nor_1137_nl;
  wire[0:0] mux_1604_nl;
  wire[0:0] mux_1603_nl;
  wire[0:0] mux_1602_nl;
  wire[0:0] mux_1601_nl;
  wire[0:0] nor_1138_nl;
  wire[0:0] nor_1139_nl;
  wire[0:0] mux_1600_nl;
  wire[0:0] nor_1140_nl;
  wire[0:0] nor_1141_nl;
  wire[0:0] mux_1599_nl;
  wire[0:0] mux_1598_nl;
  wire[0:0] nor_1142_nl;
  wire[0:0] nor_1143_nl;
  wire[0:0] mux_1597_nl;
  wire[0:0] nor_1144_nl;
  wire[0:0] nor_1145_nl;
  wire[0:0] mux_1596_nl;
  wire[0:0] mux_1595_nl;
  wire[0:0] mux_1594_nl;
  wire[0:0] nor_1146_nl;
  wire[0:0] nor_1147_nl;
  wire[0:0] mux_1593_nl;
  wire[0:0] nor_1148_nl;
  wire[0:0] nor_1149_nl;
  wire[0:0] mux_1592_nl;
  wire[0:0] mux_1591_nl;
  wire[0:0] nor_1150_nl;
  wire[0:0] nor_1151_nl;
  wire[0:0] mux_1590_nl;
  wire[0:0] nor_1152_nl;
  wire[0:0] nor_1153_nl;
  wire[0:0] mux_1650_nl;
  wire[0:0] mux_1649_nl;
  wire[0:0] mux_1648_nl;
  wire[0:0] nor_1101_nl;
  wire[0:0] mux_1647_nl;
  wire[0:0] mux_1646_nl;
  wire[0:0] nor_1102_nl;
  wire[0:0] nor_1103_nl;
  wire[0:0] nor_1104_nl;
  wire[0:0] mux_1645_nl;
  wire[0:0] mux_1644_nl;
  wire[0:0] mux_1643_nl;
  wire[0:0] nor_1105_nl;
  wire[0:0] nor_1106_nl;
  wire[0:0] nor_1107_nl;
  wire[0:0] nor_1108_nl;
  wire[0:0] mux_1642_nl;
  wire[0:0] mux_1641_nl;
  wire[0:0] mux_1640_nl;
  wire[0:0] nor_1109_nl;
  wire[0:0] mux_1639_nl;
  wire[0:0] nor_1110_nl;
  wire[0:0] nor_1111_nl;
  wire[0:0] nor_1112_nl;
  wire[0:0] mux_1638_nl;
  wire[0:0] nor_1113_nl;
  wire[0:0] mux_1637_nl;
  wire[0:0] mux_1636_nl;
  wire[0:0] nor_1114_nl;
  wire[0:0] nor_1115_nl;
  wire[0:0] nor_1116_nl;
  wire[0:0] mux_1635_nl;
  wire[0:0] mux_1634_nl;
  wire[0:0] mux_1633_nl;
  wire[0:0] and_525_nl;
  wire[0:0] mux_1632_nl;
  wire[0:0] nor_1117_nl;
  wire[0:0] nor_1118_nl;
  wire[0:0] nor_1119_nl;
  wire[0:0] mux_1631_nl;
  wire[0:0] or_1561_nl;
  wire[0:0] or_1559_nl;
  wire[0:0] mux_1630_nl;
  wire[0:0] nor_1120_nl;
  wire[0:0] mux_1629_nl;
  wire[0:0] or_1557_nl;
  wire[0:0] or_1555_nl;
  wire[0:0] and_526_nl;
  wire[0:0] mux_1627_nl;
  wire[0:0] nor_1123_nl;
  wire[0:0] mux_1626_nl;
  wire[0:0] mux_1625_nl;
  wire[0:0] or_1551_nl;
  wire[0:0] or_1549_nl;
  wire[0:0] mux_1624_nl;
  wire[0:0] or_1548_nl;
  wire[0:0] or_1546_nl;
  wire[0:0] and_527_nl;
  wire[0:0] mux_1623_nl;
  wire[0:0] mux_1622_nl;
  wire[0:0] nor_1124_nl;
  wire[0:0] nor_1125_nl;
  wire[0:0] mux_1621_nl;
  wire[0:0] nor_1126_nl;
  wire[0:0] nor_1127_nl;
  wire[0:0] nor_1071_nl;
  wire[0:0] mux_1681_nl;
  wire[0:0] mux_1680_nl;
  wire[0:0] and_524_nl;
  wire[0:0] mux_1679_nl;
  wire[0:0] nor_1072_nl;
  wire[0:0] mux_1676_nl;
  wire[0:0] mux_1675_nl;
  wire[0:0] nor_1073_nl;
  wire[0:0] nor_1074_nl;
  wire[0:0] mux_1674_nl;
  wire[0:0] nor_1075_nl;
  wire[0:0] nor_1076_nl;
  wire[0:0] mux_1673_nl;
  wire[0:0] mux_1672_nl;
  wire[0:0] mux_1671_nl;
  wire[0:0] nor_1077_nl;
  wire[0:0] nor_1078_nl;
  wire[0:0] mux_1670_nl;
  wire[0:0] nor_1079_nl;
  wire[0:0] nor_1080_nl;
  wire[0:0] mux_1669_nl;
  wire[0:0] mux_1668_nl;
  wire[0:0] nor_1081_nl;
  wire[0:0] nor_1082_nl;
  wire[0:0] mux_1667_nl;
  wire[0:0] nor_1083_nl;
  wire[0:0] nor_1084_nl;
  wire[0:0] mux_1666_nl;
  wire[0:0] mux_1665_nl;
  wire[0:0] mux_1664_nl;
  wire[0:0] mux_1663_nl;
  wire[0:0] nor_1085_nl;
  wire[0:0] mux_1662_nl;
  wire[0:0] nor_1088_nl;
  wire[0:0] mux_1661_nl;
  wire[0:0] mux_1660_nl;
  wire[0:0] nor_1089_nl;
  wire[0:0] mux_1659_nl;
  wire[0:0] nor_1092_nl;
  wire[0:0] mux_1658_nl;
  wire[0:0] mux_1657_nl;
  wire[0:0] mux_1656_nl;
  wire[0:0] nor_1093_nl;
  wire[0:0] nor_1094_nl;
  wire[0:0] mux_1655_nl;
  wire[0:0] nor_1095_nl;
  wire[0:0] nor_1096_nl;
  wire[0:0] mux_1654_nl;
  wire[0:0] mux_1653_nl;
  wire[0:0] nor_1097_nl;
  wire[0:0] nor_1098_nl;
  wire[0:0] mux_1652_nl;
  wire[0:0] nor_1099_nl;
  wire[0:0] nor_1100_nl;
  wire[0:0] mux_1713_nl;
  wire[0:0] mux_1712_nl;
  wire[0:0] mux_1711_nl;
  wire[0:0] mux_1710_nl;
  wire[0:0] nor_1039_nl;
  wire[0:0] nor_1040_nl;
  wire[0:0] mux_1709_nl;
  wire[0:0] nor_1041_nl;
  wire[0:0] nor_1042_nl;
  wire[0:0] mux_1708_nl;
  wire[0:0] mux_1707_nl;
  wire[0:0] nor_1043_nl;
  wire[0:0] nor_1044_nl;
  wire[0:0] nor_1045_nl;
  wire[0:0] mux_1706_nl;
  wire[0:0] mux_1705_nl;
  wire[0:0] mux_1704_nl;
  wire[0:0] nor_1046_nl;
  wire[0:0] nor_1047_nl;
  wire[0:0] mux_1703_nl;
  wire[0:0] nor_1048_nl;
  wire[0:0] nor_1049_nl;
  wire[0:0] mux_1702_nl;
  wire[0:0] mux_1701_nl;
  wire[0:0] nor_1050_nl;
  wire[0:0] nor_1051_nl;
  wire[0:0] mux_1700_nl;
  wire[0:0] mux_1699_nl;
  wire[0:0] nor_1052_nl;
  wire[0:0] nor_1053_nl;
  wire[0:0] nor_1054_nl;
  wire[0:0] and_520_nl;
  wire[0:0] mux_1698_nl;
  wire[0:0] mux_1697_nl;
  wire[0:0] mux_1696_nl;
  wire[0:0] mux_1695_nl;
  wire[0:0] and_521_nl;
  wire[0:0] mux_1694_nl;
  wire[0:0] nor_1057_nl;
  wire[0:0] nor_1058_nl;
  wire[0:0] mux_1693_nl;
  wire[0:0] mux_1692_nl;
  wire[0:0] and_522_nl;
  wire[0:0] mux_1689_nl;
  wire[0:0] mux_1688_nl;
  wire[0:0] mux_1687_nl;
  wire[0:0] nor_1063_nl;
  wire[0:0] nor_1064_nl;
  wire[0:0] mux_1686_nl;
  wire[0:0] nor_1065_nl;
  wire[0:0] nor_1066_nl;
  wire[0:0] mux_1685_nl;
  wire[0:0] mux_1684_nl;
  wire[0:0] nor_1067_nl;
  wire[0:0] nor_1068_nl;
  wire[0:0] mux_1683_nl;
  wire[0:0] nor_1069_nl;
  wire[0:0] nor_1070_nl;
  wire[0:0] nor_1010_nl;
  wire[0:0] mux_1744_nl;
  wire[0:0] mux_1743_nl;
  wire[0:0] nor_1011_nl;
  wire[0:0] mux_1742_nl;
  wire[0:0] nand_63_nl;
  wire[0:0] mux_1739_nl;
  wire[0:0] mux_1738_nl;
  wire[0:0] or_1728_nl;
  wire[0:0] or_1726_nl;
  wire[0:0] mux_1737_nl;
  wire[0:0] or_1724_nl;
  wire[0:0] or_1723_nl;
  wire[0:0] mux_1736_nl;
  wire[0:0] mux_1735_nl;
  wire[0:0] mux_1734_nl;
  wire[0:0] nor_1015_nl;
  wire[0:0] nor_1016_nl;
  wire[0:0] mux_1733_nl;
  wire[0:0] nor_1017_nl;
  wire[0:0] nor_1018_nl;
  wire[0:0] mux_1732_nl;
  wire[0:0] mux_1731_nl;
  wire[0:0] nor_1019_nl;
  wire[0:0] nor_1020_nl;
  wire[0:0] mux_1730_nl;
  wire[0:0] nor_1021_nl;
  wire[0:0] nor_1022_nl;
  wire[0:0] mux_1729_nl;
  wire[0:0] mux_1728_nl;
  wire[0:0] mux_1727_nl;
  wire[0:0] mux_1726_nl;
  wire[0:0] nor_1023_nl;
  wire[0:0] nor_1024_nl;
  wire[0:0] mux_1725_nl;
  wire[0:0] nor_1025_nl;
  wire[0:0] nor_1026_nl;
  wire[0:0] mux_1724_nl;
  wire[0:0] mux_1723_nl;
  wire[0:0] nor_1027_nl;
  wire[0:0] nor_1028_nl;
  wire[0:0] mux_1722_nl;
  wire[0:0] nor_1029_nl;
  wire[0:0] nor_1030_nl;
  wire[0:0] mux_1721_nl;
  wire[0:0] mux_1720_nl;
  wire[0:0] mux_1719_nl;
  wire[0:0] nor_1031_nl;
  wire[0:0] nor_1032_nl;
  wire[0:0] mux_1718_nl;
  wire[0:0] nor_1033_nl;
  wire[0:0] nor_1034_nl;
  wire[0:0] mux_1717_nl;
  wire[0:0] mux_1716_nl;
  wire[0:0] nor_1035_nl;
  wire[0:0] nor_1036_nl;
  wire[0:0] mux_1715_nl;
  wire[0:0] nor_1037_nl;
  wire[0:0] nor_1038_nl;
  wire[0:0] mux_1775_nl;
  wire[0:0] mux_1774_nl;
  wire[0:0] mux_1773_nl;
  wire[0:0] nor_983_nl;
  wire[0:0] mux_1772_nl;
  wire[0:0] mux_1771_nl;
  wire[0:0] nor_984_nl;
  wire[0:0] nor_985_nl;
  wire[0:0] nor_986_nl;
  wire[0:0] mux_1770_nl;
  wire[0:0] mux_1769_nl;
  wire[0:0] mux_1768_nl;
  wire[0:0] nor_987_nl;
  wire[0:0] nor_988_nl;
  wire[0:0] nor_989_nl;
  wire[0:0] nor_990_nl;
  wire[0:0] mux_1767_nl;
  wire[0:0] mux_1766_nl;
  wire[0:0] mux_1765_nl;
  wire[0:0] nor_991_nl;
  wire[0:0] mux_1764_nl;
  wire[0:0] nor_992_nl;
  wire[0:0] nor_993_nl;
  wire[0:0] nor_994_nl;
  wire[0:0] mux_1763_nl;
  wire[0:0] nor_995_nl;
  wire[0:0] mux_1762_nl;
  wire[0:0] mux_1761_nl;
  wire[0:0] nor_996_nl;
  wire[0:0] nor_997_nl;
  wire[0:0] nor_998_nl;
  wire[0:0] mux_1760_nl;
  wire[0:0] mux_1759_nl;
  wire[0:0] mux_1758_nl;
  wire[0:0] and_517_nl;
  wire[0:0] mux_1757_nl;
  wire[0:0] nor_999_nl;
  wire[0:0] nor_1000_nl;
  wire[0:0] nor_1001_nl;
  wire[0:0] mux_1756_nl;
  wire[0:0] or_1755_nl;
  wire[0:0] or_1753_nl;
  wire[0:0] mux_1755_nl;
  wire[0:0] nor_1002_nl;
  wire[0:0] mux_1754_nl;
  wire[0:0] or_1751_nl;
  wire[0:0] or_1749_nl;
  wire[0:0] and_518_nl;
  wire[0:0] mux_1752_nl;
  wire[0:0] nor_1005_nl;
  wire[0:0] mux_1751_nl;
  wire[0:0] mux_1750_nl;
  wire[0:0] or_1745_nl;
  wire[0:0] or_1743_nl;
  wire[0:0] mux_1749_nl;
  wire[0:0] or_1742_nl;
  wire[0:0] or_1740_nl;
  wire[0:0] and_519_nl;
  wire[0:0] mux_1748_nl;
  wire[0:0] mux_1747_nl;
  wire[0:0] nor_1006_nl;
  wire[0:0] nor_1007_nl;
  wire[0:0] mux_1746_nl;
  wire[0:0] nor_1008_nl;
  wire[0:0] nor_1009_nl;
  wire[0:0] nor_954_nl;
  wire[0:0] mux_1806_nl;
  wire[0:0] mux_1805_nl;
  wire[0:0] and_512_nl;
  wire[0:0] mux_1804_nl;
  wire[0:0] and_513_nl;
  wire[0:0] mux_1801_nl;
  wire[0:0] mux_1800_nl;
  wire[0:0] nor_958_nl;
  wire[0:0] nor_959_nl;
  wire[0:0] mux_1799_nl;
  wire[0:0] nor_960_nl;
  wire[0:0] nor_961_nl;
  wire[0:0] mux_1798_nl;
  wire[0:0] mux_1797_nl;
  wire[0:0] mux_1796_nl;
  wire[0:0] nor_962_nl;
  wire[0:0] nor_963_nl;
  wire[0:0] mux_1795_nl;
  wire[0:0] and_514_nl;
  wire[0:0] nor_964_nl;
  wire[0:0] mux_1794_nl;
  wire[0:0] mux_1793_nl;
  wire[0:0] and_841_nl;
  wire[0:0] nor_966_nl;
  wire[0:0] mux_1792_nl;
  wire[0:0] nor_967_nl;
  wire[0:0] nor_968_nl;
  wire[0:0] mux_1791_nl;
  wire[0:0] mux_1790_nl;
  wire[0:0] mux_1789_nl;
  wire[0:0] mux_1788_nl;
  wire[0:0] nor_969_nl;
  wire[0:0] mux_1787_nl;
  wire[0:0] nor_971_nl;
  wire[0:0] mux_1786_nl;
  wire[0:0] mux_1785_nl;
  wire[0:0] and_851_nl;
  wire[0:0] mux_1784_nl;
  wire[0:0] nor_975_nl;
  wire[0:0] mux_1783_nl;
  wire[0:0] mux_1782_nl;
  wire[0:0] mux_1781_nl;
  wire[0:0] nor_976_nl;
  wire[0:0] nor_977_nl;
  wire[0:0] mux_1780_nl;
  wire[0:0] and_516_nl;
  wire[0:0] nor_978_nl;
  wire[0:0] mux_1779_nl;
  wire[0:0] mux_1778_nl;
  wire[0:0] and_869_nl;
  wire[0:0] nor_980_nl;
  wire[0:0] mux_1777_nl;
  wire[0:0] nor_981_nl;
  wire[0:0] nor_982_nl;
  wire[0:0] mux_1838_nl;
  wire[0:0] mux_1837_nl;
  wire[0:0] mux_1836_nl;
  wire[0:0] mux_1835_nl;
  wire[0:0] nor_925_nl;
  wire[0:0] nor_926_nl;
  wire[0:0] mux_1834_nl;
  wire[0:0] nor_927_nl;
  wire[0:0] nor_928_nl;
  wire[0:0] mux_1833_nl;
  wire[0:0] mux_1832_nl;
  wire[0:0] nor_929_nl;
  wire[0:0] nor_930_nl;
  wire[0:0] nor_931_nl;
  wire[0:0] mux_1831_nl;
  wire[0:0] mux_1830_nl;
  wire[0:0] mux_1829_nl;
  wire[0:0] nor_932_nl;
  wire[0:0] and_850_nl;
  wire[0:0] mux_1828_nl;
  wire[0:0] and_857_nl;
  wire[0:0] nor_935_nl;
  wire[0:0] mux_1827_nl;
  wire[0:0] mux_1826_nl;
  wire[0:0] and_867_nl;
  wire[0:0] and_868_nl;
  wire[0:0] mux_1825_nl;
  wire[0:0] mux_1824_nl;
  wire[0:0] nor_938_nl;
  wire[0:0] nor_939_nl;
  wire[0:0] nor_940_nl;
  wire[0:0] and_505_nl;
  wire[0:0] mux_1823_nl;
  wire[0:0] mux_1822_nl;
  wire[0:0] mux_1821_nl;
  wire[0:0] mux_1820_nl;
  wire[0:0] and_507_nl;
  wire[0:0] mux_1819_nl;
  wire[0:0] nor_942_nl;
  wire[0:0] nor_943_nl;
  wire[0:0] mux_1818_nl;
  wire[0:0] mux_1817_nl;
  wire[0:0] and_508_nl;
  wire[0:0] mux_1814_nl;
  wire[0:0] mux_1813_nl;
  wire[0:0] mux_1812_nl;
  wire[0:0] nor_948_nl;
  wire[0:0] nor_949_nl;
  wire[0:0] mux_1811_nl;
  wire[0:0] nor_950_nl;
  wire[0:0] nor_951_nl;
  wire[0:0] mux_1810_nl;
  wire[0:0] mux_1809_nl;
  wire[0:0] and_510_nl;
  wire[0:0] nor_952_nl;
  wire[0:0] mux_1808_nl;
  wire[0:0] and_511_nl;
  wire[0:0] nor_953_nl;
  wire[0:0] nor_899_nl;
  wire[0:0] mux_1869_nl;
  wire[0:0] mux_1868_nl;
  wire[0:0] nor_900_nl;
  wire[0:0] mux_1867_nl;
  wire[0:0] or_1925_nl;
  wire[0:0] mux_1864_nl;
  wire[0:0] mux_1863_nl;
  wire[0:0] or_1919_nl;
  wire[0:0] or_1918_nl;
  wire[0:0] mux_1862_nl;
  wire[0:0] or_1916_nl;
  wire[0:0] or_1915_nl;
  wire[0:0] mux_1861_nl;
  wire[0:0] mux_1860_nl;
  wire[0:0] mux_1859_nl;
  wire[0:0] nor_901_nl;
  wire[0:0] nor_902_nl;
  wire[0:0] mux_1858_nl;
  wire[0:0] nor_903_nl;
  wire[0:0] nor_904_nl;
  wire[0:0] mux_1857_nl;
  wire[0:0] mux_1856_nl;
  wire[0:0] nor_905_nl;
  wire[0:0] nor_906_nl;
  wire[0:0] mux_1855_nl;
  wire[0:0] nor_907_nl;
  wire[0:0] nor_908_nl;
  wire[0:0] mux_1854_nl;
  wire[0:0] mux_1853_nl;
  wire[0:0] mux_1852_nl;
  wire[0:0] mux_1851_nl;
  wire[0:0] nor_909_nl;
  wire[0:0] nor_910_nl;
  wire[0:0] mux_1850_nl;
  wire[0:0] nor_911_nl;
  wire[0:0] nor_912_nl;
  wire[0:0] mux_1849_nl;
  wire[0:0] mux_1848_nl;
  wire[0:0] nor_913_nl;
  wire[0:0] nor_914_nl;
  wire[0:0] mux_1847_nl;
  wire[0:0] nor_915_nl;
  wire[0:0] nor_916_nl;
  wire[0:0] mux_1846_nl;
  wire[0:0] mux_1845_nl;
  wire[0:0] mux_1844_nl;
  wire[0:0] nor_917_nl;
  wire[0:0] nor_918_nl;
  wire[0:0] mux_1843_nl;
  wire[0:0] nor_919_nl;
  wire[0:0] nor_920_nl;
  wire[0:0] mux_1842_nl;
  wire[0:0] mux_1841_nl;
  wire[0:0] nor_921_nl;
  wire[0:0] nor_922_nl;
  wire[0:0] mux_1840_nl;
  wire[0:0] nor_923_nl;
  wire[0:0] nor_924_nl;
  wire[0:0] mux_1900_nl;
  wire[0:0] mux_1899_nl;
  wire[0:0] mux_1898_nl;
  wire[0:0] nor_873_nl;
  wire[0:0] mux_1897_nl;
  wire[0:0] mux_1896_nl;
  wire[0:0] nor_874_nl;
  wire[0:0] nor_875_nl;
  wire[0:0] nor_876_nl;
  wire[0:0] mux_1895_nl;
  wire[0:0] mux_1894_nl;
  wire[0:0] mux_1893_nl;
  wire[0:0] nor_877_nl;
  wire[0:0] nor_878_nl;
  wire[0:0] nor_879_nl;
  wire[0:0] nor_880_nl;
  wire[0:0] mux_1892_nl;
  wire[0:0] mux_1891_nl;
  wire[0:0] mux_1890_nl;
  wire[0:0] nor_881_nl;
  wire[0:0] mux_1889_nl;
  wire[0:0] nor_882_nl;
  wire[0:0] nor_883_nl;
  wire[0:0] nor_884_nl;
  wire[0:0] mux_1888_nl;
  wire[0:0] nor_885_nl;
  wire[0:0] mux_1887_nl;
  wire[0:0] mux_1886_nl;
  wire[0:0] nor_886_nl;
  wire[0:0] nor_887_nl;
  wire[0:0] nor_888_nl;
  wire[0:0] mux_1885_nl;
  wire[0:0] mux_1884_nl;
  wire[0:0] mux_1883_nl;
  wire[0:0] and_501_nl;
  wire[0:0] mux_1882_nl;
  wire[0:0] nor_889_nl;
  wire[0:0] nor_890_nl;
  wire[0:0] nor_891_nl;
  wire[0:0] mux_1881_nl;
  wire[0:0] or_1947_nl;
  wire[0:0] or_1945_nl;
  wire[0:0] mux_1880_nl;
  wire[0:0] nor_892_nl;
  wire[0:0] mux_1879_nl;
  wire[0:0] or_1943_nl;
  wire[0:0] or_1941_nl;
  wire[0:0] and_502_nl;
  wire[0:0] mux_1877_nl;
  wire[0:0] nor_894_nl;
  wire[0:0] mux_1876_nl;
  wire[0:0] mux_1875_nl;
  wire[0:0] or_1937_nl;
  wire[0:0] or_1935_nl;
  wire[0:0] mux_1874_nl;
  wire[0:0] or_1934_nl;
  wire[0:0] or_1932_nl;
  wire[0:0] and_504_nl;
  wire[0:0] mux_1873_nl;
  wire[0:0] mux_1872_nl;
  wire[0:0] nor_895_nl;
  wire[0:0] nor_896_nl;
  wire[0:0] mux_1871_nl;
  wire[0:0] nor_897_nl;
  wire[0:0] nor_898_nl;
  wire[0:0] nor_846_nl;
  wire[0:0] mux_1931_nl;
  wire[0:0] mux_1930_nl;
  wire[0:0] and_497_nl;
  wire[0:0] mux_1929_nl;
  wire[0:0] nor_847_nl;
  wire[0:0] mux_1926_nl;
  wire[0:0] mux_1925_nl;
  wire[0:0] nor_848_nl;
  wire[0:0] nor_849_nl;
  wire[0:0] mux_1924_nl;
  wire[0:0] nor_850_nl;
  wire[0:0] nor_851_nl;
  wire[0:0] mux_1923_nl;
  wire[0:0] mux_1922_nl;
  wire[0:0] mux_1921_nl;
  wire[0:0] nor_852_nl;
  wire[0:0] nor_853_nl;
  wire[0:0] mux_1920_nl;
  wire[0:0] and_498_nl;
  wire[0:0] nor_854_nl;
  wire[0:0] mux_1919_nl;
  wire[0:0] mux_1918_nl;
  wire[0:0] and_840_nl;
  wire[0:0] nor_856_nl;
  wire[0:0] mux_1917_nl;
  wire[0:0] nor_857_nl;
  wire[0:0] nor_858_nl;
  wire[0:0] mux_1916_nl;
  wire[0:0] mux_1915_nl;
  wire[0:0] mux_1914_nl;
  wire[0:0] mux_1913_nl;
  wire[0:0] nor_859_nl;
  wire[0:0] mux_1912_nl;
  wire[0:0] nor_861_nl;
  wire[0:0] mux_1911_nl;
  wire[0:0] mux_1910_nl;
  wire[0:0] and_849_nl;
  wire[0:0] mux_1909_nl;
  wire[0:0] nor_865_nl;
  wire[0:0] mux_1908_nl;
  wire[0:0] mux_1907_nl;
  wire[0:0] mux_1906_nl;
  wire[0:0] nor_866_nl;
  wire[0:0] nor_867_nl;
  wire[0:0] mux_1905_nl;
  wire[0:0] and_500_nl;
  wire[0:0] nor_868_nl;
  wire[0:0] mux_1904_nl;
  wire[0:0] mux_1903_nl;
  wire[0:0] and_866_nl;
  wire[0:0] nor_870_nl;
  wire[0:0] mux_1902_nl;
  wire[0:0] nor_871_nl;
  wire[0:0] nor_872_nl;
  wire[0:0] mux_1963_nl;
  wire[0:0] mux_1962_nl;
  wire[0:0] mux_1961_nl;
  wire[0:0] mux_1960_nl;
  wire[0:0] nor_818_nl;
  wire[0:0] nor_819_nl;
  wire[0:0] mux_1959_nl;
  wire[0:0] nor_820_nl;
  wire[0:0] nor_821_nl;
  wire[0:0] mux_1958_nl;
  wire[0:0] mux_1957_nl;
  wire[0:0] nor_822_nl;
  wire[0:0] nor_823_nl;
  wire[0:0] nor_824_nl;
  wire[0:0] mux_1956_nl;
  wire[0:0] mux_1955_nl;
  wire[0:0] mux_1954_nl;
  wire[0:0] nor_825_nl;
  wire[0:0] and_848_nl;
  wire[0:0] mux_1953_nl;
  wire[0:0] and_856_nl;
  wire[0:0] nor_828_nl;
  wire[0:0] mux_1952_nl;
  wire[0:0] mux_1951_nl;
  wire[0:0] and_864_nl;
  wire[0:0] and_865_nl;
  wire[0:0] mux_1950_nl;
  wire[0:0] mux_1949_nl;
  wire[0:0] nor_831_nl;
  wire[0:0] nor_832_nl;
  wire[0:0] nor_833_nl;
  wire[0:0] and_489_nl;
  wire[0:0] mux_1948_nl;
  wire[0:0] mux_1947_nl;
  wire[0:0] mux_1946_nl;
  wire[0:0] mux_1945_nl;
  wire[0:0] and_491_nl;
  wire[0:0] mux_1944_nl;
  wire[0:0] nor_835_nl;
  wire[0:0] nor_836_nl;
  wire[0:0] mux_1943_nl;
  wire[0:0] mux_1942_nl;
  wire[0:0] and_492_nl;
  wire[0:0] mux_1939_nl;
  wire[0:0] mux_1938_nl;
  wire[0:0] mux_1937_nl;
  wire[0:0] nor_840_nl;
  wire[0:0] nor_841_nl;
  wire[0:0] mux_1936_nl;
  wire[0:0] nor_842_nl;
  wire[0:0] nor_843_nl;
  wire[0:0] mux_1935_nl;
  wire[0:0] mux_1934_nl;
  wire[0:0] and_495_nl;
  wire[0:0] nor_844_nl;
  wire[0:0] mux_1933_nl;
  wire[0:0] and_496_nl;
  wire[0:0] nor_845_nl;
  wire[0:0] nor_792_nl;
  wire[0:0] mux_1994_nl;
  wire[0:0] mux_1993_nl;
  wire[0:0] nor_793_nl;
  wire[0:0] mux_1992_nl;
  wire[0:0] nand_79_nl;
  wire[0:0] mux_1989_nl;
  wire[0:0] mux_1988_nl;
  wire[0:0] nand_156_nl;
  wire[0:0] or_2109_nl;
  wire[0:0] mux_1987_nl;
  wire[0:0] nand_158_nl;
  wire[0:0] or_2106_nl;
  wire[0:0] mux_1986_nl;
  wire[0:0] mux_1985_nl;
  wire[0:0] mux_1984_nl;
  wire[0:0] nor_797_nl;
  wire[0:0] nor_798_nl;
  wire[0:0] mux_1983_nl;
  wire[0:0] and_486_nl;
  wire[0:0] nor_799_nl;
  wire[0:0] mux_1982_nl;
  wire[0:0] mux_1981_nl;
  wire[0:0] and_839_nl;
  wire[0:0] nor_801_nl;
  wire[0:0] mux_1980_nl;
  wire[0:0] nor_802_nl;
  wire[0:0] nor_803_nl;
  wire[0:0] mux_1979_nl;
  wire[0:0] mux_1978_nl;
  wire[0:0] mux_1977_nl;
  wire[0:0] mux_1976_nl;
  wire[0:0] nor_804_nl;
  wire[0:0] nor_805_nl;
  wire[0:0] mux_1975_nl;
  wire[0:0] and_487_nl;
  wire[0:0] nor_806_nl;
  wire[0:0] mux_1974_nl;
  wire[0:0] mux_1973_nl;
  wire[0:0] and_847_nl;
  wire[0:0] nor_808_nl;
  wire[0:0] mux_1972_nl;
  wire[0:0] nor_809_nl;
  wire[0:0] nor_810_nl;
  wire[0:0] mux_1971_nl;
  wire[0:0] mux_1970_nl;
  wire[0:0] mux_1969_nl;
  wire[0:0] nor_811_nl;
  wire[0:0] nor_812_nl;
  wire[0:0] mux_1968_nl;
  wire[0:0] and_488_nl;
  wire[0:0] nor_813_nl;
  wire[0:0] mux_1967_nl;
  wire[0:0] mux_1966_nl;
  wire[0:0] and_863_nl;
  wire[0:0] nor_815_nl;
  wire[0:0] mux_1965_nl;
  wire[0:0] nor_816_nl;
  wire[0:0] nor_817_nl;
  wire[0:0] mux_2025_nl;
  wire[0:0] mux_2024_nl;
  wire[0:0] mux_2023_nl;
  wire[0:0] nor_769_nl;
  wire[0:0] mux_2022_nl;
  wire[0:0] mux_2021_nl;
  wire[0:0] nor_770_nl;
  wire[0:0] nor_771_nl;
  wire[0:0] nor_772_nl;
  wire[0:0] mux_2020_nl;
  wire[0:0] mux_2019_nl;
  wire[0:0] mux_2018_nl;
  wire[0:0] nor_773_nl;
  wire[0:0] nor_774_nl;
  wire[0:0] nor_775_nl;
  wire[0:0] nor_776_nl;
  wire[0:0] mux_2017_nl;
  wire[0:0] mux_2016_nl;
  wire[0:0] mux_2015_nl;
  wire[0:0] nor_777_nl;
  wire[0:0] mux_2014_nl;
  wire[0:0] nor_778_nl;
  wire[0:0] nor_779_nl;
  wire[0:0] nor_780_nl;
  wire[0:0] mux_2013_nl;
  wire[0:0] nor_781_nl;
  wire[0:0] mux_2012_nl;
  wire[0:0] mux_2011_nl;
  wire[0:0] nor_782_nl;
  wire[0:0] nor_783_nl;
  wire[0:0] nor_784_nl;
  wire[0:0] mux_2010_nl;
  wire[0:0] mux_2009_nl;
  wire[0:0] mux_2008_nl;
  wire[0:0] and_479_nl;
  wire[0:0] mux_2007_nl;
  wire[0:0] nor_785_nl;
  wire[0:0] and_480_nl;
  wire[0:0] nor_786_nl;
  wire[0:0] mux_2006_nl;
  wire[0:0] or_2136_nl;
  wire[0:0] nand_149_nl;
  wire[0:0] mux_2005_nl;
  wire[0:0] nor_787_nl;
  wire[0:0] mux_2004_nl;
  wire[0:0] or_2132_nl;
  wire[0:0] nand_150_nl;
  wire[0:0] and_481_nl;
  wire[0:0] mux_2002_nl;
  wire[0:0] nor_789_nl;
  wire[0:0] mux_2001_nl;
  wire[0:0] mux_2000_nl;
  wire[0:0] or_2126_nl;
  wire[0:0] nand_151_nl;
  wire[0:0] mux_1999_nl;
  wire[0:0] or_2123_nl;
  wire[0:0] nand_152_nl;
  wire[0:0] and_483_nl;
  wire[0:0] mux_1998_nl;
  wire[0:0] mux_1997_nl;
  wire[0:0] and_484_nl;
  wire[0:0] nor_790_nl;
  wire[0:0] mux_1996_nl;
  wire[0:0] and_485_nl;
  wire[0:0] nor_791_nl;
  wire[0:0] nor_751_nl;
  wire[0:0] mux_2056_nl;
  wire[0:0] mux_2055_nl;
  wire[0:0] and_463_nl;
  wire[0:0] mux_2054_nl;
  wire[0:0] and_464_nl;
  wire[0:0] mux_2051_nl;
  wire[0:0] mux_2050_nl;
  wire[0:0] and_465_nl;
  wire[0:0] nor_755_nl;
  wire[0:0] mux_2049_nl;
  wire[0:0] and_466_nl;
  wire[0:0] nor_756_nl;
  wire[0:0] mux_2048_nl;
  wire[0:0] mux_2047_nl;
  wire[0:0] mux_2046_nl;
  wire[0:0] and_467_nl;
  wire[0:0] nor_757_nl;
  wire[0:0] mux_2045_nl;
  wire[0:0] and_468_nl;
  wire[0:0] and_469_nl;
  wire[0:0] mux_2044_nl;
  wire[0:0] mux_2043_nl;
  wire[0:0] and_838_nl;
  wire[0:0] and_844_nl;
  wire[0:0] mux_2042_nl;
  wire[0:0] and_470_nl;
  wire[0:0] nor_760_nl;
  wire[0:0] mux_2041_nl;
  wire[0:0] mux_2040_nl;
  wire[0:0] mux_2039_nl;
  wire[0:0] mux_2038_nl;
  wire[0:0] and_471_nl;
  wire[0:0] mux_2037_nl;
  wire[0:0] and_473_nl;
  wire[0:0] mux_2036_nl;
  wire[0:0] mux_2035_nl;
  wire[0:0] and_846_nl;
  wire[0:0] mux_2034_nl;
  wire[0:0] nor_764_nl;
  wire[0:0] mux_2033_nl;
  wire[0:0] mux_2032_nl;
  wire[0:0] mux_2031_nl;
  wire[0:0] and_475_nl;
  wire[0:0] nor_765_nl;
  wire[0:0] mux_2030_nl;
  wire[0:0] and_476_nl;
  wire[0:0] and_477_nl;
  wire[0:0] mux_2029_nl;
  wire[0:0] mux_2028_nl;
  wire[0:0] and_861_nl;
  wire[0:0] and_862_nl;
  wire[0:0] mux_2027_nl;
  wire[0:0] and_478_nl;
  wire[0:0] nor_768_nl;
  wire[0:0] mux_2088_nl;
  wire[0:0] mux_2087_nl;
  wire[0:0] mux_2086_nl;
  wire[0:0] mux_2085_nl;
  wire[0:0] nor_731_nl;
  wire[0:0] nor_732_nl;
  wire[0:0] mux_2084_nl;
  wire[0:0] nor_733_nl;
  wire[0:0] nor_734_nl;
  wire[0:0] mux_2083_nl;
  wire[0:0] mux_2082_nl;
  wire[0:0] nor_735_nl;
  wire[0:0] nor_736_nl;
  wire[0:0] nor_737_nl;
  wire[0:0] mux_2081_nl;
  wire[0:0] mux_2080_nl;
  wire[0:0] mux_2079_nl;
  wire[0:0] and_447_nl;
  wire[0:0] and_845_nl;
  wire[0:0] mux_2078_nl;
  wire[0:0] and_854_nl;
  wire[0:0] nor_740_nl;
  wire[0:0] mux_2077_nl;
  wire[0:0] mux_2076_nl;
  wire[0:0] and_859_nl;
  wire[0:0] and_860_nl;
  wire[0:0] mux_2075_nl;
  wire[0:0] mux_2074_nl;
  wire[0:0] and_448_nl;
  wire[0:0] nor_743_nl;
  wire[0:0] nor_744_nl;
  wire[0:0] and_449_nl;
  wire[0:0] mux_2073_nl;
  wire[0:0] mux_2072_nl;
  wire[0:0] mux_2071_nl;
  wire[0:0] mux_2070_nl;
  wire[0:0] and_451_nl;
  wire[0:0] mux_2069_nl;
  wire[0:0] and_833_nl;
  wire[0:0] and_452_nl;
  wire[0:0] mux_2068_nl;
  wire[0:0] mux_2067_nl;
  wire[0:0] and_454_nl;
  wire[0:0] mux_2064_nl;
  wire[0:0] mux_2063_nl;
  wire[0:0] mux_2062_nl;
  wire[0:0] and_837_nl;
  wire[0:0] and_457_nl;
  wire[0:0] mux_2061_nl;
  wire[0:0] and_843_nl;
  wire[0:0] and_458_nl;
  wire[0:0] mux_2060_nl;
  wire[0:0] mux_2059_nl;
  wire[0:0] and_459_nl;
  wire[0:0] and_460_nl;
  wire[0:0] mux_2058_nl;
  wire[0:0] and_461_nl;
  wire[0:0] and_462_nl;
  wire[5:0] COMP_LOOP_1_tmp_mul_nl;
  wire[11:0] nl_COMP_LOOP_1_tmp_mul_nl;
  wire[0:0] mux_2097_nl;
  wire[0:0] mux_2096_nl;
  wire[0:0] or_2260_nl;
  wire[0:0] mux_2095_nl;
  wire[0:0] mux_2094_nl;
  wire[0:0] or_2257_nl;
  wire[0:0] mux_2093_nl;
  wire[0:0] mux_2092_nl;
  wire[0:0] mux_2091_nl;
  wire[0:0] or_2255_nl;
  wire[0:0] mux_2090_nl;
  wire[0:0] or_2254_nl;
  wire[0:0] or_2253_nl;
  wire[0:0] mux_2104_nl;
  wire[0:0] mux_2103_nl;
  wire[0:0] mux_2102_nl;
  wire[0:0] nor_723_nl;
  wire[0:0] mux_2115_nl;
  wire[0:0] mux_2114_nl;
  wire[0:0] mux_2113_nl;
  wire[0:0] mux_2112_nl;
  wire[0:0] nor_711_nl;
  wire[0:0] and_445_nl;
  wire[0:0] mux_2122_nl;
  wire[0:0] mux_2121_nl;
  wire[0:0] mux_2120_nl;
  wire[0:0] nor_703_nl;
  wire[0:0] nor_692_nl;
  wire[0:0] mux_2135_nl;
  wire[0:0] mux_2134_nl;
  wire[0:0] mux_2133_nl;
  wire[0:0] nor_689_nl;
  wire[0:0] nor_690_nl;
  wire[0:0] mux_2129_nl;
  wire[0:0] mux_2127_nl;
  wire[0:0] nor_696_nl;
  wire[0:0] mux_2142_nl;
  wire[0:0] mux_2141_nl;
  wire[0:0] mux_2140_nl;
  wire[0:0] nor_681_nl;
  wire[0:0] mux_2153_nl;
  wire[0:0] mux_2152_nl;
  wire[0:0] mux_2151_nl;
  wire[0:0] mux_2150_nl;
  wire[0:0] nor_669_nl;
  wire[0:0] and_443_nl;
  wire[0:0] mux_2160_nl;
  wire[0:0] mux_2159_nl;
  wire[0:0] mux_2158_nl;
  wire[0:0] nor_661_nl;
  wire[0:0] nor_650_nl;
  wire[0:0] mux_2174_nl;
  wire[0:0] mux_2173_nl;
  wire[0:0] mux_2172_nl;
  wire[0:0] nor_646_nl;
  wire[0:0] mux_2171_nl;
  wire[0:0] nor_648_nl;
  wire[0:0] mux_2167_nl;
  wire[0:0] mux_2165_nl;
  wire[0:0] nor_654_nl;
  wire[0:0] mux_2181_nl;
  wire[0:0] mux_2180_nl;
  wire[0:0] mux_2179_nl;
  wire[0:0] nor_638_nl;
  wire[0:0] mux_2192_nl;
  wire[0:0] mux_2191_nl;
  wire[0:0] mux_2190_nl;
  wire[0:0] mux_2189_nl;
  wire[0:0] nor_626_nl;
  wire[0:0] and_441_nl;
  wire[0:0] mux_2199_nl;
  wire[0:0] mux_2198_nl;
  wire[0:0] mux_2197_nl;
  wire[0:0] nor_618_nl;
  wire[0:0] nor_607_nl;
  wire[0:0] mux_2212_nl;
  wire[0:0] mux_2211_nl;
  wire[0:0] mux_2210_nl;
  wire[0:0] nor_604_nl;
  wire[0:0] nor_605_nl;
  wire[0:0] mux_2206_nl;
  wire[0:0] mux_2204_nl;
  wire[0:0] nor_611_nl;
  wire[0:0] mux_2219_nl;
  wire[0:0] mux_2218_nl;
  wire[0:0] mux_2217_nl;
  wire[0:0] nor_596_nl;
  wire[0:0] mux_2230_nl;
  wire[0:0] mux_2229_nl;
  wire[0:0] mux_2228_nl;
  wire[0:0] mux_2227_nl;
  wire[0:0] and_434_nl;
  wire[0:0] and_435_nl;
  wire[0:0] mux_2237_nl;
  wire[0:0] mux_2236_nl;
  wire[0:0] mux_2235_nl;
  wire[0:0] and_426_nl;
  wire[11:0] acc_nl;
  wire[12:0] nl_acc_nl;
  wire[10:0] COMP_LOOP_mux_358_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_nand_1_nl;
  wire[9:0] COMP_LOOP_mux_359_nl;
  wire[53:0] COMP_LOOP_and_260_nl;
  wire[53:0] COMP_LOOP_mux1h_710_nl;
  wire[0:0] COMP_LOOP_and_261_nl;
  wire[0:0] COMP_LOOP_mux1h_711_nl;
  wire[0:0] COMP_LOOP_and_262_nl;
  wire[0:0] COMP_LOOP_mux1h_712_nl;
  wire[7:0] COMP_LOOP_mux1h_713_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_983_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_984_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_985_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_986_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_987_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_988_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_989_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_990_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_991_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_992_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_993_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_994_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_995_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_996_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_997_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_998_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_999_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1000_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1001_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1002_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1003_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1004_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1005_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1006_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1007_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1008_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1009_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1010_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1011_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1012_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1013_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1014_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1015_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1016_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1017_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1018_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1019_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1020_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1021_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1022_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1023_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1024_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1025_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1026_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1027_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1028_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1029_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1030_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1031_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1032_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1033_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1034_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1035_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1036_nl;
  wire[0:0] COMP_LOOP_and_263_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_mux_8_nl;
  wire[0:0] COMP_LOOP_and_264_nl;
  wire[0:0] COMP_LOOP_mux1h_714_nl;
  wire[3:0] COMP_LOOP_mux1h_715_nl;
  wire[0:0] COMP_LOOP_or_61_nl;
  wire[0:0] COMP_LOOP_mux1h_716_nl;
  wire[0:0] COMP_LOOP_or_62_nl;
  wire[0:0] COMP_LOOP_mux1h_717_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_2_nl;
  wire[0:0] COMP_LOOP_mux_360_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_3_nl;
  wire[3:0] STAGE_LOOP_mux_4_nl;
  wire[0:0] COMP_LOOP_mux1h_718_nl;
  wire[0:0] COMP_LOOP_mux1h_719_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1037_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1038_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1039_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1040_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1041_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1042_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1043_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1044_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1045_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1046_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1047_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1048_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1049_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1050_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1051_nl;
  wire[0:0] COMP_LOOP_mux1h_720_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1052_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1053_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1054_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1055_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1056_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1057_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1058_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1059_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1060_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1061_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1062_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1063_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1064_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1065_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1066_nl;
  wire[0:0] COMP_LOOP_mux1h_721_nl;
  wire[0:0] COMP_LOOP_mux1h_722_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1067_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1068_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1069_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1070_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1071_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1072_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1073_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1074_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1075_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1076_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1077_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1078_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1079_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1080_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1081_nl;
  wire[0:0] COMP_LOOP_mux1h_723_nl;
  wire[0:0] COMP_LOOP_mux1h_724_nl;
  wire[0:0] COMP_LOOP_mux1h_725_nl;
  wire[0:0] COMP_LOOP_mux1h_726_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1082_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1083_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1084_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1085_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1086_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1087_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1088_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1089_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1090_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1091_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1092_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1093_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1094_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1095_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1096_nl;
  wire[0:0] COMP_LOOP_mux1h_727_nl;
  wire[0:0] COMP_LOOP_mux1h_728_nl;
  wire[0:0] COMP_LOOP_mux1h_729_nl;
  wire[0:0] COMP_LOOP_mux1h_730_nl;
  wire[0:0] COMP_LOOP_mux1h_731_nl;
  wire[0:0] COMP_LOOP_mux1h_732_nl;
  wire[0:0] COMP_LOOP_mux1h_733_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[64:0] acc_3_nl;
  wire[65:0] nl_acc_3_nl;
  wire[63:0] COMP_LOOP_COMP_LOOP_mux_10_nl;
  wire[0:0] mux_2274_nl;
  wire[0:0] mux_2273_nl;
  wire[0:0] mux_2272_nl;
  wire[0:0] mux_2271_nl;
  wire[0:0] mux_2270_nl;
  wire[0:0] and_423_nl;
  wire[0:0] nor_587_nl;
  wire[0:0] mux_2269_nl;
  wire[0:0] mux_2266_nl;
  wire[0:0] mux_2262_nl;
  wire[0:0] mux_2261_nl;
  wire[0:0] or_2438_nl;
  wire[0:0] mux_2260_nl;
  wire[0:0] or_2437_nl;
  wire[0:0] mux_2259_nl;
  wire[0:0] mux_2258_nl;
  wire[0:0] nand_97_nl;
  wire [63:0] nl_COMP_LOOP_1_modulo_cmp_base_rsc_dat;
  assign COMP_LOOP_COMP_LOOP_mux_10_nl = MUX_v_64_2_2((~ COMP_LOOP_10_acc_8_itm),
      (~ z_out_7), COMP_LOOP_or_18_itm);
  assign nl_acc_3_nl = ({COMP_LOOP_mux_361_cse , 1'b1}) + ({COMP_LOOP_COMP_LOOP_mux_10_nl
      , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[64:0];
  assign and_423_nl = (fsm_output[3]) & (fsm_output[8]) & (fsm_output[0]) & (fsm_output[5]);
  assign nor_587_nl = ~((fsm_output[3]) | (fsm_output[8]) | not_tmp_676);
  assign mux_2270_nl = MUX_s_1_2_2(and_423_nl, nor_587_nl, fsm_output[4]);
  assign mux_2271_nl = MUX_s_1_2_2(mux_2270_nl, mux_tmp_2249, fsm_output[6]);
  assign mux_2269_nl = MUX_s_1_2_2((~ mux_tmp_2249), mux_tmp_2245, fsm_output[6]);
  assign mux_2272_nl = MUX_s_1_2_2((~ mux_2271_nl), mux_2269_nl, fsm_output[1]);
  assign mux_2273_nl = MUX_s_1_2_2(mux_2272_nl, mux_tmp_2246, fsm_output[7]);
  assign or_2438_nl = (fsm_output[4]) | mux_tmp_2238;
  assign or_2437_nl = (~ (fsm_output[3])) | (fsm_output[8]) | not_tmp_676;
  assign mux_2260_nl = MUX_s_1_2_2(mux_tmp_2237, or_2437_nl, fsm_output[4]);
  assign mux_2261_nl = MUX_s_1_2_2(or_2438_nl, mux_2260_nl, fsm_output[6]);
  assign mux_2258_nl = MUX_s_1_2_2(mux_tmp_2237, mux_tmp_2238, fsm_output[4]);
  assign nand_97_nl = ~((fsm_output[4]) & (~ mux_tmp_2237));
  assign mux_2259_nl = MUX_s_1_2_2(mux_2258_nl, nand_97_nl, fsm_output[6]);
  assign mux_2262_nl = MUX_s_1_2_2(mux_2261_nl, mux_2259_nl, fsm_output[1]);
  assign mux_2266_nl = MUX_s_1_2_2(mux_tmp_2246, mux_2262_nl, fsm_output[7]);
  assign mux_2274_nl = MUX_s_1_2_2(mux_2273_nl, mux_2266_nl, fsm_output[2]);
  assign nl_COMP_LOOP_1_modulo_cmp_base_rsc_dat = MUX_v_64_2_2(COMP_LOOP_10_acc_8_itm,
      (readslicef_65_64_1(acc_3_nl)), mux_2274_nl);
  wire [63:0] nl_COMP_LOOP_1_modulo_cmp_m_rsc_dat;
  assign nl_COMP_LOOP_1_modulo_cmp_m_rsc_dat = p_sva;
  wire[0:0] mux_2293_nl;
  wire[0:0] mux_2292_nl;
  wire[0:0] mux_2291_nl;
  wire[0:0] mux_2290_nl;
  wire[0:0] or_2456_nl;
  wire[0:0] mux_2289_nl;
  wire[0:0] or_2661_nl;
  wire[0:0] mux_2288_nl;
  wire[0:0] mux_2287_nl;
  wire[0:0] mux_2286_nl;
  wire[0:0] nand_98_nl;
  wire[0:0] mux_2285_nl;
  wire[0:0] mux_2284_nl;
  wire[0:0] mux_2282_nl;
  wire[0:0] or_2453_nl;
  wire[0:0] mux_2281_nl;
  wire[0:0] mux_2280_nl;
  wire[0:0] mux_2279_nl;
  wire[0:0] or_2450_nl;
  wire [0:0] nl_COMP_LOOP_1_modulo_cmp_ccs_ccore_start_rsc_dat;
  assign or_2456_nl = (fsm_output[3]) | mux_tmp_2258;
  assign mux_2290_nl = MUX_s_1_2_2(or_2456_nl, mux_tmp_2257, and_421_cse);
  assign or_2661_nl = (fsm_output[0]) | (~ (fsm_output[3])) | mux_tmp_2259;
  assign mux_2289_nl = MUX_s_1_2_2(or_2661_nl, or_tmp_2279, fsm_output[5]);
  assign mux_2291_nl = MUX_s_1_2_2(mux_2290_nl, mux_2289_nl, fsm_output[4]);
  assign mux_2286_nl = MUX_s_1_2_2(or_tmp_2277, mux_tmp_2257, fsm_output[0]);
  assign nand_98_nl = ~((fsm_output[3]) & (~ mux_tmp_2256));
  assign mux_2287_nl = MUX_s_1_2_2(mux_2286_nl, nand_98_nl, fsm_output[5]);
  assign mux_2288_nl = MUX_s_1_2_2(mux_tmp_2264, mux_2287_nl, fsm_output[4]);
  assign mux_2292_nl = MUX_s_1_2_2(mux_2291_nl, mux_2288_nl, fsm_output[6]);
  assign or_2453_nl = (fsm_output[5]) | (fsm_output[0]);
  assign mux_2282_nl = MUX_s_1_2_2(or_tmp_2277, mux_tmp_2257, or_2453_nl);
  assign mux_2284_nl = MUX_s_1_2_2(mux_tmp_2264, mux_2282_nl, fsm_output[4]);
  assign mux_2279_nl = MUX_s_1_2_2(mux_tmp_2259, mux_tmp_2258, fsm_output[3]);
  assign mux_2280_nl = MUX_s_1_2_2(or_tmp_2277, mux_2279_nl, and_421_cse);
  assign or_2450_nl = (fsm_output[5]) | (fsm_output[0]) | mux_tmp_2257;
  assign mux_2281_nl = MUX_s_1_2_2(mux_2280_nl, or_2450_nl, fsm_output[4]);
  assign mux_2285_nl = MUX_s_1_2_2(mux_2284_nl, mux_2281_nl, fsm_output[6]);
  assign mux_2293_nl = MUX_s_1_2_2(mux_2292_nl, mux_2285_nl, fsm_output[1]);
  assign nl_COMP_LOOP_1_modulo_cmp_ccs_ccore_start_rsc_dat = ~ mux_2293_nl;
  wire[0:0] and_884_nl;
  wire [3:0] nl_COMP_LOOP_9_tmp_lshift_rg_s;
  assign and_884_nl = (fsm_output==9'b000000010);
  assign nl_COMP_LOOP_9_tmp_lshift_rg_s = MUX_v_4_2_2(STAGE_LOOP_i_3_0_sva, z_out_4,
      and_884_nl);
  wire[0:0] and_897_nl;
  wire [3:0] nl_COMP_LOOP_2_tmp_lshift_rg_s;
  assign and_897_nl = (fsm_output==9'b000000010);
  assign nl_COMP_LOOP_2_tmp_lshift_rg_s = MUX_v_4_2_2(COMP_LOOP_1_tmp_acc_cse_sva,
      z_out_4, and_897_nl);
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_31_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_31_tr0 = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_62_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_62_tr0 = ~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_93_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_93_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_124_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_124_tr0 = ~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_155_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_155_tr0 = ~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_186_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_186_tr0 = ~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_217_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_217_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_248_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_248_tr0 = ~ COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_279_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_279_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_310_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_310_tr0 = ~ COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_341_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_341_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_372_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_372_tr0 = ~ COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_403_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_403_tr0 = ~ COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_434_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_434_tr0 = ~ COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_465_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_465_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_496_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_496_tr0 = ~ COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0 = z_out_2[10];
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0 = ~ STAGE_LOOP_acc_itm_4_1;
  ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd64)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_15_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_14_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_13_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_12_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_11_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_10_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_9_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_8_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_7_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_6_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_5_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_4_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_3_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_2_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_1_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_15_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_14_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_13_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_12_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_11_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_10_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_9_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_8_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_7_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_6_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_5_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_4_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_3_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_2_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_1_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_0_lz)
    );
  modulo  COMP_LOOP_1_modulo_cmp (
      .base_rsc_dat(nl_COMP_LOOP_1_modulo_cmp_base_rsc_dat[63:0]),
      .m_rsc_dat(nl_COMP_LOOP_1_modulo_cmp_m_rsc_dat[63:0]),
      .return_rsc_z(COMP_LOOP_1_modulo_cmp_return_rsc_z),
      .ccs_ccore_start_rsc_dat(nl_COMP_LOOP_1_modulo_cmp_ccs_ccore_start_rsc_dat[0:0]),
      .ccs_ccore_clk(clk),
      .ccs_ccore_srst(rst),
      .ccs_ccore_en(COMP_LOOP_1_modulo_cmp_ccs_ccore_en)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd6)) COMP_LOOP_1_tmp_lshift_rg (
      .a(1'b1),
      .s(z_out_4),
      .z(COMP_LOOP_1_tmp_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) COMP_LOOP_9_tmp_lshift_rg (
      .a(1'b1),
      .s(nl_COMP_LOOP_9_tmp_lshift_rg_s[3:0]),
      .z(z_out)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd10)) COMP_LOOP_2_tmp_lshift_rg (
      .a(1'b1),
      .s(nl_COMP_LOOP_2_tmp_lshift_rg_s[3:0]),
      .z(z_out_1)
    );
  inPlaceNTT_DIF_core_wait_dp inPlaceNTT_DIF_core_wait_dp_inst (
      .ensig_cgo_iro(mux_2255_rmff),
      .ensig_cgo(reg_ensig_cgo_cse),
      .COMP_LOOP_1_modulo_cmp_ccs_ccore_en(COMP_LOOP_1_modulo_cmp_ccs_ccore_en)
    );
  inPlaceNTT_DIF_core_core_fsm inPlaceNTT_DIF_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .COMP_LOOP_C_31_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_31_tr0[0:0]),
      .COMP_LOOP_C_62_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_62_tr0[0:0]),
      .COMP_LOOP_C_93_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_93_tr0[0:0]),
      .COMP_LOOP_C_124_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_124_tr0[0:0]),
      .COMP_LOOP_C_155_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_155_tr0[0:0]),
      .COMP_LOOP_C_186_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_186_tr0[0:0]),
      .COMP_LOOP_C_217_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_217_tr0[0:0]),
      .COMP_LOOP_C_248_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_248_tr0[0:0]),
      .COMP_LOOP_C_279_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_279_tr0[0:0]),
      .COMP_LOOP_C_310_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_310_tr0[0:0]),
      .COMP_LOOP_C_341_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_341_tr0[0:0]),
      .COMP_LOOP_C_372_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_372_tr0[0:0]),
      .COMP_LOOP_C_403_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_403_tr0[0:0]),
      .COMP_LOOP_C_434_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_434_tr0[0:0]),
      .COMP_LOOP_C_465_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_465_tr0[0:0]),
      .COMP_LOOP_C_496_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_496_tr0[0:0]),
      .VEC_LOOP_C_0_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0[0:0]),
      .STAGE_LOOP_C_1_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0[0:0])
    );
  assign nor_1589_nl = ~((VEC_LOOP_j_10_0_sva_9_0[2]) | (COMP_LOOP_acc_16_psp_sva[0])
      | (~ COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm) | (VEC_LOOP_j_10_0_sva_9_0[0]) |
      (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_1590_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00)
      | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) | (fsm_output[7]) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign mux_1128_cse = MUX_s_1_2_2(nor_1589_nl, nor_1590_nl, fsm_output[2]);
  assign nor_346_cse = ~((VEC_LOOP_j_10_0_sva_9_0[1]) | (~ (fsm_output[5])));
  assign nor_1554_cse = ~((COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b0001) | (fsm_output[7])
      | not_tmp_395);
  assign nand_271_cse = ~((fsm_output[2]) & (fsm_output[7]) & (fsm_output[6]) & (fsm_output[8]));
  assign nand_272_cse = ~((COMP_LOOP_acc_1_cse_sva[0]) & (fsm_output[8:6]==3'b111));
  assign nor_1528_cse = ~((COMP_LOOP_acc_16_psp_sva[0]) | (~ COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b011));
  assign nor_1529_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b001));
  assign mux_1190_nl = MUX_s_1_2_2(nor_1528_cse, nor_1529_nl, fsm_output[2]);
  assign nor_1530_nl = ~((~ (fsm_output[2])) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00)
      | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) | (fsm_output[8:6]!=3'b001));
  assign mux_1191_cse = MUX_s_1_2_2(mux_1190_nl, nor_1530_nl, VEC_LOOP_j_10_0_sva_9_0[2]);
  assign nor_351_cse = ~((VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01));
  assign nor_1523_cse = ~((COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b011));
  assign nor_1526_cse = ~((COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b100));
  assign nor_1527_cse = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b010));
  assign nand_265_cse = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[1]) & (fsm_output[7])
      & (fsm_output[4]) & (fsm_output[8]));
  assign nor_1435_cse = ~((COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b0011) | (fsm_output[7])
      | not_tmp_395);
  assign nor_1402_cse = ~((COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b011));
  assign nor_1405_cse = ~((COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b100));
  assign nor_1406_cse = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b010));
  assign nor_1352_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[2])) | (COMP_LOOP_acc_16_psp_sva[0])
      | (~ COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm) | (VEC_LOOP_j_10_0_sva_9_0[0]) |
      (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_1353_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01)
      | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) | (fsm_output[7]) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign mux_1378_cse = MUX_s_1_2_2(nor_1352_nl, nor_1353_nl, fsm_output[2]);
  assign nor_1317_cse = ~((COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b0101) | (fsm_output[7])
      | not_tmp_395);
  assign nor_1286_cse = ~((COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b011));
  assign nor_1289_cse = ~((COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b100));
  assign nor_1290_cse = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b010));
  assign nor_1291_nl = ~((~ (fsm_output[2])) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01)
      | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) | (fsm_output[8:6]!=3'b001));
  assign nor_1293_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b001));
  assign mux_1440_nl = MUX_s_1_2_2(nor_1528_cse, nor_1293_nl, fsm_output[2]);
  assign mux_1441_cse = MUX_s_1_2_2(nor_1291_nl, mux_1440_nl, VEC_LOOP_j_10_0_sva_9_0[2]);
  assign nor_1200_cse = ~((COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b0111) | (fsm_output[7])
      | not_tmp_395);
  assign nand_226_cse = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:0]==4'b0111));
  assign and_529_cse = (COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]==4'b0111) & (fsm_output[8:6]==3'b011);
  assign nor_1173_cse = ~((COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b0111) | (fsm_output[8:6]!=3'b100));
  assign nor_1174_cse = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0111) | (fsm_output[8:6]!=3'b010));
  assign nand_219_cse = ~((COMP_LOOP_acc_10_cse_10_1_sva[3]) & (fsm_output[7]) &
      (fsm_output[4]) & (fsm_output[8]));
  assign nor_1121_nl = ~((VEC_LOOP_j_10_0_sva_9_0[2]) | (~ (COMP_LOOP_acc_16_psp_sva[0]))
      | (~ COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm) | (VEC_LOOP_j_10_0_sva_9_0[0]) |
      (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_1122_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10)
      | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) | (fsm_output[7]) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign mux_1628_cse = MUX_s_1_2_2(nor_1121_nl, nor_1122_nl, fsm_output[2]);
  assign nor_1086_cse = ~((COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b1001) | (fsm_output[7])
      | not_tmp_395);
  assign nand_211_cse = ~((COMP_LOOP_acc_10_cse_10_1_sva[3]) & (fsm_output[2]) &
      (fsm_output[7]) & (fsm_output[6]) & (fsm_output[8]));
  assign nand_212_cse = ~((COMP_LOOP_acc_1_cse_sva[3]) & (COMP_LOOP_acc_1_cse_sva[0])
      & (fsm_output[8:6]==3'b111));
  assign and_523_cse = (COMP_LOOP_acc_16_psp_sva[0]) & COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[8:6]==3'b011);
  assign nor_1061_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b001));
  assign mux_1690_nl = MUX_s_1_2_2(and_523_cse, nor_1061_nl, fsm_output[2]);
  assign nor_1062_nl = ~((~ (fsm_output[2])) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10)
      | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) | (fsm_output[8:6]!=3'b001));
  assign mux_1691_cse = MUX_s_1_2_2(mux_1690_nl, nor_1062_nl, VEC_LOOP_j_10_0_sva_9_0[2]);
  assign nor_1056_cse = ~((COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b011));
  assign nor_1059_cse = ~((COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b100));
  assign nor_1060_cse = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b010));
  assign nor_970_cse = ~((COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b1011) | (fsm_output[7])
      | not_tmp_395);
  assign and_506_cse = (COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]==4'b1011) & (fsm_output[8:6]==3'b011);
  assign nor_944_cse = ~((COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b1011) | (fsm_output[8:6]!=3'b100));
  assign nor_945_cse = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b1011) | (fsm_output[8:6]!=3'b010));
  assign and_503_nl = (VEC_LOOP_j_10_0_sva_9_0[2]) & (COMP_LOOP_acc_16_psp_sva[0])
      & COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm & (~ (VEC_LOOP_j_10_0_sva_9_0[0])) &
      (fsm_output[7]) & (fsm_output[4]) & (~ (fsm_output[8]));
  assign nor_893_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11)
      | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) | (fsm_output[7]) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign mux_1878_cse = MUX_s_1_2_2(and_503_nl, nor_893_nl, fsm_output[2]);
  assign nor_860_cse = ~((COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b1101) | (fsm_output[7])
      | not_tmp_395);
  assign and_490_cse = (COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]==4'b1101) & (fsm_output[8:6]==3'b011);
  assign nor_837_cse = ~((COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b1101) | (fsm_output[8:6]!=3'b100));
  assign nor_838_cse = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b1101) | (fsm_output[8:6]!=3'b010));
  assign nand_170_cse = ~((COMP_LOOP_acc_1_cse_sva[2]) & (COMP_LOOP_acc_1_cse_sva[3])
      & (COMP_LOOP_acc_1_cse_sva[0]) & (fsm_output[8:6]==3'b111));
  assign and_493_nl = (fsm_output[2]) & (COMP_LOOP_acc_13_psp_sva[1:0]==2'b11) &
      COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm & (fsm_output[8:6]==3'b001);
  assign nor_839_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b001));
  assign mux_1940_nl = MUX_s_1_2_2(and_523_cse, nor_839_nl, fsm_output[2]);
  assign mux_1941_cse = MUX_s_1_2_2(and_493_nl, mux_1940_nl, VEC_LOOP_j_10_0_sva_9_0[2]);
  assign nor_761_cse = ~((~((COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]==4'b1111) & (~
      (fsm_output[7])))) | not_tmp_395);
  assign and_450_cse = (COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b011);
  assign and_836_cse = (COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b100);
  assign and_453_cse = (COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b010);
  assign or_2259_cse_1 = (fsm_output[3:2]!=2'b00);
  assign nand_122_cse = ~((z_out_3[0]) & (fsm_output[4]));
  assign nand_121_cse = ~((z_out_3[1:0]==2'b11) & (fsm_output[4]));
  assign mux_2251_nl = MUX_s_1_2_2((~ mux_tmp_2224), mux_955_cse, fsm_output[7]);
  assign mux_2252_nl = MUX_s_1_2_2(mux_2251_nl, mux_965_cse, fsm_output[0]);
  assign mux_2253_nl = MUX_s_1_2_2(mux_tmp_2229, (~ mux_2252_nl), fsm_output[5]);
  assign mux_2254_nl = MUX_s_1_2_2(mux_952_cse, mux_2253_nl, fsm_output[6]);
  assign mux_2245_nl = MUX_s_1_2_2(mux_tmp_2225, mux_949_cse, fsm_output[0]);
  assign mux_2249_nl = MUX_s_1_2_2(mux_tmp_2229, mux_2245_nl, fsm_output[5]);
  assign mux_2242_nl = MUX_s_1_2_2(mux_949_cse, (~ mux_965_cse), fsm_output[5]);
  assign mux_2250_nl = MUX_s_1_2_2(mux_2249_nl, mux_2242_nl, fsm_output[6]);
  assign mux_2255_rmff = MUX_s_1_2_2(mux_2254_nl, mux_2250_nl, fsm_output[1]);
  assign and_421_cse = (fsm_output[5]) & (fsm_output[0]);
  assign nor_1624_cse = ~((fsm_output[3:2]!=2'b00));
  assign and_1189_cse = (fsm_output[1:0]==2'b11);
  assign nand_324_cse = ~((fsm_output[8:6]==3'b111));
  assign and_831_cse = (fsm_output[3:1]==3'b111);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_nor_cse = ~((z_out_3[3:0]!=4'b0000));
  assign COMP_LOOP_tmp_nor_cse = ~((z_out_3[3:1]!=3'b000));
  assign COMP_LOOP_tmp_nor_1_cse = ~((z_out_3[3]) | (z_out_3[2]) | (z_out_3[0]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_cse = (z_out_3[3:0]==4'b0011);
  assign COMP_LOOP_tmp_nor_3_cse = ~((z_out_3[3]) | (z_out_3[1]) | (z_out_3[0]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_cse = (z_out_3[3:0]==4'b0101);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_cse = (z_out_3[3:0]==4'b0110);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_cse = (z_out_3[3:0]==4'b0111);
  assign COMP_LOOP_tmp_nor_6_cse = ~((z_out_3[2:0]!=3'b000));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_cse = (z_out_3[3:0]==4'b1001);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_cse = (z_out_3[3:0]==4'b1010);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_cse = (z_out_3[3:0]==4'b1011);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse = (z_out_3[3:0]==4'b1100);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse = (z_out_3[3:0]==4'b1101);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse = (z_out_3[3:0]==4'b1110);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse = (z_out_3[3:0]==4'b1111);
  assign nor_1767_cse = ~((fsm_output[5]) | (fsm_output[0]));
  assign and_407_cse = (fsm_output[4:3]==2'b11);
  assign and_733_cse = (fsm_output[8:7]==2'b11);
  assign or_2729_cse = (fsm_output[6]) | (fsm_output[1]) | (fsm_output[7]) | (fsm_output[2]);
  assign and_728_cse = or_2729_cse & (fsm_output[8]);
  assign and_712_cse = (fsm_output[0]) & (fsm_output[3]);
  assign or_432_cse = (fsm_output[2:1]!=2'b00);
  assign and_674_cse = (fsm_output[2:1]==2'b11);
  assign and_675_cse = (fsm_output[4]) & (fsm_output[8]);
  assign or_2697_cse = (fsm_output[6]) | (fsm_output[2]);
  assign nand_301_cse = ~((fsm_output[7]) & (fsm_output[4]) & (fsm_output[8]));
  assign nor_298_nl = ~((fsm_output[3:2]!=2'b10));
  assign mux_955_cse = MUX_s_1_2_2(and_675_cse, (fsm_output[4]), nor_298_nl);
  assign or_611_cse = (fsm_output[2]) | mux_tmp_929;
  assign nor_1642_nl = ~((fsm_output[4]) | (fsm_output[8]));
  assign mux_951_nl = MUX_s_1_2_2(nor_1642_nl, and_675_cse, fsm_output[3]);
  assign or_614_nl = (fsm_output[2]) | (~ mux_951_nl);
  assign mux_952_cse = MUX_s_1_2_2(or_614_nl, nand_tmp_13, fsm_output[7]);
  assign mux_949_cse = MUX_s_1_2_2(nand_tmp_13, or_611_cse, fsm_output[7]);
  assign mux_965_cse = MUX_s_1_2_2((~ nand_tmp_13), mux_955_cse, fsm_output[7]);
  assign COMP_LOOP_tmp_or_1_cse = and_dcpl_62 | and_dcpl_189 | and_dcpl_181 | and_dcpl_190
      | and_dcpl_183 | and_dcpl_191 | and_dcpl_184 | and_dcpl_192;
  assign COMP_LOOP_tmp_or_2_cse = and_dcpl_62 | and_dcpl_65 | and_dcpl_181 | and_dcpl_190
      | and_dcpl_183 | and_dcpl_191 | and_dcpl_184 | and_dcpl_192;
  assign COMP_LOOP_or_27_cse = and_dcpl_181 | and_dcpl_190 | and_dcpl_183 | and_dcpl_191
      | and_dcpl_184 | and_dcpl_192;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_17_cse = (z_out_3[2:0]==3'b011);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_19_cse = (z_out_3[2:0]==3'b101);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_20_cse = (z_out_3[2:0]==3'b110);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_21_cse = (z_out_3[2:0]==3'b111);
  assign COMP_LOOP_or_31_cse = and_dcpl_195 | and_dcpl_197 | and_dcpl_198;
  assign COMP_LOOP_or_23_cse = and_dcpl_189 | and_dcpl_181 | and_dcpl_190 | and_dcpl_183
      | and_dcpl_191 | and_dcpl_184 | and_dcpl_192;
  assign nor_1630_cse = ~((fsm_output[8:7]!=2'b00));
  assign and_1191_cse = (COMP_LOOP_10_tmp_mul_idiv_sva[1]) & COMP_LOOP_tmp_nor_14_itm;
  assign and_1190_cse = (COMP_LOOP_10_tmp_mul_idiv_sva[2]) & COMP_LOOP_tmp_nor_16_itm;
  assign and_314_m1c = and_dcpl_51 & and_dcpl_111;
  assign COMP_LOOP_tmp_or_29_cse = COMP_LOOP_tmp_COMP_LOOP_tmp_and_155 | COMP_LOOP_tmp_COMP_LOOP_tmp_and_157
      | COMP_LOOP_tmp_COMP_LOOP_tmp_and_159;
  assign COMP_LOOP_tmp_or_19_cse = and_dcpl_65 | and_dcpl_195 | and_dcpl_197 | and_dcpl_198;
  assign nor_572_cse = ~((fsm_output[7:6]!=2'b00));
  assign or_2589_cse = (fsm_output[5:4]!=2'b00);
  assign COMP_LOOP_tmp_or_21_cse = and_dcpl_189 | and_dcpl_195 | and_dcpl_197 | and_dcpl_198;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_nor_14_cse = ~((COMP_LOOP_13_tmp_mul_idiv_sva[1:0]!=2'b00));
  assign and_570_cse = (fsm_output[3:2]==2'b11);
  assign or_2612_cse = (fsm_output[3:0]!=4'b0000);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_nor_16_rgt = ~((COMP_LOOP_5_tmp_mul_idiv_sva[1:0]!=2'b00)
      | nor_1798_tmp);
  assign COMP_LOOP_tmp_and_14_rgt = (COMP_LOOP_5_tmp_mul_idiv_sva[1:0]==2'b01) &
      (~ nor_1798_tmp);
  assign COMP_LOOP_tmp_and_15_rgt = (COMP_LOOP_5_tmp_mul_idiv_sva[1:0]==2'b10) &
      (~ nor_1798_tmp);
  assign COMP_LOOP_tmp_and_16_rgt = (COMP_LOOP_5_tmp_mul_idiv_sva[1:0]==2'b11) &
      (~ nor_1798_tmp);
  assign mux_228_cse = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[6]);
  assign or_2621_cse = and_570_cse | (fsm_output[7:6]!=2'b00);
  assign mux_464_cse = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), fsm_output[7]);
  assign mux_559_cse = MUX_s_1_2_2(mux_464_cse, and_733_cse, fsm_output[6]);
  assign or_455_cse = (fsm_output[8:7]!=2'b00);
  assign or_454_cse = (fsm_output[8:7]!=2'b01);
  assign or_2626_cse = ((fsm_output[3:0]==4'b1111)) | (fsm_output[6]);
  assign and_655_cse = (((fsm_output[6]) & (fsm_output[1]) & (fsm_output[2])) | (fsm_output[7]))
      & (fsm_output[8]);
  assign nl_COMP_LOOP_1_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_4_sva_5_0
      , 4'b0000}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_1_acc_10_nl = nl_COMP_LOOP_1_acc_10_nl[10:0];
  assign COMP_LOOP_1_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_1_acc_10_nl);
  assign nl_COMP_LOOP_acc_13_psp_sva_1 = (VEC_LOOP_j_10_0_sva_9_0[9:2]) + ({COMP_LOOP_k_10_4_sva_5_0
      , 2'b01});
  assign COMP_LOOP_acc_13_psp_sva_1 = nl_COMP_LOOP_acc_13_psp_sva_1[7:0];
  assign nl_COMP_LOOP_acc_1_cse_4_sva_1 = VEC_LOOP_j_10_0_sva_9_0 + ({COMP_LOOP_k_10_4_sva_5_0
      , 4'b0011});
  assign COMP_LOOP_acc_1_cse_4_sva_1 = nl_COMP_LOOP_acc_1_cse_4_sva_1[9:0];
  assign nl_COMP_LOOP_acc_1_cse_2_sva_1 = VEC_LOOP_j_10_0_sva_9_0 + ({COMP_LOOP_k_10_4_sva_5_0
      , 4'b0001});
  assign COMP_LOOP_acc_1_cse_2_sva_1 = nl_COMP_LOOP_acc_1_cse_2_sva_1[9:0];
  assign nl_COMP_LOOP_2_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_4_sva_5_0
      , 4'b0001}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_2_acc_10_nl = nl_COMP_LOOP_2_acc_10_nl[10:0];
  assign COMP_LOOP_2_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_2_acc_10_nl);
  assign nl_COMP_LOOP_3_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_4_sva_5_0
      , 4'b0010}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_3_acc_10_nl = nl_COMP_LOOP_3_acc_10_nl[10:0];
  assign COMP_LOOP_3_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_3_acc_10_nl);
  assign nl_COMP_LOOP_4_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_4_sva_5_0
      , 4'b0011}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_4_acc_10_nl = nl_COMP_LOOP_4_acc_10_nl[10:0];
  assign COMP_LOOP_4_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_4_acc_10_nl);
  assign nl_COMP_LOOP_5_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_4_sva_5_0
      , 4'b0100}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_5_acc_10_nl = nl_COMP_LOOP_5_acc_10_nl[10:0];
  assign COMP_LOOP_5_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_5_acc_10_nl);
  assign nl_COMP_LOOP_6_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_4_sva_5_0
      , 4'b0101}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_6_acc_10_nl = nl_COMP_LOOP_6_acc_10_nl[10:0];
  assign COMP_LOOP_6_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_6_acc_10_nl);
  assign nl_COMP_LOOP_7_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_4_sva_5_0
      , 4'b0110}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_7_acc_10_nl = nl_COMP_LOOP_7_acc_10_nl[10:0];
  assign COMP_LOOP_7_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_7_acc_10_nl);
  assign nl_COMP_LOOP_8_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_4_sva_5_0
      , 4'b0111}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_8_acc_10_nl = nl_COMP_LOOP_8_acc_10_nl[10:0];
  assign COMP_LOOP_8_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_8_acc_10_nl);
  assign nl_COMP_LOOP_9_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_4_sva_5_0
      , 4'b1000}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_9_acc_10_nl = nl_COMP_LOOP_9_acc_10_nl[10:0];
  assign COMP_LOOP_9_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_9_acc_10_nl);
  assign nl_COMP_LOOP_10_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_4_sva_5_0
      , 4'b1001}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_10_acc_10_nl = nl_COMP_LOOP_10_acc_10_nl[10:0];
  assign COMP_LOOP_10_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_10_acc_10_nl);
  assign nl_COMP_LOOP_11_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_4_sva_5_0
      , 4'b1010}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_11_acc_10_nl = nl_COMP_LOOP_11_acc_10_nl[10:0];
  assign COMP_LOOP_11_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_11_acc_10_nl);
  assign nl_COMP_LOOP_12_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_4_sva_5_0
      , 4'b1011}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_12_acc_10_nl = nl_COMP_LOOP_12_acc_10_nl[10:0];
  assign COMP_LOOP_12_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_12_acc_10_nl);
  assign nl_COMP_LOOP_13_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_4_sva_5_0
      , 4'b1100}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_13_acc_10_nl = nl_COMP_LOOP_13_acc_10_nl[10:0];
  assign COMP_LOOP_13_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_13_acc_10_nl);
  assign nl_COMP_LOOP_14_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_4_sva_5_0
      , 4'b1101}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_14_acc_10_nl = nl_COMP_LOOP_14_acc_10_nl[10:0];
  assign COMP_LOOP_14_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_14_acc_10_nl);
  assign nl_COMP_LOOP_15_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_4_sva_5_0
      , 4'b1110}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_15_acc_10_nl = nl_COMP_LOOP_15_acc_10_nl[10:0];
  assign COMP_LOOP_15_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_15_acc_10_nl);
  assign nl_COMP_LOOP_16_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_4_sva_5_0
      , 4'b1111}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_16_acc_10_nl = nl_COMP_LOOP_16_acc_10_nl[10:0];
  assign COMP_LOOP_16_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_16_acc_10_nl);
  assign nl_COMP_LOOP_k_10_4_sva_2 = conv_u2u_6_7(COMP_LOOP_k_10_4_sva_5_0) + 7'b0000001;
  assign COMP_LOOP_k_10_4_sva_2 = nl_COMP_LOOP_k_10_4_sva_2[6:0];
  assign COMP_LOOP_tmp_mux1h_4_itm_mx0w3 = MUX1HOT_v_64_16_2(twiddle_rsc_0_0_i_q_d,
      tmp_33_sva_1, tmp_33_sva_2, tmp_33_sva_3, tmp_33_sva_4, tmp_33_sva_5, tmp_33_sva_6,
      tmp_33_sva_7, tmp_33_sva_8, tmp_33_sva_9, tmp_33_sva_10, tmp_33_sva_11, tmp_33_sva_12,
      tmp_33_sva_13, tmp_33_sva_14, tmp_33_sva_15, {COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_itm
      , COMP_LOOP_tmp_COMP_LOOP_tmp_and_167 , and_1191_cse , COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm
      , and_1190_cse , COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm , COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm
      , COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm , COMP_LOOP_tmp_COMP_LOOP_tmp_and_161
      , COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm , COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm
      , COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm , COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm
      , COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm , COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm
      , COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm});
  assign nor_1792_cse = ~((COMP_LOOP_11_tmp_mul_idiv_sva[2:1]!=2'b00));
  assign and_313_nl = (COMP_LOOP_11_tmp_mul_idiv_sva[2:1]==2'b10);
  assign tmp_33_sva_13_mx0w1 = MUX1HOT_v_64_3_2(twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_4_i_q_d,
      twiddle_rsc_0_8_i_q_d, {nor_1792_cse , (COMP_LOOP_11_tmp_mul_idiv_sva[1]) ,
      and_313_nl});
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_155 = (COMP_LOOP_11_tmp_mul_idiv_sva[0])
      & nor_1792_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_157 = (COMP_LOOP_11_tmp_mul_idiv_sva[2:0]==3'b010);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_159 = (COMP_LOOP_11_tmp_mul_idiv_sva[2:0]==3'b100);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_161 = (COMP_LOOP_10_tmp_mul_idiv_sva[3])
      & COMP_LOOP_tmp_nor_19_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_167 = (COMP_LOOP_10_tmp_mul_idiv_sva[0])
      & COMP_LOOP_tmp_nor_13_itm;
  assign or_dcpl_5 = COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm;
  assign and_dcpl_5 = nor_1630_cse & (~ (fsm_output[6]));
  assign or_36_cse = (fsm_output[3:1]!=3'b000);
  assign nor_tmp_10 = (fsm_output[3]) & (fsm_output[2]) & (fsm_output[1]) & (fsm_output[6]);
  assign or_tmp_29 = and_674_cse | (fsm_output[6]);
  assign nor_tmp_47 = (fsm_output[7:6]==2'b11);
  assign or_2732_cse = (fsm_output[7:6]!=2'b00);
  assign nor_tmp_115 = or_2732_cse & (fsm_output[8]);
  assign mux_tmp_439 = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), or_2732_cse);
  assign mux_tmp_538 = MUX_s_1_2_2(mux_tmp_439, nor_tmp_115, and_674_cse);
  assign or_610_cse = (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_tmp_929 = MUX_s_1_2_2((~ and_675_cse), or_610_cse, fsm_output[3]);
  assign nand_tmp_13 = ~((fsm_output[2]) & (~ mux_tmp_929));
  assign and_dcpl_45 = ~((fsm_output[5:4]!=2'b00));
  assign and_dcpl_46 = ~((fsm_output[3]) | (fsm_output[0]));
  assign and_dcpl_47 = and_dcpl_46 & and_dcpl_45;
  assign and_dcpl_48 = ~((fsm_output[2:1]!=2'b00));
  assign and_dcpl_51 = and_dcpl_5 & and_dcpl_48;
  assign and_dcpl_53 = (fsm_output[5:4]==2'b11);
  assign and_dcpl_54 = and_dcpl_46 & and_dcpl_53;
  assign and_dcpl_55 = (fsm_output[2:1]==2'b10);
  assign and_dcpl_57 = and_733_cse & (fsm_output[6]);
  assign and_dcpl_58 = and_dcpl_57 & and_dcpl_55;
  assign nor_tmp_339 = or_2259_cse_1 & (fsm_output[8:6]==3'b111);
  assign and_565_nl = (fsm_output[2]) & (fsm_output[1]) & (fsm_output[6]) & (fsm_output[7])
      & (fsm_output[8]);
  assign mux_1080_nl = MUX_s_1_2_2(and_565_nl, and_dcpl_57, fsm_output[3]);
  assign mux_tmp_1062 = MUX_s_1_2_2(mux_1080_nl, nor_tmp_339, fsm_output[0]);
  assign or_714_nl = (~ (fsm_output[4])) | (fsm_output[0]) | (~((fsm_output[1]) &
      (fsm_output[6])));
  assign mux_1083_nl = MUX_s_1_2_2((fsm_output[6]), (~ (fsm_output[6])), fsm_output[1]);
  assign nand_22_nl = ~((fsm_output[4]) & (fsm_output[0]) & mux_1083_nl);
  assign mux_tmp_1065 = MUX_s_1_2_2(or_714_nl, nand_22_nl, fsm_output[5]);
  assign nand_23_nl = ~((fsm_output[7]) & (~ mux_tmp_1065));
  assign or_712_nl = (fsm_output[5]) | (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[1])
      | (fsm_output[6]);
  assign mux_1085_nl = MUX_s_1_2_2(mux_tmp_1065, or_712_nl, fsm_output[7]);
  assign mux_tmp_1067 = MUX_s_1_2_2(nand_23_nl, mux_1085_nl, fsm_output[2]);
  assign and_dcpl_60 = (fsm_output[2:1]==2'b01);
  assign and_dcpl_61 = and_dcpl_5 & and_dcpl_60;
  assign and_dcpl_62 = and_dcpl_61 & and_dcpl_47;
  assign and_dcpl_63 = (~ (fsm_output[3])) & (fsm_output[0]);
  assign and_dcpl_64 = and_dcpl_63 & and_dcpl_45;
  assign and_dcpl_65 = and_dcpl_61 & and_dcpl_64;
  assign and_dcpl_66 = (fsm_output[5:4]==2'b10);
  assign and_dcpl_67 = and_dcpl_63 & and_dcpl_66;
  assign and_dcpl_69 = and_dcpl_46 & and_dcpl_66;
  assign and_dcpl_70 = and_dcpl_61 & and_dcpl_69;
  assign and_dcpl_71 = nor_1630_cse & (fsm_output[6]);
  assign and_dcpl_72 = and_dcpl_71 & and_dcpl_48;
  assign and_dcpl_74 = and_dcpl_72 & and_dcpl_64;
  assign and_dcpl_75 = (fsm_output[5:4]==2'b01);
  assign and_dcpl_77 = and_712_cse & and_dcpl_75;
  assign and_dcpl_79 = and_dcpl_71 & and_674_cse;
  assign and_dcpl_81 = and_dcpl_72 & and_dcpl_69;
  assign and_dcpl_82 = (fsm_output[3]) & (~ (fsm_output[0]));
  assign and_dcpl_83 = and_dcpl_82 & and_dcpl_53;
  assign and_dcpl_85 = and_712_cse & and_dcpl_53;
  assign and_dcpl_86 = and_dcpl_79 & and_dcpl_85;
  assign and_dcpl_87 = (fsm_output[8:7]==2'b01);
  assign and_dcpl_88 = and_dcpl_87 & (~ (fsm_output[6]));
  assign and_dcpl_89 = and_dcpl_88 & and_dcpl_55;
  assign and_dcpl_91 = and_dcpl_82 & and_dcpl_75;
  assign and_dcpl_92 = and_dcpl_88 & and_674_cse;
  assign and_dcpl_93 = and_dcpl_92 & and_dcpl_91;
  assign and_dcpl_95 = and_dcpl_89 & and_dcpl_85;
  assign and_dcpl_96 = and_dcpl_87 & (fsm_output[6]);
  assign and_dcpl_97 = and_dcpl_96 & and_dcpl_60;
  assign and_dcpl_99 = and_dcpl_96 & and_dcpl_55;
  assign and_dcpl_100 = and_dcpl_99 & and_dcpl_91;
  assign and_dcpl_102 = and_dcpl_97 & and_dcpl_85;
  assign and_dcpl_103 = (fsm_output[8:7]==2'b10);
  assign and_dcpl_104 = and_dcpl_103 & (~ (fsm_output[6]));
  assign and_dcpl_105 = and_dcpl_104 & and_dcpl_48;
  assign and_dcpl_107 = and_dcpl_104 & and_dcpl_60;
  assign and_dcpl_108 = and_dcpl_107 & and_dcpl_91;
  assign and_dcpl_110 = and_dcpl_105 & and_dcpl_85;
  assign and_dcpl_111 = and_dcpl_63 & and_dcpl_75;
  assign and_dcpl_112 = and_dcpl_103 & (fsm_output[6]);
  assign and_dcpl_113 = and_dcpl_112 & and_674_cse;
  assign and_dcpl_115 = and_dcpl_112 & and_dcpl_48;
  assign and_dcpl_116 = and_dcpl_115 & and_dcpl_91;
  assign and_dcpl_118 = and_dcpl_63 & and_dcpl_53;
  assign and_dcpl_119 = and_dcpl_113 & and_dcpl_118;
  assign and_dcpl_120 = and_733_cse & (~ (fsm_output[6]));
  assign and_dcpl_121 = and_dcpl_120 & and_dcpl_55;
  assign and_dcpl_123 = and_dcpl_46 & and_dcpl_75;
  assign and_dcpl_124 = and_dcpl_120 & and_674_cse;
  assign and_dcpl_125 = and_dcpl_124 & and_dcpl_123;
  assign and_dcpl_127 = and_dcpl_121 & and_dcpl_118;
  assign and_dcpl_128 = and_dcpl_57 & and_dcpl_60;
  assign and_dcpl_130 = and_dcpl_58 & and_dcpl_123;
  assign and_dcpl_131 = and_dcpl_5 & and_674_cse;
  assign and_dcpl_136 = and_dcpl_71 & and_dcpl_55;
  assign and_dcpl_141 = and_dcpl_88 & and_dcpl_60;
  assign and_dcpl_146 = and_dcpl_96 & and_dcpl_48;
  assign and_dcpl_151 = and_dcpl_104 & and_674_cse;
  assign and_dcpl_156 = and_dcpl_112 & and_dcpl_55;
  assign and_dcpl_161 = and_dcpl_120 & and_dcpl_60;
  assign and_dcpl_166 = and_dcpl_57 & and_dcpl_48;
  assign not_tmp_395 = ~((fsm_output[6]) & (fsm_output[8]));
  assign or_762_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8]));
  assign or_760_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_10_0_sva_9_0[2])
      | (fsm_output[8:6]!=3'b100);
  assign or_758_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (fsm_output[8:6]!=3'b010);
  assign mux_1115_nl = MUX_s_1_2_2(or_760_nl, or_758_nl, fsm_output[2]);
  assign mux_1116_cse = MUX_s_1_2_2(or_762_nl, mux_1115_nl, fsm_output[3]);
  assign not_tmp_399 = ~((fsm_output[4]) & (fsm_output[8]));
  assign nor_1479_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign nor_1480_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_10_0_sva_9_0[2])
      | (fsm_output[8:6]!=3'b100));
  assign nor_1481_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (fsm_output[8:6]!=3'b010));
  assign mux_1240_nl = MUX_s_1_2_2(nor_1480_nl, nor_1481_nl, fsm_output[2]);
  assign mux_1241_cse = MUX_s_1_2_2(nor_1479_nl, mux_1240_nl, fsm_output[3]);
  assign nand_268_cse = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[1]) & (fsm_output[8:6]==3'b111));
  assign nand_261_cse = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[1:0]==2'b11) & (fsm_output[8:6]==3'b111));
  assign or_1150_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8]));
  assign or_1148_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (~ (VEC_LOOP_j_10_0_sva_9_0[2]))
      | (fsm_output[8:6]!=3'b100);
  assign or_1146_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (fsm_output[8:6]!=3'b010);
  assign mux_1365_nl = MUX_s_1_2_2(or_1148_nl, or_1146_nl, fsm_output[2]);
  assign mux_1366_cse = MUX_s_1_2_2(or_1150_nl, mux_1365_nl, fsm_output[3]);
  assign nor_1242_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign nor_1243_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) | (~ (VEC_LOOP_j_10_0_sva_9_0[2]))
      | (fsm_output[8:6]!=3'b100));
  assign nor_1244_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (fsm_output[8:6]!=3'b010));
  assign mux_1490_nl = MUX_s_1_2_2(nor_1243_nl, nor_1244_nl, fsm_output[2]);
  assign mux_1491_cse = MUX_s_1_2_2(nor_1242_nl, mux_1490_nl, fsm_output[3]);
  assign or_1538_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8]));
  assign or_1536_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_10_0_sva_9_0[2])
      | (fsm_output[8:6]!=3'b100);
  assign or_1534_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (fsm_output[8:6]!=3'b010);
  assign mux_1615_nl = MUX_s_1_2_2(or_1536_nl, or_1534_nl, fsm_output[2]);
  assign mux_1616_cse = MUX_s_1_2_2(or_1538_nl, mux_1615_nl, fsm_output[3]);
  assign nand_222_cse = ~((COMP_LOOP_acc_20_psp_sva[2]) & (fsm_output[8:6]==3'b111));
  assign nand_223_cse = ~((COMP_LOOP_acc_10_cse_10_1_sva[3]) & (fsm_output[8:6]==3'b111));
  assign nor_1012_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign nor_1013_nl = ~((~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_10_0_sva_9_0[2])
      | (fsm_output[8:6]!=3'b100));
  assign nor_1014_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (fsm_output[8:6]!=3'b010));
  assign mux_1740_nl = MUX_s_1_2_2(nor_1013_nl, nor_1014_nl, fsm_output[2]);
  assign mux_1741_cse = MUX_s_1_2_2(nor_1012_nl, mux_1740_nl, fsm_output[3]);
  assign nand_322_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]==2'b11) & (fsm_output[2])
      & (fsm_output[7]) & (~ (fsm_output[6])) & (fsm_output[8]));
  assign or_1922_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (~ (VEC_LOOP_j_10_0_sva_9_0[2]))
      | (fsm_output[8:6]!=3'b100);
  assign or_1920_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (fsm_output[8:6]!=3'b010);
  assign mux_1865_nl = MUX_s_1_2_2(or_1922_nl, or_1920_nl, fsm_output[2]);
  assign mux_1866_cse = MUX_s_1_2_2(nand_322_nl, mux_1865_nl, fsm_output[3]);
  assign nand_184_cse = ~((COMP_LOOP_acc_20_psp_sva[2:1]==2'b11) & (fsm_output[8:6]==3'b111));
  assign nand_185_cse = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:2]==2'b11) & (fsm_output[8:6]==3'b111));
  assign and_835_nl = (COMP_LOOP_acc_19_psp_sva[1:0]==2'b11) & (fsm_output[2]) &
      (fsm_output[7]) & (~ (fsm_output[6])) & (fsm_output[8]);
  assign nor_795_nl = ~((~ (COMP_LOOP_acc_16_psp_sva[0])) | (~ (VEC_LOOP_j_10_0_sva_9_0[2]))
      | (fsm_output[8:6]!=3'b100));
  assign nor_796_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (fsm_output[8:6]!=3'b010));
  assign mux_1990_nl = MUX_s_1_2_2(nor_795_nl, nor_796_nl, fsm_output[2]);
  assign mux_1991_cse = MUX_s_1_2_2(and_835_nl, mux_1990_nl, fsm_output[3]);
  assign nand_157_cse = ~((COMP_LOOP_acc_17_psp_sva[2:0]==3'b111) & (~ (fsm_output[7])));
  assign and_dcpl_171 = (fsm_output[0]) & (~ (fsm_output[5]));
  assign and_dcpl_175 = (or_36_cse ^ (fsm_output[4])) & (~ (fsm_output[8])) & nor_572_cse
      & and_dcpl_171;
  assign and_dcpl_180 = (or_2259_cse_1 ^ (fsm_output[4])) & nor_1630_cse & (~ (fsm_output[6]))
      & (~ (fsm_output[1])) & nor_1767_cse;
  assign and_dcpl_181 = and_dcpl_131 & and_dcpl_47;
  assign and_dcpl_182 = and_dcpl_82 & and_dcpl_45;
  assign and_dcpl_183 = and_dcpl_61 & and_dcpl_182;
  assign and_dcpl_184 = and_dcpl_131 & and_dcpl_182;
  assign and_dcpl_186 = nor_1630_cse & (fsm_output[6:5]==2'b00);
  assign or_tmp_2077 = (fsm_output[4]) | (COMP_LOOP_10_tmp_mul_idiv_sva[3:0]!=4'b0000);
  assign and_dcpl_188 = and_dcpl_5 & and_dcpl_55;
  assign and_dcpl_189 = and_dcpl_188 & and_dcpl_47;
  assign and_dcpl_190 = and_dcpl_51 & and_dcpl_182;
  assign and_dcpl_191 = and_dcpl_188 & and_dcpl_182;
  assign and_dcpl_192 = and_dcpl_51 & and_dcpl_123;
  assign and_dcpl_193 = and_dcpl_5 & nor_1767_cse;
  assign and_dcpl_195 = and_dcpl_131 & and_dcpl_64;
  assign and_dcpl_196 = and_712_cse & and_dcpl_45;
  assign and_dcpl_197 = and_dcpl_61 & and_dcpl_196;
  assign and_dcpl_198 = and_dcpl_131 & and_dcpl_196;
  assign and_dcpl_202 = and_dcpl_188 & and_dcpl_196;
  assign and_dcpl_207 = and_dcpl_51 & and_dcpl_196;
  assign or_2430_nl = (fsm_output[3]) | (fsm_output[4]) | (fsm_output[8]);
  assign mux_tmp_2224 = MUX_s_1_2_2(or_2430_nl, mux_tmp_929, fsm_output[2]);
  assign mux_tmp_2225 = MUX_s_1_2_2(mux_tmp_2224, or_611_cse, fsm_output[7]);
  assign mux_tmp_2229 = MUX_s_1_2_2(mux_952_cse, mux_tmp_2225, fsm_output[0]);
  assign or_tmp_2258 = (fsm_output[8]) | (fsm_output[0]) | (fsm_output[5]);
  assign or_2434_nl = (~ (fsm_output[8])) | (fsm_output[0]) | (fsm_output[5]);
  assign mux_tmp_2237 = MUX_s_1_2_2(or_2434_nl, or_tmp_2258, fsm_output[3]);
  assign not_tmp_676 = ~((fsm_output[0]) & (fsm_output[5]));
  assign nor_tmp_480 = (fsm_output[8]) & (fsm_output[0]) & (fsm_output[5]);
  assign or_2435_nl = (fsm_output[8]) | not_tmp_676;
  assign mux_tmp_2238 = MUX_s_1_2_2((~ nor_tmp_480), or_2435_nl, fsm_output[3]);
  assign or_tmp_2266 = (~ (fsm_output[3])) | (~ (fsm_output[8])) | (fsm_output[0])
      | (fsm_output[5]);
  assign mux_2263_nl = MUX_s_1_2_2((~ (fsm_output[5])), (fsm_output[5]), fsm_output[0]);
  assign or_2443_nl = (fsm_output[3]) | (fsm_output[8]) | mux_2263_nl;
  assign mux_tmp_2245 = MUX_s_1_2_2(or_2443_nl, or_tmp_2266, fsm_output[4]);
  assign or_2444_nl = (fsm_output[6]) | mux_tmp_2245;
  assign or_2440_nl = (~ (fsm_output[6])) | (fsm_output[4]) | mux_tmp_2238;
  assign mux_tmp_2246 = MUX_s_1_2_2(or_2444_nl, or_2440_nl, fsm_output[1]);
  assign mux_2267_nl = MUX_s_1_2_2((~ or_tmp_2258), nor_tmp_480, fsm_output[3]);
  assign mux_tmp_2249 = MUX_s_1_2_2((~ or_tmp_2266), mux_2267_nl, fsm_output[4]);
  assign and_dcpl_220 = and_dcpl_61 & and_dcpl_67;
  assign and_dcpl_222 = and_dcpl_71 & and_dcpl_60 & and_dcpl_47;
  assign and_dcpl_223 = and_dcpl_72 & and_dcpl_67;
  assign and_dcpl_225 = and_dcpl_88 & and_dcpl_48 & and_dcpl_47;
  assign and_dcpl_226 = and_dcpl_92 & and_dcpl_77;
  assign and_dcpl_227 = and_dcpl_92 & and_dcpl_83;
  assign and_dcpl_228 = and_dcpl_99 & and_dcpl_77;
  assign and_dcpl_229 = and_dcpl_99 & and_dcpl_83;
  assign and_dcpl_230 = and_dcpl_107 & and_dcpl_77;
  assign and_dcpl_231 = and_dcpl_107 & and_dcpl_83;
  assign and_dcpl_232 = and_dcpl_115 & and_dcpl_77;
  assign and_dcpl_233 = and_dcpl_115 & and_dcpl_83;
  assign and_dcpl_234 = and_dcpl_124 & and_dcpl_111;
  assign and_dcpl_235 = and_dcpl_124 & and_dcpl_54;
  assign and_dcpl_236 = and_dcpl_58 & and_dcpl_111;
  assign or_tmp_2274 = (fsm_output[8:7]!=2'b10);
  assign mux_tmp_2256 = MUX_s_1_2_2(or_tmp_2274, or_454_cse, fsm_output[2]);
  assign nand_114_nl = ~((fsm_output[2]) & (fsm_output[7]) & (fsm_output[8]));
  assign mux_tmp_2257 = MUX_s_1_2_2(nand_114_nl, mux_tmp_2256, fsm_output[3]);
  assign mux_tmp_2258 = MUX_s_1_2_2(or_454_cse, or_455_cse, fsm_output[2]);
  assign nand_113_nl = ~((fsm_output[8:7]==2'b11));
  assign mux_tmp_2259 = MUX_s_1_2_2(nand_113_nl, or_tmp_2274, fsm_output[2]);
  assign or_tmp_2277 = (fsm_output[3]) | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[8]);
  assign or_tmp_2279 = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[2]) |
      (fsm_output[7]) | (fsm_output[8]);
  assign or_2455_nl = (fsm_output[0]) | mux_tmp_2257;
  assign mux_tmp_2264 = MUX_s_1_2_2(or_2455_nl, or_tmp_2279, fsm_output[5]);
  assign or_dcpl_182 = or_455_cse | (fsm_output[6]);
  assign or_dcpl_183 = or_dcpl_182 | (fsm_output[2:1]!=2'b01);
  assign or_dcpl_184 = or_dcpl_183 | (fsm_output[3]) | (fsm_output[0]) | or_2589_cse;
  assign or_2482_nl = (fsm_output[3]) | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[7])
      | (fsm_output[8]);
  assign or_2481_nl = (fsm_output[3]) | (fsm_output[2]) | (fsm_output[1]) | (fsm_output[6])
      | (fsm_output[7]) | (fsm_output[8]);
  assign mux_tmp_2282 = MUX_s_1_2_2(or_2482_nl, or_2481_nl, fsm_output[0]);
  assign mux_2302_nl = MUX_s_1_2_2((~ mux_tmp_2282), nor_tmp_339, fsm_output[4]);
  assign mux_2303_itm = MUX_s_1_2_2(mux_2302_nl, and_dcpl_57, fsm_output[5]);
  assign nor_tmp_489 = (and_570_cse | (fsm_output[6])) & (fsm_output[7]);
  assign mux_2306_nl = MUX_s_1_2_2(mux_228_cse, nor_tmp_47, or_2259_cse_1);
  assign mux_2305_nl = MUX_s_1_2_2(mux_228_cse, nor_tmp_47, or_36_cse);
  assign mux_tmp_2288 = MUX_s_1_2_2(mux_2306_nl, mux_2305_nl, fsm_output[0]);
  assign and_416_nl = (fsm_output[3]) & (fsm_output[2]) & (fsm_output[6]);
  assign mux_tmp_2291 = MUX_s_1_2_2(nor_tmp_10, and_416_nl, fsm_output[0]);
  assign or_2487_cse = (fsm_output[3]) | (fsm_output[2]) | (fsm_output[6]);
  assign or_2486_cse = (fsm_output[3]) | (fsm_output[2]) | (fsm_output[1]) | (fsm_output[6]);
  assign mux_tmp_2292 = MUX_s_1_2_2(or_2487_cse, or_2486_cse, fsm_output[0]);
  assign not_tmp_703 = ~((fsm_output[4]) | mux_tmp_2292);
  assign mux_22_nl = MUX_s_1_2_2(or_2259_cse_1, or_36_cse, fsm_output[0]);
  assign or_tmp_2300 = (fsm_output[4]) | mux_22_nl;
  assign or_dcpl_190 = (fsm_output[5:3]!=3'b000);
  assign and_dcpl_248 = (or_tmp_2300 ^ (fsm_output[5])) & and_dcpl_5;
  assign or_2497_nl = (fsm_output[1]) | (~ (fsm_output[6]));
  assign mux_2323_nl = MUX_s_1_2_2(or_2497_nl, (fsm_output[6]), or_2259_cse_1);
  assign mux_61_nl = MUX_s_1_2_2((~ (fsm_output[6])), (fsm_output[6]), or_36_cse);
  assign mux_2324_nl = MUX_s_1_2_2(mux_2323_nl, mux_61_nl, fsm_output[0]);
  assign mux_2325_nl = MUX_s_1_2_2(mux_2324_nl, (fsm_output[6]), or_2589_cse);
  assign and_dcpl_252 = (~ mux_2325_nl) & nor_1630_cse;
  assign and_411_nl = ((fsm_output[4:0]!=5'b00000)) & (fsm_output[6]);
  assign mux_2328_nl = MUX_s_1_2_2(not_tmp_703, and_411_nl, fsm_output[5]);
  assign and_dcpl_255 = (~ mux_2328_nl) & nor_1630_cse;
  assign nor_tmp_499 = ((fsm_output[2]) | (fsm_output[1]) | (fsm_output[6])) & (fsm_output[7]);
  assign mux_2329_nl = MUX_s_1_2_2(nor_tmp_47, nor_tmp_499, fsm_output[3]);
  assign mux_tmp_2311 = MUX_s_1_2_2(nor_tmp_489, mux_2329_nl, fsm_output[0]);
  assign and_dcpl_258 = (or_2697_cse | and_1189_cse | or_dcpl_190) & nor_1630_cse;
  assign mux_tmp_2318 = MUX_s_1_2_2(mux_tmp_2288, nor_tmp_47, fsm_output[4]);
  assign and_403_nl = or_2626_cse & (fsm_output[7]);
  assign mux_2342_nl = MUX_s_1_2_2(mux_tmp_2288, and_403_nl, fsm_output[4]);
  assign mux_2343_nl = MUX_s_1_2_2(mux_2342_nl, (fsm_output[7]), fsm_output[5]);
  assign and_dcpl_262 = ~(mux_2343_nl | (fsm_output[8]));
  assign nor_tmp_507 = or_432_cse & (fsm_output[7:6]==2'b11);
  assign and_tmp_28 = (fsm_output[3]) & nor_tmp_507;
  assign or_2507_nl = (fsm_output[3]) | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[7]);
  assign or_2506_nl = (fsm_output[3]) | (fsm_output[2]) | (fsm_output[1]) | (fsm_output[6])
      | (fsm_output[7]);
  assign mux_tmp_2325 = MUX_s_1_2_2(or_2507_nl, or_2506_nl, fsm_output[0]);
  assign and_401_nl = (fsm_output[3]) & (fsm_output[6]) & (fsm_output[7]);
  assign mux_tmp_2328 = MUX_s_1_2_2(and_tmp_28, and_401_nl, fsm_output[0]);
  assign nor_tmp_509 = (fsm_output[3]) & (fsm_output[2]) & (fsm_output[6]) & (fsm_output[7]);
  assign and_398_nl = (((fsm_output[4:1]==4'b1111)) | (fsm_output[6])) & (fsm_output[7]);
  assign mux_2353_nl = MUX_s_1_2_2(mux_tmp_2318, and_398_nl, fsm_output[5]);
  assign and_dcpl_266 = ~(mux_2353_nl | (fsm_output[8]));
  assign not_tmp_727 = ~((fsm_output[4]) | mux_tmp_2325);
  assign and_396_nl = (fsm_output[3]) & (fsm_output[2]) & (fsm_output[1]) & (fsm_output[6])
      & (fsm_output[7]);
  assign mux_2357_nl = MUX_s_1_2_2(and_396_nl, nor_tmp_509, fsm_output[0]);
  assign mux_2358_nl = MUX_s_1_2_2((~ mux_tmp_2325), mux_2357_nl, fsm_output[4]);
  assign mux_2359_nl = MUX_s_1_2_2(mux_2358_nl, nor_tmp_47, fsm_output[5]);
  assign and_dcpl_270 = ~(mux_2359_nl | (fsm_output[8]));
  assign nor_tmp_515 = ((fsm_output[3]) | (fsm_output[6]) | (fsm_output[7])) & (fsm_output[8]);
  assign mux_2362_nl = MUX_s_1_2_2(mux_tmp_439, nor_tmp_115, or_2259_cse_1);
  assign mux_2361_nl = MUX_s_1_2_2(mux_tmp_439, nor_tmp_115, or_36_cse);
  assign mux_tmp_2344 = MUX_s_1_2_2(mux_2362_nl, mux_2361_nl, fsm_output[0]);
  assign and_566_nl = (and_674_cse | (fsm_output[7:6]!=2'b00)) & (fsm_output[8]);
  assign mux_tmp_2347 = MUX_s_1_2_2(and_566_nl, (fsm_output[8]), fsm_output[3]);
  assign mux_tmp_2348 = MUX_s_1_2_2(nor_tmp_515, mux_tmp_2347, fsm_output[0]);
  assign mux_tmp_2351 = MUX_s_1_2_2(nor_tmp_115, and_728_cse, fsm_output[3]);
  assign and_392_nl = (fsm_output[4]) & (fsm_output[3]) & (fsm_output[2]) & (fsm_output[6])
      & (fsm_output[7]);
  assign mux_2374_nl = MUX_s_1_2_2(not_tmp_727, and_392_nl, fsm_output[5]);
  assign and_dcpl_271 = ~(mux_2374_nl | (fsm_output[8]));
  assign mux_tmp_2357 = MUX_s_1_2_2(mux_tmp_2344, nor_tmp_115, fsm_output[4]);
  assign and_388_nl = or_2621_cse & (fsm_output[8]);
  assign mux_2381_nl = MUX_s_1_2_2(and_388_nl, mux_tmp_2351, fsm_output[0]);
  assign mux_2382_nl = MUX_s_1_2_2(mux_tmp_2344, mux_2381_nl, fsm_output[4]);
  assign mux_2383_itm = MUX_s_1_2_2(mux_2382_nl, (fsm_output[8]), fsm_output[5]);
  assign mux_tmp_2365 = MUX_s_1_2_2(and_655_cse, nor_tmp_115, fsm_output[3]);
  assign mux_2387_nl = MUX_s_1_2_2(mux_464_cse, and_733_cse, or_2487_cse);
  assign mux_2386_nl = MUX_s_1_2_2(mux_464_cse, and_733_cse, or_2486_cse);
  assign mux_tmp_2369 = MUX_s_1_2_2(mux_2387_nl, mux_2386_nl, fsm_output[0]);
  assign nor_tmp_528 = ((or_2259_cse_1 & (fsm_output[6])) | (fsm_output[7])) & (fsm_output[8]);
  assign nor_tmp_530 = (((fsm_output[3]) & (fsm_output[6])) | (fsm_output[7])) &
      (fsm_output[8]);
  assign mux_2397_nl = MUX_s_1_2_2(nor_tmp_115, and_728_cse, and_407_cse);
  assign mux_2398_itm = MUX_s_1_2_2(mux_tmp_2357, mux_2397_nl, fsm_output[5]);
  assign mux_tmp_2384 = MUX_s_1_2_2(mux_tmp_2369, and_733_cse, fsm_output[4]);
  assign and_376_nl = ((or_432_cse & (fsm_output[6])) | (fsm_output[7])) & (fsm_output[8]);
  assign mux_2407_nl = MUX_s_1_2_2(and_733_cse, and_376_nl, fsm_output[3]);
  assign mux_2408_nl = MUX_s_1_2_2(mux_2407_nl, nor_tmp_530, fsm_output[0]);
  assign mux_2409_nl = MUX_s_1_2_2(mux_tmp_2369, mux_2408_nl, fsm_output[4]);
  assign mux_2410_itm = MUX_s_1_2_2(mux_2409_nl, nor_tmp_115, fsm_output[5]);
  assign nor_tmp_537 = or_2487_cse & (fsm_output[8:7]==2'b11);
  assign mux_tmp_2392 = MUX_s_1_2_2(nor_1630_cse, and_733_cse, fsm_output[6]);
  assign mux_2413_nl = MUX_s_1_2_2(mux_tmp_2392, and_dcpl_57, or_2259_cse_1);
  assign mux_2412_nl = MUX_s_1_2_2(mux_tmp_2392, and_dcpl_57, or_36_cse);
  assign mux_tmp_2395 = MUX_s_1_2_2(mux_2413_nl, mux_2412_nl, fsm_output[0]);
  assign nor_tmp_538 = or_2486_cse & (fsm_output[8:7]==2'b11);
  assign and_372_nl = or_tmp_29 & (fsm_output[8:7]==2'b11);
  assign mux_tmp_2401 = MUX_s_1_2_2(and_372_nl, and_733_cse, fsm_output[3]);
  assign and_370_nl = (((fsm_output[3]) & (fsm_output[4]) & (fsm_output[6])) | (fsm_output[7]))
      & (fsm_output[8]);
  assign mux_2424_itm = MUX_s_1_2_2(mux_tmp_2384, and_370_nl, fsm_output[5]);
  assign nor_tmp_544 = (fsm_output[4]) & (fsm_output[5]) & (fsm_output[7]) & (fsm_output[8]);
  assign mux_tmp_2410 = MUX_s_1_2_2(mux_tmp_2395, and_dcpl_57, fsm_output[4]);
  assign or_2635_cse = (fsm_output[3]) | (fsm_output[6]);
  assign and_366_nl = or_2635_cse & (fsm_output[8:7]==2'b11);
  assign mux_2433_nl = MUX_s_1_2_2(and_366_nl, mux_tmp_2401, fsm_output[0]);
  assign mux_2434_nl = MUX_s_1_2_2(mux_tmp_2395, mux_2433_nl, fsm_output[4]);
  assign mux_2435_itm = MUX_s_1_2_2(mux_2434_nl, and_733_cse, fsm_output[5]);
  assign nor_tmp_547 = or_36_cse & (fsm_output[8:6]==3'b111);
  assign nor_tmp_548 = or_2612_cse & (fsm_output[8:6]==3'b111);
  assign mux_2440_nl = MUX_s_1_2_2(nor_tmp_339, nor_tmp_547, fsm_output[0]);
  assign mux_2441_nl = MUX_s_1_2_2((~ mux_tmp_2282), mux_2440_nl, fsm_output[4]);
  assign mux_2442_itm = MUX_s_1_2_2(mux_2441_nl, and_dcpl_57, fsm_output[5]);
  assign mux_2443_nl = MUX_s_1_2_2(and_dcpl_57, mux_tmp_2401, fsm_output[4]);
  assign mux_2444_itm = MUX_s_1_2_2(mux_tmp_2410, mux_2443_nl, fsm_output[5]);
  assign not_tmp_762 = ~((fsm_output[4]) | mux_tmp_2282);
  assign mux_2448_nl = MUX_s_1_2_2((~ mux_tmp_2282), mux_tmp_1062, fsm_output[4]);
  assign mux_2449_itm = MUX_s_1_2_2(mux_2448_nl, and_dcpl_57, fsm_output[5]);
  assign or_dcpl_207 = (fsm_output[3]) | (~ (fsm_output[0])) | or_2589_cse;
  assign and_dcpl_277 = nor_1630_cse & (~ (fsm_output[6])) & (fsm_output[1]) & (fsm_output[2])
      & (~ (fsm_output[0])) & and_dcpl_45;
  assign or_tmp_2358 = (~ (fsm_output[8])) | (fsm_output[4]);
  assign or_427_nl = (fsm_output[4]) | (fsm_output[8]);
  assign mux_tmp_2447 = MUX_s_1_2_2(or_tmp_2358, or_427_nl, fsm_output[3]);
  assign nand_tmp_100 = ~((fsm_output[7]) & (~ mux_tmp_2447));
  assign mux_2468_nl = MUX_s_1_2_2(or_610_cse, or_tmp_2358, fsm_output[3]);
  assign or_2571_nl = (fsm_output[7]) | mux_2468_nl;
  assign mux_tmp_2450 = MUX_s_1_2_2(or_2571_nl, nand_tmp_100, fsm_output[2]);
  assign or_tmp_2362 = (fsm_output[6]) | mux_tmp_2450;
  assign and_dcpl_286 = and_dcpl_82 & and_dcpl_66;
  assign or_tmp_2384 = (fsm_output[3]) | or_tmp_29;
  assign STAGE_LOOP_i_3_0_sva_mx0c1 = and_dcpl_58 & and_dcpl_54;
  assign VEC_LOOP_j_10_0_sva_9_0_mx0c0 = and_dcpl_51 & and_dcpl_64;
  assign and_361_nl = (fsm_output[1]) & (fsm_output[6]) & (fsm_output[7]) & (fsm_output[8]);
  assign nor_577_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[8]));
  assign mux_2465_cse = MUX_s_1_2_2(and_361_nl, nor_577_nl, fsm_output[4]);
  assign COMP_LOOP_10_acc_8_itm_mx0c2 = mux_2465_cse & nor_1624_cse & and_dcpl_171;
  assign nand_103_nl = ~((fsm_output[6]) & (~ mux_tmp_2450));
  assign mux_2471_nl = MUX_s_1_2_2(nand_103_nl, or_tmp_2362, fsm_output[1]);
  assign nor_576_nl = ~((fsm_output[5]) | mux_2471_nl);
  assign or_2569_nl = (fsm_output[7]) | mux_tmp_2447;
  assign mux_2467_nl = MUX_s_1_2_2(nand_tmp_100, or_2569_nl, fsm_output[2]);
  assign nand_101_nl = ~((fsm_output[6]) & (~ mux_2467_nl));
  assign mux_2470_nl = MUX_s_1_2_2(or_tmp_2362, nand_101_nl, fsm_output[1]);
  assign and_360_nl = (fsm_output[5]) & (~ mux_2470_nl);
  assign COMP_LOOP_10_acc_8_itm_mx0c3 = MUX_s_1_2_2(nor_576_nl, and_360_nl, fsm_output[0]);
  assign COMP_LOOP_10_acc_8_itm_mx0c6 = and_dcpl_51 & and_dcpl_54;
  assign COMP_LOOP_10_acc_8_itm_mx0c9 = and_dcpl_79 & and_dcpl_196;
  assign COMP_LOOP_10_acc_8_itm_mx0c12 = and_dcpl_79 & and_dcpl_286;
  assign COMP_LOOP_10_acc_8_itm_mx0c15 = and_dcpl_89 & and_dcpl_196;
  assign COMP_LOOP_10_acc_8_itm_mx0c18 = and_dcpl_89 & and_dcpl_286;
  assign COMP_LOOP_10_acc_8_itm_mx0c21 = and_dcpl_97 & and_dcpl_196;
  assign COMP_LOOP_10_acc_8_itm_mx0c24 = and_dcpl_97 & and_dcpl_286;
  assign COMP_LOOP_10_acc_8_itm_mx0c27 = and_dcpl_105 & and_dcpl_196;
  assign COMP_LOOP_10_acc_8_itm_mx0c30 = and_dcpl_105 & and_dcpl_286;
  assign COMP_LOOP_10_acc_8_itm_mx0c33 = and_dcpl_113 & and_dcpl_64;
  assign COMP_LOOP_10_acc_8_itm_mx0c36 = and_dcpl_113 & and_dcpl_69;
  assign COMP_LOOP_10_acc_8_itm_mx0c39 = and_dcpl_121 & and_dcpl_64;
  assign COMP_LOOP_10_acc_8_itm_mx0c42 = and_dcpl_121 & and_dcpl_69;
  assign COMP_LOOP_10_acc_8_itm_mx0c47 = and_dcpl_128 & and_dcpl_69;
  assign nl_STAGE_LOOP_acc_nl = ({1'b1 , (~ z_out_4)}) + 5'b00001;
  assign STAGE_LOOP_acc_nl = nl_STAGE_LOOP_acc_nl[4:0];
  assign STAGE_LOOP_acc_itm_4_1 = readslicef_5_1_4(STAGE_LOOP_acc_nl);
  assign or_44_nl = (fsm_output[3]) | and_674_cse;
  assign mux_27_nl = MUX_s_1_2_2(or_44_nl, or_2259_cse_1, fsm_output[0]);
  assign nor_575_nl = ~((fsm_output[4]) | mux_27_nl);
  assign mux_2498_nl = MUX_s_1_2_2(nor_575_nl, (fsm_output[4]), fsm_output[5]);
  assign and_332_tmp = (~ mux_2498_nl) & and_dcpl_5;
  assign nand_107_nl = ~((fsm_output[2]) & (fsm_output[1]) & (fsm_output[6]));
  assign mux_2507_nl = MUX_s_1_2_2(or_tmp_29, nand_107_nl, fsm_output[3]);
  assign mux_2508_nl = MUX_s_1_2_2(or_tmp_2384, mux_2507_nl, fsm_output[0]);
  assign mux_2509_nl = MUX_s_1_2_2(mux_2508_nl, (~ (fsm_output[6])), or_2589_cse);
  assign and_341_tmp = mux_2509_nl & nor_1630_cse;
  assign mux_2511_nl = MUX_s_1_2_2(or_2635_cse, or_tmp_2384, fsm_output[0]);
  assign nor_570_nl = ~((fsm_output[4]) | mux_2511_nl);
  assign mux_2510_nl = MUX_s_1_2_2(nor_tmp_10, (fsm_output[6]), fsm_output[4]);
  assign mux_2512_nl = MUX_s_1_2_2(nor_570_nl, mux_2510_nl, fsm_output[5]);
  assign and_342_tmp = (~ mux_2512_nl) & nor_1630_cse;
  assign and_354_nl = or_tmp_29 & (fsm_output[7]);
  assign mux_2523_nl = MUX_s_1_2_2(mux_228_cse, and_354_nl, fsm_output[3]);
  assign and_356_nl = or_2697_cse & (fsm_output[7]);
  assign mux_2522_nl = MUX_s_1_2_2(mux_228_cse, and_356_nl, fsm_output[3]);
  assign mux_2524_nl = MUX_s_1_2_2(mux_2523_nl, mux_2522_nl, fsm_output[0]);
  assign mux_2525_nl = MUX_s_1_2_2(mux_2524_nl, (fsm_output[7]), or_2589_cse);
  assign nor_1798_tmp = ~(mux_2525_nl | (fsm_output[8]));
  assign nor_1750_nl = ~((fsm_output[6]) | (fsm_output[1]) | (fsm_output[7]));
  assign mux_234_nl = MUX_s_1_2_2(nor_1750_nl, nor_tmp_47, fsm_output[2]);
  assign mux_2536_nl = MUX_s_1_2_2(nor_572_cse, mux_234_nl, fsm_output[3]);
  assign mux_232_nl = MUX_s_1_2_2(nor_572_cse, nor_tmp_47, or_432_cse);
  assign mux_233_nl = MUX_s_1_2_2(nor_572_cse, mux_232_nl, fsm_output[3]);
  assign mux_2537_nl = MUX_s_1_2_2(mux_2536_nl, mux_233_nl, fsm_output[0]);
  assign mux_2538_nl = MUX_s_1_2_2(mux_2537_nl, nor_tmp_47, or_2589_cse);
  assign nor_1796_tmp = ~(mux_2538_nl | (fsm_output[8]));
  assign or_715_nl = (fsm_output[2]) | (fsm_output[7]) | (~ (fsm_output[5])) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[6]);
  assign mux_1088_nl = MUX_s_1_2_2(or_715_nl, mux_tmp_1067, fsm_output[8]);
  assign or_711_nl = (fsm_output[2]) | (fsm_output[7]) | (fsm_output[5]) | (~ (fsm_output[4]))
      | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[6]);
  assign mux_1087_nl = MUX_s_1_2_2(mux_tmp_1067, or_711_nl, fsm_output[8]);
  assign mux_1089_nl = MUX_s_1_2_2(mux_1088_nl, mux_1087_nl, fsm_output[3]);
  assign vec_rsc_0_0_i_d_d_pff = MUX_v_64_2_2(COMP_LOOP_10_acc_8_itm, COMP_LOOP_1_modulo_cmp_return_rsc_z,
      mux_1089_nl);
  assign and_94_nl = and_dcpl_51 & and_dcpl_67;
  assign and_99_nl = and_dcpl_72 & and_dcpl_47;
  assign and_106_nl = and_dcpl_79 & and_dcpl_77;
  assign and_110_nl = and_dcpl_79 & and_dcpl_83;
  assign and_116_nl = and_dcpl_89 & and_dcpl_77;
  assign and_120_nl = and_dcpl_89 & and_dcpl_83;
  assign and_124_nl = and_dcpl_97 & and_dcpl_77;
  assign and_127_nl = and_dcpl_97 & and_dcpl_83;
  assign and_132_nl = and_dcpl_105 & and_dcpl_77;
  assign and_135_nl = and_dcpl_105 & and_dcpl_83;
  assign and_140_nl = and_dcpl_113 & and_dcpl_111;
  assign and_143_nl = and_dcpl_113 & and_dcpl_54;
  assign and_148_nl = and_dcpl_121 & and_dcpl_111;
  assign and_152_nl = and_dcpl_121 & and_dcpl_54;
  assign and_155_nl = and_dcpl_128 & and_dcpl_111;
  assign vec_rsc_0_0_i_radr_d_pff = MUX1HOT_v_6_32_2((COMP_LOOP_1_acc_10_itm_10_1_1[9:4]),
      COMP_LOOP_acc_psp_sva, (COMP_LOOP_acc_1_cse_2_sva[9:4]), (COMP_LOOP_acc_10_cse_10_1_2_sva[9:4]),
      (COMP_LOOP_acc_11_psp_sva[8:3]), (COMP_LOOP_acc_10_cse_10_1_3_sva[9:4]), (COMP_LOOP_acc_1_cse_4_sva[9:4]),
      (COMP_LOOP_acc_10_cse_10_1_4_sva[9:4]), (COMP_LOOP_acc_13_psp_sva[7:2]), (COMP_LOOP_acc_10_cse_10_1_5_sva[9:4]),
      (COMP_LOOP_acc_1_cse_6_sva[9:4]), (COMP_LOOP_acc_10_cse_10_1_6_sva[9:4]), (COMP_LOOP_acc_14_psp_sva[8:3]),
      (COMP_LOOP_acc_10_cse_10_1_7_sva[9:4]), (COMP_LOOP_acc_1_cse_8_sva[9:4]), (COMP_LOOP_acc_10_cse_10_1_8_sva[9:4]),
      (COMP_LOOP_acc_16_psp_sva[6:1]), (COMP_LOOP_acc_10_cse_10_1_9_sva[9:4]), (COMP_LOOP_acc_1_cse_10_sva[9:4]),
      (COMP_LOOP_acc_10_cse_10_1_10_sva[9:4]), (COMP_LOOP_acc_17_psp_sva[8:3]), (COMP_LOOP_acc_10_cse_10_1_11_sva[9:4]),
      (COMP_LOOP_acc_1_cse_12_sva[9:4]), (COMP_LOOP_acc_10_cse_10_1_12_sva[9:4]),
      (COMP_LOOP_acc_19_psp_sva[7:2]), (COMP_LOOP_acc_10_cse_10_1_13_sva[9:4]), (COMP_LOOP_acc_1_cse_14_sva[9:4]),
      (COMP_LOOP_acc_10_cse_10_1_14_sva[9:4]), (COMP_LOOP_acc_20_psp_sva[8:3]), (COMP_LOOP_acc_10_cse_10_1_15_sva[9:4]),
      (COMP_LOOP_acc_1_cse_sva[9:4]), (COMP_LOOP_acc_10_cse_10_1_sva[9:4]), {and_dcpl_62
      , and_dcpl_65 , and_94_nl , and_dcpl_70 , and_99_nl , and_dcpl_74 , and_106_nl
      , and_dcpl_81 , and_110_nl , and_dcpl_86 , and_116_nl , and_dcpl_93 , and_120_nl
      , and_dcpl_95 , and_124_nl , and_dcpl_100 , and_127_nl , and_dcpl_102 , and_132_nl
      , and_dcpl_108 , and_135_nl , and_dcpl_110 , and_140_nl , and_dcpl_116 , and_143_nl
      , and_dcpl_119 , and_148_nl , and_dcpl_125 , and_152_nl , and_dcpl_127 , and_155_nl
      , and_dcpl_130});
  assign and_158_nl = and_dcpl_131 & and_dcpl_77;
  assign and_159_nl = and_dcpl_51 & and_dcpl_69;
  assign and_160_nl = and_dcpl_131 & and_dcpl_83;
  assign and_161_nl = and_dcpl_131 & and_dcpl_85;
  assign and_163_nl = and_dcpl_136 & and_dcpl_77;
  assign and_164_nl = and_dcpl_79 & and_dcpl_91;
  assign and_165_nl = and_dcpl_136 & and_dcpl_83;
  assign and_166_nl = and_dcpl_136 & and_dcpl_85;
  assign and_168_nl = and_dcpl_141 & and_dcpl_77;
  assign and_169_nl = and_dcpl_89 & and_dcpl_91;
  assign and_170_nl = and_dcpl_141 & and_dcpl_83;
  assign and_171_nl = and_dcpl_141 & and_dcpl_85;
  assign and_173_nl = and_dcpl_146 & and_dcpl_77;
  assign and_174_nl = and_dcpl_97 & and_dcpl_91;
  assign and_175_nl = and_dcpl_146 & and_dcpl_83;
  assign and_176_nl = and_dcpl_146 & and_dcpl_85;
  assign and_178_nl = and_dcpl_151 & and_dcpl_111;
  assign and_179_nl = and_dcpl_105 & and_dcpl_91;
  assign and_180_nl = and_dcpl_151 & and_dcpl_54;
  assign and_181_nl = and_dcpl_151 & and_dcpl_118;
  assign and_183_nl = and_dcpl_156 & and_dcpl_111;
  assign and_184_nl = and_dcpl_113 & and_dcpl_123;
  assign and_185_nl = and_dcpl_156 & and_dcpl_54;
  assign and_186_nl = and_dcpl_156 & and_dcpl_118;
  assign and_188_nl = and_dcpl_161 & and_dcpl_111;
  assign and_189_nl = and_dcpl_121 & and_dcpl_123;
  assign and_190_nl = and_dcpl_161 & and_dcpl_54;
  assign and_191_nl = and_dcpl_161 & and_dcpl_118;
  assign and_193_nl = and_dcpl_166 & and_dcpl_111;
  assign and_194_nl = and_dcpl_128 & and_dcpl_123;
  assign and_195_nl = and_dcpl_166 & and_dcpl_54;
  assign and_196_nl = and_dcpl_166 & and_dcpl_118;
  assign vec_rsc_0_0_i_wadr_d_pff = MUX1HOT_v_6_32_2((COMP_LOOP_acc_10_cse_10_1_1_sva[9:4]),
      COMP_LOOP_acc_psp_sva, (COMP_LOOP_acc_10_cse_10_1_2_sva[9:4]), (COMP_LOOP_acc_1_cse_2_sva[9:4]),
      (COMP_LOOP_acc_10_cse_10_1_3_sva[9:4]), (COMP_LOOP_acc_11_psp_sva[8:3]), (COMP_LOOP_acc_10_cse_10_1_4_sva[9:4]),
      (COMP_LOOP_acc_1_cse_4_sva[9:4]), (COMP_LOOP_acc_10_cse_10_1_5_sva[9:4]), (COMP_LOOP_acc_13_psp_sva[7:2]),
      (COMP_LOOP_acc_10_cse_10_1_6_sva[9:4]), (COMP_LOOP_acc_1_cse_6_sva[9:4]), (COMP_LOOP_acc_10_cse_10_1_7_sva[9:4]),
      (COMP_LOOP_acc_14_psp_sva[8:3]), (COMP_LOOP_acc_10_cse_10_1_8_sva[9:4]), (COMP_LOOP_acc_1_cse_8_sva[9:4]),
      (COMP_LOOP_acc_10_cse_10_1_9_sva[9:4]), (COMP_LOOP_acc_16_psp_sva[6:1]), (COMP_LOOP_acc_10_cse_10_1_10_sva[9:4]),
      (COMP_LOOP_acc_1_cse_10_sva[9:4]), (COMP_LOOP_acc_10_cse_10_1_11_sva[9:4]),
      (COMP_LOOP_acc_17_psp_sva[8:3]), (COMP_LOOP_acc_10_cse_10_1_12_sva[9:4]), (COMP_LOOP_acc_1_cse_12_sva[9:4]),
      (COMP_LOOP_acc_10_cse_10_1_13_sva[9:4]), (COMP_LOOP_acc_19_psp_sva[7:2]), (COMP_LOOP_acc_10_cse_10_1_14_sva[9:4]),
      (COMP_LOOP_acc_1_cse_14_sva[9:4]), (COMP_LOOP_acc_10_cse_10_1_15_sva[9:4]),
      (COMP_LOOP_acc_20_psp_sva[8:3]), (COMP_LOOP_acc_10_cse_10_1_sva[9:4]), (COMP_LOOP_acc_1_cse_sva[9:4]),
      {and_158_nl , and_159_nl , and_160_nl , and_161_nl , and_163_nl , and_164_nl
      , and_165_nl , and_166_nl , and_168_nl , and_169_nl , and_170_nl , and_171_nl
      , and_173_nl , and_174_nl , and_175_nl , and_176_nl , and_178_nl , and_179_nl
      , and_180_nl , and_181_nl , and_183_nl , and_184_nl , and_185_nl , and_186_nl
      , and_188_nl , and_189_nl , and_190_nl , and_191_nl , and_193_nl , and_194_nl
      , and_195_nl , and_196_nl});
  assign nor_1596_nl = ~((~ (fsm_output[5])) | (VEC_LOOP_j_10_0_sva_9_0[3]) | (fsm_output[0])
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[1]) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | (fsm_output[3:2]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2]) | (fsm_output[8:6]!=3'b000));
  assign or_763_nl = (VEC_LOOP_j_10_0_sva_9_0[1]) | mux_1116_cse;
  assign or_757_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000) | nand_324_cse;
  assign or_755_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b000) | (fsm_output[7]) |
      not_tmp_395;
  assign mux_1113_nl = MUX_s_1_2_2(or_757_nl, or_755_nl, fsm_output[2]);
  assign or_753_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000) | (fsm_output[8:6]!=3'b011);
  assign or_752_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000) | (fsm_output[8:6]!=3'b001);
  assign mux_1112_nl = MUX_s_1_2_2(or_753_nl, or_752_nl, fsm_output[2]);
  assign mux_1114_nl = MUX_s_1_2_2(mux_1113_nl, mux_1112_nl, fsm_output[3]);
  assign mux_1117_nl = MUX_s_1_2_2(or_763_nl, mux_1114_nl, fsm_output[1]);
  assign nor_1597_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1117_nl);
  assign nor_1598_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]!=4'b0000) | nand_324_cse);
  assign nor_1599_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b0000) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1109_nl = MUX_s_1_2_2(nor_1598_nl, nor_1599_nl, fsm_output[2]);
  assign nor_1600_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b011));
  assign nor_1601_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b001));
  assign mux_1108_nl = MUX_s_1_2_2(nor_1600_nl, nor_1601_nl, fsm_output[2]);
  assign mux_1110_nl = MUX_s_1_2_2(mux_1109_nl, mux_1108_nl, fsm_output[3]);
  assign nor_1602_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b110));
  assign nor_1603_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b100));
  assign mux_1106_nl = MUX_s_1_2_2(nor_1602_nl, nor_1603_nl, fsm_output[2]);
  assign nor_1604_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b010));
  assign nor_1605_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b000));
  assign mux_1105_nl = MUX_s_1_2_2(nor_1604_nl, nor_1605_nl, fsm_output[2]);
  assign mux_1107_nl = MUX_s_1_2_2(mux_1106_nl, mux_1105_nl, fsm_output[3]);
  assign mux_1111_nl = MUX_s_1_2_2(mux_1110_nl, mux_1107_nl, fsm_output[1]);
  assign mux_1118_nl = MUX_s_1_2_2(nor_1597_nl, mux_1111_nl, fsm_output[0]);
  assign nor_1606_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:0]!=4'b0000) | nand_324_cse);
  assign nor_1607_nl = ~((COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b0000) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1101_nl = MUX_s_1_2_2(nor_1606_nl, nor_1607_nl, fsm_output[2]);
  assign nor_1608_nl = ~((COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b011));
  assign nor_1609_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b001));
  assign mux_1100_nl = MUX_s_1_2_2(nor_1608_nl, nor_1609_nl, fsm_output[2]);
  assign mux_1102_nl = MUX_s_1_2_2(mux_1101_nl, mux_1100_nl, fsm_output[3]);
  assign nor_1610_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b110));
  assign nor_1611_nl = ~((COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b100));
  assign mux_1098_nl = MUX_s_1_2_2(nor_1610_nl, nor_1611_nl, fsm_output[2]);
  assign nor_1612_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b010));
  assign nor_1613_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b000));
  assign mux_1097_nl = MUX_s_1_2_2(nor_1612_nl, nor_1613_nl, fsm_output[2]);
  assign mux_1099_nl = MUX_s_1_2_2(mux_1098_nl, mux_1097_nl, fsm_output[3]);
  assign mux_1103_nl = MUX_s_1_2_2(mux_1102_nl, mux_1099_nl, fsm_output[1]);
  assign nor_1614_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0000) | nand_324_cse);
  assign nor_1615_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0000) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1094_nl = MUX_s_1_2_2(nor_1614_nl, nor_1615_nl, fsm_output[2]);
  assign nor_1616_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b011));
  assign nor_1617_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b001));
  assign mux_1093_nl = MUX_s_1_2_2(nor_1616_nl, nor_1617_nl, fsm_output[2]);
  assign mux_1095_nl = MUX_s_1_2_2(mux_1094_nl, mux_1093_nl, fsm_output[3]);
  assign nor_1618_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b110));
  assign nor_1619_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b100));
  assign mux_1091_nl = MUX_s_1_2_2(nor_1618_nl, nor_1619_nl, fsm_output[2]);
  assign nor_1620_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b010));
  assign nor_1621_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0000) | (fsm_output[8:6]!=3'b000));
  assign mux_1090_nl = MUX_s_1_2_2(nor_1620_nl, nor_1621_nl, fsm_output[2]);
  assign mux_1092_nl = MUX_s_1_2_2(mux_1091_nl, mux_1090_nl, fsm_output[3]);
  assign mux_1096_nl = MUX_s_1_2_2(mux_1095_nl, mux_1092_nl, fsm_output[1]);
  assign mux_1104_nl = MUX_s_1_2_2(mux_1103_nl, mux_1096_nl, fsm_output[0]);
  assign mux_1119_nl = MUX_s_1_2_2(mux_1118_nl, mux_1104_nl, fsm_output[5]);
  assign vec_rsc_0_0_i_we_d_pff = MUX_s_1_2_2(nor_1596_nl, mux_1119_nl, fsm_output[4]);
  assign nor_1569_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[2])) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000) | (~ COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm)
      | nand_301_cse);
  assign nor_1570_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1571_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:0]!=4'b0000) | nand_301_cse);
  assign mux_1146_nl = MUX_s_1_2_2(nor_1570_nl, nor_1571_nl, fsm_output[2]);
  assign nor_1572_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b0000) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1147_nl = MUX_s_1_2_2(mux_1146_nl, nor_1572_nl, fsm_output[5]);
  assign mux_1148_nl = MUX_s_1_2_2(nor_1569_nl, mux_1147_nl, fsm_output[6]);
  assign nor_1573_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b0000) | (fsm_output[7])
      | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1574_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b0000) | nand_301_cse);
  assign mux_1143_nl = MUX_s_1_2_2(nor_1573_nl, nor_1574_nl, fsm_output[2]);
  assign nor_1575_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b0000) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1144_nl = MUX_s_1_2_2(mux_1143_nl, nor_1575_nl, fsm_output[5]);
  assign nor_1576_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1]) | (~ (fsm_output[5])) | (~
      (fsm_output[2])) | (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (~ COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | not_tmp_399);
  assign mux_1145_nl = MUX_s_1_2_2(mux_1144_nl, nor_1576_nl, fsm_output[6]);
  assign mux_1149_nl = MUX_s_1_2_2(mux_1148_nl, mux_1145_nl, fsm_output[1]);
  assign nor_1577_nl = ~((~ (fsm_output[2])) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0000)
      | (~ COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm) | nand_301_cse);
  assign nor_1578_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0000)
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1579_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]!=4'b0000) | nand_301_cse);
  assign mux_1139_nl = MUX_s_1_2_2(nor_1578_nl, nor_1579_nl, fsm_output[2]);
  assign mux_1140_nl = MUX_s_1_2_2(nor_1577_nl, mux_1139_nl, fsm_output[5]);
  assign nor_1580_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b0000) | (fsm_output[5])
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1141_nl = MUX_s_1_2_2(mux_1140_nl, nor_1580_nl, fsm_output[6]);
  assign nor_1581_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1]) | (VEC_LOOP_j_10_0_sva_9_0[3])
      | (fsm_output[5]) | (fsm_output[2]) | (VEC_LOOP_j_10_0_sva_9_0[2]) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1582_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) | (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0000)
      | nand_301_cse);
  assign nor_1583_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm)
      | (fsm_output[7]) | not_tmp_399);
  assign mux_1136_nl = MUX_s_1_2_2(nor_1582_nl, nor_1583_nl, fsm_output[2]);
  assign nor_1584_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b0000) | (~ (fsm_output[2]))
      | (fsm_output[7]) | not_tmp_399);
  assign mux_1137_nl = MUX_s_1_2_2(mux_1136_nl, nor_1584_nl, fsm_output[5]);
  assign mux_1138_nl = MUX_s_1_2_2(nor_1581_nl, mux_1137_nl, fsm_output[6]);
  assign mux_1142_nl = MUX_s_1_2_2(mux_1141_nl, mux_1138_nl, fsm_output[1]);
  assign mux_1150_nl = MUX_s_1_2_2(mux_1149_nl, mux_1142_nl, fsm_output[0]);
  assign nor_1585_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b000) | (~ COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | not_tmp_399);
  assign nor_1586_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[7])) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign mux_1132_nl = MUX_s_1_2_2(nor_1585_nl, nor_1586_nl, fsm_output[2]);
  assign and_561_nl = (fsm_output[5]) & mux_1132_nl;
  assign or_785_nl = (COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b0000) | (fsm_output[7])
      | not_tmp_399;
  assign or_783_nl = (COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b0000) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1131_nl = MUX_s_1_2_2(or_785_nl, or_783_nl, fsm_output[2]);
  assign nor_1587_nl = ~((fsm_output[5]) | mux_1131_nl);
  assign mux_1133_nl = MUX_s_1_2_2(and_561_nl, nor_1587_nl, fsm_output[6]);
  assign or_781_nl = (COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b0000) | (fsm_output[7])
      | not_tmp_399;
  assign or_779_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0000) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1129_nl = MUX_s_1_2_2(or_781_nl, or_779_nl, fsm_output[2]);
  assign nor_1588_nl = ~((fsm_output[5]) | mux_1129_nl);
  assign and_562_nl = nor_346_cse & mux_1128_cse;
  assign mux_1130_nl = MUX_s_1_2_2(nor_1588_nl, and_562_nl, fsm_output[6]);
  assign mux_1134_nl = MUX_s_1_2_2(mux_1133_nl, mux_1130_nl, fsm_output[1]);
  assign or_775_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0000) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7]) | not_tmp_399;
  assign or_773_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0000) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1125_nl = MUX_s_1_2_2(or_775_nl, or_773_nl, fsm_output[2]);
  assign or_772_nl = (COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b0000) | (fsm_output[7])
      | not_tmp_399;
  assign or_770_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0000) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1124_nl = MUX_s_1_2_2(or_772_nl, or_770_nl, fsm_output[2]);
  assign mux_1126_nl = MUX_s_1_2_2(mux_1125_nl, mux_1124_nl, fsm_output[5]);
  assign nor_1591_nl = ~((fsm_output[6]) | mux_1126_nl);
  assign nor_1592_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_1593_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7]) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_1122_nl = MUX_s_1_2_2(nor_1592_nl, nor_1593_nl, fsm_output[2]);
  assign nor_1594_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b0000) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_1595_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0000) | (fsm_output[7])
      | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_1121_nl = MUX_s_1_2_2(nor_1594_nl, nor_1595_nl, fsm_output[2]);
  assign mux_1123_nl = MUX_s_1_2_2(mux_1122_nl, mux_1121_nl, fsm_output[5]);
  assign and_563_nl = (fsm_output[6]) & mux_1123_nl;
  assign mux_1127_nl = MUX_s_1_2_2(nor_1591_nl, and_563_nl, fsm_output[1]);
  assign mux_1135_nl = MUX_s_1_2_2(mux_1134_nl, mux_1127_nl, fsm_output[0]);
  assign vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1150_nl,
      mux_1135_nl, fsm_output[3]);
  assign nor_1539_nl = ~((~ (fsm_output[5])) | (VEC_LOOP_j_10_0_sva_9_0[3]) | (fsm_output[0])
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (fsm_output[1]) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | (fsm_output[3:2]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2]) | (fsm_output[8:6]!=3'b000));
  assign nor_1540_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1]) | mux_1116_cse);
  assign nor_1541_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000) | nand_324_cse);
  assign nor_1542_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b000) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1175_nl = MUX_s_1_2_2(nor_1541_nl, nor_1542_nl, fsm_output[2]);
  assign nor_1543_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000) | (fsm_output[8:6]!=3'b011));
  assign nor_1544_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000) | (fsm_output[8:6]!=3'b001));
  assign mux_1174_nl = MUX_s_1_2_2(nor_1543_nl, nor_1544_nl, fsm_output[2]);
  assign mux_1176_nl = MUX_s_1_2_2(mux_1175_nl, mux_1174_nl, fsm_output[3]);
  assign mux_1179_nl = MUX_s_1_2_2(nor_1540_nl, mux_1176_nl, fsm_output[1]);
  assign and_560_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1179_nl;
  assign nor_1545_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]!=4'b0001) | nand_324_cse);
  assign nor_1546_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b0001) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1171_nl = MUX_s_1_2_2(nor_1545_nl, nor_1546_nl, fsm_output[2]);
  assign nor_1547_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b011));
  assign nor_1548_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b001));
  assign mux_1170_nl = MUX_s_1_2_2(nor_1547_nl, nor_1548_nl, fsm_output[2]);
  assign mux_1172_nl = MUX_s_1_2_2(mux_1171_nl, mux_1170_nl, fsm_output[3]);
  assign nor_1549_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b110));
  assign nor_1550_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b100));
  assign mux_1168_nl = MUX_s_1_2_2(nor_1549_nl, nor_1550_nl, fsm_output[2]);
  assign nor_1551_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b010));
  assign nor_1552_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b000));
  assign mux_1167_nl = MUX_s_1_2_2(nor_1551_nl, nor_1552_nl, fsm_output[2]);
  assign mux_1169_nl = MUX_s_1_2_2(mux_1168_nl, mux_1167_nl, fsm_output[3]);
  assign mux_1173_nl = MUX_s_1_2_2(mux_1172_nl, mux_1169_nl, fsm_output[1]);
  assign mux_1180_nl = MUX_s_1_2_2(and_560_nl, mux_1173_nl, fsm_output[0]);
  assign nor_1553_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:0]!=4'b0001) | nand_324_cse);
  assign mux_1163_nl = MUX_s_1_2_2(nor_1553_nl, nor_1554_cse, fsm_output[2]);
  assign nor_1556_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b001));
  assign mux_1162_nl = MUX_s_1_2_2(nor_1523_cse, nor_1556_nl, fsm_output[2]);
  assign mux_1164_nl = MUX_s_1_2_2(mux_1163_nl, mux_1162_nl, fsm_output[3]);
  assign nor_1557_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b110));
  assign mux_1160_nl = MUX_s_1_2_2(nor_1557_nl, nor_1526_cse, fsm_output[2]);
  assign nor_1560_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b000));
  assign mux_1159_nl = MUX_s_1_2_2(nor_1527_cse, nor_1560_nl, fsm_output[2]);
  assign mux_1161_nl = MUX_s_1_2_2(mux_1160_nl, mux_1159_nl, fsm_output[3]);
  assign mux_1165_nl = MUX_s_1_2_2(mux_1164_nl, mux_1161_nl, fsm_output[1]);
  assign nor_1561_nl = ~((COMP_LOOP_acc_1_cse_sva[3:1]!=3'b000) | nand_272_cse);
  assign nor_1562_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0001) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1156_nl = MUX_s_1_2_2(nor_1561_nl, nor_1562_nl, fsm_output[2]);
  assign nor_1563_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b011));
  assign nor_1564_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b001));
  assign mux_1155_nl = MUX_s_1_2_2(nor_1563_nl, nor_1564_nl, fsm_output[2]);
  assign mux_1157_nl = MUX_s_1_2_2(mux_1156_nl, mux_1155_nl, fsm_output[3]);
  assign nor_1565_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b110));
  assign nor_1566_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b100));
  assign mux_1153_nl = MUX_s_1_2_2(nor_1565_nl, nor_1566_nl, fsm_output[2]);
  assign nor_1567_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b010));
  assign nor_1568_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b000));
  assign mux_1152_nl = MUX_s_1_2_2(nor_1567_nl, nor_1568_nl, fsm_output[2]);
  assign mux_1154_nl = MUX_s_1_2_2(mux_1153_nl, mux_1152_nl, fsm_output[3]);
  assign mux_1158_nl = MUX_s_1_2_2(mux_1157_nl, mux_1154_nl, fsm_output[1]);
  assign mux_1166_nl = MUX_s_1_2_2(mux_1165_nl, mux_1158_nl, fsm_output[0]);
  assign mux_1181_nl = MUX_s_1_2_2(mux_1180_nl, mux_1166_nl, fsm_output[5]);
  assign vec_rsc_0_1_i_we_d_pff = MUX_s_1_2_2(nor_1539_nl, mux_1181_nl, fsm_output[4]);
  assign nor_1506_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000)
      | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) | (fsm_output[2]) | (fsm_output[7])
      | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_1507_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b0001) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_1210_nl = MUX_s_1_2_2(nor_1506_nl, nor_1507_nl, fsm_output[5]);
  assign nor_1508_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b0001) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign nor_1509_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b0001) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1209_nl = MUX_s_1_2_2(nor_1508_nl, nor_1509_nl, fsm_output[5]);
  assign mux_1211_nl = MUX_s_1_2_2(mux_1210_nl, mux_1209_nl, fsm_output[1]);
  assign nor_1510_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b0001) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_1511_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0001)
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1207_nl = MUX_s_1_2_2(nor_1510_nl, nor_1511_nl, fsm_output[5]);
  assign nor_1512_nl = ~((VEC_LOOP_j_10_0_sva_9_0[3]) | (fsm_output[5]) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1208_nl = MUX_s_1_2_2(mux_1207_nl, nor_1512_nl, fsm_output[1]);
  assign mux_1212_nl = MUX_s_1_2_2(mux_1211_nl, mux_1208_nl, fsm_output[0]);
  assign nor_1513_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:0]!=4'b0001) | nand_271_cse);
  assign nor_1514_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[2])) |
      (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000) | (~ COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b110));
  assign mux_1204_nl = MUX_s_1_2_2(nor_1513_nl, nor_1514_nl, fsm_output[5]);
  assign nor_1515_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b0001) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign nor_1516_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (~ (fsm_output[2]))
      | (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (~ COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1203_nl = MUX_s_1_2_2(nor_1515_nl, nor_1516_nl, fsm_output[5]);
  assign mux_1205_nl = MUX_s_1_2_2(mux_1204_nl, mux_1203_nl, fsm_output[1]);
  assign nor_1517_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0001) | (~ COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm)
      | (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign nor_1518_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]!=4'b0001) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign mux_1201_nl = MUX_s_1_2_2(nor_1517_nl, nor_1518_nl, fsm_output[5]);
  assign nor_1519_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) | (COMP_LOOP_acc_1_cse_sva[3:1]!=3'b000)
      | nand_272_cse);
  assign nor_1520_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm)
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1199_nl = MUX_s_1_2_2(nor_1519_nl, nor_1520_nl, fsm_output[2]);
  assign nor_1521_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b0001) | (~ (fsm_output[2]))
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1200_nl = MUX_s_1_2_2(mux_1199_nl, nor_1521_nl, fsm_output[5]);
  assign mux_1202_nl = MUX_s_1_2_2(mux_1201_nl, mux_1200_nl, fsm_output[1]);
  assign mux_1206_nl = MUX_s_1_2_2(mux_1205_nl, mux_1202_nl, fsm_output[0]);
  assign mux_1213_nl = MUX_s_1_2_2(mux_1212_nl, mux_1206_nl, fsm_output[4]);
  assign mux_1195_nl = MUX_s_1_2_2(nor_1554_cse, nor_1523_cse, fsm_output[2]);
  assign nor_1524_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b000) | (~ COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b100));
  assign nor_1525_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b010));
  assign mux_1194_nl = MUX_s_1_2_2(nor_1524_nl, nor_1525_nl, fsm_output[2]);
  assign and_558_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1194_nl;
  assign mux_1196_nl = MUX_s_1_2_2(mux_1195_nl, and_558_nl, fsm_output[5]);
  assign mux_1192_nl = MUX_s_1_2_2(nor_1526_cse, nor_1527_cse, fsm_output[2]);
  assign and_559_nl = nor_351_cse & mux_1191_cse;
  assign mux_1193_nl = MUX_s_1_2_2(mux_1192_nl, and_559_nl, fsm_output[5]);
  assign mux_1197_nl = MUX_s_1_2_2(mux_1196_nl, mux_1193_nl, fsm_output[1]);
  assign nor_1531_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0001) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b100));
  assign nor_1532_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0001) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b010));
  assign mux_1187_nl = MUX_s_1_2_2(nor_1531_nl, nor_1532_nl, fsm_output[2]);
  assign nor_1533_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b100));
  assign nor_1534_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b010));
  assign mux_1186_nl = MUX_s_1_2_2(nor_1533_nl, nor_1534_nl, fsm_output[2]);
  assign mux_1188_nl = MUX_s_1_2_2(mux_1187_nl, mux_1186_nl, fsm_output[5]);
  assign nor_1535_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | (fsm_output[8:6]!=3'b011));
  assign nor_1536_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[8:6]!=3'b001));
  assign mux_1184_nl = MUX_s_1_2_2(nor_1535_nl, nor_1536_nl, fsm_output[2]);
  assign nor_1537_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b011));
  assign nor_1538_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0001) | (fsm_output[8:6]!=3'b001));
  assign mux_1183_nl = MUX_s_1_2_2(nor_1537_nl, nor_1538_nl, fsm_output[2]);
  assign mux_1185_nl = MUX_s_1_2_2(mux_1184_nl, mux_1183_nl, fsm_output[5]);
  assign mux_1189_nl = MUX_s_1_2_2(mux_1188_nl, mux_1185_nl, fsm_output[1]);
  assign mux_1198_nl = MUX_s_1_2_2(mux_1197_nl, mux_1189_nl, fsm_output[0]);
  assign and_557_nl = (fsm_output[4]) & mux_1198_nl;
  assign vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1213_nl,
      and_557_nl, fsm_output[3]);
  assign nor_1477_nl = ~((~ (fsm_output[5])) | (VEC_LOOP_j_10_0_sva_9_0[3]) | (fsm_output[0])
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[1]) | (~ (VEC_LOOP_j_10_0_sva_9_0[1]))
      | (fsm_output[3:2]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2]) | (fsm_output[8:6]!=3'b000));
  assign nand_31_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1]) & mux_1241_cse);
  assign or_952_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001) | nand_324_cse;
  assign or_950_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b001) | (fsm_output[7]) |
      not_tmp_395;
  assign mux_1238_nl = MUX_s_1_2_2(or_952_nl, or_950_nl, fsm_output[2]);
  assign or_948_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001) | (fsm_output[8:6]!=3'b011);
  assign or_947_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001) | (fsm_output[8:6]!=3'b001);
  assign mux_1237_nl = MUX_s_1_2_2(or_948_nl, or_947_nl, fsm_output[2]);
  assign mux_1239_nl = MUX_s_1_2_2(mux_1238_nl, mux_1237_nl, fsm_output[3]);
  assign mux_1242_nl = MUX_s_1_2_2(nand_31_nl, mux_1239_nl, fsm_output[1]);
  assign nor_1478_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1242_nl);
  assign nor_1482_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[2]) | (COMP_LOOP_acc_10_cse_10_1_15_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_15_sva[0]) | nand_268_cse);
  assign nor_1483_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b0010) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1234_nl = MUX_s_1_2_2(nor_1482_nl, nor_1483_nl, fsm_output[2]);
  assign nor_1484_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b011));
  assign nor_1485_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b001));
  assign mux_1233_nl = MUX_s_1_2_2(nor_1484_nl, nor_1485_nl, fsm_output[2]);
  assign mux_1235_nl = MUX_s_1_2_2(mux_1234_nl, mux_1233_nl, fsm_output[3]);
  assign nor_1486_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b110));
  assign nor_1487_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b100));
  assign mux_1231_nl = MUX_s_1_2_2(nor_1486_nl, nor_1487_nl, fsm_output[2]);
  assign nor_1488_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b010));
  assign nor_1489_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b000));
  assign mux_1230_nl = MUX_s_1_2_2(nor_1488_nl, nor_1489_nl, fsm_output[2]);
  assign mux_1232_nl = MUX_s_1_2_2(mux_1231_nl, mux_1230_nl, fsm_output[3]);
  assign mux_1236_nl = MUX_s_1_2_2(mux_1235_nl, mux_1232_nl, fsm_output[1]);
  assign mux_1243_nl = MUX_s_1_2_2(nor_1478_nl, mux_1236_nl, fsm_output[0]);
  assign nor_1490_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:0]!=4'b0010) | nand_324_cse);
  assign nor_1491_nl = ~((COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b0010) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1226_nl = MUX_s_1_2_2(nor_1490_nl, nor_1491_nl, fsm_output[2]);
  assign nor_1492_nl = ~((COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b011));
  assign nor_1493_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b001));
  assign mux_1225_nl = MUX_s_1_2_2(nor_1492_nl, nor_1493_nl, fsm_output[2]);
  assign mux_1227_nl = MUX_s_1_2_2(mux_1226_nl, mux_1225_nl, fsm_output[3]);
  assign nor_1494_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b110));
  assign nor_1495_nl = ~((COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b100));
  assign mux_1223_nl = MUX_s_1_2_2(nor_1494_nl, nor_1495_nl, fsm_output[2]);
  assign nor_1496_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b010));
  assign nor_1497_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b000));
  assign mux_1222_nl = MUX_s_1_2_2(nor_1496_nl, nor_1497_nl, fsm_output[2]);
  assign mux_1224_nl = MUX_s_1_2_2(mux_1223_nl, mux_1222_nl, fsm_output[3]);
  assign mux_1228_nl = MUX_s_1_2_2(mux_1227_nl, mux_1224_nl, fsm_output[1]);
  assign nor_1498_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0010) | nand_324_cse);
  assign nor_1499_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0010) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1219_nl = MUX_s_1_2_2(nor_1498_nl, nor_1499_nl, fsm_output[2]);
  assign nor_1500_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b011));
  assign nor_1501_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b001));
  assign mux_1218_nl = MUX_s_1_2_2(nor_1500_nl, nor_1501_nl, fsm_output[2]);
  assign mux_1220_nl = MUX_s_1_2_2(mux_1219_nl, mux_1218_nl, fsm_output[3]);
  assign nor_1502_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b110));
  assign nor_1503_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b100));
  assign mux_1216_nl = MUX_s_1_2_2(nor_1502_nl, nor_1503_nl, fsm_output[2]);
  assign nor_1504_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b010));
  assign nor_1505_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0010) | (fsm_output[8:6]!=3'b000));
  assign mux_1215_nl = MUX_s_1_2_2(nor_1504_nl, nor_1505_nl, fsm_output[2]);
  assign mux_1217_nl = MUX_s_1_2_2(mux_1216_nl, mux_1215_nl, fsm_output[3]);
  assign mux_1221_nl = MUX_s_1_2_2(mux_1220_nl, mux_1217_nl, fsm_output[1]);
  assign mux_1229_nl = MUX_s_1_2_2(mux_1228_nl, mux_1221_nl, fsm_output[0]);
  assign mux_1244_nl = MUX_s_1_2_2(mux_1243_nl, mux_1229_nl, fsm_output[5]);
  assign vec_rsc_0_2_i_we_d_pff = MUX_s_1_2_2(nor_1477_nl, mux_1244_nl, fsm_output[4]);
  assign nor_1450_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[2])) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001) | (~ COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm)
      | nand_301_cse);
  assign nor_1451_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1452_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:0]!=4'b0010) | nand_301_cse);
  assign mux_1271_nl = MUX_s_1_2_2(nor_1451_nl, nor_1452_nl, fsm_output[2]);
  assign nor_1453_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b0010) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1272_nl = MUX_s_1_2_2(mux_1271_nl, nor_1453_nl, fsm_output[5]);
  assign mux_1273_nl = MUX_s_1_2_2(nor_1450_nl, mux_1272_nl, fsm_output[6]);
  assign nor_1454_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b0010) | (fsm_output[7])
      | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1455_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b0010) | nand_301_cse);
  assign mux_1268_nl = MUX_s_1_2_2(nor_1454_nl, nor_1455_nl, fsm_output[2]);
  assign nor_1456_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b0010) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1269_nl = MUX_s_1_2_2(mux_1268_nl, nor_1456_nl, fsm_output[5]);
  assign nor_1457_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[1])) | (~ (fsm_output[5])) |
      (~ (fsm_output[2])) | (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (~ COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | not_tmp_399);
  assign mux_1270_nl = MUX_s_1_2_2(mux_1269_nl, nor_1457_nl, fsm_output[6]);
  assign mux_1274_nl = MUX_s_1_2_2(mux_1273_nl, mux_1270_nl, fsm_output[1]);
  assign nor_1458_nl = ~((~ (fsm_output[2])) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0010)
      | (~ COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm) | nand_301_cse);
  assign nor_1459_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0010)
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1460_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[2]) | (COMP_LOOP_acc_10_cse_10_1_15_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_15_sva[0]) | nand_265_cse);
  assign mux_1264_nl = MUX_s_1_2_2(nor_1459_nl, nor_1460_nl, fsm_output[2]);
  assign mux_1265_nl = MUX_s_1_2_2(nor_1458_nl, mux_1264_nl, fsm_output[5]);
  assign nor_1461_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b0010) | (fsm_output[5])
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1266_nl = MUX_s_1_2_2(mux_1265_nl, nor_1461_nl, fsm_output[6]);
  assign nor_1462_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[1])) | (VEC_LOOP_j_10_0_sva_9_0[3])
      | (fsm_output[5]) | (fsm_output[2]) | (VEC_LOOP_j_10_0_sva_9_0[2]) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1463_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) | (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0010)
      | nand_301_cse);
  assign nor_1464_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm)
      | (fsm_output[7]) | not_tmp_399);
  assign mux_1261_nl = MUX_s_1_2_2(nor_1463_nl, nor_1464_nl, fsm_output[2]);
  assign nor_1465_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b0010) | (~ (fsm_output[2]))
      | (fsm_output[7]) | not_tmp_399);
  assign mux_1262_nl = MUX_s_1_2_2(mux_1261_nl, nor_1465_nl, fsm_output[5]);
  assign mux_1263_nl = MUX_s_1_2_2(nor_1462_nl, mux_1262_nl, fsm_output[6]);
  assign mux_1267_nl = MUX_s_1_2_2(mux_1266_nl, mux_1263_nl, fsm_output[1]);
  assign mux_1275_nl = MUX_s_1_2_2(mux_1274_nl, mux_1267_nl, fsm_output[0]);
  assign nor_1466_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b001) | (~ COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | not_tmp_399);
  assign nor_1467_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[7])) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign mux_1257_nl = MUX_s_1_2_2(nor_1466_nl, nor_1467_nl, fsm_output[2]);
  assign and_554_nl = (fsm_output[5]) & mux_1257_nl;
  assign or_979_nl = (COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b0010) | (fsm_output[7])
      | not_tmp_399;
  assign or_977_nl = (COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b0010) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1256_nl = MUX_s_1_2_2(or_979_nl, or_977_nl, fsm_output[2]);
  assign nor_1468_nl = ~((fsm_output[5]) | mux_1256_nl);
  assign mux_1258_nl = MUX_s_1_2_2(and_554_nl, nor_1468_nl, fsm_output[6]);
  assign or_975_nl = (COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b0010) | (fsm_output[7])
      | not_tmp_399;
  assign or_973_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0010) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1254_nl = MUX_s_1_2_2(or_975_nl, or_973_nl, fsm_output[2]);
  assign nor_1469_nl = ~((fsm_output[5]) | mux_1254_nl);
  assign and_555_nl = (VEC_LOOP_j_10_0_sva_9_0[1]) & (fsm_output[5]) & mux_1128_cse;
  assign mux_1255_nl = MUX_s_1_2_2(nor_1469_nl, and_555_nl, fsm_output[6]);
  assign mux_1259_nl = MUX_s_1_2_2(mux_1258_nl, mux_1255_nl, fsm_output[1]);
  assign or_969_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0010) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7]) | not_tmp_399;
  assign or_967_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0010) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1250_nl = MUX_s_1_2_2(or_969_nl, or_967_nl, fsm_output[2]);
  assign or_966_nl = (COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b0010) | (fsm_output[7])
      | not_tmp_399;
  assign or_964_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0010) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1249_nl = MUX_s_1_2_2(or_966_nl, or_964_nl, fsm_output[2]);
  assign mux_1251_nl = MUX_s_1_2_2(mux_1250_nl, mux_1249_nl, fsm_output[5]);
  assign nor_1472_nl = ~((fsm_output[6]) | mux_1251_nl);
  assign nor_1473_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_1474_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7]) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_1247_nl = MUX_s_1_2_2(nor_1473_nl, nor_1474_nl, fsm_output[2]);
  assign nor_1475_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b0010) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_1476_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0010) | (fsm_output[7])
      | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_1246_nl = MUX_s_1_2_2(nor_1475_nl, nor_1476_nl, fsm_output[2]);
  assign mux_1248_nl = MUX_s_1_2_2(mux_1247_nl, mux_1246_nl, fsm_output[5]);
  assign and_556_nl = (fsm_output[6]) & mux_1248_nl;
  assign mux_1252_nl = MUX_s_1_2_2(nor_1472_nl, and_556_nl, fsm_output[1]);
  assign mux_1260_nl = MUX_s_1_2_2(mux_1259_nl, mux_1252_nl, fsm_output[0]);
  assign vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1275_nl,
      mux_1260_nl, fsm_output[3]);
  assign nor_1418_nl = ~((~ (fsm_output[5])) | (VEC_LOOP_j_10_0_sva_9_0[3]) | (fsm_output[0])
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (fsm_output[1]) | (~ (VEC_LOOP_j_10_0_sva_9_0[1]))
      | (fsm_output[3:2]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2]) | (fsm_output[8:6]!=3'b000));
  assign and_553_nl = (VEC_LOOP_j_10_0_sva_9_0[1]) & mux_1241_cse;
  assign nor_1422_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001) | nand_324_cse);
  assign nor_1423_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b001) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1300_nl = MUX_s_1_2_2(nor_1422_nl, nor_1423_nl, fsm_output[2]);
  assign nor_1424_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001) | (fsm_output[8:6]!=3'b011));
  assign nor_1425_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001) | (fsm_output[8:6]!=3'b001));
  assign mux_1299_nl = MUX_s_1_2_2(nor_1424_nl, nor_1425_nl, fsm_output[2]);
  assign mux_1301_nl = MUX_s_1_2_2(mux_1300_nl, mux_1299_nl, fsm_output[3]);
  assign mux_1304_nl = MUX_s_1_2_2(and_553_nl, mux_1301_nl, fsm_output[1]);
  assign and_552_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1304_nl;
  assign nor_1426_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:2]!=2'b00) | nand_261_cse);
  assign nor_1427_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b0011) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1296_nl = MUX_s_1_2_2(nor_1426_nl, nor_1427_nl, fsm_output[2]);
  assign nor_1428_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b011));
  assign nor_1429_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b001));
  assign mux_1295_nl = MUX_s_1_2_2(nor_1428_nl, nor_1429_nl, fsm_output[2]);
  assign mux_1297_nl = MUX_s_1_2_2(mux_1296_nl, mux_1295_nl, fsm_output[3]);
  assign nor_1430_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b110));
  assign nor_1431_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b100));
  assign mux_1293_nl = MUX_s_1_2_2(nor_1430_nl, nor_1431_nl, fsm_output[2]);
  assign nor_1432_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b010));
  assign nor_1433_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b000));
  assign mux_1292_nl = MUX_s_1_2_2(nor_1432_nl, nor_1433_nl, fsm_output[2]);
  assign mux_1294_nl = MUX_s_1_2_2(mux_1293_nl, mux_1292_nl, fsm_output[3]);
  assign mux_1298_nl = MUX_s_1_2_2(mux_1297_nl, mux_1294_nl, fsm_output[1]);
  assign mux_1305_nl = MUX_s_1_2_2(and_552_nl, mux_1298_nl, fsm_output[0]);
  assign nor_1434_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:0]!=4'b0011) | nand_324_cse);
  assign mux_1288_nl = MUX_s_1_2_2(nor_1434_nl, nor_1435_cse, fsm_output[2]);
  assign nor_1437_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b001));
  assign mux_1287_nl = MUX_s_1_2_2(nor_1402_cse, nor_1437_nl, fsm_output[2]);
  assign mux_1289_nl = MUX_s_1_2_2(mux_1288_nl, mux_1287_nl, fsm_output[3]);
  assign nor_1438_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b110));
  assign mux_1285_nl = MUX_s_1_2_2(nor_1438_nl, nor_1405_cse, fsm_output[2]);
  assign nor_1441_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b000));
  assign mux_1284_nl = MUX_s_1_2_2(nor_1406_cse, nor_1441_nl, fsm_output[2]);
  assign mux_1286_nl = MUX_s_1_2_2(mux_1285_nl, mux_1284_nl, fsm_output[3]);
  assign mux_1290_nl = MUX_s_1_2_2(mux_1289_nl, mux_1286_nl, fsm_output[1]);
  assign nor_1442_nl = ~((COMP_LOOP_acc_1_cse_sva[3:1]!=3'b001) | nand_272_cse);
  assign nor_1443_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0011) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1281_nl = MUX_s_1_2_2(nor_1442_nl, nor_1443_nl, fsm_output[2]);
  assign nor_1444_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b011));
  assign nor_1445_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b001));
  assign mux_1280_nl = MUX_s_1_2_2(nor_1444_nl, nor_1445_nl, fsm_output[2]);
  assign mux_1282_nl = MUX_s_1_2_2(mux_1281_nl, mux_1280_nl, fsm_output[3]);
  assign nor_1446_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b110));
  assign nor_1447_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b100));
  assign mux_1278_nl = MUX_s_1_2_2(nor_1446_nl, nor_1447_nl, fsm_output[2]);
  assign nor_1448_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b010));
  assign nor_1449_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b000));
  assign mux_1277_nl = MUX_s_1_2_2(nor_1448_nl, nor_1449_nl, fsm_output[2]);
  assign mux_1279_nl = MUX_s_1_2_2(mux_1278_nl, mux_1277_nl, fsm_output[3]);
  assign mux_1283_nl = MUX_s_1_2_2(mux_1282_nl, mux_1279_nl, fsm_output[1]);
  assign mux_1291_nl = MUX_s_1_2_2(mux_1290_nl, mux_1283_nl, fsm_output[0]);
  assign mux_1306_nl = MUX_s_1_2_2(mux_1305_nl, mux_1291_nl, fsm_output[5]);
  assign vec_rsc_0_3_i_we_d_pff = MUX_s_1_2_2(nor_1418_nl, mux_1306_nl, fsm_output[4]);
  assign nor_1385_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001)
      | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) | (fsm_output[2]) | (fsm_output[7])
      | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_1386_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b0011) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_1335_nl = MUX_s_1_2_2(nor_1385_nl, nor_1386_nl, fsm_output[5]);
  assign nor_1387_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b0011) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign nor_1388_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b0011) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1334_nl = MUX_s_1_2_2(nor_1387_nl, nor_1388_nl, fsm_output[5]);
  assign mux_1336_nl = MUX_s_1_2_2(mux_1335_nl, mux_1334_nl, fsm_output[1]);
  assign nor_1389_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b0011) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_1390_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0011)
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1332_nl = MUX_s_1_2_2(nor_1389_nl, nor_1390_nl, fsm_output[5]);
  assign nor_1391_nl = ~((VEC_LOOP_j_10_0_sva_9_0[3]) | (fsm_output[5]) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1333_nl = MUX_s_1_2_2(mux_1332_nl, nor_1391_nl, fsm_output[1]);
  assign mux_1337_nl = MUX_s_1_2_2(mux_1336_nl, mux_1333_nl, fsm_output[0]);
  assign nor_1392_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:0]!=4'b0011) | nand_271_cse);
  assign nor_1393_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[2])) |
      (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001) | (~ COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b110));
  assign mux_1329_nl = MUX_s_1_2_2(nor_1392_nl, nor_1393_nl, fsm_output[5]);
  assign nor_1394_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b0011) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign nor_1395_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b11) | (~ (fsm_output[2]))
      | (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (~ COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1328_nl = MUX_s_1_2_2(nor_1394_nl, nor_1395_nl, fsm_output[5]);
  assign mux_1330_nl = MUX_s_1_2_2(mux_1329_nl, mux_1328_nl, fsm_output[1]);
  assign nor_1396_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0011) | (~ COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm)
      | (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign nor_1397_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]!=4'b0011) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign mux_1326_nl = MUX_s_1_2_2(nor_1396_nl, nor_1397_nl, fsm_output[5]);
  assign nor_1398_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) | (COMP_LOOP_acc_1_cse_sva[3:1]!=3'b001)
      | nand_272_cse);
  assign nor_1399_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm)
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1324_nl = MUX_s_1_2_2(nor_1398_nl, nor_1399_nl, fsm_output[2]);
  assign nor_1400_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b0011) | (~ (fsm_output[2]))
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1325_nl = MUX_s_1_2_2(mux_1324_nl, nor_1400_nl, fsm_output[5]);
  assign mux_1327_nl = MUX_s_1_2_2(mux_1326_nl, mux_1325_nl, fsm_output[1]);
  assign mux_1331_nl = MUX_s_1_2_2(mux_1330_nl, mux_1327_nl, fsm_output[0]);
  assign mux_1338_nl = MUX_s_1_2_2(mux_1337_nl, mux_1331_nl, fsm_output[4]);
  assign mux_1320_nl = MUX_s_1_2_2(nor_1435_cse, nor_1402_cse, fsm_output[2]);
  assign nor_1403_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b001) | (~ COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b100));
  assign nor_1404_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b010));
  assign mux_1319_nl = MUX_s_1_2_2(nor_1403_nl, nor_1404_nl, fsm_output[2]);
  assign and_550_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1319_nl;
  assign mux_1321_nl = MUX_s_1_2_2(mux_1320_nl, and_550_nl, fsm_output[5]);
  assign mux_1317_nl = MUX_s_1_2_2(nor_1405_cse, nor_1406_cse, fsm_output[2]);
  assign and_551_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & mux_1191_cse;
  assign mux_1318_nl = MUX_s_1_2_2(mux_1317_nl, and_551_nl, fsm_output[5]);
  assign mux_1322_nl = MUX_s_1_2_2(mux_1321_nl, mux_1318_nl, fsm_output[1]);
  assign nor_1410_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0011) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b100));
  assign nor_1411_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0011) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b010));
  assign mux_1312_nl = MUX_s_1_2_2(nor_1410_nl, nor_1411_nl, fsm_output[2]);
  assign nor_1412_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b100));
  assign nor_1413_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b010));
  assign mux_1311_nl = MUX_s_1_2_2(nor_1412_nl, nor_1413_nl, fsm_output[2]);
  assign mux_1313_nl = MUX_s_1_2_2(mux_1312_nl, mux_1311_nl, fsm_output[5]);
  assign nor_1414_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | (fsm_output[8:6]!=3'b011));
  assign nor_1415_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[8:6]!=3'b001));
  assign mux_1309_nl = MUX_s_1_2_2(nor_1414_nl, nor_1415_nl, fsm_output[2]);
  assign nor_1416_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b011));
  assign nor_1417_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0011) | (fsm_output[8:6]!=3'b001));
  assign mux_1308_nl = MUX_s_1_2_2(nor_1416_nl, nor_1417_nl, fsm_output[2]);
  assign mux_1310_nl = MUX_s_1_2_2(mux_1309_nl, mux_1308_nl, fsm_output[5]);
  assign mux_1314_nl = MUX_s_1_2_2(mux_1313_nl, mux_1310_nl, fsm_output[1]);
  assign mux_1323_nl = MUX_s_1_2_2(mux_1322_nl, mux_1314_nl, fsm_output[0]);
  assign and_549_nl = (fsm_output[4]) & mux_1323_nl;
  assign vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1338_nl,
      and_549_nl, fsm_output[3]);
  assign nor_1359_nl = ~((~ (fsm_output[5])) | (VEC_LOOP_j_10_0_sva_9_0[3]) | (fsm_output[0])
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[1]) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | (fsm_output[3:2]!=2'b00) | (~ (VEC_LOOP_j_10_0_sva_9_0[2])) | (fsm_output[8:6]!=3'b000));
  assign or_1151_nl = (VEC_LOOP_j_10_0_sva_9_0[1]) | mux_1366_cse;
  assign or_1145_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010) | nand_324_cse;
  assign or_1143_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b010) | (fsm_output[7]) |
      not_tmp_395;
  assign mux_1363_nl = MUX_s_1_2_2(or_1145_nl, or_1143_nl, fsm_output[2]);
  assign or_1141_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010) | (fsm_output[8:6]!=3'b011);
  assign or_1140_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010) | (fsm_output[8:6]!=3'b001);
  assign mux_1362_nl = MUX_s_1_2_2(or_1141_nl, or_1140_nl, fsm_output[2]);
  assign mux_1364_nl = MUX_s_1_2_2(mux_1363_nl, mux_1362_nl, fsm_output[3]);
  assign mux_1367_nl = MUX_s_1_2_2(or_1151_nl, mux_1364_nl, fsm_output[1]);
  assign nor_1360_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1367_nl);
  assign nor_1361_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]!=4'b0100) | nand_324_cse);
  assign nor_1362_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b0100) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1359_nl = MUX_s_1_2_2(nor_1361_nl, nor_1362_nl, fsm_output[2]);
  assign nor_1363_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b011));
  assign nor_1364_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b001));
  assign mux_1358_nl = MUX_s_1_2_2(nor_1363_nl, nor_1364_nl, fsm_output[2]);
  assign mux_1360_nl = MUX_s_1_2_2(mux_1359_nl, mux_1358_nl, fsm_output[3]);
  assign nor_1365_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b110));
  assign nor_1366_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b100));
  assign mux_1356_nl = MUX_s_1_2_2(nor_1365_nl, nor_1366_nl, fsm_output[2]);
  assign nor_1367_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b010));
  assign nor_1368_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b000));
  assign mux_1355_nl = MUX_s_1_2_2(nor_1367_nl, nor_1368_nl, fsm_output[2]);
  assign mux_1357_nl = MUX_s_1_2_2(mux_1356_nl, mux_1355_nl, fsm_output[3]);
  assign mux_1361_nl = MUX_s_1_2_2(mux_1360_nl, mux_1357_nl, fsm_output[1]);
  assign mux_1368_nl = MUX_s_1_2_2(nor_1360_nl, mux_1361_nl, fsm_output[0]);
  assign nor_1369_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:0]!=4'b0100) | nand_324_cse);
  assign nor_1370_nl = ~((COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b0100) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1351_nl = MUX_s_1_2_2(nor_1369_nl, nor_1370_nl, fsm_output[2]);
  assign nor_1371_nl = ~((COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b011));
  assign nor_1372_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b001));
  assign mux_1350_nl = MUX_s_1_2_2(nor_1371_nl, nor_1372_nl, fsm_output[2]);
  assign mux_1352_nl = MUX_s_1_2_2(mux_1351_nl, mux_1350_nl, fsm_output[3]);
  assign nor_1373_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b110));
  assign nor_1374_nl = ~((COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b100));
  assign mux_1348_nl = MUX_s_1_2_2(nor_1373_nl, nor_1374_nl, fsm_output[2]);
  assign nor_1375_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b010));
  assign nor_1376_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b000));
  assign mux_1347_nl = MUX_s_1_2_2(nor_1375_nl, nor_1376_nl, fsm_output[2]);
  assign mux_1349_nl = MUX_s_1_2_2(mux_1348_nl, mux_1347_nl, fsm_output[3]);
  assign mux_1353_nl = MUX_s_1_2_2(mux_1352_nl, mux_1349_nl, fsm_output[1]);
  assign nor_1377_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0100) | nand_324_cse);
  assign nor_1378_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0100) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1344_nl = MUX_s_1_2_2(nor_1377_nl, nor_1378_nl, fsm_output[2]);
  assign nor_1379_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b011));
  assign nor_1380_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b001));
  assign mux_1343_nl = MUX_s_1_2_2(nor_1379_nl, nor_1380_nl, fsm_output[2]);
  assign mux_1345_nl = MUX_s_1_2_2(mux_1344_nl, mux_1343_nl, fsm_output[3]);
  assign nor_1381_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b110));
  assign nor_1382_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b100));
  assign mux_1341_nl = MUX_s_1_2_2(nor_1381_nl, nor_1382_nl, fsm_output[2]);
  assign nor_1383_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b010));
  assign nor_1384_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0100) | (fsm_output[8:6]!=3'b000));
  assign mux_1340_nl = MUX_s_1_2_2(nor_1383_nl, nor_1384_nl, fsm_output[2]);
  assign mux_1342_nl = MUX_s_1_2_2(mux_1341_nl, mux_1340_nl, fsm_output[3]);
  assign mux_1346_nl = MUX_s_1_2_2(mux_1345_nl, mux_1342_nl, fsm_output[1]);
  assign mux_1354_nl = MUX_s_1_2_2(mux_1353_nl, mux_1346_nl, fsm_output[0]);
  assign mux_1369_nl = MUX_s_1_2_2(mux_1368_nl, mux_1354_nl, fsm_output[5]);
  assign vec_rsc_0_4_i_we_d_pff = MUX_s_1_2_2(nor_1359_nl, mux_1369_nl, fsm_output[4]);
  assign nor_1332_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[2])) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010) | (~ COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm)
      | nand_301_cse);
  assign nor_1333_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1334_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:0]!=4'b0100) | nand_301_cse);
  assign mux_1396_nl = MUX_s_1_2_2(nor_1333_nl, nor_1334_nl, fsm_output[2]);
  assign nor_1335_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b0100) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1397_nl = MUX_s_1_2_2(mux_1396_nl, nor_1335_nl, fsm_output[5]);
  assign mux_1398_nl = MUX_s_1_2_2(nor_1332_nl, mux_1397_nl, fsm_output[6]);
  assign nor_1336_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b0100) | (fsm_output[7])
      | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1337_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b0100) | nand_301_cse);
  assign mux_1393_nl = MUX_s_1_2_2(nor_1336_nl, nor_1337_nl, fsm_output[2]);
  assign nor_1338_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b0100) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1394_nl = MUX_s_1_2_2(mux_1393_nl, nor_1338_nl, fsm_output[5]);
  assign nor_1339_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1]) | (~ (fsm_output[5])) | (~
      (fsm_output[2])) | (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (~ COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | not_tmp_399);
  assign mux_1395_nl = MUX_s_1_2_2(mux_1394_nl, nor_1339_nl, fsm_output[6]);
  assign mux_1399_nl = MUX_s_1_2_2(mux_1398_nl, mux_1395_nl, fsm_output[1]);
  assign nor_1340_nl = ~((~ (fsm_output[2])) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0100)
      | (~ COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm) | nand_301_cse);
  assign nor_1341_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0100)
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1342_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]!=4'b0100) | nand_301_cse);
  assign mux_1389_nl = MUX_s_1_2_2(nor_1341_nl, nor_1342_nl, fsm_output[2]);
  assign mux_1390_nl = MUX_s_1_2_2(nor_1340_nl, mux_1389_nl, fsm_output[5]);
  assign nor_1343_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b0100) | (fsm_output[5])
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1391_nl = MUX_s_1_2_2(mux_1390_nl, nor_1343_nl, fsm_output[6]);
  assign nor_1344_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1]) | (VEC_LOOP_j_10_0_sva_9_0[3])
      | (fsm_output[5]) | (fsm_output[2]) | (~ (VEC_LOOP_j_10_0_sva_9_0[2])) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1345_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) | (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0100)
      | nand_301_cse);
  assign nor_1346_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm)
      | (fsm_output[7]) | not_tmp_399);
  assign mux_1386_nl = MUX_s_1_2_2(nor_1345_nl, nor_1346_nl, fsm_output[2]);
  assign nor_1347_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b0100) | (~ (fsm_output[2]))
      | (fsm_output[7]) | not_tmp_399);
  assign mux_1387_nl = MUX_s_1_2_2(mux_1386_nl, nor_1347_nl, fsm_output[5]);
  assign mux_1388_nl = MUX_s_1_2_2(nor_1344_nl, mux_1387_nl, fsm_output[6]);
  assign mux_1392_nl = MUX_s_1_2_2(mux_1391_nl, mux_1388_nl, fsm_output[1]);
  assign mux_1400_nl = MUX_s_1_2_2(mux_1399_nl, mux_1392_nl, fsm_output[0]);
  assign nor_1348_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b010) | (~ COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | not_tmp_399);
  assign nor_1349_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[7])) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign mux_1382_nl = MUX_s_1_2_2(nor_1348_nl, nor_1349_nl, fsm_output[2]);
  assign and_546_nl = (fsm_output[5]) & mux_1382_nl;
  assign or_1173_nl = (COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b0100) | (fsm_output[7])
      | not_tmp_399;
  assign or_1171_nl = (COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b0100) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1381_nl = MUX_s_1_2_2(or_1173_nl, or_1171_nl, fsm_output[2]);
  assign nor_1350_nl = ~((fsm_output[5]) | mux_1381_nl);
  assign mux_1383_nl = MUX_s_1_2_2(and_546_nl, nor_1350_nl, fsm_output[6]);
  assign or_1169_nl = (COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b0100) | (fsm_output[7])
      | not_tmp_399;
  assign or_1167_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0100) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1379_nl = MUX_s_1_2_2(or_1169_nl, or_1167_nl, fsm_output[2]);
  assign nor_1351_nl = ~((fsm_output[5]) | mux_1379_nl);
  assign and_547_nl = nor_346_cse & mux_1378_cse;
  assign mux_1380_nl = MUX_s_1_2_2(nor_1351_nl, and_547_nl, fsm_output[6]);
  assign mux_1384_nl = MUX_s_1_2_2(mux_1383_nl, mux_1380_nl, fsm_output[1]);
  assign or_1163_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0100) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7]) | not_tmp_399;
  assign or_1161_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0100) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1375_nl = MUX_s_1_2_2(or_1163_nl, or_1161_nl, fsm_output[2]);
  assign or_1160_nl = (COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b0100) | (fsm_output[7])
      | not_tmp_399;
  assign or_1158_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0100) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1374_nl = MUX_s_1_2_2(or_1160_nl, or_1158_nl, fsm_output[2]);
  assign mux_1376_nl = MUX_s_1_2_2(mux_1375_nl, mux_1374_nl, fsm_output[5]);
  assign nor_1354_nl = ~((fsm_output[6]) | mux_1376_nl);
  assign nor_1355_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_1356_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7]) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_1372_nl = MUX_s_1_2_2(nor_1355_nl, nor_1356_nl, fsm_output[2]);
  assign nor_1357_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b0100) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_1358_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0100) | (fsm_output[7])
      | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_1371_nl = MUX_s_1_2_2(nor_1357_nl, nor_1358_nl, fsm_output[2]);
  assign mux_1373_nl = MUX_s_1_2_2(mux_1372_nl, mux_1371_nl, fsm_output[5]);
  assign and_548_nl = (fsm_output[6]) & mux_1373_nl;
  assign mux_1377_nl = MUX_s_1_2_2(nor_1354_nl, and_548_nl, fsm_output[1]);
  assign mux_1385_nl = MUX_s_1_2_2(mux_1384_nl, mux_1377_nl, fsm_output[0]);
  assign vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1400_nl,
      mux_1385_nl, fsm_output[3]);
  assign nor_1302_nl = ~((~ (fsm_output[5])) | (VEC_LOOP_j_10_0_sva_9_0[3]) | (fsm_output[0])
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (fsm_output[1]) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | (fsm_output[3:2]!=2'b00) | (~ (VEC_LOOP_j_10_0_sva_9_0[2])) | (fsm_output[8:6]!=3'b000));
  assign nor_1303_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1]) | mux_1366_cse);
  assign nor_1304_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010) | nand_324_cse);
  assign nor_1305_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b010) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1425_nl = MUX_s_1_2_2(nor_1304_nl, nor_1305_nl, fsm_output[2]);
  assign nor_1306_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010) | (fsm_output[8:6]!=3'b011));
  assign nor_1307_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010) | (fsm_output[8:6]!=3'b001));
  assign mux_1424_nl = MUX_s_1_2_2(nor_1306_nl, nor_1307_nl, fsm_output[2]);
  assign mux_1426_nl = MUX_s_1_2_2(mux_1425_nl, mux_1424_nl, fsm_output[3]);
  assign mux_1429_nl = MUX_s_1_2_2(nor_1303_nl, mux_1426_nl, fsm_output[1]);
  assign and_545_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1429_nl;
  assign nor_1308_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]!=4'b0101) | nand_324_cse);
  assign nor_1309_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b0101) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1421_nl = MUX_s_1_2_2(nor_1308_nl, nor_1309_nl, fsm_output[2]);
  assign nor_1310_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b011));
  assign nor_1311_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b001));
  assign mux_1420_nl = MUX_s_1_2_2(nor_1310_nl, nor_1311_nl, fsm_output[2]);
  assign mux_1422_nl = MUX_s_1_2_2(mux_1421_nl, mux_1420_nl, fsm_output[3]);
  assign nor_1312_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b110));
  assign nor_1313_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b100));
  assign mux_1418_nl = MUX_s_1_2_2(nor_1312_nl, nor_1313_nl, fsm_output[2]);
  assign nor_1314_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b010));
  assign nor_1315_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b000));
  assign mux_1417_nl = MUX_s_1_2_2(nor_1314_nl, nor_1315_nl, fsm_output[2]);
  assign mux_1419_nl = MUX_s_1_2_2(mux_1418_nl, mux_1417_nl, fsm_output[3]);
  assign mux_1423_nl = MUX_s_1_2_2(mux_1422_nl, mux_1419_nl, fsm_output[1]);
  assign mux_1430_nl = MUX_s_1_2_2(and_545_nl, mux_1423_nl, fsm_output[0]);
  assign nor_1316_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:0]!=4'b0101) | nand_324_cse);
  assign mux_1413_nl = MUX_s_1_2_2(nor_1316_nl, nor_1317_cse, fsm_output[2]);
  assign nor_1319_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b001));
  assign mux_1412_nl = MUX_s_1_2_2(nor_1286_cse, nor_1319_nl, fsm_output[2]);
  assign mux_1414_nl = MUX_s_1_2_2(mux_1413_nl, mux_1412_nl, fsm_output[3]);
  assign nor_1320_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b110));
  assign mux_1410_nl = MUX_s_1_2_2(nor_1320_nl, nor_1289_cse, fsm_output[2]);
  assign nor_1323_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b000));
  assign mux_1409_nl = MUX_s_1_2_2(nor_1290_cse, nor_1323_nl, fsm_output[2]);
  assign mux_1411_nl = MUX_s_1_2_2(mux_1410_nl, mux_1409_nl, fsm_output[3]);
  assign mux_1415_nl = MUX_s_1_2_2(mux_1414_nl, mux_1411_nl, fsm_output[1]);
  assign nor_1324_nl = ~((COMP_LOOP_acc_1_cse_sva[3:1]!=3'b010) | nand_272_cse);
  assign nor_1325_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0101) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1406_nl = MUX_s_1_2_2(nor_1324_nl, nor_1325_nl, fsm_output[2]);
  assign nor_1326_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b011));
  assign nor_1327_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b001));
  assign mux_1405_nl = MUX_s_1_2_2(nor_1326_nl, nor_1327_nl, fsm_output[2]);
  assign mux_1407_nl = MUX_s_1_2_2(mux_1406_nl, mux_1405_nl, fsm_output[3]);
  assign nor_1328_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b110));
  assign nor_1329_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b100));
  assign mux_1403_nl = MUX_s_1_2_2(nor_1328_nl, nor_1329_nl, fsm_output[2]);
  assign nor_1330_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b010));
  assign nor_1331_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b000));
  assign mux_1402_nl = MUX_s_1_2_2(nor_1330_nl, nor_1331_nl, fsm_output[2]);
  assign mux_1404_nl = MUX_s_1_2_2(mux_1403_nl, mux_1402_nl, fsm_output[3]);
  assign mux_1408_nl = MUX_s_1_2_2(mux_1407_nl, mux_1404_nl, fsm_output[1]);
  assign mux_1416_nl = MUX_s_1_2_2(mux_1415_nl, mux_1408_nl, fsm_output[0]);
  assign mux_1431_nl = MUX_s_1_2_2(mux_1430_nl, mux_1416_nl, fsm_output[5]);
  assign vec_rsc_0_5_i_we_d_pff = MUX_s_1_2_2(nor_1302_nl, mux_1431_nl, fsm_output[4]);
  assign nor_1269_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010)
      | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) | (fsm_output[2]) | (fsm_output[7])
      | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_1270_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b0101) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_1460_nl = MUX_s_1_2_2(nor_1269_nl, nor_1270_nl, fsm_output[5]);
  assign nor_1271_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b0101) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign nor_1272_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b0101) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1459_nl = MUX_s_1_2_2(nor_1271_nl, nor_1272_nl, fsm_output[5]);
  assign mux_1461_nl = MUX_s_1_2_2(mux_1460_nl, mux_1459_nl, fsm_output[1]);
  assign nor_1273_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b0101) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_1274_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0101)
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1457_nl = MUX_s_1_2_2(nor_1273_nl, nor_1274_nl, fsm_output[5]);
  assign nor_1275_nl = ~((VEC_LOOP_j_10_0_sva_9_0[3]) | (fsm_output[5]) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1458_nl = MUX_s_1_2_2(mux_1457_nl, nor_1275_nl, fsm_output[1]);
  assign mux_1462_nl = MUX_s_1_2_2(mux_1461_nl, mux_1458_nl, fsm_output[0]);
  assign nor_1276_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:0]!=4'b0101) | nand_271_cse);
  assign nor_1277_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[2])) |
      (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010) | (~ COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b110));
  assign mux_1454_nl = MUX_s_1_2_2(nor_1276_nl, nor_1277_nl, fsm_output[5]);
  assign nor_1278_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b0101) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign nor_1279_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (~ (fsm_output[2]))
      | (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (~ COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1453_nl = MUX_s_1_2_2(nor_1278_nl, nor_1279_nl, fsm_output[5]);
  assign mux_1455_nl = MUX_s_1_2_2(mux_1454_nl, mux_1453_nl, fsm_output[1]);
  assign nor_1280_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0101) | (~ COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm)
      | (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign nor_1281_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]!=4'b0101) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign mux_1451_nl = MUX_s_1_2_2(nor_1280_nl, nor_1281_nl, fsm_output[5]);
  assign nor_1282_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) | (COMP_LOOP_acc_1_cse_sva[3:1]!=3'b010)
      | nand_272_cse);
  assign nor_1283_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm)
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1449_nl = MUX_s_1_2_2(nor_1282_nl, nor_1283_nl, fsm_output[2]);
  assign nor_1284_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b0101) | (~ (fsm_output[2]))
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1450_nl = MUX_s_1_2_2(mux_1449_nl, nor_1284_nl, fsm_output[5]);
  assign mux_1452_nl = MUX_s_1_2_2(mux_1451_nl, mux_1450_nl, fsm_output[1]);
  assign mux_1456_nl = MUX_s_1_2_2(mux_1455_nl, mux_1452_nl, fsm_output[0]);
  assign mux_1463_nl = MUX_s_1_2_2(mux_1462_nl, mux_1456_nl, fsm_output[4]);
  assign mux_1445_nl = MUX_s_1_2_2(nor_1317_cse, nor_1286_cse, fsm_output[2]);
  assign nor_1287_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b010) | (~ COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b100));
  assign nor_1288_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b010));
  assign mux_1444_nl = MUX_s_1_2_2(nor_1287_nl, nor_1288_nl, fsm_output[2]);
  assign and_543_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1444_nl;
  assign mux_1446_nl = MUX_s_1_2_2(mux_1445_nl, and_543_nl, fsm_output[5]);
  assign mux_1442_nl = MUX_s_1_2_2(nor_1289_cse, nor_1290_cse, fsm_output[2]);
  assign and_544_nl = nor_351_cse & mux_1441_cse;
  assign mux_1443_nl = MUX_s_1_2_2(mux_1442_nl, and_544_nl, fsm_output[5]);
  assign mux_1447_nl = MUX_s_1_2_2(mux_1446_nl, mux_1443_nl, fsm_output[1]);
  assign nor_1294_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0101) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b100));
  assign nor_1295_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0101) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b010));
  assign mux_1437_nl = MUX_s_1_2_2(nor_1294_nl, nor_1295_nl, fsm_output[2]);
  assign nor_1296_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b100));
  assign nor_1297_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b010));
  assign mux_1436_nl = MUX_s_1_2_2(nor_1296_nl, nor_1297_nl, fsm_output[2]);
  assign mux_1438_nl = MUX_s_1_2_2(mux_1437_nl, mux_1436_nl, fsm_output[5]);
  assign nor_1298_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | (fsm_output[8:6]!=3'b011));
  assign nor_1299_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[8:6]!=3'b001));
  assign mux_1434_nl = MUX_s_1_2_2(nor_1298_nl, nor_1299_nl, fsm_output[2]);
  assign nor_1300_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b011));
  assign nor_1301_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0101) | (fsm_output[8:6]!=3'b001));
  assign mux_1433_nl = MUX_s_1_2_2(nor_1300_nl, nor_1301_nl, fsm_output[2]);
  assign mux_1435_nl = MUX_s_1_2_2(mux_1434_nl, mux_1433_nl, fsm_output[5]);
  assign mux_1439_nl = MUX_s_1_2_2(mux_1438_nl, mux_1435_nl, fsm_output[1]);
  assign mux_1448_nl = MUX_s_1_2_2(mux_1447_nl, mux_1439_nl, fsm_output[0]);
  assign and_542_nl = (fsm_output[4]) & mux_1448_nl;
  assign vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1463_nl,
      and_542_nl, fsm_output[3]);
  assign nor_1240_nl = ~((~ (fsm_output[5])) | (VEC_LOOP_j_10_0_sva_9_0[3]) | (fsm_output[0])
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[1]) | (~ (VEC_LOOP_j_10_0_sva_9_0[1]))
      | (fsm_output[3:2]!=2'b00) | (~ (VEC_LOOP_j_10_0_sva_9_0[2])) | (fsm_output[8:6]!=3'b000));
  assign nand_47_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1]) & mux_1491_cse);
  assign or_1340_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b011) | nand_324_cse;
  assign or_1338_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b011) | (fsm_output[7]) |
      not_tmp_395;
  assign mux_1488_nl = MUX_s_1_2_2(or_1340_nl, or_1338_nl, fsm_output[2]);
  assign or_1336_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b011) | (fsm_output[8:6]!=3'b011);
  assign or_1335_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b011) | (fsm_output[8:6]!=3'b001);
  assign mux_1487_nl = MUX_s_1_2_2(or_1336_nl, or_1335_nl, fsm_output[2]);
  assign mux_1489_nl = MUX_s_1_2_2(mux_1488_nl, mux_1487_nl, fsm_output[3]);
  assign mux_1492_nl = MUX_s_1_2_2(nand_47_nl, mux_1489_nl, fsm_output[1]);
  assign nor_1241_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1492_nl);
  assign nor_1245_nl = ~((~ (COMP_LOOP_acc_10_cse_10_1_15_sva[2])) | (COMP_LOOP_acc_10_cse_10_1_15_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_15_sva[0]) | nand_268_cse);
  assign nor_1246_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b0110) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1484_nl = MUX_s_1_2_2(nor_1245_nl, nor_1246_nl, fsm_output[2]);
  assign nor_1247_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b011));
  assign nor_1248_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b001));
  assign mux_1483_nl = MUX_s_1_2_2(nor_1247_nl, nor_1248_nl, fsm_output[2]);
  assign mux_1485_nl = MUX_s_1_2_2(mux_1484_nl, mux_1483_nl, fsm_output[3]);
  assign nor_1249_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b110));
  assign nor_1250_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b100));
  assign mux_1481_nl = MUX_s_1_2_2(nor_1249_nl, nor_1250_nl, fsm_output[2]);
  assign nor_1251_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b010));
  assign nor_1252_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b000));
  assign mux_1480_nl = MUX_s_1_2_2(nor_1251_nl, nor_1252_nl, fsm_output[2]);
  assign mux_1482_nl = MUX_s_1_2_2(mux_1481_nl, mux_1480_nl, fsm_output[3]);
  assign mux_1486_nl = MUX_s_1_2_2(mux_1485_nl, mux_1482_nl, fsm_output[1]);
  assign mux_1493_nl = MUX_s_1_2_2(nor_1241_nl, mux_1486_nl, fsm_output[0]);
  assign nor_1253_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:0]!=4'b0110) | nand_324_cse);
  assign nor_1254_nl = ~((COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b0110) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1476_nl = MUX_s_1_2_2(nor_1253_nl, nor_1254_nl, fsm_output[2]);
  assign nor_1255_nl = ~((COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b011));
  assign nor_1256_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b001));
  assign mux_1475_nl = MUX_s_1_2_2(nor_1255_nl, nor_1256_nl, fsm_output[2]);
  assign mux_1477_nl = MUX_s_1_2_2(mux_1476_nl, mux_1475_nl, fsm_output[3]);
  assign nor_1257_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b110));
  assign nor_1258_nl = ~((COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b100));
  assign mux_1473_nl = MUX_s_1_2_2(nor_1257_nl, nor_1258_nl, fsm_output[2]);
  assign nor_1259_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b010));
  assign nor_1260_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b000));
  assign mux_1472_nl = MUX_s_1_2_2(nor_1259_nl, nor_1260_nl, fsm_output[2]);
  assign mux_1474_nl = MUX_s_1_2_2(mux_1473_nl, mux_1472_nl, fsm_output[3]);
  assign mux_1478_nl = MUX_s_1_2_2(mux_1477_nl, mux_1474_nl, fsm_output[1]);
  assign nor_1261_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0110) | nand_324_cse);
  assign nor_1262_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0110) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1469_nl = MUX_s_1_2_2(nor_1261_nl, nor_1262_nl, fsm_output[2]);
  assign nor_1263_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b011));
  assign nor_1264_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b001));
  assign mux_1468_nl = MUX_s_1_2_2(nor_1263_nl, nor_1264_nl, fsm_output[2]);
  assign mux_1470_nl = MUX_s_1_2_2(mux_1469_nl, mux_1468_nl, fsm_output[3]);
  assign nor_1265_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b110));
  assign nor_1266_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b100));
  assign mux_1466_nl = MUX_s_1_2_2(nor_1265_nl, nor_1266_nl, fsm_output[2]);
  assign nor_1267_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b010));
  assign nor_1268_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0110) | (fsm_output[8:6]!=3'b000));
  assign mux_1465_nl = MUX_s_1_2_2(nor_1267_nl, nor_1268_nl, fsm_output[2]);
  assign mux_1467_nl = MUX_s_1_2_2(mux_1466_nl, mux_1465_nl, fsm_output[3]);
  assign mux_1471_nl = MUX_s_1_2_2(mux_1470_nl, mux_1467_nl, fsm_output[1]);
  assign mux_1479_nl = MUX_s_1_2_2(mux_1478_nl, mux_1471_nl, fsm_output[0]);
  assign mux_1494_nl = MUX_s_1_2_2(mux_1493_nl, mux_1479_nl, fsm_output[5]);
  assign vec_rsc_0_6_i_we_d_pff = MUX_s_1_2_2(nor_1240_nl, mux_1494_nl, fsm_output[4]);
  assign nor_1213_nl = ~((~((fsm_output[5]) & (fsm_output[2]) & (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      & (COMP_LOOP_acc_20_psp_sva[2:0]==3'b011) & COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm))
      | nand_301_cse);
  assign nor_1214_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b011) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1215_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:0]!=4'b0110) | nand_301_cse);
  assign mux_1521_nl = MUX_s_1_2_2(nor_1214_nl, nor_1215_nl, fsm_output[2]);
  assign nor_1216_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b0110) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1522_nl = MUX_s_1_2_2(mux_1521_nl, nor_1216_nl, fsm_output[5]);
  assign mux_1523_nl = MUX_s_1_2_2(nor_1213_nl, mux_1522_nl, fsm_output[6]);
  assign nor_1217_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b0110) | (fsm_output[7])
      | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1218_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b0110) | nand_301_cse);
  assign mux_1518_nl = MUX_s_1_2_2(nor_1217_nl, nor_1218_nl, fsm_output[2]);
  assign nor_1219_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b0110) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1519_nl = MUX_s_1_2_2(mux_1518_nl, nor_1219_nl, fsm_output[5]);
  assign nor_1220_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[1])) | (~ (fsm_output[5])) |
      (~ (fsm_output[2])) | (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (~ COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | not_tmp_399);
  assign mux_1520_nl = MUX_s_1_2_2(mux_1519_nl, nor_1220_nl, fsm_output[6]);
  assign mux_1524_nl = MUX_s_1_2_2(mux_1523_nl, mux_1520_nl, fsm_output[1]);
  assign nor_1221_nl = ~((~ (fsm_output[2])) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0110)
      | (~ COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm) | nand_301_cse);
  assign nor_1222_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0110)
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1223_nl = ~((~ (COMP_LOOP_acc_10_cse_10_1_15_sva[2])) | (COMP_LOOP_acc_10_cse_10_1_15_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_15_sva[0]) | nand_265_cse);
  assign mux_1514_nl = MUX_s_1_2_2(nor_1222_nl, nor_1223_nl, fsm_output[2]);
  assign mux_1515_nl = MUX_s_1_2_2(nor_1221_nl, mux_1514_nl, fsm_output[5]);
  assign nor_1224_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b0110) | (fsm_output[5])
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1516_nl = MUX_s_1_2_2(mux_1515_nl, nor_1224_nl, fsm_output[6]);
  assign nor_1225_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[1])) | (VEC_LOOP_j_10_0_sva_9_0[3])
      | (fsm_output[5]) | (fsm_output[2]) | (~ (VEC_LOOP_j_10_0_sva_9_0[2])) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1226_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) | (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0110)
      | nand_301_cse);
  assign nor_1227_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm)
      | (fsm_output[7]) | not_tmp_399);
  assign mux_1511_nl = MUX_s_1_2_2(nor_1226_nl, nor_1227_nl, fsm_output[2]);
  assign nor_1228_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b0110) | (~ (fsm_output[2]))
      | (fsm_output[7]) | not_tmp_399);
  assign mux_1512_nl = MUX_s_1_2_2(mux_1511_nl, nor_1228_nl, fsm_output[5]);
  assign mux_1513_nl = MUX_s_1_2_2(nor_1225_nl, mux_1512_nl, fsm_output[6]);
  assign mux_1517_nl = MUX_s_1_2_2(mux_1516_nl, mux_1513_nl, fsm_output[1]);
  assign mux_1525_nl = MUX_s_1_2_2(mux_1524_nl, mux_1517_nl, fsm_output[0]);
  assign nor_1229_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b011) | (~ COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | not_tmp_399);
  assign nor_1230_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b011) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[7])) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign mux_1507_nl = MUX_s_1_2_2(nor_1229_nl, nor_1230_nl, fsm_output[2]);
  assign and_539_nl = (fsm_output[5]) & mux_1507_nl;
  assign or_1367_nl = (COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b0110) | (fsm_output[7])
      | not_tmp_399;
  assign or_1365_nl = (COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b0110) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1506_nl = MUX_s_1_2_2(or_1367_nl, or_1365_nl, fsm_output[2]);
  assign nor_1231_nl = ~((fsm_output[5]) | mux_1506_nl);
  assign mux_1508_nl = MUX_s_1_2_2(and_539_nl, nor_1231_nl, fsm_output[6]);
  assign or_1363_nl = (COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b0110) | (fsm_output[7])
      | not_tmp_399;
  assign or_1361_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0110) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1504_nl = MUX_s_1_2_2(or_1363_nl, or_1361_nl, fsm_output[2]);
  assign nor_1232_nl = ~((fsm_output[5]) | mux_1504_nl);
  assign and_540_nl = (VEC_LOOP_j_10_0_sva_9_0[1]) & (fsm_output[5]) & mux_1378_cse;
  assign mux_1505_nl = MUX_s_1_2_2(nor_1232_nl, and_540_nl, fsm_output[6]);
  assign mux_1509_nl = MUX_s_1_2_2(mux_1508_nl, mux_1505_nl, fsm_output[1]);
  assign or_1357_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0110) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7]) | not_tmp_399;
  assign or_1355_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0110) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1500_nl = MUX_s_1_2_2(or_1357_nl, or_1355_nl, fsm_output[2]);
  assign or_1354_nl = (COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b0110) | (fsm_output[7])
      | not_tmp_399;
  assign or_1352_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0110) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1499_nl = MUX_s_1_2_2(or_1354_nl, or_1352_nl, fsm_output[2]);
  assign mux_1501_nl = MUX_s_1_2_2(mux_1500_nl, mux_1499_nl, fsm_output[5]);
  assign nor_1235_nl = ~((fsm_output[6]) | mux_1501_nl);
  assign nor_1236_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_1237_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7]) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_1497_nl = MUX_s_1_2_2(nor_1236_nl, nor_1237_nl, fsm_output[2]);
  assign nor_1238_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b0110) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_1239_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0110) | (fsm_output[7])
      | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_1496_nl = MUX_s_1_2_2(nor_1238_nl, nor_1239_nl, fsm_output[2]);
  assign mux_1498_nl = MUX_s_1_2_2(mux_1497_nl, mux_1496_nl, fsm_output[5]);
  assign and_541_nl = (fsm_output[6]) & mux_1498_nl;
  assign mux_1502_nl = MUX_s_1_2_2(nor_1235_nl, and_541_nl, fsm_output[1]);
  assign mux_1510_nl = MUX_s_1_2_2(mux_1509_nl, mux_1502_nl, fsm_output[0]);
  assign vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1525_nl,
      mux_1510_nl, fsm_output[3]);
  assign nor_1184_nl = ~((~ (fsm_output[5])) | (VEC_LOOP_j_10_0_sva_9_0[3]) | (fsm_output[0])
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (fsm_output[1]) | (~ (VEC_LOOP_j_10_0_sva_9_0[1]))
      | (fsm_output[3:2]!=2'b00) | (~ (VEC_LOOP_j_10_0_sva_9_0[2])) | (fsm_output[8:6]!=3'b000));
  assign and_535_nl = (VEC_LOOP_j_10_0_sva_9_0[1]) & mux_1491_cse;
  assign nor_1188_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b011) | nand_324_cse);
  assign nor_1189_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b011) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1550_nl = MUX_s_1_2_2(nor_1188_nl, nor_1189_nl, fsm_output[2]);
  assign nor_1190_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b011) | (fsm_output[8:6]!=3'b011));
  assign nor_1191_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b011) | (fsm_output[8:6]!=3'b001));
  assign mux_1549_nl = MUX_s_1_2_2(nor_1190_nl, nor_1191_nl, fsm_output[2]);
  assign mux_1551_nl = MUX_s_1_2_2(mux_1550_nl, mux_1549_nl, fsm_output[3]);
  assign mux_1554_nl = MUX_s_1_2_2(and_535_nl, mux_1551_nl, fsm_output[1]);
  assign and_534_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1554_nl;
  assign nor_1192_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:2]!=2'b01) | nand_261_cse);
  assign nor_1193_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b0111) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1546_nl = MUX_s_1_2_2(nor_1192_nl, nor_1193_nl, fsm_output[2]);
  assign and_536_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]==4'b0111) & (fsm_output[8:6]==3'b011);
  assign nor_1194_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b0111) | (fsm_output[8:6]!=3'b001));
  assign mux_1545_nl = MUX_s_1_2_2(and_536_nl, nor_1194_nl, fsm_output[2]);
  assign mux_1547_nl = MUX_s_1_2_2(mux_1546_nl, mux_1545_nl, fsm_output[3]);
  assign and_842_nl = (COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]==4'b0111) & (fsm_output[8:6]==3'b110);
  assign nor_1196_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b0111) | (fsm_output[8:6]!=3'b100));
  assign mux_1543_nl = MUX_s_1_2_2(and_842_nl, nor_1196_nl, fsm_output[2]);
  assign nor_1197_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0111) | (fsm_output[8:6]!=3'b010));
  assign nor_1198_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[3:0]!=4'b0111) | (fsm_output[8:6]!=3'b000));
  assign mux_1542_nl = MUX_s_1_2_2(nor_1197_nl, nor_1198_nl, fsm_output[2]);
  assign mux_1544_nl = MUX_s_1_2_2(mux_1543_nl, mux_1542_nl, fsm_output[3]);
  assign mux_1548_nl = MUX_s_1_2_2(mux_1547_nl, mux_1544_nl, fsm_output[1]);
  assign mux_1555_nl = MUX_s_1_2_2(and_534_nl, mux_1548_nl, fsm_output[0]);
  assign nor_1199_nl = ~(nand_226_cse | nand_324_cse);
  assign mux_1538_nl = MUX_s_1_2_2(nor_1199_nl, nor_1200_cse, fsm_output[2]);
  assign nor_1201_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b0111) | (fsm_output[8:6]!=3'b001));
  assign mux_1537_nl = MUX_s_1_2_2(and_529_cse, nor_1201_nl, fsm_output[2]);
  assign mux_1539_nl = MUX_s_1_2_2(mux_1538_nl, mux_1537_nl, fsm_output[3]);
  assign and_853_nl = (COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]==4'b0111) & (fsm_output[8:6]==3'b110);
  assign mux_1535_nl = MUX_s_1_2_2(and_853_nl, nor_1173_cse, fsm_output[2]);
  assign nor_1205_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b0111) | (fsm_output[8:6]!=3'b000));
  assign mux_1534_nl = MUX_s_1_2_2(nor_1174_cse, nor_1205_nl, fsm_output[2]);
  assign mux_1536_nl = MUX_s_1_2_2(mux_1535_nl, mux_1534_nl, fsm_output[3]);
  assign mux_1540_nl = MUX_s_1_2_2(mux_1539_nl, mux_1536_nl, fsm_output[1]);
  assign nor_1206_nl = ~((COMP_LOOP_acc_1_cse_sva[3:1]!=3'b011) | nand_272_cse);
  assign nor_1207_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0111) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1531_nl = MUX_s_1_2_2(nor_1206_nl, nor_1207_nl, fsm_output[2]);
  assign and_538_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b0111) & (fsm_output[8:6]==3'b011);
  assign nor_1208_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0111) | (fsm_output[8:6]!=3'b001));
  assign mux_1530_nl = MUX_s_1_2_2(and_538_nl, nor_1208_nl, fsm_output[2]);
  assign mux_1532_nl = MUX_s_1_2_2(mux_1531_nl, mux_1530_nl, fsm_output[3]);
  assign and_872_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b0111) & (fsm_output[8:6]==3'b110);
  assign nor_1210_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0111) | (fsm_output[8:6]!=3'b100));
  assign mux_1528_nl = MUX_s_1_2_2(and_872_nl, nor_1210_nl, fsm_output[2]);
  assign nor_1211_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0111) | (fsm_output[8:6]!=3'b010));
  assign nor_1212_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0111) | (fsm_output[8:6]!=3'b000));
  assign mux_1527_nl = MUX_s_1_2_2(nor_1211_nl, nor_1212_nl, fsm_output[2]);
  assign mux_1529_nl = MUX_s_1_2_2(mux_1528_nl, mux_1527_nl, fsm_output[3]);
  assign mux_1533_nl = MUX_s_1_2_2(mux_1532_nl, mux_1529_nl, fsm_output[1]);
  assign mux_1541_nl = MUX_s_1_2_2(mux_1540_nl, mux_1533_nl, fsm_output[0]);
  assign mux_1556_nl = MUX_s_1_2_2(mux_1555_nl, mux_1541_nl, fsm_output[5]);
  assign vec_rsc_0_7_i_we_d_pff = MUX_s_1_2_2(nor_1184_nl, mux_1556_nl, fsm_output[4]);
  assign nor_1154_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b011)
      | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) | (fsm_output[2]) | (fsm_output[7])
      | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_1155_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b0111) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_1585_nl = MUX_s_1_2_2(nor_1154_nl, nor_1155_nl, fsm_output[5]);
  assign nor_1156_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b0111) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign nor_1157_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b0111) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1584_nl = MUX_s_1_2_2(nor_1156_nl, nor_1157_nl, fsm_output[5]);
  assign mux_1586_nl = MUX_s_1_2_2(mux_1585_nl, mux_1584_nl, fsm_output[1]);
  assign nor_1158_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b0111) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_1159_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0111)
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1582_nl = MUX_s_1_2_2(nor_1158_nl, nor_1159_nl, fsm_output[5]);
  assign nor_1160_nl = ~((VEC_LOOP_j_10_0_sva_9_0[3]) | (fsm_output[5]) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1583_nl = MUX_s_1_2_2(mux_1582_nl, nor_1160_nl, fsm_output[1]);
  assign mux_1587_nl = MUX_s_1_2_2(mux_1586_nl, mux_1583_nl, fsm_output[0]);
  assign nor_1161_nl = ~(nand_226_cse | nand_271_cse);
  assign and_852_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (fsm_output[2]) & (COMP_LOOP_acc_20_psp_sva[2:0]==3'b011)
      & COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm & (fsm_output[8:6]==3'b110);
  assign mux_1579_nl = MUX_s_1_2_2(nor_1161_nl, and_852_nl, fsm_output[5]);
  assign and_858_nl = (COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]==4'b0111) & (fsm_output[2])
      & (fsm_output[7]) & (~ (fsm_output[6])) & (fsm_output[8]);
  assign nor_1164_nl = ~((~((VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & (fsm_output[2])
      & (COMP_LOOP_acc_19_psp_sva[1:0]==2'b01) & COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm
      & (~ (fsm_output[7])))) | not_tmp_395);
  assign mux_1578_nl = MUX_s_1_2_2(and_858_nl, nor_1164_nl, fsm_output[5]);
  assign mux_1580_nl = MUX_s_1_2_2(mux_1579_nl, mux_1578_nl, fsm_output[1]);
  assign and_870_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b0111) & COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[2]) & (fsm_output[7]) & (~ (fsm_output[6])) & (fsm_output[8]);
  assign and_871_nl = (COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]==4'b0111) & (fsm_output[2])
      & (fsm_output[7]) & (~ (fsm_output[6])) & (fsm_output[8]);
  assign mux_1576_nl = MUX_s_1_2_2(and_870_nl, and_871_nl, fsm_output[5]);
  assign nor_1167_nl = ~((~(COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm & (COMP_LOOP_acc_1_cse_sva[3:1]==3'b011)))
      | nand_272_cse);
  assign nor_1168_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0111) | (~ COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm)
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1574_nl = MUX_s_1_2_2(nor_1167_nl, nor_1168_nl, fsm_output[2]);
  assign nor_1169_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b0111) | (~ (fsm_output[2]))
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1575_nl = MUX_s_1_2_2(mux_1574_nl, nor_1169_nl, fsm_output[5]);
  assign mux_1577_nl = MUX_s_1_2_2(mux_1576_nl, mux_1575_nl, fsm_output[1]);
  assign mux_1581_nl = MUX_s_1_2_2(mux_1580_nl, mux_1577_nl, fsm_output[0]);
  assign mux_1588_nl = MUX_s_1_2_2(mux_1587_nl, mux_1581_nl, fsm_output[4]);
  assign mux_1570_nl = MUX_s_1_2_2(nor_1200_cse, and_529_cse, fsm_output[2]);
  assign nor_1171_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b011) | (~ COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b100));
  assign nor_1172_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b011) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b010));
  assign mux_1569_nl = MUX_s_1_2_2(nor_1171_nl, nor_1172_nl, fsm_output[2]);
  assign and_530_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1569_nl;
  assign mux_1571_nl = MUX_s_1_2_2(mux_1570_nl, and_530_nl, fsm_output[5]);
  assign mux_1567_nl = MUX_s_1_2_2(nor_1173_cse, nor_1174_cse, fsm_output[2]);
  assign and_531_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & mux_1441_cse;
  assign mux_1568_nl = MUX_s_1_2_2(mux_1567_nl, and_531_nl, fsm_output[5]);
  assign mux_1572_nl = MUX_s_1_2_2(mux_1571_nl, mux_1568_nl, fsm_output[1]);
  assign nor_1178_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0111) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b100));
  assign nor_1179_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0111) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b010));
  assign mux_1562_nl = MUX_s_1_2_2(nor_1178_nl, nor_1179_nl, fsm_output[2]);
  assign nor_1180_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b0111) | (fsm_output[8:6]!=3'b100));
  assign nor_1181_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0111) | (fsm_output[8:6]!=3'b010));
  assign mux_1561_nl = MUX_s_1_2_2(nor_1180_nl, nor_1181_nl, fsm_output[2]);
  assign mux_1563_nl = MUX_s_1_2_2(mux_1562_nl, mux_1561_nl, fsm_output[5]);
  assign and_532_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b0111) & COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm
      & (fsm_output[8:6]==3'b011);
  assign nor_1182_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0111) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[8:6]!=3'b001));
  assign mux_1559_nl = MUX_s_1_2_2(and_532_nl, nor_1182_nl, fsm_output[2]);
  assign and_533_nl = (COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]==4'b0111) & (fsm_output[8:6]==3'b011);
  assign nor_1183_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0111) | (fsm_output[8:6]!=3'b001));
  assign mux_1558_nl = MUX_s_1_2_2(and_533_nl, nor_1183_nl, fsm_output[2]);
  assign mux_1560_nl = MUX_s_1_2_2(mux_1559_nl, mux_1558_nl, fsm_output[5]);
  assign mux_1564_nl = MUX_s_1_2_2(mux_1563_nl, mux_1560_nl, fsm_output[1]);
  assign mux_1573_nl = MUX_s_1_2_2(mux_1572_nl, mux_1564_nl, fsm_output[0]);
  assign and_528_nl = (fsm_output[4]) & mux_1573_nl;
  assign vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1588_nl,
      and_528_nl, fsm_output[3]);
  assign nor_1128_nl = ~((~ (fsm_output[5])) | (~ (VEC_LOOP_j_10_0_sva_9_0[3])) |
      (fsm_output[0]) | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[1]) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | (fsm_output[3:2]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2]) | (fsm_output[8:6]!=3'b000));
  assign or_1539_nl = (VEC_LOOP_j_10_0_sva_9_0[1]) | mux_1616_cse;
  assign or_1533_nl = (COMP_LOOP_acc_20_psp_sva[1:0]!=2'b00) | nand_222_cse;
  assign or_1531_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b100) | (fsm_output[7]) |
      not_tmp_395;
  assign mux_1613_nl = MUX_s_1_2_2(or_1533_nl, or_1531_nl, fsm_output[2]);
  assign or_1529_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100) | (fsm_output[8:6]!=3'b011);
  assign or_1528_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100) | (fsm_output[8:6]!=3'b001);
  assign mux_1612_nl = MUX_s_1_2_2(or_1529_nl, or_1528_nl, fsm_output[2]);
  assign mux_1614_nl = MUX_s_1_2_2(mux_1613_nl, mux_1612_nl, fsm_output[3]);
  assign mux_1617_nl = MUX_s_1_2_2(or_1539_nl, mux_1614_nl, fsm_output[1]);
  assign nor_1129_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1617_nl);
  assign nor_1130_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]!=4'b1000) | nand_324_cse);
  assign nor_1131_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b1000) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1609_nl = MUX_s_1_2_2(nor_1130_nl, nor_1131_nl, fsm_output[2]);
  assign nor_1132_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b011));
  assign nor_1133_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b001));
  assign mux_1608_nl = MUX_s_1_2_2(nor_1132_nl, nor_1133_nl, fsm_output[2]);
  assign mux_1610_nl = MUX_s_1_2_2(mux_1609_nl, mux_1608_nl, fsm_output[3]);
  assign nor_1134_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b110));
  assign nor_1135_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b100));
  assign mux_1606_nl = MUX_s_1_2_2(nor_1134_nl, nor_1135_nl, fsm_output[2]);
  assign nor_1136_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b010));
  assign nor_1137_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b000));
  assign mux_1605_nl = MUX_s_1_2_2(nor_1136_nl, nor_1137_nl, fsm_output[2]);
  assign mux_1607_nl = MUX_s_1_2_2(mux_1606_nl, mux_1605_nl, fsm_output[3]);
  assign mux_1611_nl = MUX_s_1_2_2(mux_1610_nl, mux_1607_nl, fsm_output[1]);
  assign mux_1618_nl = MUX_s_1_2_2(nor_1129_nl, mux_1611_nl, fsm_output[0]);
  assign nor_1138_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[2:0]!=3'b000) | nand_223_cse);
  assign nor_1139_nl = ~((COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b1000) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1601_nl = MUX_s_1_2_2(nor_1138_nl, nor_1139_nl, fsm_output[2]);
  assign nor_1140_nl = ~((COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b011));
  assign nor_1141_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b001));
  assign mux_1600_nl = MUX_s_1_2_2(nor_1140_nl, nor_1141_nl, fsm_output[2]);
  assign mux_1602_nl = MUX_s_1_2_2(mux_1601_nl, mux_1600_nl, fsm_output[3]);
  assign nor_1142_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b110));
  assign nor_1143_nl = ~((COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b100));
  assign mux_1598_nl = MUX_s_1_2_2(nor_1142_nl, nor_1143_nl, fsm_output[2]);
  assign nor_1144_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b010));
  assign nor_1145_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b000));
  assign mux_1597_nl = MUX_s_1_2_2(nor_1144_nl, nor_1145_nl, fsm_output[2]);
  assign mux_1599_nl = MUX_s_1_2_2(mux_1598_nl, mux_1597_nl, fsm_output[3]);
  assign mux_1603_nl = MUX_s_1_2_2(mux_1602_nl, mux_1599_nl, fsm_output[1]);
  assign nor_1146_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1000) | nand_324_cse);
  assign nor_1147_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1000) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1594_nl = MUX_s_1_2_2(nor_1146_nl, nor_1147_nl, fsm_output[2]);
  assign nor_1148_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b011));
  assign nor_1149_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b001));
  assign mux_1593_nl = MUX_s_1_2_2(nor_1148_nl, nor_1149_nl, fsm_output[2]);
  assign mux_1595_nl = MUX_s_1_2_2(mux_1594_nl, mux_1593_nl, fsm_output[3]);
  assign nor_1150_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b110));
  assign nor_1151_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b100));
  assign mux_1591_nl = MUX_s_1_2_2(nor_1150_nl, nor_1151_nl, fsm_output[2]);
  assign nor_1152_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b010));
  assign nor_1153_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1000) | (fsm_output[8:6]!=3'b000));
  assign mux_1590_nl = MUX_s_1_2_2(nor_1152_nl, nor_1153_nl, fsm_output[2]);
  assign mux_1592_nl = MUX_s_1_2_2(mux_1591_nl, mux_1590_nl, fsm_output[3]);
  assign mux_1596_nl = MUX_s_1_2_2(mux_1595_nl, mux_1592_nl, fsm_output[1]);
  assign mux_1604_nl = MUX_s_1_2_2(mux_1603_nl, mux_1596_nl, fsm_output[0]);
  assign mux_1619_nl = MUX_s_1_2_2(mux_1618_nl, mux_1604_nl, fsm_output[5]);
  assign vec_rsc_0_8_i_we_d_pff = MUX_s_1_2_2(nor_1128_nl, mux_1619_nl, fsm_output[4]);
  assign nor_1101_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[2])) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b100) | (~ COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm)
      | nand_301_cse);
  assign nor_1102_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1103_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[2:0]!=3'b000) | nand_219_cse);
  assign mux_1646_nl = MUX_s_1_2_2(nor_1102_nl, nor_1103_nl, fsm_output[2]);
  assign nor_1104_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b1000) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1647_nl = MUX_s_1_2_2(mux_1646_nl, nor_1104_nl, fsm_output[5]);
  assign mux_1648_nl = MUX_s_1_2_2(nor_1101_nl, mux_1647_nl, fsm_output[6]);
  assign nor_1105_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b1000) | (fsm_output[7])
      | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1106_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b1000) | nand_301_cse);
  assign mux_1643_nl = MUX_s_1_2_2(nor_1105_nl, nor_1106_nl, fsm_output[2]);
  assign nor_1107_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b1000) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1644_nl = MUX_s_1_2_2(mux_1643_nl, nor_1107_nl, fsm_output[5]);
  assign nor_1108_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1]) | (~ (fsm_output[5])) | (~
      (fsm_output[2])) | (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (~ COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | not_tmp_399);
  assign mux_1645_nl = MUX_s_1_2_2(mux_1644_nl, nor_1108_nl, fsm_output[6]);
  assign mux_1649_nl = MUX_s_1_2_2(mux_1648_nl, mux_1645_nl, fsm_output[1]);
  assign nor_1109_nl = ~((~ (fsm_output[2])) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1000)
      | (~ COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm) | nand_301_cse);
  assign nor_1110_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1000)
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1111_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]!=4'b1000) | nand_301_cse);
  assign mux_1639_nl = MUX_s_1_2_2(nor_1110_nl, nor_1111_nl, fsm_output[2]);
  assign mux_1640_nl = MUX_s_1_2_2(nor_1109_nl, mux_1639_nl, fsm_output[5]);
  assign nor_1112_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b1000) | (fsm_output[5])
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1641_nl = MUX_s_1_2_2(mux_1640_nl, nor_1112_nl, fsm_output[6]);
  assign nor_1113_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1]) | (~ (VEC_LOOP_j_10_0_sva_9_0[3]))
      | (fsm_output[5]) | (fsm_output[2]) | (VEC_LOOP_j_10_0_sva_9_0[2]) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_1114_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) | (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1000)
      | nand_301_cse);
  assign nor_1115_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm)
      | (fsm_output[7]) | not_tmp_399);
  assign mux_1636_nl = MUX_s_1_2_2(nor_1114_nl, nor_1115_nl, fsm_output[2]);
  assign nor_1116_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b1000) | (~ (fsm_output[2]))
      | (fsm_output[7]) | not_tmp_399);
  assign mux_1637_nl = MUX_s_1_2_2(mux_1636_nl, nor_1116_nl, fsm_output[5]);
  assign mux_1638_nl = MUX_s_1_2_2(nor_1113_nl, mux_1637_nl, fsm_output[6]);
  assign mux_1642_nl = MUX_s_1_2_2(mux_1641_nl, mux_1638_nl, fsm_output[1]);
  assign mux_1650_nl = MUX_s_1_2_2(mux_1649_nl, mux_1642_nl, fsm_output[0]);
  assign nor_1117_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b100) | (~ COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | not_tmp_399);
  assign nor_1118_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[7])) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign mux_1632_nl = MUX_s_1_2_2(nor_1117_nl, nor_1118_nl, fsm_output[2]);
  assign and_525_nl = (fsm_output[5]) & mux_1632_nl;
  assign or_1561_nl = (COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b1000) | (fsm_output[7])
      | not_tmp_399;
  assign or_1559_nl = (COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b1000) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1631_nl = MUX_s_1_2_2(or_1561_nl, or_1559_nl, fsm_output[2]);
  assign nor_1119_nl = ~((fsm_output[5]) | mux_1631_nl);
  assign mux_1633_nl = MUX_s_1_2_2(and_525_nl, nor_1119_nl, fsm_output[6]);
  assign or_1557_nl = (COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b1000) | (fsm_output[7])
      | not_tmp_399;
  assign or_1555_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b1000) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1629_nl = MUX_s_1_2_2(or_1557_nl, or_1555_nl, fsm_output[2]);
  assign nor_1120_nl = ~((fsm_output[5]) | mux_1629_nl);
  assign and_526_nl = nor_346_cse & mux_1628_cse;
  assign mux_1630_nl = MUX_s_1_2_2(nor_1120_nl, and_526_nl, fsm_output[6]);
  assign mux_1634_nl = MUX_s_1_2_2(mux_1633_nl, mux_1630_nl, fsm_output[1]);
  assign or_1551_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1000) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7]) | not_tmp_399;
  assign or_1549_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1000) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1625_nl = MUX_s_1_2_2(or_1551_nl, or_1549_nl, fsm_output[2]);
  assign or_1548_nl = (COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b1000) | (fsm_output[7])
      | not_tmp_399;
  assign or_1546_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b1000) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1624_nl = MUX_s_1_2_2(or_1548_nl, or_1546_nl, fsm_output[2]);
  assign mux_1626_nl = MUX_s_1_2_2(mux_1625_nl, mux_1624_nl, fsm_output[5]);
  assign nor_1123_nl = ~((fsm_output[6]) | mux_1626_nl);
  assign nor_1124_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_1125_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7]) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_1622_nl = MUX_s_1_2_2(nor_1124_nl, nor_1125_nl, fsm_output[2]);
  assign nor_1126_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b1000) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_1127_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b1000) | (fsm_output[7])
      | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_1621_nl = MUX_s_1_2_2(nor_1126_nl, nor_1127_nl, fsm_output[2]);
  assign mux_1623_nl = MUX_s_1_2_2(mux_1622_nl, mux_1621_nl, fsm_output[5]);
  assign and_527_nl = (fsm_output[6]) & mux_1623_nl;
  assign mux_1627_nl = MUX_s_1_2_2(nor_1123_nl, and_527_nl, fsm_output[1]);
  assign mux_1635_nl = MUX_s_1_2_2(mux_1634_nl, mux_1627_nl, fsm_output[0]);
  assign vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1650_nl,
      mux_1635_nl, fsm_output[3]);
  assign nor_1071_nl = ~((~ (fsm_output[5])) | (~ (VEC_LOOP_j_10_0_sva_9_0[3])) |
      (fsm_output[0]) | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (fsm_output[1]) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | (fsm_output[3:2]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2]) | (fsm_output[8:6]!=3'b000));
  assign nor_1072_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1]) | mux_1616_cse);
  assign nor_1073_nl = ~((COMP_LOOP_acc_20_psp_sva[1:0]!=2'b00) | nand_222_cse);
  assign nor_1074_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b100) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1675_nl = MUX_s_1_2_2(nor_1073_nl, nor_1074_nl, fsm_output[2]);
  assign nor_1075_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100) | (fsm_output[8:6]!=3'b011));
  assign nor_1076_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100) | (fsm_output[8:6]!=3'b001));
  assign mux_1674_nl = MUX_s_1_2_2(nor_1075_nl, nor_1076_nl, fsm_output[2]);
  assign mux_1676_nl = MUX_s_1_2_2(mux_1675_nl, mux_1674_nl, fsm_output[3]);
  assign mux_1679_nl = MUX_s_1_2_2(nor_1072_nl, mux_1676_nl, fsm_output[1]);
  assign and_524_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1679_nl;
  assign nor_1077_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]!=4'b1001) | nand_324_cse);
  assign nor_1078_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b1001) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1671_nl = MUX_s_1_2_2(nor_1077_nl, nor_1078_nl, fsm_output[2]);
  assign nor_1079_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b011));
  assign nor_1080_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b001));
  assign mux_1670_nl = MUX_s_1_2_2(nor_1079_nl, nor_1080_nl, fsm_output[2]);
  assign mux_1672_nl = MUX_s_1_2_2(mux_1671_nl, mux_1670_nl, fsm_output[3]);
  assign nor_1081_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b110));
  assign nor_1082_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b100));
  assign mux_1668_nl = MUX_s_1_2_2(nor_1081_nl, nor_1082_nl, fsm_output[2]);
  assign nor_1083_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b010));
  assign nor_1084_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b000));
  assign mux_1667_nl = MUX_s_1_2_2(nor_1083_nl, nor_1084_nl, fsm_output[2]);
  assign mux_1669_nl = MUX_s_1_2_2(mux_1668_nl, mux_1667_nl, fsm_output[3]);
  assign mux_1673_nl = MUX_s_1_2_2(mux_1672_nl, mux_1669_nl, fsm_output[1]);
  assign mux_1680_nl = MUX_s_1_2_2(and_524_nl, mux_1673_nl, fsm_output[0]);
  assign nor_1085_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[2:0]!=3'b001) | nand_223_cse);
  assign mux_1663_nl = MUX_s_1_2_2(nor_1085_nl, nor_1086_cse, fsm_output[2]);
  assign nor_1088_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b001));
  assign mux_1662_nl = MUX_s_1_2_2(nor_1056_cse, nor_1088_nl, fsm_output[2]);
  assign mux_1664_nl = MUX_s_1_2_2(mux_1663_nl, mux_1662_nl, fsm_output[3]);
  assign nor_1089_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b110));
  assign mux_1660_nl = MUX_s_1_2_2(nor_1089_nl, nor_1059_cse, fsm_output[2]);
  assign nor_1092_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b000));
  assign mux_1659_nl = MUX_s_1_2_2(nor_1060_cse, nor_1092_nl, fsm_output[2]);
  assign mux_1661_nl = MUX_s_1_2_2(mux_1660_nl, mux_1659_nl, fsm_output[3]);
  assign mux_1665_nl = MUX_s_1_2_2(mux_1664_nl, mux_1661_nl, fsm_output[1]);
  assign nor_1093_nl = ~((COMP_LOOP_acc_1_cse_sva[2:1]!=2'b00) | nand_212_cse);
  assign nor_1094_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1001) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1656_nl = MUX_s_1_2_2(nor_1093_nl, nor_1094_nl, fsm_output[2]);
  assign nor_1095_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b011));
  assign nor_1096_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b001));
  assign mux_1655_nl = MUX_s_1_2_2(nor_1095_nl, nor_1096_nl, fsm_output[2]);
  assign mux_1657_nl = MUX_s_1_2_2(mux_1656_nl, mux_1655_nl, fsm_output[3]);
  assign nor_1097_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b110));
  assign nor_1098_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b100));
  assign mux_1653_nl = MUX_s_1_2_2(nor_1097_nl, nor_1098_nl, fsm_output[2]);
  assign nor_1099_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b010));
  assign nor_1100_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b000));
  assign mux_1652_nl = MUX_s_1_2_2(nor_1099_nl, nor_1100_nl, fsm_output[2]);
  assign mux_1654_nl = MUX_s_1_2_2(mux_1653_nl, mux_1652_nl, fsm_output[3]);
  assign mux_1658_nl = MUX_s_1_2_2(mux_1657_nl, mux_1654_nl, fsm_output[1]);
  assign mux_1666_nl = MUX_s_1_2_2(mux_1665_nl, mux_1658_nl, fsm_output[0]);
  assign mux_1681_nl = MUX_s_1_2_2(mux_1680_nl, mux_1666_nl, fsm_output[5]);
  assign vec_rsc_0_9_i_we_d_pff = MUX_s_1_2_2(nor_1071_nl, mux_1681_nl, fsm_output[4]);
  assign nor_1039_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100)
      | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) | (fsm_output[2]) | (fsm_output[7])
      | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_1040_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b1001) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_1710_nl = MUX_s_1_2_2(nor_1039_nl, nor_1040_nl, fsm_output[5]);
  assign nor_1041_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b1001) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign nor_1042_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b1001) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1709_nl = MUX_s_1_2_2(nor_1041_nl, nor_1042_nl, fsm_output[5]);
  assign mux_1711_nl = MUX_s_1_2_2(mux_1710_nl, mux_1709_nl, fsm_output[1]);
  assign nor_1043_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b1001) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_1044_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1001)
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1707_nl = MUX_s_1_2_2(nor_1043_nl, nor_1044_nl, fsm_output[5]);
  assign nor_1045_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[3])) | (fsm_output[5]) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1708_nl = MUX_s_1_2_2(mux_1707_nl, nor_1045_nl, fsm_output[1]);
  assign mux_1712_nl = MUX_s_1_2_2(mux_1711_nl, mux_1708_nl, fsm_output[0]);
  assign nor_1046_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[2:0]!=3'b001) | nand_211_cse);
  assign nor_1047_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[2])) |
      (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b100) | (~ COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b110));
  assign mux_1704_nl = MUX_s_1_2_2(nor_1046_nl, nor_1047_nl, fsm_output[5]);
  assign nor_1048_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b1001) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign nor_1049_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (~ (fsm_output[2]))
      | (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (~ COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1703_nl = MUX_s_1_2_2(nor_1048_nl, nor_1049_nl, fsm_output[5]);
  assign mux_1705_nl = MUX_s_1_2_2(mux_1704_nl, mux_1703_nl, fsm_output[1]);
  assign nor_1050_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1001) | (~ COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm)
      | (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign nor_1051_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]!=4'b1001) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign mux_1701_nl = MUX_s_1_2_2(nor_1050_nl, nor_1051_nl, fsm_output[5]);
  assign nor_1052_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) | (COMP_LOOP_acc_1_cse_sva[2:1]!=2'b00)
      | nand_212_cse);
  assign nor_1053_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm)
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1699_nl = MUX_s_1_2_2(nor_1052_nl, nor_1053_nl, fsm_output[2]);
  assign nor_1054_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b1001) | (~ (fsm_output[2]))
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1700_nl = MUX_s_1_2_2(mux_1699_nl, nor_1054_nl, fsm_output[5]);
  assign mux_1702_nl = MUX_s_1_2_2(mux_1701_nl, mux_1700_nl, fsm_output[1]);
  assign mux_1706_nl = MUX_s_1_2_2(mux_1705_nl, mux_1702_nl, fsm_output[0]);
  assign mux_1713_nl = MUX_s_1_2_2(mux_1712_nl, mux_1706_nl, fsm_output[4]);
  assign mux_1695_nl = MUX_s_1_2_2(nor_1086_cse, nor_1056_cse, fsm_output[2]);
  assign nor_1057_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b100) | (~ COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b100));
  assign nor_1058_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b010));
  assign mux_1694_nl = MUX_s_1_2_2(nor_1057_nl, nor_1058_nl, fsm_output[2]);
  assign and_521_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1694_nl;
  assign mux_1696_nl = MUX_s_1_2_2(mux_1695_nl, and_521_nl, fsm_output[5]);
  assign mux_1692_nl = MUX_s_1_2_2(nor_1059_cse, nor_1060_cse, fsm_output[2]);
  assign and_522_nl = nor_351_cse & mux_1691_cse;
  assign mux_1693_nl = MUX_s_1_2_2(mux_1692_nl, and_522_nl, fsm_output[5]);
  assign mux_1697_nl = MUX_s_1_2_2(mux_1696_nl, mux_1693_nl, fsm_output[1]);
  assign nor_1063_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1001) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b100));
  assign nor_1064_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1001) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b010));
  assign mux_1687_nl = MUX_s_1_2_2(nor_1063_nl, nor_1064_nl, fsm_output[2]);
  assign nor_1065_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b100));
  assign nor_1066_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b010));
  assign mux_1686_nl = MUX_s_1_2_2(nor_1065_nl, nor_1066_nl, fsm_output[2]);
  assign mux_1688_nl = MUX_s_1_2_2(mux_1687_nl, mux_1686_nl, fsm_output[5]);
  assign nor_1067_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | (fsm_output[8:6]!=3'b011));
  assign nor_1068_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[8:6]!=3'b001));
  assign mux_1684_nl = MUX_s_1_2_2(nor_1067_nl, nor_1068_nl, fsm_output[2]);
  assign nor_1069_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b011));
  assign nor_1070_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b1001) | (fsm_output[8:6]!=3'b001));
  assign mux_1683_nl = MUX_s_1_2_2(nor_1069_nl, nor_1070_nl, fsm_output[2]);
  assign mux_1685_nl = MUX_s_1_2_2(mux_1684_nl, mux_1683_nl, fsm_output[5]);
  assign mux_1689_nl = MUX_s_1_2_2(mux_1688_nl, mux_1685_nl, fsm_output[1]);
  assign mux_1698_nl = MUX_s_1_2_2(mux_1697_nl, mux_1689_nl, fsm_output[0]);
  assign and_520_nl = (fsm_output[4]) & mux_1698_nl;
  assign vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1713_nl,
      and_520_nl, fsm_output[3]);
  assign nor_1010_nl = ~((~ (fsm_output[5])) | (~ (VEC_LOOP_j_10_0_sva_9_0[3])) |
      (fsm_output[0]) | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[1]) | (~ (VEC_LOOP_j_10_0_sva_9_0[1]))
      | (fsm_output[3:2]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2]) | (fsm_output[8:6]!=3'b000));
  assign nand_63_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1]) & mux_1741_cse);
  assign or_1728_nl = (COMP_LOOP_acc_20_psp_sva[1:0]!=2'b01) | nand_222_cse;
  assign or_1726_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b101) | (fsm_output[7]) |
      not_tmp_395;
  assign mux_1738_nl = MUX_s_1_2_2(or_1728_nl, or_1726_nl, fsm_output[2]);
  assign or_1724_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b101) | (fsm_output[8:6]!=3'b011);
  assign or_1723_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b101) | (fsm_output[8:6]!=3'b001);
  assign mux_1737_nl = MUX_s_1_2_2(or_1724_nl, or_1723_nl, fsm_output[2]);
  assign mux_1739_nl = MUX_s_1_2_2(mux_1738_nl, mux_1737_nl, fsm_output[3]);
  assign mux_1742_nl = MUX_s_1_2_2(nand_63_nl, mux_1739_nl, fsm_output[1]);
  assign nor_1011_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1742_nl);
  assign nor_1015_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[2]) | (~ (COMP_LOOP_acc_10_cse_10_1_15_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_15_sva[0]) | nand_268_cse);
  assign nor_1016_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b1010) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1734_nl = MUX_s_1_2_2(nor_1015_nl, nor_1016_nl, fsm_output[2]);
  assign nor_1017_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b011));
  assign nor_1018_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b001));
  assign mux_1733_nl = MUX_s_1_2_2(nor_1017_nl, nor_1018_nl, fsm_output[2]);
  assign mux_1735_nl = MUX_s_1_2_2(mux_1734_nl, mux_1733_nl, fsm_output[3]);
  assign nor_1019_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b110));
  assign nor_1020_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b100));
  assign mux_1731_nl = MUX_s_1_2_2(nor_1019_nl, nor_1020_nl, fsm_output[2]);
  assign nor_1021_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b010));
  assign nor_1022_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b000));
  assign mux_1730_nl = MUX_s_1_2_2(nor_1021_nl, nor_1022_nl, fsm_output[2]);
  assign mux_1732_nl = MUX_s_1_2_2(mux_1731_nl, mux_1730_nl, fsm_output[3]);
  assign mux_1736_nl = MUX_s_1_2_2(mux_1735_nl, mux_1732_nl, fsm_output[1]);
  assign mux_1743_nl = MUX_s_1_2_2(nor_1011_nl, mux_1736_nl, fsm_output[0]);
  assign nor_1023_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[2:0]!=3'b010) | nand_223_cse);
  assign nor_1024_nl = ~((COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b1010) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1726_nl = MUX_s_1_2_2(nor_1023_nl, nor_1024_nl, fsm_output[2]);
  assign nor_1025_nl = ~((COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b011));
  assign nor_1026_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b001));
  assign mux_1725_nl = MUX_s_1_2_2(nor_1025_nl, nor_1026_nl, fsm_output[2]);
  assign mux_1727_nl = MUX_s_1_2_2(mux_1726_nl, mux_1725_nl, fsm_output[3]);
  assign nor_1027_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b110));
  assign nor_1028_nl = ~((COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b100));
  assign mux_1723_nl = MUX_s_1_2_2(nor_1027_nl, nor_1028_nl, fsm_output[2]);
  assign nor_1029_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b010));
  assign nor_1030_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b000));
  assign mux_1722_nl = MUX_s_1_2_2(nor_1029_nl, nor_1030_nl, fsm_output[2]);
  assign mux_1724_nl = MUX_s_1_2_2(mux_1723_nl, mux_1722_nl, fsm_output[3]);
  assign mux_1728_nl = MUX_s_1_2_2(mux_1727_nl, mux_1724_nl, fsm_output[1]);
  assign nor_1031_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1010) | nand_324_cse);
  assign nor_1032_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1010) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1719_nl = MUX_s_1_2_2(nor_1031_nl, nor_1032_nl, fsm_output[2]);
  assign nor_1033_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b011));
  assign nor_1034_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b001));
  assign mux_1718_nl = MUX_s_1_2_2(nor_1033_nl, nor_1034_nl, fsm_output[2]);
  assign mux_1720_nl = MUX_s_1_2_2(mux_1719_nl, mux_1718_nl, fsm_output[3]);
  assign nor_1035_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b110));
  assign nor_1036_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b100));
  assign mux_1716_nl = MUX_s_1_2_2(nor_1035_nl, nor_1036_nl, fsm_output[2]);
  assign nor_1037_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b010));
  assign nor_1038_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1010) | (fsm_output[8:6]!=3'b000));
  assign mux_1715_nl = MUX_s_1_2_2(nor_1037_nl, nor_1038_nl, fsm_output[2]);
  assign mux_1717_nl = MUX_s_1_2_2(mux_1716_nl, mux_1715_nl, fsm_output[3]);
  assign mux_1721_nl = MUX_s_1_2_2(mux_1720_nl, mux_1717_nl, fsm_output[1]);
  assign mux_1729_nl = MUX_s_1_2_2(mux_1728_nl, mux_1721_nl, fsm_output[0]);
  assign mux_1744_nl = MUX_s_1_2_2(mux_1743_nl, mux_1729_nl, fsm_output[5]);
  assign vec_rsc_0_10_i_we_d_pff = MUX_s_1_2_2(nor_1010_nl, mux_1744_nl, fsm_output[4]);
  assign nor_983_nl = ~((~((fsm_output[5]) & (fsm_output[2]) & (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      & (COMP_LOOP_acc_20_psp_sva[2:0]==3'b101) & COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm))
      | nand_301_cse);
  assign nor_984_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b101) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_985_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[2:0]!=3'b010) | nand_219_cse);
  assign mux_1771_nl = MUX_s_1_2_2(nor_984_nl, nor_985_nl, fsm_output[2]);
  assign nor_986_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b1010) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1772_nl = MUX_s_1_2_2(mux_1771_nl, nor_986_nl, fsm_output[5]);
  assign mux_1773_nl = MUX_s_1_2_2(nor_983_nl, mux_1772_nl, fsm_output[6]);
  assign nor_987_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b1010) | (fsm_output[7])
      | (fsm_output[4]) | (fsm_output[8]));
  assign nor_988_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b1010) | nand_301_cse);
  assign mux_1768_nl = MUX_s_1_2_2(nor_987_nl, nor_988_nl, fsm_output[2]);
  assign nor_989_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b1010) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1769_nl = MUX_s_1_2_2(mux_1768_nl, nor_989_nl, fsm_output[5]);
  assign nor_990_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[1])) | (~ (fsm_output[5])) |
      (~ (fsm_output[2])) | (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (~ COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | not_tmp_399);
  assign mux_1770_nl = MUX_s_1_2_2(mux_1769_nl, nor_990_nl, fsm_output[6]);
  assign mux_1774_nl = MUX_s_1_2_2(mux_1773_nl, mux_1770_nl, fsm_output[1]);
  assign nor_991_nl = ~((~ (fsm_output[2])) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1010)
      | (~ COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm) | nand_301_cse);
  assign nor_992_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1010)
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_993_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[2]) | (~ (COMP_LOOP_acc_10_cse_10_1_15_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_15_sva[0]) | nand_265_cse);
  assign mux_1764_nl = MUX_s_1_2_2(nor_992_nl, nor_993_nl, fsm_output[2]);
  assign mux_1765_nl = MUX_s_1_2_2(nor_991_nl, mux_1764_nl, fsm_output[5]);
  assign nor_994_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b1010) | (fsm_output[5])
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1766_nl = MUX_s_1_2_2(mux_1765_nl, nor_994_nl, fsm_output[6]);
  assign nor_995_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[1])) | (~ (VEC_LOOP_j_10_0_sva_9_0[3]))
      | (fsm_output[5]) | (fsm_output[2]) | (VEC_LOOP_j_10_0_sva_9_0[2]) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_996_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) | (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1010)
      | nand_301_cse);
  assign nor_997_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm)
      | (fsm_output[7]) | not_tmp_399);
  assign mux_1761_nl = MUX_s_1_2_2(nor_996_nl, nor_997_nl, fsm_output[2]);
  assign nor_998_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b1010) | (~ (fsm_output[2]))
      | (fsm_output[7]) | not_tmp_399);
  assign mux_1762_nl = MUX_s_1_2_2(mux_1761_nl, nor_998_nl, fsm_output[5]);
  assign mux_1763_nl = MUX_s_1_2_2(nor_995_nl, mux_1762_nl, fsm_output[6]);
  assign mux_1767_nl = MUX_s_1_2_2(mux_1766_nl, mux_1763_nl, fsm_output[1]);
  assign mux_1775_nl = MUX_s_1_2_2(mux_1774_nl, mux_1767_nl, fsm_output[0]);
  assign nor_999_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b101) | (~ COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | not_tmp_399);
  assign nor_1000_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b101) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[7])) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign mux_1757_nl = MUX_s_1_2_2(nor_999_nl, nor_1000_nl, fsm_output[2]);
  assign and_517_nl = (fsm_output[5]) & mux_1757_nl;
  assign or_1755_nl = (COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b1010) | (fsm_output[7])
      | not_tmp_399;
  assign or_1753_nl = (COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b1010) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1756_nl = MUX_s_1_2_2(or_1755_nl, or_1753_nl, fsm_output[2]);
  assign nor_1001_nl = ~((fsm_output[5]) | mux_1756_nl);
  assign mux_1758_nl = MUX_s_1_2_2(and_517_nl, nor_1001_nl, fsm_output[6]);
  assign or_1751_nl = (COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b1010) | (fsm_output[7])
      | not_tmp_399;
  assign or_1749_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b1010) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1754_nl = MUX_s_1_2_2(or_1751_nl, or_1749_nl, fsm_output[2]);
  assign nor_1002_nl = ~((fsm_output[5]) | mux_1754_nl);
  assign and_518_nl = (VEC_LOOP_j_10_0_sva_9_0[1]) & (fsm_output[5]) & mux_1628_cse;
  assign mux_1755_nl = MUX_s_1_2_2(nor_1002_nl, and_518_nl, fsm_output[6]);
  assign mux_1759_nl = MUX_s_1_2_2(mux_1758_nl, mux_1755_nl, fsm_output[1]);
  assign or_1745_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1010) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7]) | not_tmp_399;
  assign or_1743_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1010) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1750_nl = MUX_s_1_2_2(or_1745_nl, or_1743_nl, fsm_output[2]);
  assign or_1742_nl = (COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b1010) | (fsm_output[7])
      | not_tmp_399;
  assign or_1740_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b1010) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1749_nl = MUX_s_1_2_2(or_1742_nl, or_1740_nl, fsm_output[2]);
  assign mux_1751_nl = MUX_s_1_2_2(mux_1750_nl, mux_1749_nl, fsm_output[5]);
  assign nor_1005_nl = ~((fsm_output[6]) | mux_1751_nl);
  assign nor_1006_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_1007_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7]) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_1747_nl = MUX_s_1_2_2(nor_1006_nl, nor_1007_nl, fsm_output[2]);
  assign nor_1008_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b1010) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_1009_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b1010) | (fsm_output[7])
      | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_1746_nl = MUX_s_1_2_2(nor_1008_nl, nor_1009_nl, fsm_output[2]);
  assign mux_1748_nl = MUX_s_1_2_2(mux_1747_nl, mux_1746_nl, fsm_output[5]);
  assign and_519_nl = (fsm_output[6]) & mux_1748_nl;
  assign mux_1752_nl = MUX_s_1_2_2(nor_1005_nl, and_519_nl, fsm_output[1]);
  assign mux_1760_nl = MUX_s_1_2_2(mux_1759_nl, mux_1752_nl, fsm_output[0]);
  assign vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1775_nl,
      mux_1760_nl, fsm_output[3]);
  assign nor_954_nl = ~((~ (fsm_output[5])) | (~ (VEC_LOOP_j_10_0_sva_9_0[3])) |
      (fsm_output[0]) | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (fsm_output[1]) | (~ (VEC_LOOP_j_10_0_sva_9_0[1]))
      | (fsm_output[3:2]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2]) | (fsm_output[8:6]!=3'b000));
  assign and_513_nl = (VEC_LOOP_j_10_0_sva_9_0[1]) & mux_1741_cse;
  assign nor_958_nl = ~((COMP_LOOP_acc_20_psp_sva[1:0]!=2'b01) | nand_222_cse);
  assign nor_959_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b101) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1800_nl = MUX_s_1_2_2(nor_958_nl, nor_959_nl, fsm_output[2]);
  assign nor_960_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b101) | (fsm_output[8:6]!=3'b011));
  assign nor_961_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b101) | (fsm_output[8:6]!=3'b001));
  assign mux_1799_nl = MUX_s_1_2_2(nor_960_nl, nor_961_nl, fsm_output[2]);
  assign mux_1801_nl = MUX_s_1_2_2(mux_1800_nl, mux_1799_nl, fsm_output[3]);
  assign mux_1804_nl = MUX_s_1_2_2(and_513_nl, mux_1801_nl, fsm_output[1]);
  assign and_512_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1804_nl;
  assign nor_962_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[2]) | (~((COMP_LOOP_acc_10_cse_10_1_15_sva[3])
      & (COMP_LOOP_acc_10_cse_10_1_15_sva[0]) & (COMP_LOOP_acc_10_cse_10_1_15_sva[1])
      & (fsm_output[8:6]==3'b111))));
  assign nor_963_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b1011) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1796_nl = MUX_s_1_2_2(nor_962_nl, nor_963_nl, fsm_output[2]);
  assign and_514_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]==4'b1011) & (fsm_output[8:6]==3'b011);
  assign nor_964_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b1011) | (fsm_output[8:6]!=3'b001));
  assign mux_1795_nl = MUX_s_1_2_2(and_514_nl, nor_964_nl, fsm_output[2]);
  assign mux_1797_nl = MUX_s_1_2_2(mux_1796_nl, mux_1795_nl, fsm_output[3]);
  assign and_841_nl = (COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]==4'b1011) & (fsm_output[8:6]==3'b110);
  assign nor_966_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b1011) | (fsm_output[8:6]!=3'b100));
  assign mux_1793_nl = MUX_s_1_2_2(and_841_nl, nor_966_nl, fsm_output[2]);
  assign nor_967_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b1011) | (fsm_output[8:6]!=3'b010));
  assign nor_968_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[3:0]!=4'b1011) | (fsm_output[8:6]!=3'b000));
  assign mux_1792_nl = MUX_s_1_2_2(nor_967_nl, nor_968_nl, fsm_output[2]);
  assign mux_1794_nl = MUX_s_1_2_2(mux_1793_nl, mux_1792_nl, fsm_output[3]);
  assign mux_1798_nl = MUX_s_1_2_2(mux_1797_nl, mux_1794_nl, fsm_output[1]);
  assign mux_1805_nl = MUX_s_1_2_2(and_512_nl, mux_1798_nl, fsm_output[0]);
  assign nor_969_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[2:0]!=3'b011) | nand_223_cse);
  assign mux_1788_nl = MUX_s_1_2_2(nor_969_nl, nor_970_cse, fsm_output[2]);
  assign nor_971_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b1011) | (fsm_output[8:6]!=3'b001));
  assign mux_1787_nl = MUX_s_1_2_2(and_506_cse, nor_971_nl, fsm_output[2]);
  assign mux_1789_nl = MUX_s_1_2_2(mux_1788_nl, mux_1787_nl, fsm_output[3]);
  assign and_851_nl = (COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]==4'b1011) & (fsm_output[8:6]==3'b110);
  assign mux_1785_nl = MUX_s_1_2_2(and_851_nl, nor_944_cse, fsm_output[2]);
  assign nor_975_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b1011) | (fsm_output[8:6]!=3'b000));
  assign mux_1784_nl = MUX_s_1_2_2(nor_945_cse, nor_975_nl, fsm_output[2]);
  assign mux_1786_nl = MUX_s_1_2_2(mux_1785_nl, mux_1784_nl, fsm_output[3]);
  assign mux_1790_nl = MUX_s_1_2_2(mux_1789_nl, mux_1786_nl, fsm_output[1]);
  assign nor_976_nl = ~((COMP_LOOP_acc_1_cse_sva[2:1]!=2'b01) | nand_212_cse);
  assign nor_977_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1011) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1781_nl = MUX_s_1_2_2(nor_976_nl, nor_977_nl, fsm_output[2]);
  assign and_516_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b1011) & (fsm_output[8:6]==3'b011);
  assign nor_978_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1011) | (fsm_output[8:6]!=3'b001));
  assign mux_1780_nl = MUX_s_1_2_2(and_516_nl, nor_978_nl, fsm_output[2]);
  assign mux_1782_nl = MUX_s_1_2_2(mux_1781_nl, mux_1780_nl, fsm_output[3]);
  assign and_869_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1011) & (fsm_output[8:6]==3'b110);
  assign nor_980_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1011) | (fsm_output[8:6]!=3'b100));
  assign mux_1778_nl = MUX_s_1_2_2(and_869_nl, nor_980_nl, fsm_output[2]);
  assign nor_981_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1011) | (fsm_output[8:6]!=3'b010));
  assign nor_982_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1011) | (fsm_output[8:6]!=3'b000));
  assign mux_1777_nl = MUX_s_1_2_2(nor_981_nl, nor_982_nl, fsm_output[2]);
  assign mux_1779_nl = MUX_s_1_2_2(mux_1778_nl, mux_1777_nl, fsm_output[3]);
  assign mux_1783_nl = MUX_s_1_2_2(mux_1782_nl, mux_1779_nl, fsm_output[1]);
  assign mux_1791_nl = MUX_s_1_2_2(mux_1790_nl, mux_1783_nl, fsm_output[0]);
  assign mux_1806_nl = MUX_s_1_2_2(mux_1805_nl, mux_1791_nl, fsm_output[5]);
  assign vec_rsc_0_11_i_we_d_pff = MUX_s_1_2_2(nor_954_nl, mux_1806_nl, fsm_output[4]);
  assign nor_925_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b101)
      | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) | (fsm_output[2]) | (fsm_output[7])
      | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_926_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b1011) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_1835_nl = MUX_s_1_2_2(nor_925_nl, nor_926_nl, fsm_output[5]);
  assign nor_927_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b1011) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign nor_928_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b1011) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1834_nl = MUX_s_1_2_2(nor_927_nl, nor_928_nl, fsm_output[5]);
  assign mux_1836_nl = MUX_s_1_2_2(mux_1835_nl, mux_1834_nl, fsm_output[1]);
  assign nor_929_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b1011) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_930_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1011)
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1832_nl = MUX_s_1_2_2(nor_929_nl, nor_930_nl, fsm_output[5]);
  assign nor_931_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[3])) | (fsm_output[5]) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1833_nl = MUX_s_1_2_2(mux_1832_nl, nor_931_nl, fsm_output[1]);
  assign mux_1837_nl = MUX_s_1_2_2(mux_1836_nl, mux_1833_nl, fsm_output[0]);
  assign nor_932_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[2:0]!=3'b011) | nand_211_cse);
  assign and_850_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (fsm_output[2]) & (COMP_LOOP_acc_20_psp_sva[2:0]==3'b101)
      & COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm & (fsm_output[8:6]==3'b110);
  assign mux_1829_nl = MUX_s_1_2_2(nor_932_nl, and_850_nl, fsm_output[5]);
  assign and_857_nl = (COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]==4'b1011) & (fsm_output[2])
      & (fsm_output[7]) & (~ (fsm_output[6])) & (fsm_output[8]);
  assign nor_935_nl = ~((~((VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & (fsm_output[2])
      & (COMP_LOOP_acc_19_psp_sva[1:0]==2'b10) & COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm
      & (~ (fsm_output[7])))) | not_tmp_395);
  assign mux_1828_nl = MUX_s_1_2_2(and_857_nl, nor_935_nl, fsm_output[5]);
  assign mux_1830_nl = MUX_s_1_2_2(mux_1829_nl, mux_1828_nl, fsm_output[1]);
  assign and_867_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1011) & COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[2]) & (fsm_output[7]) & (~ (fsm_output[6])) & (fsm_output[8]);
  assign and_868_nl = (COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]==4'b1011) & (fsm_output[2])
      & (fsm_output[7]) & (~ (fsm_output[6])) & (fsm_output[8]);
  assign mux_1826_nl = MUX_s_1_2_2(and_867_nl, and_868_nl, fsm_output[5]);
  assign nor_938_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) | (COMP_LOOP_acc_1_cse_sva[2:1]!=2'b01)
      | nand_212_cse);
  assign nor_939_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm)
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1824_nl = MUX_s_1_2_2(nor_938_nl, nor_939_nl, fsm_output[2]);
  assign nor_940_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b1011) | (~ (fsm_output[2]))
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1825_nl = MUX_s_1_2_2(mux_1824_nl, nor_940_nl, fsm_output[5]);
  assign mux_1827_nl = MUX_s_1_2_2(mux_1826_nl, mux_1825_nl, fsm_output[1]);
  assign mux_1831_nl = MUX_s_1_2_2(mux_1830_nl, mux_1827_nl, fsm_output[0]);
  assign mux_1838_nl = MUX_s_1_2_2(mux_1837_nl, mux_1831_nl, fsm_output[4]);
  assign mux_1820_nl = MUX_s_1_2_2(nor_970_cse, and_506_cse, fsm_output[2]);
  assign nor_942_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b101) | (~ COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b100));
  assign nor_943_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b101) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b010));
  assign mux_1819_nl = MUX_s_1_2_2(nor_942_nl, nor_943_nl, fsm_output[2]);
  assign and_507_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1819_nl;
  assign mux_1821_nl = MUX_s_1_2_2(mux_1820_nl, and_507_nl, fsm_output[5]);
  assign mux_1817_nl = MUX_s_1_2_2(nor_944_cse, nor_945_cse, fsm_output[2]);
  assign and_508_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & mux_1691_cse;
  assign mux_1818_nl = MUX_s_1_2_2(mux_1817_nl, and_508_nl, fsm_output[5]);
  assign mux_1822_nl = MUX_s_1_2_2(mux_1821_nl, mux_1818_nl, fsm_output[1]);
  assign nor_948_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1011) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b100));
  assign nor_949_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1011) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b010));
  assign mux_1812_nl = MUX_s_1_2_2(nor_948_nl, nor_949_nl, fsm_output[2]);
  assign nor_950_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b1011) | (fsm_output[8:6]!=3'b100));
  assign nor_951_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b1011) | (fsm_output[8:6]!=3'b010));
  assign mux_1811_nl = MUX_s_1_2_2(nor_950_nl, nor_951_nl, fsm_output[2]);
  assign mux_1813_nl = MUX_s_1_2_2(mux_1812_nl, mux_1811_nl, fsm_output[5]);
  assign and_510_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b1011) & COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm
      & (fsm_output[8:6]==3'b011);
  assign nor_952_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[8:6]!=3'b001));
  assign mux_1809_nl = MUX_s_1_2_2(and_510_nl, nor_952_nl, fsm_output[2]);
  assign and_511_nl = (COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]==4'b1011) & (fsm_output[8:6]==3'b011);
  assign nor_953_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b1011) | (fsm_output[8:6]!=3'b001));
  assign mux_1808_nl = MUX_s_1_2_2(and_511_nl, nor_953_nl, fsm_output[2]);
  assign mux_1810_nl = MUX_s_1_2_2(mux_1809_nl, mux_1808_nl, fsm_output[5]);
  assign mux_1814_nl = MUX_s_1_2_2(mux_1813_nl, mux_1810_nl, fsm_output[1]);
  assign mux_1823_nl = MUX_s_1_2_2(mux_1822_nl, mux_1814_nl, fsm_output[0]);
  assign and_505_nl = (fsm_output[4]) & mux_1823_nl;
  assign vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1838_nl,
      and_505_nl, fsm_output[3]);
  assign nor_899_nl = ~((~ (fsm_output[5])) | (~ (VEC_LOOP_j_10_0_sva_9_0[3])) |
      (fsm_output[0]) | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[1]) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | (fsm_output[3:2]!=2'b00) | (~ (VEC_LOOP_j_10_0_sva_9_0[2])) | (fsm_output[8:6]!=3'b000));
  assign or_1925_nl = (VEC_LOOP_j_10_0_sva_9_0[1]) | mux_1866_cse;
  assign or_1919_nl = (COMP_LOOP_acc_20_psp_sva[0]) | nand_184_cse;
  assign or_1918_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b110) | (fsm_output[7]) |
      not_tmp_395;
  assign mux_1863_nl = MUX_s_1_2_2(or_1919_nl, or_1918_nl, fsm_output[2]);
  assign or_1916_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b110) | (fsm_output[8:6]!=3'b011);
  assign or_1915_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b110) | (fsm_output[8:6]!=3'b001);
  assign mux_1862_nl = MUX_s_1_2_2(or_1916_nl, or_1915_nl, fsm_output[2]);
  assign mux_1864_nl = MUX_s_1_2_2(mux_1863_nl, mux_1862_nl, fsm_output[3]);
  assign mux_1867_nl = MUX_s_1_2_2(or_1925_nl, mux_1864_nl, fsm_output[1]);
  assign nor_900_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1867_nl);
  assign nor_901_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]!=4'b1100) | nand_324_cse);
  assign nor_902_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b1100) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1859_nl = MUX_s_1_2_2(nor_901_nl, nor_902_nl, fsm_output[2]);
  assign nor_903_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b011));
  assign nor_904_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b001));
  assign mux_1858_nl = MUX_s_1_2_2(nor_903_nl, nor_904_nl, fsm_output[2]);
  assign mux_1860_nl = MUX_s_1_2_2(mux_1859_nl, mux_1858_nl, fsm_output[3]);
  assign nor_905_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b110));
  assign nor_906_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b100));
  assign mux_1856_nl = MUX_s_1_2_2(nor_905_nl, nor_906_nl, fsm_output[2]);
  assign nor_907_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b010));
  assign nor_908_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b000));
  assign mux_1855_nl = MUX_s_1_2_2(nor_907_nl, nor_908_nl, fsm_output[2]);
  assign mux_1857_nl = MUX_s_1_2_2(mux_1856_nl, mux_1855_nl, fsm_output[3]);
  assign mux_1861_nl = MUX_s_1_2_2(mux_1860_nl, mux_1857_nl, fsm_output[1]);
  assign mux_1868_nl = MUX_s_1_2_2(nor_900_nl, mux_1861_nl, fsm_output[0]);
  assign nor_909_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[1:0]!=2'b00) | nand_185_cse);
  assign nor_910_nl = ~((COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b1100) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1851_nl = MUX_s_1_2_2(nor_909_nl, nor_910_nl, fsm_output[2]);
  assign nor_911_nl = ~((COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b011));
  assign nor_912_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b001));
  assign mux_1850_nl = MUX_s_1_2_2(nor_911_nl, nor_912_nl, fsm_output[2]);
  assign mux_1852_nl = MUX_s_1_2_2(mux_1851_nl, mux_1850_nl, fsm_output[3]);
  assign nor_913_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b110));
  assign nor_914_nl = ~((COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b100));
  assign mux_1848_nl = MUX_s_1_2_2(nor_913_nl, nor_914_nl, fsm_output[2]);
  assign nor_915_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b010));
  assign nor_916_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b000));
  assign mux_1847_nl = MUX_s_1_2_2(nor_915_nl, nor_916_nl, fsm_output[2]);
  assign mux_1849_nl = MUX_s_1_2_2(mux_1848_nl, mux_1847_nl, fsm_output[3]);
  assign mux_1853_nl = MUX_s_1_2_2(mux_1852_nl, mux_1849_nl, fsm_output[1]);
  assign nor_917_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1100) | nand_324_cse);
  assign nor_918_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1100) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1844_nl = MUX_s_1_2_2(nor_917_nl, nor_918_nl, fsm_output[2]);
  assign nor_919_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b011));
  assign nor_920_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b001));
  assign mux_1843_nl = MUX_s_1_2_2(nor_919_nl, nor_920_nl, fsm_output[2]);
  assign mux_1845_nl = MUX_s_1_2_2(mux_1844_nl, mux_1843_nl, fsm_output[3]);
  assign nor_921_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b110));
  assign nor_922_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b100));
  assign mux_1841_nl = MUX_s_1_2_2(nor_921_nl, nor_922_nl, fsm_output[2]);
  assign nor_923_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b010));
  assign nor_924_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1100) | (fsm_output[8:6]!=3'b000));
  assign mux_1840_nl = MUX_s_1_2_2(nor_923_nl, nor_924_nl, fsm_output[2]);
  assign mux_1842_nl = MUX_s_1_2_2(mux_1841_nl, mux_1840_nl, fsm_output[3]);
  assign mux_1846_nl = MUX_s_1_2_2(mux_1845_nl, mux_1842_nl, fsm_output[1]);
  assign mux_1854_nl = MUX_s_1_2_2(mux_1853_nl, mux_1846_nl, fsm_output[0]);
  assign mux_1869_nl = MUX_s_1_2_2(mux_1868_nl, mux_1854_nl, fsm_output[5]);
  assign vec_rsc_0_12_i_we_d_pff = MUX_s_1_2_2(nor_899_nl, mux_1869_nl, fsm_output[4]);
  assign nor_873_nl = ~((~((fsm_output[5]) & (fsm_output[2]) & (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      & (COMP_LOOP_acc_20_psp_sva[2:0]==3'b110) & COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm))
      | nand_301_cse);
  assign nor_874_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b110) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_875_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[1:0]!=2'b00) | (~((COMP_LOOP_acc_10_cse_10_1_sva[3:2]==2'b11)
      & (fsm_output[7]) & (fsm_output[4]) & (fsm_output[8]))));
  assign mux_1896_nl = MUX_s_1_2_2(nor_874_nl, nor_875_nl, fsm_output[2]);
  assign nor_876_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b1100) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1897_nl = MUX_s_1_2_2(mux_1896_nl, nor_876_nl, fsm_output[5]);
  assign mux_1898_nl = MUX_s_1_2_2(nor_873_nl, mux_1897_nl, fsm_output[6]);
  assign nor_877_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b1100) | (fsm_output[7])
      | (fsm_output[4]) | (fsm_output[8]));
  assign nor_878_nl = ~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]!=4'b1100) | nand_301_cse);
  assign mux_1893_nl = MUX_s_1_2_2(nor_877_nl, nor_878_nl, fsm_output[2]);
  assign nor_879_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b1100) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1894_nl = MUX_s_1_2_2(mux_1893_nl, nor_879_nl, fsm_output[5]);
  assign nor_880_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1]) | (~ (fsm_output[5])) | (~ (fsm_output[2]))
      | (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (~ COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | not_tmp_399);
  assign mux_1895_nl = MUX_s_1_2_2(mux_1894_nl, nor_880_nl, fsm_output[6]);
  assign mux_1899_nl = MUX_s_1_2_2(mux_1898_nl, mux_1895_nl, fsm_output[1]);
  assign nor_881_nl = ~((~ (fsm_output[2])) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1100)
      | (~ COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm) | nand_301_cse);
  assign nor_882_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1100)
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_883_nl = ~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]!=4'b1100) | nand_301_cse);
  assign mux_1889_nl = MUX_s_1_2_2(nor_882_nl, nor_883_nl, fsm_output[2]);
  assign mux_1890_nl = MUX_s_1_2_2(nor_881_nl, mux_1889_nl, fsm_output[5]);
  assign nor_884_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b1100) | (fsm_output[5])
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_1891_nl = MUX_s_1_2_2(mux_1890_nl, nor_884_nl, fsm_output[6]);
  assign nor_885_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1]) | (~ (VEC_LOOP_j_10_0_sva_9_0[3]))
      | (fsm_output[5]) | (fsm_output[2]) | (~ (VEC_LOOP_j_10_0_sva_9_0[2])) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_886_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) | (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1100)
      | nand_301_cse);
  assign nor_887_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm)
      | (fsm_output[7]) | not_tmp_399);
  assign mux_1886_nl = MUX_s_1_2_2(nor_886_nl, nor_887_nl, fsm_output[2]);
  assign nor_888_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b1100) | (~ (fsm_output[2]))
      | (fsm_output[7]) | not_tmp_399);
  assign mux_1887_nl = MUX_s_1_2_2(mux_1886_nl, nor_888_nl, fsm_output[5]);
  assign mux_1888_nl = MUX_s_1_2_2(nor_885_nl, mux_1887_nl, fsm_output[6]);
  assign mux_1892_nl = MUX_s_1_2_2(mux_1891_nl, mux_1888_nl, fsm_output[1]);
  assign mux_1900_nl = MUX_s_1_2_2(mux_1899_nl, mux_1892_nl, fsm_output[0]);
  assign nor_889_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b110) | (~ COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | not_tmp_399);
  assign nor_890_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b110) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[7])) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign mux_1882_nl = MUX_s_1_2_2(nor_889_nl, nor_890_nl, fsm_output[2]);
  assign and_501_nl = (fsm_output[5]) & mux_1882_nl;
  assign or_1947_nl = (COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b1100) | (fsm_output[7])
      | not_tmp_399;
  assign or_1945_nl = (COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]!=4'b1100) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1881_nl = MUX_s_1_2_2(or_1947_nl, or_1945_nl, fsm_output[2]);
  assign nor_891_nl = ~((fsm_output[5]) | mux_1881_nl);
  assign mux_1883_nl = MUX_s_1_2_2(and_501_nl, nor_891_nl, fsm_output[6]);
  assign or_1943_nl = (COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b1100) | (fsm_output[7])
      | not_tmp_399;
  assign or_1941_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b1100) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1879_nl = MUX_s_1_2_2(or_1943_nl, or_1941_nl, fsm_output[2]);
  assign nor_892_nl = ~((fsm_output[5]) | mux_1879_nl);
  assign and_502_nl = nor_346_cse & mux_1878_cse;
  assign mux_1880_nl = MUX_s_1_2_2(nor_892_nl, and_502_nl, fsm_output[6]);
  assign mux_1884_nl = MUX_s_1_2_2(mux_1883_nl, mux_1880_nl, fsm_output[1]);
  assign or_1937_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1100) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7]) | not_tmp_399;
  assign or_1935_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1100) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1875_nl = MUX_s_1_2_2(or_1937_nl, or_1935_nl, fsm_output[2]);
  assign or_1934_nl = (COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b1100) | (fsm_output[7])
      | not_tmp_399;
  assign or_1932_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b1100) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1874_nl = MUX_s_1_2_2(or_1934_nl, or_1932_nl, fsm_output[2]);
  assign mux_1876_nl = MUX_s_1_2_2(mux_1875_nl, mux_1874_nl, fsm_output[5]);
  assign nor_894_nl = ~((fsm_output[6]) | mux_1876_nl);
  assign nor_895_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | (~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_896_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7]) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_1872_nl = MUX_s_1_2_2(nor_895_nl, nor_896_nl, fsm_output[2]);
  assign nor_897_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b1100) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_898_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b1100) | (fsm_output[7])
      | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_1871_nl = MUX_s_1_2_2(nor_897_nl, nor_898_nl, fsm_output[2]);
  assign mux_1873_nl = MUX_s_1_2_2(mux_1872_nl, mux_1871_nl, fsm_output[5]);
  assign and_504_nl = (fsm_output[6]) & mux_1873_nl;
  assign mux_1877_nl = MUX_s_1_2_2(nor_894_nl, and_504_nl, fsm_output[1]);
  assign mux_1885_nl = MUX_s_1_2_2(mux_1884_nl, mux_1877_nl, fsm_output[0]);
  assign vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1900_nl,
      mux_1885_nl, fsm_output[3]);
  assign nor_846_nl = ~((~ (fsm_output[5])) | (~ (VEC_LOOP_j_10_0_sva_9_0[3])) |
      (fsm_output[0]) | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (fsm_output[1]) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | (fsm_output[3:2]!=2'b00) | (~ (VEC_LOOP_j_10_0_sva_9_0[2])) | (fsm_output[8:6]!=3'b000));
  assign nor_847_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1]) | mux_1866_cse);
  assign nor_848_nl = ~((COMP_LOOP_acc_20_psp_sva[0]) | nand_184_cse);
  assign nor_849_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b110) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1925_nl = MUX_s_1_2_2(nor_848_nl, nor_849_nl, fsm_output[2]);
  assign nor_850_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b110) | (fsm_output[8:6]!=3'b011));
  assign nor_851_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b110) | (fsm_output[8:6]!=3'b001));
  assign mux_1924_nl = MUX_s_1_2_2(nor_850_nl, nor_851_nl, fsm_output[2]);
  assign mux_1926_nl = MUX_s_1_2_2(mux_1925_nl, mux_1924_nl, fsm_output[3]);
  assign mux_1929_nl = MUX_s_1_2_2(nor_847_nl, mux_1926_nl, fsm_output[1]);
  assign and_497_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1929_nl;
  assign nor_852_nl = ~((~((COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]==4'b1101))) | nand_324_cse);
  assign nor_853_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b1101) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1921_nl = MUX_s_1_2_2(nor_852_nl, nor_853_nl, fsm_output[2]);
  assign and_498_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]==4'b1101) & (fsm_output[8:6]==3'b011);
  assign nor_854_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b1101) | (fsm_output[8:6]!=3'b001));
  assign mux_1920_nl = MUX_s_1_2_2(and_498_nl, nor_854_nl, fsm_output[2]);
  assign mux_1922_nl = MUX_s_1_2_2(mux_1921_nl, mux_1920_nl, fsm_output[3]);
  assign and_840_nl = (COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]==4'b1101) & (fsm_output[8:6]==3'b110);
  assign nor_856_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b1101) | (fsm_output[8:6]!=3'b100));
  assign mux_1918_nl = MUX_s_1_2_2(and_840_nl, nor_856_nl, fsm_output[2]);
  assign nor_857_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b1101) | (fsm_output[8:6]!=3'b010));
  assign nor_858_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[3:0]!=4'b1101) | (fsm_output[8:6]!=3'b000));
  assign mux_1917_nl = MUX_s_1_2_2(nor_857_nl, nor_858_nl, fsm_output[2]);
  assign mux_1919_nl = MUX_s_1_2_2(mux_1918_nl, mux_1917_nl, fsm_output[3]);
  assign mux_1923_nl = MUX_s_1_2_2(mux_1922_nl, mux_1919_nl, fsm_output[1]);
  assign mux_1930_nl = MUX_s_1_2_2(and_497_nl, mux_1923_nl, fsm_output[0]);
  assign nor_859_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[1:0]!=2'b01) | nand_185_cse);
  assign mux_1913_nl = MUX_s_1_2_2(nor_859_nl, nor_860_cse, fsm_output[2]);
  assign nor_861_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b1101) | (fsm_output[8:6]!=3'b001));
  assign mux_1912_nl = MUX_s_1_2_2(and_490_cse, nor_861_nl, fsm_output[2]);
  assign mux_1914_nl = MUX_s_1_2_2(mux_1913_nl, mux_1912_nl, fsm_output[3]);
  assign and_849_nl = (COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]==4'b1101) & (fsm_output[8:6]==3'b110);
  assign mux_1910_nl = MUX_s_1_2_2(and_849_nl, nor_837_cse, fsm_output[2]);
  assign nor_865_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b1101) | (fsm_output[8:6]!=3'b000));
  assign mux_1909_nl = MUX_s_1_2_2(nor_838_cse, nor_865_nl, fsm_output[2]);
  assign mux_1911_nl = MUX_s_1_2_2(mux_1910_nl, mux_1909_nl, fsm_output[3]);
  assign mux_1915_nl = MUX_s_1_2_2(mux_1914_nl, mux_1911_nl, fsm_output[1]);
  assign nor_866_nl = ~((COMP_LOOP_acc_1_cse_sva[1]) | nand_170_cse);
  assign nor_867_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1101) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1906_nl = MUX_s_1_2_2(nor_866_nl, nor_867_nl, fsm_output[2]);
  assign and_500_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b1101) & (fsm_output[8:6]==3'b011);
  assign nor_868_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1101) | (fsm_output[8:6]!=3'b001));
  assign mux_1905_nl = MUX_s_1_2_2(and_500_nl, nor_868_nl, fsm_output[2]);
  assign mux_1907_nl = MUX_s_1_2_2(mux_1906_nl, mux_1905_nl, fsm_output[3]);
  assign and_866_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1101) & (fsm_output[8:6]==3'b110);
  assign nor_870_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1101) | (fsm_output[8:6]!=3'b100));
  assign mux_1903_nl = MUX_s_1_2_2(and_866_nl, nor_870_nl, fsm_output[2]);
  assign nor_871_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1101) | (fsm_output[8:6]!=3'b010));
  assign nor_872_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1101) | (fsm_output[8:6]!=3'b000));
  assign mux_1902_nl = MUX_s_1_2_2(nor_871_nl, nor_872_nl, fsm_output[2]);
  assign mux_1904_nl = MUX_s_1_2_2(mux_1903_nl, mux_1902_nl, fsm_output[3]);
  assign mux_1908_nl = MUX_s_1_2_2(mux_1907_nl, mux_1904_nl, fsm_output[1]);
  assign mux_1916_nl = MUX_s_1_2_2(mux_1915_nl, mux_1908_nl, fsm_output[0]);
  assign mux_1931_nl = MUX_s_1_2_2(mux_1930_nl, mux_1916_nl, fsm_output[5]);
  assign vec_rsc_0_13_i_we_d_pff = MUX_s_1_2_2(nor_846_nl, mux_1931_nl, fsm_output[4]);
  assign nor_818_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b110)
      | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) | (fsm_output[2]) | (fsm_output[7])
      | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_819_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b1101) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_1960_nl = MUX_s_1_2_2(nor_818_nl, nor_819_nl, fsm_output[5]);
  assign nor_820_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b1101) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign nor_821_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b1101) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1959_nl = MUX_s_1_2_2(nor_820_nl, nor_821_nl, fsm_output[5]);
  assign mux_1961_nl = MUX_s_1_2_2(mux_1960_nl, mux_1959_nl, fsm_output[1]);
  assign nor_822_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b1101) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_823_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1101)
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1957_nl = MUX_s_1_2_2(nor_822_nl, nor_823_nl, fsm_output[5]);
  assign nor_824_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[3])) | (fsm_output[5]) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_1958_nl = MUX_s_1_2_2(mux_1957_nl, nor_824_nl, fsm_output[1]);
  assign mux_1962_nl = MUX_s_1_2_2(mux_1961_nl, mux_1958_nl, fsm_output[0]);
  assign nor_825_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[1:0]!=2'b01) | (~((COMP_LOOP_acc_10_cse_10_1_sva[3:2]==2'b11)
      & (fsm_output[2]) & (fsm_output[7]) & (fsm_output[6]) & (fsm_output[8]))));
  assign and_848_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (fsm_output[2]) & (COMP_LOOP_acc_20_psp_sva[2:0]==3'b110)
      & COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm & (fsm_output[8:6]==3'b110);
  assign mux_1954_nl = MUX_s_1_2_2(nor_825_nl, and_848_nl, fsm_output[5]);
  assign and_856_nl = (COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]==4'b1101) & (fsm_output[2])
      & (fsm_output[7]) & (~ (fsm_output[6])) & (fsm_output[8]);
  assign nor_828_nl = ~((~((VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b01) & (fsm_output[2])
      & (COMP_LOOP_acc_19_psp_sva[1:0]==2'b11) & COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm
      & (~ (fsm_output[7])))) | not_tmp_395);
  assign mux_1953_nl = MUX_s_1_2_2(and_856_nl, nor_828_nl, fsm_output[5]);
  assign mux_1955_nl = MUX_s_1_2_2(mux_1954_nl, mux_1953_nl, fsm_output[1]);
  assign and_864_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1101) & COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[2]) & (fsm_output[7]) & (~ (fsm_output[6])) & (fsm_output[8]);
  assign and_865_nl = (COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]==4'b1101) & (fsm_output[2])
      & (fsm_output[7]) & (~ (fsm_output[6])) & (fsm_output[8]);
  assign mux_1951_nl = MUX_s_1_2_2(and_864_nl, and_865_nl, fsm_output[5]);
  assign nor_831_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) | (COMP_LOOP_acc_1_cse_sva[1])
      | nand_170_cse);
  assign nor_832_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm)
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1949_nl = MUX_s_1_2_2(nor_831_nl, nor_832_nl, fsm_output[2]);
  assign nor_833_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b1101) | (~ (fsm_output[2]))
      | (fsm_output[7]) | not_tmp_395);
  assign mux_1950_nl = MUX_s_1_2_2(mux_1949_nl, nor_833_nl, fsm_output[5]);
  assign mux_1952_nl = MUX_s_1_2_2(mux_1951_nl, mux_1950_nl, fsm_output[1]);
  assign mux_1956_nl = MUX_s_1_2_2(mux_1955_nl, mux_1952_nl, fsm_output[0]);
  assign mux_1963_nl = MUX_s_1_2_2(mux_1962_nl, mux_1956_nl, fsm_output[4]);
  assign mux_1945_nl = MUX_s_1_2_2(nor_860_cse, and_490_cse, fsm_output[2]);
  assign nor_835_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b110) | (~ COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b100));
  assign nor_836_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]!=3'b110) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b010));
  assign mux_1944_nl = MUX_s_1_2_2(nor_835_nl, nor_836_nl, fsm_output[2]);
  assign and_491_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1944_nl;
  assign mux_1946_nl = MUX_s_1_2_2(mux_1945_nl, and_491_nl, fsm_output[5]);
  assign mux_1942_nl = MUX_s_1_2_2(nor_837_cse, nor_838_cse, fsm_output[2]);
  assign and_492_nl = nor_351_cse & mux_1941_cse;
  assign mux_1943_nl = MUX_s_1_2_2(mux_1942_nl, and_492_nl, fsm_output[5]);
  assign mux_1947_nl = MUX_s_1_2_2(mux_1946_nl, mux_1943_nl, fsm_output[1]);
  assign nor_840_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1101) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b100));
  assign nor_841_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1101) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[8:6]!=3'b010));
  assign mux_1937_nl = MUX_s_1_2_2(nor_840_nl, nor_841_nl, fsm_output[2]);
  assign nor_842_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b1101) | (fsm_output[8:6]!=3'b100));
  assign nor_843_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b1101) | (fsm_output[8:6]!=3'b010));
  assign mux_1936_nl = MUX_s_1_2_2(nor_842_nl, nor_843_nl, fsm_output[2]);
  assign mux_1938_nl = MUX_s_1_2_2(mux_1937_nl, mux_1936_nl, fsm_output[5]);
  assign and_495_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b1101) & COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm
      & (fsm_output[8:6]==3'b011);
  assign nor_844_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[8:6]!=3'b001));
  assign mux_1934_nl = MUX_s_1_2_2(and_495_nl, nor_844_nl, fsm_output[2]);
  assign and_496_nl = (COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]==4'b1101) & (fsm_output[8:6]==3'b011);
  assign nor_845_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b1101) | (fsm_output[8:6]!=3'b001));
  assign mux_1933_nl = MUX_s_1_2_2(and_496_nl, nor_845_nl, fsm_output[2]);
  assign mux_1935_nl = MUX_s_1_2_2(mux_1934_nl, mux_1933_nl, fsm_output[5]);
  assign mux_1939_nl = MUX_s_1_2_2(mux_1938_nl, mux_1935_nl, fsm_output[1]);
  assign mux_1948_nl = MUX_s_1_2_2(mux_1947_nl, mux_1939_nl, fsm_output[0]);
  assign and_489_nl = (fsm_output[4]) & mux_1948_nl;
  assign vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1963_nl,
      and_489_nl, fsm_output[3]);
  assign nor_792_nl = ~((~ (fsm_output[5])) | (~ (VEC_LOOP_j_10_0_sva_9_0[3])) |
      (fsm_output[0]) | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[1]) | (~ (VEC_LOOP_j_10_0_sva_9_0[1]))
      | (fsm_output[3:2]!=2'b00) | (~ (VEC_LOOP_j_10_0_sva_9_0[2])) | (fsm_output[8:6]!=3'b000));
  assign nand_79_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1]) & mux_1991_cse);
  assign nand_156_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]==3'b111) & (fsm_output[8:6]==3'b111));
  assign or_2109_nl = nand_157_cse | not_tmp_395;
  assign mux_1988_nl = MUX_s_1_2_2(nand_156_nl, or_2109_nl, fsm_output[2]);
  assign nand_158_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]==3'b111) & (fsm_output[8:6]==3'b011));
  assign or_2106_nl = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b111) | (fsm_output[8:6]!=3'b001);
  assign mux_1987_nl = MUX_s_1_2_2(nand_158_nl, or_2106_nl, fsm_output[2]);
  assign mux_1989_nl = MUX_s_1_2_2(mux_1988_nl, mux_1987_nl, fsm_output[3]);
  assign mux_1992_nl = MUX_s_1_2_2(nand_79_nl, mux_1989_nl, fsm_output[1]);
  assign nor_793_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1992_nl);
  assign nor_797_nl = ~((~ (COMP_LOOP_acc_10_cse_10_1_15_sva[2])) | (~ (COMP_LOOP_acc_10_cse_10_1_15_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_15_sva[0]) | nand_268_cse);
  assign nor_798_nl = ~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b1110) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1984_nl = MUX_s_1_2_2(nor_797_nl, nor_798_nl, fsm_output[2]);
  assign and_486_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]==4'b1110) & (fsm_output[8:6]==3'b011);
  assign nor_799_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b1110) | (fsm_output[8:6]!=3'b001));
  assign mux_1983_nl = MUX_s_1_2_2(and_486_nl, nor_799_nl, fsm_output[2]);
  assign mux_1985_nl = MUX_s_1_2_2(mux_1984_nl, mux_1983_nl, fsm_output[3]);
  assign and_839_nl = (COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]==4'b1110) & (fsm_output[8:6]==3'b110);
  assign nor_801_nl = ~((COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]!=4'b1110) | (fsm_output[8:6]!=3'b100));
  assign mux_1981_nl = MUX_s_1_2_2(and_839_nl, nor_801_nl, fsm_output[2]);
  assign nor_802_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b1110) | (fsm_output[8:6]!=3'b010));
  assign nor_803_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[3:0]!=4'b1110) | (fsm_output[8:6]!=3'b000));
  assign mux_1980_nl = MUX_s_1_2_2(nor_802_nl, nor_803_nl, fsm_output[2]);
  assign mux_1982_nl = MUX_s_1_2_2(mux_1981_nl, mux_1980_nl, fsm_output[3]);
  assign mux_1986_nl = MUX_s_1_2_2(mux_1985_nl, mux_1982_nl, fsm_output[1]);
  assign mux_1993_nl = MUX_s_1_2_2(nor_793_nl, mux_1986_nl, fsm_output[0]);
  assign nor_804_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[0]) | (~((COMP_LOOP_acc_10_cse_10_1_sva[3:1]==3'b111)
      & (fsm_output[8:6]==3'b111))));
  assign nor_805_nl = ~((COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b1110) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1976_nl = MUX_s_1_2_2(nor_804_nl, nor_805_nl, fsm_output[2]);
  assign and_487_nl = (COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]==4'b1110) & (fsm_output[8:6]==3'b011);
  assign nor_806_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b1110) | (fsm_output[8:6]!=3'b001));
  assign mux_1975_nl = MUX_s_1_2_2(and_487_nl, nor_806_nl, fsm_output[2]);
  assign mux_1977_nl = MUX_s_1_2_2(mux_1976_nl, mux_1975_nl, fsm_output[3]);
  assign and_847_nl = (COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]==4'b1110) & (fsm_output[8:6]==3'b110);
  assign nor_808_nl = ~((COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b1110) | (fsm_output[8:6]!=3'b100));
  assign mux_1973_nl = MUX_s_1_2_2(and_847_nl, nor_808_nl, fsm_output[2]);
  assign nor_809_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b1110) | (fsm_output[8:6]!=3'b010));
  assign nor_810_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b1110) | (fsm_output[8:6]!=3'b000));
  assign mux_1972_nl = MUX_s_1_2_2(nor_809_nl, nor_810_nl, fsm_output[2]);
  assign mux_1974_nl = MUX_s_1_2_2(mux_1973_nl, mux_1972_nl, fsm_output[3]);
  assign mux_1978_nl = MUX_s_1_2_2(mux_1977_nl, mux_1974_nl, fsm_output[1]);
  assign nor_811_nl = ~((~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1110))) | nand_324_cse);
  assign nor_812_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1110) | (fsm_output[7])
      | not_tmp_395);
  assign mux_1969_nl = MUX_s_1_2_2(nor_811_nl, nor_812_nl, fsm_output[2]);
  assign and_488_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b1110) & (fsm_output[8:6]==3'b011);
  assign nor_813_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1110) | (fsm_output[8:6]!=3'b001));
  assign mux_1968_nl = MUX_s_1_2_2(and_488_nl, nor_813_nl, fsm_output[2]);
  assign mux_1970_nl = MUX_s_1_2_2(mux_1969_nl, mux_1968_nl, fsm_output[3]);
  assign and_863_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1110) & (fsm_output[8:6]==3'b110);
  assign nor_815_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1110) | (fsm_output[8:6]!=3'b100));
  assign mux_1966_nl = MUX_s_1_2_2(and_863_nl, nor_815_nl, fsm_output[2]);
  assign nor_816_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1110) | (fsm_output[8:6]!=3'b010));
  assign nor_817_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1110) | (fsm_output[8:6]!=3'b000));
  assign mux_1965_nl = MUX_s_1_2_2(nor_816_nl, nor_817_nl, fsm_output[2]);
  assign mux_1967_nl = MUX_s_1_2_2(mux_1966_nl, mux_1965_nl, fsm_output[3]);
  assign mux_1971_nl = MUX_s_1_2_2(mux_1970_nl, mux_1967_nl, fsm_output[1]);
  assign mux_1979_nl = MUX_s_1_2_2(mux_1978_nl, mux_1971_nl, fsm_output[0]);
  assign mux_1994_nl = MUX_s_1_2_2(mux_1993_nl, mux_1979_nl, fsm_output[5]);
  assign vec_rsc_0_14_i_we_d_pff = MUX_s_1_2_2(nor_792_nl, mux_1994_nl, fsm_output[4]);
  assign nor_769_nl = ~((~((fsm_output[5]) & (fsm_output[2]) & (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      & (COMP_LOOP_acc_20_psp_sva[2:0]==3'b111) & COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm))
      | nand_301_cse);
  assign nor_770_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b111) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_771_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[0]) | (~((COMP_LOOP_acc_10_cse_10_1_sva[3:1]==3'b111)
      & (fsm_output[7]) & (fsm_output[4]) & (fsm_output[8]))));
  assign mux_2021_nl = MUX_s_1_2_2(nor_770_nl, nor_771_nl, fsm_output[2]);
  assign nor_772_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b1110) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_2022_nl = MUX_s_1_2_2(mux_2021_nl, nor_772_nl, fsm_output[5]);
  assign mux_2023_nl = MUX_s_1_2_2(nor_769_nl, mux_2022_nl, fsm_output[6]);
  assign nor_773_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b1110) | (fsm_output[7])
      | (fsm_output[4]) | (fsm_output[8]));
  assign nor_774_nl = ~((~((COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]==4'b1110))) | nand_301_cse);
  assign mux_2018_nl = MUX_s_1_2_2(nor_773_nl, nor_774_nl, fsm_output[2]);
  assign nor_775_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b1110) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_2019_nl = MUX_s_1_2_2(mux_2018_nl, nor_775_nl, fsm_output[5]);
  assign nor_776_nl = ~((~((VEC_LOOP_j_10_0_sva_9_0[1]) & (fsm_output[5]) & (fsm_output[2])
      & (COMP_LOOP_acc_19_psp_sva[1:0]==2'b11) & COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm
      & (~ (VEC_LOOP_j_10_0_sva_9_0[0])) & (~ (fsm_output[7])))) | not_tmp_399);
  assign mux_2020_nl = MUX_s_1_2_2(mux_2019_nl, nor_776_nl, fsm_output[6]);
  assign mux_2024_nl = MUX_s_1_2_2(mux_2023_nl, mux_2020_nl, fsm_output[1]);
  assign nor_777_nl = ~((~((fsm_output[2]) & (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1110)
      & COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm)) | nand_301_cse);
  assign nor_778_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1110)
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_779_nl = ~((~ (COMP_LOOP_acc_10_cse_10_1_15_sva[2])) | (~ (COMP_LOOP_acc_10_cse_10_1_15_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_15_sva[0]) | nand_265_cse);
  assign mux_2014_nl = MUX_s_1_2_2(nor_778_nl, nor_779_nl, fsm_output[2]);
  assign mux_2015_nl = MUX_s_1_2_2(nor_777_nl, mux_2014_nl, fsm_output[5]);
  assign nor_780_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b1110) | (fsm_output[5])
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_2016_nl = MUX_s_1_2_2(mux_2015_nl, nor_780_nl, fsm_output[6]);
  assign nor_781_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[1])) | (~ (VEC_LOOP_j_10_0_sva_9_0[3]))
      | (fsm_output[5]) | (fsm_output[2]) | (~ (VEC_LOOP_j_10_0_sva_9_0[2])) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[7]) | (fsm_output[4]) | (fsm_output[8]));
  assign nor_782_nl = ~((~(COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm & (COMP_LOOP_acc_1_cse_sva[3:0]==4'b1110)))
      | nand_301_cse);
  assign nor_783_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm)
      | (fsm_output[7]) | not_tmp_399);
  assign mux_2011_nl = MUX_s_1_2_2(nor_782_nl, nor_783_nl, fsm_output[2]);
  assign nor_784_nl = ~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]!=4'b1110) | (~ (fsm_output[2]))
      | (fsm_output[7]) | not_tmp_399);
  assign mux_2012_nl = MUX_s_1_2_2(mux_2011_nl, nor_784_nl, fsm_output[5]);
  assign mux_2013_nl = MUX_s_1_2_2(nor_781_nl, mux_2012_nl, fsm_output[6]);
  assign mux_2017_nl = MUX_s_1_2_2(mux_2016_nl, mux_2013_nl, fsm_output[1]);
  assign mux_2025_nl = MUX_s_1_2_2(mux_2024_nl, mux_2017_nl, fsm_output[0]);
  assign nor_785_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]!=3'b111) | (~ COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (fsm_output[7]) | not_tmp_399);
  assign and_480_nl = (COMP_LOOP_acc_14_psp_sva[2:0]==3'b111) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm
      & (~ (VEC_LOOP_j_10_0_sva_9_0[0])) & (fsm_output[7]) & (fsm_output[4]) & (~
      (fsm_output[8]));
  assign mux_2007_nl = MUX_s_1_2_2(nor_785_nl, and_480_nl, fsm_output[2]);
  assign and_479_nl = (fsm_output[5]) & mux_2007_nl;
  assign or_2136_nl = (COMP_LOOP_acc_10_cse_10_1_12_sva[3:0]!=4'b1110) | (fsm_output[7])
      | not_tmp_399;
  assign nand_149_nl = ~((COMP_LOOP_acc_10_cse_10_1_8_sva[3:0]==4'b1110) & (fsm_output[7])
      & (fsm_output[4]) & (~ (fsm_output[8])));
  assign mux_2006_nl = MUX_s_1_2_2(or_2136_nl, nand_149_nl, fsm_output[2]);
  assign nor_786_nl = ~((fsm_output[5]) | mux_2006_nl);
  assign mux_2008_nl = MUX_s_1_2_2(and_479_nl, nor_786_nl, fsm_output[6]);
  assign or_2132_nl = (COMP_LOOP_acc_10_cse_10_1_10_sva[3:0]!=4'b1110) | (fsm_output[7])
      | not_tmp_399;
  assign nand_150_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]==4'b1110) & (fsm_output[7])
      & (fsm_output[4]) & (~ (fsm_output[8])));
  assign mux_2004_nl = MUX_s_1_2_2(or_2132_nl, nand_150_nl, fsm_output[2]);
  assign nor_787_nl = ~((fsm_output[5]) | mux_2004_nl);
  assign and_481_nl = (VEC_LOOP_j_10_0_sva_9_0[1]) & (fsm_output[5]) & mux_1878_cse;
  assign mux_2005_nl = MUX_s_1_2_2(nor_787_nl, and_481_nl, fsm_output[6]);
  assign mux_2009_nl = MUX_s_1_2_2(mux_2008_nl, mux_2005_nl, fsm_output[1]);
  assign or_2126_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1110) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7]) | not_tmp_399;
  assign nand_151_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1110) & COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[7]) & (fsm_output[4]) & (~ (fsm_output[8])));
  assign mux_2000_nl = MUX_s_1_2_2(or_2126_nl, nand_151_nl, fsm_output[2]);
  assign or_2123_nl = (COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]!=4'b1110) | (fsm_output[7])
      | not_tmp_399;
  assign nand_152_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]==4'b1110) & (fsm_output[7])
      & (fsm_output[4]) & (~ (fsm_output[8])));
  assign mux_1999_nl = MUX_s_1_2_2(or_2123_nl, nand_152_nl, fsm_output[2]);
  assign mux_2001_nl = MUX_s_1_2_2(mux_2000_nl, mux_1999_nl, fsm_output[5]);
  assign nor_789_nl = ~((fsm_output[6]) | mux_2001_nl);
  assign and_484_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b1110) & COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm
      & (fsm_output[7]) & (fsm_output[4]) & (~ (fsm_output[8]));
  assign nor_790_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7]) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_1997_nl = MUX_s_1_2_2(and_484_nl, nor_790_nl, fsm_output[2]);
  assign and_485_nl = (COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]==4'b1110) & (fsm_output[7])
      & (fsm_output[4]) & (~ (fsm_output[8]));
  assign nor_791_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b1110) | (fsm_output[7])
      | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_1996_nl = MUX_s_1_2_2(and_485_nl, nor_791_nl, fsm_output[2]);
  assign mux_1998_nl = MUX_s_1_2_2(mux_1997_nl, mux_1996_nl, fsm_output[5]);
  assign and_483_nl = (fsm_output[6]) & mux_1998_nl;
  assign mux_2002_nl = MUX_s_1_2_2(nor_789_nl, and_483_nl, fsm_output[1]);
  assign mux_2010_nl = MUX_s_1_2_2(mux_2009_nl, mux_2002_nl, fsm_output[0]);
  assign vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_2025_nl,
      mux_2010_nl, fsm_output[3]);
  assign nor_751_nl = ~((~ (fsm_output[5])) | (~ (VEC_LOOP_j_10_0_sva_9_0[3])) |
      (fsm_output[0]) | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (fsm_output[1]) | (~ (VEC_LOOP_j_10_0_sva_9_0[1]))
      | (fsm_output[3:2]!=2'b00) | (~ (VEC_LOOP_j_10_0_sva_9_0[2])) | (fsm_output[8:6]!=3'b000));
  assign and_464_nl = (VEC_LOOP_j_10_0_sva_9_0[1]) & mux_1991_cse;
  assign and_465_nl = (COMP_LOOP_acc_20_psp_sva[2:0]==3'b111) & (fsm_output[8:6]==3'b111);
  assign nor_755_nl = ~(nand_157_cse | not_tmp_395);
  assign mux_2050_nl = MUX_s_1_2_2(and_465_nl, nor_755_nl, fsm_output[2]);
  assign and_466_nl = (COMP_LOOP_acc_14_psp_sva[2:0]==3'b111) & (fsm_output[8:6]==3'b011);
  assign nor_756_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b111) | (fsm_output[8:6]!=3'b001));
  assign mux_2049_nl = MUX_s_1_2_2(and_466_nl, nor_756_nl, fsm_output[2]);
  assign mux_2051_nl = MUX_s_1_2_2(mux_2050_nl, mux_2049_nl, fsm_output[3]);
  assign mux_2054_nl = MUX_s_1_2_2(and_464_nl, mux_2051_nl, fsm_output[1]);
  assign and_463_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_2054_nl;
  assign and_467_nl = (COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b111);
  assign nor_757_nl = ~((~((COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]==4'b1111) & (~
      (fsm_output[7])))) | not_tmp_395);
  assign mux_2046_nl = MUX_s_1_2_2(and_467_nl, nor_757_nl, fsm_output[2]);
  assign and_468_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b011);
  assign and_469_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b001);
  assign mux_2045_nl = MUX_s_1_2_2(and_468_nl, and_469_nl, fsm_output[2]);
  assign mux_2047_nl = MUX_s_1_2_2(mux_2046_nl, mux_2045_nl, fsm_output[3]);
  assign and_838_nl = (COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b110);
  assign and_844_nl = (COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b100);
  assign mux_2043_nl = MUX_s_1_2_2(and_838_nl, and_844_nl, fsm_output[2]);
  assign and_470_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b010);
  assign nor_760_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[3:0]!=4'b1111) | (fsm_output[8:6]!=3'b000));
  assign mux_2042_nl = MUX_s_1_2_2(and_470_nl, nor_760_nl, fsm_output[2]);
  assign mux_2044_nl = MUX_s_1_2_2(mux_2043_nl, mux_2042_nl, fsm_output[3]);
  assign mux_2048_nl = MUX_s_1_2_2(mux_2047_nl, mux_2044_nl, fsm_output[1]);
  assign mux_2055_nl = MUX_s_1_2_2(and_463_nl, mux_2048_nl, fsm_output[0]);
  assign and_471_nl = (COMP_LOOP_acc_10_cse_10_1_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b111);
  assign mux_2038_nl = MUX_s_1_2_2(and_471_nl, nor_761_cse, fsm_output[2]);
  assign and_473_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b001);
  assign mux_2037_nl = MUX_s_1_2_2(and_450_cse, and_473_nl, fsm_output[2]);
  assign mux_2039_nl = MUX_s_1_2_2(mux_2038_nl, mux_2037_nl, fsm_output[3]);
  assign and_846_nl = (COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b110);
  assign mux_2035_nl = MUX_s_1_2_2(and_846_nl, and_836_cse, fsm_output[2]);
  assign nor_764_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b1111) | (fsm_output[8:6]!=3'b000));
  assign mux_2034_nl = MUX_s_1_2_2(and_453_cse, nor_764_nl, fsm_output[2]);
  assign mux_2036_nl = MUX_s_1_2_2(mux_2035_nl, mux_2034_nl, fsm_output[3]);
  assign mux_2040_nl = MUX_s_1_2_2(mux_2039_nl, mux_2036_nl, fsm_output[1]);
  assign and_475_nl = (COMP_LOOP_acc_1_cse_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b111);
  assign nor_765_nl = ~((~((COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b1111) & (~ (fsm_output[7]))))
      | not_tmp_395);
  assign mux_2031_nl = MUX_s_1_2_2(and_475_nl, nor_765_nl, fsm_output[2]);
  assign and_476_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b011);
  assign and_477_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b001);
  assign mux_2030_nl = MUX_s_1_2_2(and_476_nl, and_477_nl, fsm_output[2]);
  assign mux_2032_nl = MUX_s_1_2_2(mux_2031_nl, mux_2030_nl, fsm_output[3]);
  assign and_861_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b110);
  assign and_862_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b100);
  assign mux_2028_nl = MUX_s_1_2_2(and_861_nl, and_862_nl, fsm_output[2]);
  assign and_478_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b010);
  assign nor_768_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1111) | (fsm_output[8:6]!=3'b000));
  assign mux_2027_nl = MUX_s_1_2_2(and_478_nl, nor_768_nl, fsm_output[2]);
  assign mux_2029_nl = MUX_s_1_2_2(mux_2028_nl, mux_2027_nl, fsm_output[3]);
  assign mux_2033_nl = MUX_s_1_2_2(mux_2032_nl, mux_2029_nl, fsm_output[1]);
  assign mux_2041_nl = MUX_s_1_2_2(mux_2040_nl, mux_2033_nl, fsm_output[0]);
  assign mux_2056_nl = MUX_s_1_2_2(mux_2055_nl, mux_2041_nl, fsm_output[5]);
  assign vec_rsc_0_15_i_we_d_pff = MUX_s_1_2_2(nor_751_nl, mux_2056_nl, fsm_output[4]);
  assign nor_731_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b111)
      | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) | (fsm_output[2]) | (fsm_output[7])
      | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_732_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[3:0]!=4'b1111) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_2085_nl = MUX_s_1_2_2(nor_731_nl, nor_732_nl, fsm_output[5]);
  assign nor_733_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b1111) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign nor_734_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[3:0]!=4'b1111) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_2084_nl = MUX_s_1_2_2(nor_733_nl, nor_734_nl, fsm_output[5]);
  assign mux_2086_nl = MUX_s_1_2_2(mux_2085_nl, mux_2084_nl, fsm_output[1]);
  assign nor_735_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[3:0]!=4'b1111) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_736_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1111)
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_2082_nl = MUX_s_1_2_2(nor_735_nl, nor_736_nl, fsm_output[5]);
  assign nor_737_nl = ~((~ (VEC_LOOP_j_10_0_sva_9_0[3])) | (fsm_output[5]) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_2083_nl = MUX_s_1_2_2(mux_2082_nl, nor_737_nl, fsm_output[1]);
  assign mux_2087_nl = MUX_s_1_2_2(mux_2086_nl, mux_2083_nl, fsm_output[0]);
  assign and_447_nl = (COMP_LOOP_acc_10_cse_10_1_sva[3:0]==4'b1111) & (fsm_output[2])
      & (fsm_output[7]) & (fsm_output[6]) & (fsm_output[8]);
  assign and_845_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (fsm_output[2]) & (COMP_LOOP_acc_20_psp_sva[2:0]==3'b111)
      & COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm & (fsm_output[8:6]==3'b110);
  assign mux_2079_nl = MUX_s_1_2_2(and_447_nl, and_845_nl, fsm_output[5]);
  assign and_854_nl = (COMP_LOOP_acc_10_cse_10_1_14_sva[3:0]==4'b1111) & (fsm_output[2])
      & (fsm_output[7]) & (~ (fsm_output[6])) & (fsm_output[8]);
  assign nor_740_nl = ~((~((VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & (fsm_output[2])
      & (COMP_LOOP_acc_19_psp_sva[1:0]==2'b11) & COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm
      & (~ (fsm_output[7])))) | not_tmp_395);
  assign mux_2078_nl = MUX_s_1_2_2(and_854_nl, nor_740_nl, fsm_output[5]);
  assign mux_2080_nl = MUX_s_1_2_2(mux_2079_nl, mux_2078_nl, fsm_output[1]);
  assign and_859_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1111) & COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[2]) & (fsm_output[7]) & (~ (fsm_output[6])) & (fsm_output[8]);
  assign and_860_nl = (COMP_LOOP_acc_10_cse_10_1_15_sva[3:0]==4'b1111) & (fsm_output[2])
      & (fsm_output[7]) & (~ (fsm_output[6])) & (fsm_output[8]);
  assign mux_2076_nl = MUX_s_1_2_2(and_859_nl, and_860_nl, fsm_output[5]);
  assign and_448_nl = COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm & (COMP_LOOP_acc_1_cse_sva[3:0]==4'b1111)
      & (fsm_output[8:6]==3'b111);
  assign nor_743_nl = ~((~((COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b1111) & COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm
      & (~ (fsm_output[7])))) | not_tmp_395);
  assign mux_2074_nl = MUX_s_1_2_2(and_448_nl, nor_743_nl, fsm_output[2]);
  assign nor_744_nl = ~((~((COMP_LOOP_acc_10_cse_10_1_13_sva[3:0]==4'b1111) & (fsm_output[2])
      & (~ (fsm_output[7])))) | not_tmp_395);
  assign mux_2075_nl = MUX_s_1_2_2(mux_2074_nl, nor_744_nl, fsm_output[5]);
  assign mux_2077_nl = MUX_s_1_2_2(mux_2076_nl, mux_2075_nl, fsm_output[1]);
  assign mux_2081_nl = MUX_s_1_2_2(mux_2080_nl, mux_2077_nl, fsm_output[0]);
  assign mux_2088_nl = MUX_s_1_2_2(mux_2087_nl, mux_2081_nl, fsm_output[4]);
  assign mux_2070_nl = MUX_s_1_2_2(nor_761_cse, and_450_cse, fsm_output[2]);
  assign and_833_nl = (COMP_LOOP_acc_17_psp_sva[2:0]==3'b111) & COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[8:6]==3'b100);
  assign and_452_nl = (COMP_LOOP_acc_14_psp_sva[2:0]==3'b111) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[8:6]==3'b010);
  assign mux_2069_nl = MUX_s_1_2_2(and_833_nl, and_452_nl, fsm_output[2]);
  assign and_451_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_2069_nl;
  assign mux_2071_nl = MUX_s_1_2_2(mux_2070_nl, and_451_nl, fsm_output[5]);
  assign mux_2067_nl = MUX_s_1_2_2(and_836_cse, and_453_cse, fsm_output[2]);
  assign and_454_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & mux_1941_cse;
  assign mux_2068_nl = MUX_s_1_2_2(mux_2067_nl, and_454_nl, fsm_output[5]);
  assign mux_2072_nl = MUX_s_1_2_2(mux_2071_nl, mux_2068_nl, fsm_output[1]);
  assign and_837_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]==4'b1111) & COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[8:6]==3'b100);
  assign and_457_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1111) & COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[8:6]==3'b010);
  assign mux_2062_nl = MUX_s_1_2_2(and_837_nl, and_457_nl, fsm_output[2]);
  assign and_843_nl = (COMP_LOOP_acc_10_cse_10_1_11_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b100);
  assign and_458_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b010);
  assign mux_2061_nl = MUX_s_1_2_2(and_843_nl, and_458_nl, fsm_output[2]);
  assign mux_2063_nl = MUX_s_1_2_2(mux_2062_nl, mux_2061_nl, fsm_output[5]);
  assign and_459_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b1111) & COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm
      & (fsm_output[8:6]==3'b011);
  assign and_460_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]==4'b1111) & COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm
      & (fsm_output[8:6]==3'b001);
  assign mux_2059_nl = MUX_s_1_2_2(and_459_nl, and_460_nl, fsm_output[2]);
  assign and_461_nl = (COMP_LOOP_acc_10_cse_10_1_9_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b011);
  assign and_462_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]==4'b1111) & (fsm_output[8:6]==3'b001);
  assign mux_2058_nl = MUX_s_1_2_2(and_461_nl, and_462_nl, fsm_output[2]);
  assign mux_2060_nl = MUX_s_1_2_2(mux_2059_nl, mux_2058_nl, fsm_output[5]);
  assign mux_2064_nl = MUX_s_1_2_2(mux_2063_nl, mux_2060_nl, fsm_output[1]);
  assign mux_2073_nl = MUX_s_1_2_2(mux_2072_nl, mux_2064_nl, fsm_output[0]);
  assign and_449_nl = (fsm_output[4]) & mux_2073_nl;
  assign vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_2088_nl,
      and_449_nl, fsm_output[3]);
  assign nl_COMP_LOOP_1_tmp_mul_nl = COMP_LOOP_1_tmp_lshift_itm * COMP_LOOP_k_10_4_sva_5_0;
  assign COMP_LOOP_1_tmp_mul_nl = nl_COMP_LOOP_1_tmp_mul_nl[5:0];
  assign twiddle_rsc_0_0_i_radr_d = MUX1HOT_v_6_6_2(COMP_LOOP_1_tmp_mul_nl, (COMP_LOOP_10_tmp_mul_idiv_sva[9:4]),
      (COMP_LOOP_11_tmp_mul_idiv_sva[8:3]), (COMP_LOOP_5_tmp_mul_idiv_sva[7:2]),
      (COMP_LOOP_9_tmp_lshift_itm[6:1]), (COMP_LOOP_13_tmp_mul_idiv_sva[7:2]), {and_dcpl_62
      , and_dcpl_175 , and_dcpl_180 , and_dcpl_181 , and_dcpl_183 , and_dcpl_184});
  assign mux_2095_nl = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), or_2259_cse_1);
  assign or_2260_nl = (COMP_LOOP_11_tmp_mul_idiv_sva[2:0]!=3'b000) | mux_2095_nl;
  assign or_2257_nl = (~ (fsm_output[4])) | (COMP_LOOP_10_tmp_mul_idiv_sva[3:0]!=4'b0000);
  assign mux_2094_nl = MUX_s_1_2_2(or_2257_nl, or_tmp_2077, or_2259_cse_1);
  assign mux_2096_nl = MUX_s_1_2_2(or_2260_nl, mux_2094_nl, fsm_output[0]);
  assign or_2255_nl = (COMP_LOOP_5_tmp_mul_idiv_sva[1:0]!=2'b00) | (fsm_output[4]);
  assign mux_2091_nl = MUX_s_1_2_2((fsm_output[4]), or_2255_nl, fsm_output[2]);
  assign or_2254_nl = (COMP_LOOP_9_tmp_lshift_itm[0]) | (fsm_output[4]);
  assign or_2253_nl = (COMP_LOOP_13_tmp_mul_idiv_sva[1:0]!=2'b00) | (fsm_output[4]);
  assign mux_2090_nl = MUX_s_1_2_2(or_2254_nl, or_2253_nl, fsm_output[2]);
  assign mux_2092_nl = MUX_s_1_2_2(mux_2091_nl, mux_2090_nl, fsm_output[3]);
  assign mux_2093_nl = MUX_s_1_2_2(mux_2092_nl, or_tmp_2077, fsm_output[0]);
  assign mux_2097_nl = MUX_s_1_2_2(mux_2096_nl, mux_2093_nl, fsm_output[1]);
  assign twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2097_nl) &
      and_dcpl_186;
  assign twiddle_rsc_0_1_i_radr_d_pff = z_out_3[9:4];
  assign nor_724_cse = ~((z_out_3[3:0]!=4'b0001) | (fsm_output[4]));
  assign nor_723_nl = ~((z_out_3[3:1]!=3'b000) | nand_122_cse);
  assign mux_2102_nl = MUX_s_1_2_2(nor_723_nl, nor_724_cse, fsm_output[1]);
  assign mux_2103_nl = MUX_s_1_2_2(mux_2102_nl, nor_724_cse, fsm_output[2]);
  assign mux_2104_nl = MUX_s_1_2_2(mux_2103_nl, nor_724_cse, fsm_output[3]);
  assign twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2104_nl & and_dcpl_193;
  assign twiddle_rsc_0_2_i_radr_d_pff = MUX_v_6_2_2((z_out_3[9:4]), (z_out_3[8:3]),
      COMP_LOOP_tmp_or_19_cse);
  assign nor_712_cse = ~((z_out_3[3:0]!=4'b0010) | (fsm_output[4]));
  assign nor_711_nl = ~((z_out_3[3:0]!=4'b0010) | (~ (fsm_output[4])));
  assign mux_2112_nl = MUX_s_1_2_2(nor_711_nl, nor_712_cse, fsm_output[2]);
  assign mux_2113_nl = MUX_s_1_2_2(mux_2112_nl, nor_712_cse, fsm_output[1]);
  assign mux_2114_nl = MUX_s_1_2_2(mux_2113_nl, nor_712_cse, fsm_output[3]);
  assign and_445_nl = (fsm_output[1]) & (~((z_out_3[2:0]!=3'b001) | (fsm_output[4])));
  assign mux_2115_nl = MUX_s_1_2_2(mux_2114_nl, and_445_nl, fsm_output[0]);
  assign twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2115_nl & and_dcpl_186;
  assign nor_704_cse = ~((z_out_3[3:0]!=4'b0011) | (fsm_output[4]));
  assign nor_703_nl = ~((z_out_3[3:2]!=2'b00) | nand_121_cse);
  assign mux_2120_nl = MUX_s_1_2_2(nor_703_nl, nor_704_cse, fsm_output[1]);
  assign mux_2121_nl = MUX_s_1_2_2(mux_2120_nl, nor_704_cse, fsm_output[2]);
  assign mux_2122_nl = MUX_s_1_2_2(mux_2121_nl, nor_704_cse, fsm_output[3]);
  assign twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2122_nl & and_dcpl_193;
  assign COMP_LOOP_tmp_or_46_cse = (and_dcpl_188 & and_dcpl_64) | and_dcpl_202;
  assign twiddle_rsc_0_4_i_radr_d_pff = MUX1HOT_v_6_3_2((z_out_3[9:4]), (z_out_3[8:3]),
      (z_out_3[7:2]), {COMP_LOOP_tmp_or_1_cse , COMP_LOOP_tmp_or_19_cse , COMP_LOOP_tmp_or_46_cse});
  assign nor_691_cse = ~((z_out_3[3:0]!=4'b0100) | (fsm_output[4]));
  assign nor_692_nl = ~((z_out_3[2:0]!=3'b010) | (fsm_output[4]));
  assign mux_2131_cse = MUX_s_1_2_2(nor_691_cse, nor_692_nl, fsm_output[0]);
  assign nor_689_nl = ~((z_out_3[3:0]!=4'b0100) | (fsm_output[0]) | (~ (fsm_output[4])));
  assign nor_690_nl = ~((fsm_output[0]) | (z_out_3[3:0]!=4'b0100) | (fsm_output[4]));
  assign mux_2133_nl = MUX_s_1_2_2(nor_689_nl, nor_690_nl, fsm_output[3]);
  assign mux_2134_nl = MUX_s_1_2_2(mux_2133_nl, mux_2131_cse, fsm_output[1]);
  assign nor_696_nl = ~((z_out_3[1:0]!=2'b01) | (fsm_output[4]));
  assign mux_2127_nl = MUX_s_1_2_2(nor_691_cse, nor_696_nl, fsm_output[0]);
  assign mux_2129_nl = MUX_s_1_2_2(mux_2127_nl, mux_2131_cse, fsm_output[1]);
  assign mux_2135_nl = MUX_s_1_2_2(mux_2134_nl, mux_2129_nl, fsm_output[2]);
  assign twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2135_nl & and_dcpl_186;
  assign nor_682_cse = ~((z_out_3[3:0]!=4'b0101) | (fsm_output[4]));
  assign nor_681_nl = ~((z_out_3[3:1]!=3'b010) | nand_122_cse);
  assign mux_2140_nl = MUX_s_1_2_2(nor_681_nl, nor_682_cse, fsm_output[1]);
  assign mux_2141_nl = MUX_s_1_2_2(mux_2140_nl, nor_682_cse, fsm_output[2]);
  assign mux_2142_nl = MUX_s_1_2_2(mux_2141_nl, nor_682_cse, fsm_output[3]);
  assign twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2142_nl & and_dcpl_193;
  assign nor_670_cse = ~((z_out_3[3:0]!=4'b0110) | (fsm_output[4]));
  assign nor_669_nl = ~((z_out_3[3:0]!=4'b0110) | (~ (fsm_output[4])));
  assign mux_2150_nl = MUX_s_1_2_2(nor_669_nl, nor_670_cse, fsm_output[2]);
  assign mux_2151_nl = MUX_s_1_2_2(mux_2150_nl, nor_670_cse, fsm_output[1]);
  assign mux_2152_nl = MUX_s_1_2_2(mux_2151_nl, nor_670_cse, fsm_output[3]);
  assign and_443_nl = (fsm_output[1]) & (~((z_out_3[2:0]!=3'b011) | (fsm_output[4])));
  assign mux_2153_nl = MUX_s_1_2_2(mux_2152_nl, and_443_nl, fsm_output[0]);
  assign twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2153_nl & and_dcpl_186;
  assign nor_662_cse = ~((z_out_3[3:0]!=4'b0111) | (fsm_output[4]));
  assign nor_661_nl = ~((z_out_3[3]) | (~((z_out_3[2:0]==3'b111) & (fsm_output[4]))));
  assign mux_2158_nl = MUX_s_1_2_2(nor_661_nl, nor_662_cse, fsm_output[1]);
  assign mux_2159_nl = MUX_s_1_2_2(mux_2158_nl, nor_662_cse, fsm_output[2]);
  assign mux_2160_nl = MUX_s_1_2_2(mux_2159_nl, nor_662_cse, fsm_output[3]);
  assign twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2160_nl & and_dcpl_193;
  assign twiddle_rsc_0_8_i_radr_d = MUX1HOT_v_6_4_2((z_out_3[9:4]), (z_out_3[8:3]),
      (z_out_3[7:2]), (z_out_3[6:1]), {COMP_LOOP_tmp_or_1_cse , COMP_LOOP_tmp_or_19_cse
      , COMP_LOOP_tmp_or_46_cse , and_dcpl_207});
  assign nor_647_cse = ~((z_out_3[3:0]!=4'b1000) | (fsm_output[4]));
  assign nor_650_nl = ~((z_out_3[2:0]!=3'b100) | (fsm_output[4]));
  assign mux_2169_cse = MUX_s_1_2_2(nor_647_cse, nor_650_nl, fsm_output[0]);
  assign nor_646_nl = ~((z_out_3[3:0]!=4'b1000) | (fsm_output[0]) | (~ (fsm_output[4])));
  assign nor_648_nl = ~((~ (z_out_3[0])) | (fsm_output[4]));
  assign mux_2171_nl = MUX_s_1_2_2(nor_647_cse, nor_648_nl, fsm_output[0]);
  assign mux_2172_nl = MUX_s_1_2_2(nor_646_nl, mux_2171_nl, fsm_output[3]);
  assign mux_2173_nl = MUX_s_1_2_2(mux_2172_nl, mux_2169_cse, fsm_output[1]);
  assign nor_654_nl = ~((z_out_3[1:0]!=2'b10) | (fsm_output[4]));
  assign mux_2165_nl = MUX_s_1_2_2(nor_647_cse, nor_654_nl, fsm_output[0]);
  assign mux_2167_nl = MUX_s_1_2_2(mux_2165_nl, mux_2169_cse, fsm_output[1]);
  assign mux_2174_nl = MUX_s_1_2_2(mux_2173_nl, mux_2167_nl, fsm_output[2]);
  assign twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2174_nl & and_dcpl_186;
  assign nor_639_cse = ~((z_out_3[3:0]!=4'b1001) | (fsm_output[4]));
  assign nor_638_nl = ~((z_out_3[3:1]!=3'b100) | nand_122_cse);
  assign mux_2179_nl = MUX_s_1_2_2(nor_638_nl, nor_639_cse, fsm_output[1]);
  assign mux_2180_nl = MUX_s_1_2_2(mux_2179_nl, nor_639_cse, fsm_output[2]);
  assign mux_2181_nl = MUX_s_1_2_2(mux_2180_nl, nor_639_cse, fsm_output[3]);
  assign twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2181_nl & and_dcpl_193;
  assign nor_627_cse = ~((z_out_3[3:0]!=4'b1010) | (fsm_output[4]));
  assign nor_626_nl = ~((z_out_3[3:0]!=4'b1010) | (~ (fsm_output[4])));
  assign mux_2189_nl = MUX_s_1_2_2(nor_626_nl, nor_627_cse, fsm_output[2]);
  assign mux_2190_nl = MUX_s_1_2_2(mux_2189_nl, nor_627_cse, fsm_output[1]);
  assign mux_2191_nl = MUX_s_1_2_2(mux_2190_nl, nor_627_cse, fsm_output[3]);
  assign and_441_nl = (fsm_output[1]) & (~((z_out_3[2:0]!=3'b101) | (fsm_output[4])));
  assign mux_2192_nl = MUX_s_1_2_2(mux_2191_nl, and_441_nl, fsm_output[0]);
  assign twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2192_nl & and_dcpl_186;
  assign nor_619_cse = ~((z_out_3[3:0]!=4'b1011) | (fsm_output[4]));
  assign nor_618_nl = ~((z_out_3[3:2]!=2'b10) | nand_121_cse);
  assign mux_2197_nl = MUX_s_1_2_2(nor_618_nl, nor_619_cse, fsm_output[1]);
  assign mux_2198_nl = MUX_s_1_2_2(mux_2197_nl, nor_619_cse, fsm_output[2]);
  assign mux_2199_nl = MUX_s_1_2_2(mux_2198_nl, nor_619_cse, fsm_output[3]);
  assign twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2199_nl & and_dcpl_193;
  assign nor_606_cse = ~((z_out_3[3:0]!=4'b1100) | (fsm_output[4]));
  assign nor_607_nl = ~((z_out_3[2:0]!=3'b110) | (fsm_output[4]));
  assign mux_2208_cse = MUX_s_1_2_2(nor_606_cse, nor_607_nl, fsm_output[0]);
  assign nor_604_nl = ~((z_out_3[3:0]!=4'b1100) | (fsm_output[0]) | (~ (fsm_output[4])));
  assign nor_605_nl = ~((fsm_output[0]) | (z_out_3[3:0]!=4'b1100) | (fsm_output[4]));
  assign mux_2210_nl = MUX_s_1_2_2(nor_604_nl, nor_605_nl, fsm_output[3]);
  assign mux_2211_nl = MUX_s_1_2_2(mux_2210_nl, mux_2208_cse, fsm_output[1]);
  assign nor_611_nl = ~((z_out_3[1:0]!=2'b11) | (fsm_output[4]));
  assign mux_2204_nl = MUX_s_1_2_2(nor_606_cse, nor_611_nl, fsm_output[0]);
  assign mux_2206_nl = MUX_s_1_2_2(mux_2204_nl, mux_2208_cse, fsm_output[1]);
  assign mux_2212_nl = MUX_s_1_2_2(mux_2211_nl, mux_2206_nl, fsm_output[2]);
  assign twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2212_nl & and_dcpl_186;
  assign nor_597_cse = ~((z_out_3[3:0]!=4'b1101) | (fsm_output[4]));
  assign nor_596_nl = ~((z_out_3[3:1]!=3'b110) | nand_122_cse);
  assign mux_2217_nl = MUX_s_1_2_2(nor_596_nl, nor_597_cse, fsm_output[1]);
  assign mux_2218_nl = MUX_s_1_2_2(mux_2217_nl, nor_597_cse, fsm_output[2]);
  assign mux_2219_nl = MUX_s_1_2_2(mux_2218_nl, nor_597_cse, fsm_output[3]);
  assign twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2219_nl & and_dcpl_193;
  assign nor_589_cse = ~((z_out_3[3:0]!=4'b1110) | (fsm_output[4]));
  assign and_434_nl = (z_out_3[3:0]==4'b1110) & (fsm_output[4]);
  assign mux_2227_nl = MUX_s_1_2_2(and_434_nl, nor_589_cse, fsm_output[2]);
  assign mux_2228_nl = MUX_s_1_2_2(mux_2227_nl, nor_589_cse, fsm_output[1]);
  assign mux_2229_nl = MUX_s_1_2_2(mux_2228_nl, nor_589_cse, fsm_output[3]);
  assign and_435_nl = (fsm_output[1]) & (z_out_3[2:0]==3'b111) & (~ (fsm_output[4]));
  assign mux_2230_nl = MUX_s_1_2_2(mux_2229_nl, and_435_nl, fsm_output[0]);
  assign twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2230_nl & and_dcpl_186;
  assign and_427_cse = (z_out_3[3:0]==4'b1111) & (~ (fsm_output[4]));
  assign and_426_nl = (z_out_3[3:0]==4'b1111) & (fsm_output[4]);
  assign mux_2235_nl = MUX_s_1_2_2(and_426_nl, and_427_cse, fsm_output[1]);
  assign mux_2236_nl = MUX_s_1_2_2(mux_2235_nl, and_427_cse, fsm_output[2]);
  assign mux_2237_nl = MUX_s_1_2_2(mux_2236_nl, and_427_cse, fsm_output[3]);
  assign twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2237_nl & and_dcpl_193;
  assign and_dcpl_356 = (fsm_output[8:6]==3'b111) & nor_1624_cse & (fsm_output[1])
      & (fsm_output[0]) & (fsm_output[4]) & (fsm_output[5]);
  assign and_dcpl_360 = mux_2465_cse & nor_1624_cse & (fsm_output[0]) & (~ (fsm_output[5]));
  assign and_dcpl_362 = ~((fsm_output[1:0]!=2'b00));
  assign and_dcpl_366 = and_dcpl_5 & nor_1624_cse;
  assign and_dcpl_367 = and_dcpl_366 & and_dcpl_362 & (fsm_output[5:4]==2'b11);
  assign and_dcpl_370 = (fsm_output[1:0]==2'b11) & and_dcpl_45;
  assign and_dcpl_373 = nor_1630_cse & (fsm_output[6]) & and_570_cse;
  assign and_dcpl_374 = and_dcpl_373 & and_dcpl_370;
  assign and_dcpl_376 = (fsm_output[1:0]==2'b10);
  assign and_dcpl_377 = and_dcpl_376 & and_dcpl_66;
  assign and_dcpl_378 = and_dcpl_373 & and_dcpl_377;
  assign and_dcpl_380 = (fsm_output[1:0]==2'b01) & and_dcpl_45;
  assign and_dcpl_383 = and_dcpl_87 & (~ (fsm_output[6])) & and_570_cse;
  assign and_dcpl_384 = and_dcpl_383 & and_dcpl_380;
  assign and_dcpl_385 = and_dcpl_362 & and_dcpl_66;
  assign and_dcpl_386 = and_dcpl_383 & and_dcpl_385;
  assign and_dcpl_387 = (fsm_output[3:2]==2'b10);
  assign and_dcpl_389 = and_dcpl_87 & (fsm_output[6]) & and_dcpl_387;
  assign and_dcpl_390 = and_dcpl_389 & and_dcpl_370;
  assign and_dcpl_391 = and_dcpl_389 & and_dcpl_377;
  assign and_dcpl_394 = and_dcpl_103 & (~ (fsm_output[6])) & and_dcpl_387;
  assign and_dcpl_395 = and_dcpl_394 & and_dcpl_380;
  assign and_dcpl_396 = and_dcpl_394 & and_dcpl_385;
  assign and_dcpl_397 = (fsm_output[3:2]==2'b01);
  assign and_dcpl_399 = and_dcpl_103 & (fsm_output[6]) & and_dcpl_397;
  assign and_dcpl_400 = and_dcpl_399 & and_dcpl_370;
  assign and_dcpl_401 = and_dcpl_399 & and_dcpl_377;
  assign and_dcpl_404 = and_733_cse & (~ (fsm_output[6])) & and_dcpl_397;
  assign and_dcpl_405 = and_dcpl_404 & and_dcpl_380;
  assign and_dcpl_406 = and_dcpl_404 & and_dcpl_385;
  assign and_dcpl_409 = and_733_cse & (fsm_output[6]) & nor_1624_cse & and_dcpl_377;
  assign and_dcpl_410 = and_dcpl_376 & and_dcpl_45;
  assign and_dcpl_411 = and_dcpl_366 & and_dcpl_410;
  assign and_dcpl_412 = and_dcpl_5 & and_dcpl_387;
  assign and_dcpl_413 = and_dcpl_412 & and_dcpl_380;
  assign and_dcpl_414 = and_dcpl_362 & and_dcpl_45;
  assign and_dcpl_415 = and_dcpl_5 & and_dcpl_397;
  assign and_dcpl_416 = and_dcpl_415 & and_dcpl_414;
  assign and_dcpl_417 = and_dcpl_415 & and_dcpl_410;
  assign and_dcpl_418 = and_dcpl_412 & and_dcpl_414;
  assign and_dcpl_419 = and_dcpl_412 & and_dcpl_410;
  assign and_dcpl_420 = and_dcpl_5 & and_570_cse;
  assign and_dcpl_421 = and_dcpl_420 & and_dcpl_414;
  assign and_dcpl_422 = and_dcpl_420 & and_dcpl_410;
  assign and_dcpl_425 = and_dcpl_366 & and_dcpl_362 & (fsm_output[5:4]==2'b01);
  assign and_dcpl_426 = and_dcpl_366 & and_dcpl_370;
  assign and_dcpl_427 = and_dcpl_415 & and_dcpl_370;
  assign and_dcpl_428 = and_dcpl_412 & and_dcpl_370;
  assign and_dcpl_429 = and_dcpl_420 & and_dcpl_370;
  assign and_dcpl_430 = and_dcpl_420 & and_dcpl_380;
  assign and_dcpl_431 = and_dcpl_415 & and_dcpl_380;
  assign and_dcpl_447 = ~((fsm_output!=9'b000000010));
  assign and_dcpl_465 = nor_1630_cse & (fsm_output[6]) & nor_1624_cse;
  assign and_1025_cse = and_dcpl_465 & and_dcpl_376 & and_dcpl_45;
  assign and_dcpl_467 = (fsm_output[1:0]==2'b01);
  assign and_1028_cse = and_dcpl_465 & and_dcpl_467 & and_dcpl_66;
  assign and_dcpl_475 = and_1189_cse & and_dcpl_75;
  assign and_dcpl_477 = and_dcpl_88 & and_570_cse;
  assign and_1037_cse = and_dcpl_477 & and_dcpl_475;
  assign and_dcpl_480 = and_dcpl_376 & and_dcpl_53;
  assign and_1040_cse = and_dcpl_477 & and_dcpl_480;
  assign and_dcpl_482 = and_dcpl_467 & and_dcpl_75;
  assign and_dcpl_484 = and_dcpl_87 & (fsm_output[6]) & and_570_cse;
  assign and_1044_cse = and_dcpl_484 & and_dcpl_482;
  assign and_dcpl_486 = and_dcpl_362 & and_dcpl_53;
  assign and_1046_cse = and_dcpl_484 & and_dcpl_486;
  assign and_1051_cse = and_dcpl_394 & and_dcpl_475;
  assign and_1052_cse = and_dcpl_394 & and_dcpl_480;
  assign and_dcpl_495 = and_dcpl_103 & (fsm_output[6]) & and_dcpl_387;
  assign and_1055_cse = and_dcpl_495 & and_dcpl_482;
  assign and_1056_cse = and_dcpl_495 & and_dcpl_486;
  assign and_1060_cse = and_dcpl_404 & and_dcpl_475;
  assign and_1061_cse = and_dcpl_404 & and_dcpl_480;
  assign and_1064_cse = and_733_cse & (fsm_output[6]) & and_dcpl_397 & and_dcpl_482;
  assign and_dcpl_571 = and_dcpl_5 & and_dcpl_397 & and_dcpl_414;
  assign and_dcpl_577 = and_dcpl_5 & nor_1624_cse & and_1189_cse & and_dcpl_66;
  assign and_dcpl_589 = and_dcpl_88 & nor_1624_cse & and_dcpl_414;
  assign COMP_LOOP_or_17_ssc = and_dcpl_360 | and_dcpl_367 | and_dcpl_374 | and_dcpl_378
      | and_dcpl_384 | and_dcpl_386 | and_dcpl_390 | and_dcpl_391 | and_dcpl_395
      | and_dcpl_396 | and_dcpl_400 | and_dcpl_401 | and_dcpl_405 | and_dcpl_406
      | and_dcpl_409;
  assign or_tmp_2410 = (fsm_output[3]) | (fsm_output[0]) | (fsm_output[2]);
  assign COMP_LOOP_nor_itm = ~(and_dcpl_411 | and_dcpl_413 | and_dcpl_416 | and_dcpl_417
      | and_dcpl_418 | and_dcpl_419 | and_dcpl_421 | and_dcpl_422 | and_dcpl_425
      | and_dcpl_426 | and_dcpl_427 | and_dcpl_428 | and_dcpl_429 | and_dcpl_430
      | and_dcpl_431);
  assign COMP_LOOP_or_40_itm = and_dcpl_416 | and_dcpl_417 | and_dcpl_418 | and_dcpl_419
      | and_dcpl_421 | and_dcpl_422 | and_dcpl_425;
  assign COMP_LOOP_nor_621_itm = ~(and_dcpl_413 | and_dcpl_426 | and_dcpl_427 | and_dcpl_428
      | and_dcpl_429 | and_dcpl_430 | and_dcpl_431);
  assign COMP_LOOP_or_41_itm = and_dcpl_411 | and_dcpl_426;
  assign COMP_LOOP_or_43_itm = and_dcpl_427 | and_dcpl_428 | and_dcpl_429;
  assign COMP_LOOP_nor_622_itm = ~(and_dcpl_413 | and_dcpl_430 | and_dcpl_431);
  assign COMP_LOOP_or_47_itm = and_dcpl_430 | and_dcpl_431;
  assign COMP_LOOP_or_52_itm = and_dcpl_411 | and_dcpl_416 | and_dcpl_417 | and_dcpl_418
      | and_dcpl_419 | and_dcpl_421 | and_dcpl_422 | and_dcpl_425;
  assign COMP_LOOP_or_54_itm = and_dcpl_426 | and_dcpl_427 | and_dcpl_428 | and_dcpl_429;
  assign COMP_LOOP_or_18_itm = (nor_1630_cse & (~ (fsm_output[6])) & nor_1624_cse
      & and_1189_cse & and_dcpl_66) | and_1025_cse | and_1028_cse | (and_dcpl_88
      & nor_1624_cse & and_dcpl_362 & and_dcpl_45) | and_1037_cse | and_1040_cse
      | and_1044_cse | and_1046_cse | and_1051_cse | and_1052_cse | and_1055_cse
      | and_1056_cse | and_1060_cse | and_1061_cse | and_1064_cse;
  always @(posedge clk) begin
    if ( (and_dcpl_51 & and_dcpl_47) | STAGE_LOOP_i_3_0_sva_mx0c1 ) begin
      STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(4'b1010, z_out_4, STAGE_LOOP_i_3_0_sva_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(nor_1871_nl, and_1183_nl, fsm_output[5]) ) begin
      p_sva <= p_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_vec_rsc_triosy_0_15_obj_ld_cse <= 1'b0;
      reg_ensig_cgo_cse <= 1'b0;
    end
    else begin
      reg_vec_rsc_triosy_0_15_obj_ld_cse <= and_dcpl_58 & and_dcpl_46 & (fsm_output[5:4]==2'b11)
          & (~ STAGE_LOOP_acc_itm_4_1);
      reg_ensig_cgo_cse <= mux_2255_rmff;
    end
  end
  always @(posedge clk) begin
    tmp_33_sva_6 <= twiddle_rsc_0_6_i_q_d;
    tmp_33_sva_8 <= twiddle_rsc_0_8_i_q_d;
    tmp_33_sva_11 <= MUX_v_64_2_2(twiddle_rsc_0_11_i_q_d, twiddle_rsc_0_12_i_q_d,
        and_dcpl_180);
    tmp_33_sva_12 <= MUX_v_64_2_2(twiddle_rsc_0_12_i_q_d, twiddle_rsc_0_14_i_q_d,
        and_dcpl_180);
    tmp_33_sva_13 <= MUX_v_64_2_2(twiddle_rsc_0_13_i_q_d, tmp_33_sva_13_mx0w1, and_dcpl_192);
    tmp_33_sva_14 <= twiddle_rsc_0_14_i_q_d;
  end
  always @(posedge clk) begin
    if ( rst ) begin
      VEC_LOOP_j_10_0_sva_9_0 <= 10'b0000000000;
    end
    else if ( VEC_LOOP_j_10_0_sva_9_0_mx0c0 | (and_dcpl_128 & and_dcpl_118) ) begin
      VEC_LOOP_j_10_0_sva_9_0 <= MUX_v_10_2_2(10'b0000000000, (z_out_2[9:0]), VEC_LOOP_j_not_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(nor_1870_nl, and_nl, fsm_output[5]) ) begin
      STAGE_LOOP_lshift_psp_sva <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_2558_nl, mux_nl, fsm_output[4]) ) begin
      COMP_LOOP_k_10_4_sva_5_0 <= MUX_v_6_2_2(6'b000000, reg_COMP_LOOP_k_10_4_ftd,
          nand_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_1_sva <= 10'b0000000000;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_acc_10_cse_10_1_1_sva <= COMP_LOOP_1_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_acc_psp_sva <= nl_COMP_LOOP_acc_psp_sva[5:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm <= z_out_2[10];
    end
  end
  always @(posedge clk) begin
    if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_2_tmp_lshift_ncse_sva <= z_out_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_9_tmp_lshift_itm <= 7'b0000000;
    end
    else if ( and_dcpl_62 | and_dcpl_207 ) begin
      COMP_LOOP_9_tmp_lshift_itm <= MUX_v_7_2_2((z_out[6:0]), (z_out_3[6:0]), and_dcpl_207);
    end
  end
  always @(posedge clk) begin
    if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_1_tmp_acc_cse_sva <= z_out_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_244_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_62_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_185_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_64_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_65_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_66_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_6_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_68_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_69_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_70_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_10_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_72_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_12_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_13_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_14_itm <= 1'b0;
    end
    else if ( mux_2303_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_itm <= ~((VEC_LOOP_j_10_0_sva_9_0[3:0]!=4'b0000));
      COMP_LOOP_COMP_LOOP_and_244_itm <= (COMP_LOOP_acc_13_psp_sva_1[0]) & (VEC_LOOP_j_10_0_sva_9_0[0])
          & (~((COMP_LOOP_acc_13_psp_sva_1[1]) | (VEC_LOOP_j_10_0_sva_9_0[1])));
      COMP_LOOP_COMP_LOOP_and_62_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b0011);
      COMP_LOOP_COMP_LOOP_and_185_itm <= (COMP_LOOP_acc_1_cse_4_sva_1[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_64_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_65_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_66_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b0111);
      COMP_LOOP_COMP_LOOP_and_6_itm <= (VEC_LOOP_j_10_0_sva_9_0[3:0]==4'b0111);
      COMP_LOOP_COMP_LOOP_and_68_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_69_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_70_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_10_itm <= (VEC_LOOP_j_10_0_sva_9_0[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_72_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_12_itm <= (VEC_LOOP_j_10_0_sva_9_0[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_13_itm <= (VEC_LOOP_j_10_0_sva_9_0[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_14_itm <= (VEC_LOOP_j_10_0_sva_9_0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_13_psp_sva <= 8'b00000000;
    end
    else if ( mux_2309_nl | (fsm_output[8]) ) begin
      COMP_LOOP_acc_13_psp_sva <= COMP_LOOP_acc_13_psp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_4_sva <= 10'b0000000000;
    end
    else if ( ~((~ mux_2312_nl) & nor_1630_cse) ) begin
      COMP_LOOP_acc_1_cse_4_sva <= COMP_LOOP_acc_1_cse_4_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_2_sva <= 10'b0000000000;
    end
    else if ( ~(mux_2314_nl & and_dcpl_5) ) begin
      COMP_LOOP_acc_1_cse_2_sva <= COMP_LOOP_acc_1_cse_2_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_2_sva <= 10'b0000000000;
    end
    else if ( ~(mux_2315_nl & and_dcpl_5) ) begin
      COMP_LOOP_acc_10_cse_10_1_2_sva <= COMP_LOOP_2_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( ~((and_1189_cse | (fsm_output[2]) | or_dcpl_190) & and_dcpl_5) ) begin
      COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_3_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_5_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_248 ) begin
      COMP_LOOP_COMP_LOOP_nor_5_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_51_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_248 ) begin
      COMP_LOOP_nor_51_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_52_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_248 ) begin
      COMP_LOOP_nor_52_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[3]) | (COMP_LOOP_2_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_77_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_248 ) begin
      COMP_LOOP_COMP_LOOP_and_77_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_54_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_248 ) begin
      COMP_LOOP_nor_54_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[3]) | (COMP_LOOP_2_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_79_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_248 ) begin
      COMP_LOOP_COMP_LOOP_and_79_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_80_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_248 ) begin
      COMP_LOOP_COMP_LOOP_and_80_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_81_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_248 ) begin
      COMP_LOOP_COMP_LOOP_and_81_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_57_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_248 ) begin
      COMP_LOOP_nor_57_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_83_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_248 ) begin
      COMP_LOOP_COMP_LOOP_and_83_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_84_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_248 ) begin
      COMP_LOOP_COMP_LOOP_and_84_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_85_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_248 ) begin
      COMP_LOOP_COMP_LOOP_and_85_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_86_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_248 ) begin
      COMP_LOOP_COMP_LOOP_and_86_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_87_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_248 ) begin
      COMP_LOOP_COMP_LOOP_and_87_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_88_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_248 ) begin
      COMP_LOOP_COMP_LOOP_and_88_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_89_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_248 ) begin
      COMP_LOOP_COMP_LOOP_and_89_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_nor_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_tmp_nor_itm <= COMP_LOOP_tmp_nor_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_nor_1_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_tmp_nor_1_itm <= COMP_LOOP_tmp_nor_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_nor_3_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_tmp_nor_3_itm <= COMP_LOOP_tmp_nor_3_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_nor_6_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_tmp_nor_6_itm <= COMP_LOOP_tmp_nor_6_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_184 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_11_psp_sva <= 9'b000000000;
    end
    else if ( ~((~ mux_2317_nl) & nor_1630_cse) ) begin
      COMP_LOOP_acc_11_psp_sva <= nl_COMP_LOOP_acc_11_psp_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_3_sva <= 10'b0000000000;
    end
    else if ( ~((~ mux_2319_nl) & nor_1630_cse) ) begin
      COMP_LOOP_acc_10_cse_10_1_3_sva <= COMP_LOOP_3_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( ~(mux_2321_nl & nor_1630_cse) ) begin
      COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm <= readslicef_9_1_8(COMP_LOOP_acc_12_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_9_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_nor_9_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_91_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_nor_91_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_92_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_nor_92_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[3]) | (COMP_LOOP_3_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_3_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_137_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_137_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_94_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_nor_94_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[3]) | (COMP_LOOP_3_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_3_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_139_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_139_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_140_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_140_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_141_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_141_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_97_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_nor_97_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_143_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_143_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_144_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_144_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_145_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_145_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_146_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_146_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_147_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_147_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_148_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_148_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_149_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_149_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_4_sva <= 10'b0000000000;
    end
    else if ( ~((~ mux_2326_nl) & nor_1630_cse) ) begin
      COMP_LOOP_acc_10_cse_10_1_4_sva <= COMP_LOOP_4_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( ~((~ mux_2327_nl) & nor_1630_cse) ) begin
      COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_5_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_13_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_255 ) begin
      COMP_LOOP_COMP_LOOP_nor_13_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_131_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_255 ) begin
      COMP_LOOP_nor_131_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_132_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_255 ) begin
      COMP_LOOP_nor_132_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[3]) | (COMP_LOOP_4_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_4_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_197_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_255 ) begin
      COMP_LOOP_COMP_LOOP_and_197_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_134_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_255 ) begin
      COMP_LOOP_nor_134_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[3]) | (COMP_LOOP_4_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_4_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_199_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_255 ) begin
      COMP_LOOP_COMP_LOOP_and_199_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_200_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_255 ) begin
      COMP_LOOP_COMP_LOOP_and_200_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_201_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_255 ) begin
      COMP_LOOP_COMP_LOOP_and_201_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_137_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_255 ) begin
      COMP_LOOP_nor_137_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_203_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_255 ) begin
      COMP_LOOP_COMP_LOOP_and_203_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_204_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_255 ) begin
      COMP_LOOP_COMP_LOOP_and_204_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_205_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_255 ) begin
      COMP_LOOP_COMP_LOOP_and_205_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_206_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_255 ) begin
      COMP_LOOP_COMP_LOOP_and_206_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_207_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_255 ) begin
      COMP_LOOP_COMP_LOOP_and_207_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_208_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_255 ) begin
      COMP_LOOP_COMP_LOOP_and_208_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_209_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_255 ) begin
      COMP_LOOP_COMP_LOOP_and_209_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_5_sva <= 10'b0000000000;
    end
    else if ( mux_2332_nl | (fsm_output[8]) ) begin
      COMP_LOOP_acc_10_cse_10_1_5_sva <= COMP_LOOP_5_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( mux_2335_nl | (fsm_output[8]) ) begin
      COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_6_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_17_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_258 ) begin
      COMP_LOOP_COMP_LOOP_nor_17_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_171_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_258 ) begin
      COMP_LOOP_nor_171_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_172_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_258 ) begin
      COMP_LOOP_nor_172_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[3]) | (COMP_LOOP_5_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_257_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_258 ) begin
      COMP_LOOP_COMP_LOOP_and_257_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_174_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_258 ) begin
      COMP_LOOP_nor_174_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[3]) | (COMP_LOOP_5_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_259_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_258 ) begin
      COMP_LOOP_COMP_LOOP_and_259_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_260_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_258 ) begin
      COMP_LOOP_COMP_LOOP_and_260_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_261_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_258 ) begin
      COMP_LOOP_COMP_LOOP_and_261_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_177_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_258 ) begin
      COMP_LOOP_nor_177_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_263_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_258 ) begin
      COMP_LOOP_COMP_LOOP_and_263_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_264_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_258 ) begin
      COMP_LOOP_COMP_LOOP_and_264_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_265_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_258 ) begin
      COMP_LOOP_COMP_LOOP_and_265_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_266_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_258 ) begin
      COMP_LOOP_COMP_LOOP_and_266_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_267_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_258 ) begin
      COMP_LOOP_COMP_LOOP_and_267_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_268_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_258 ) begin
      COMP_LOOP_COMP_LOOP_and_268_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_269_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_258 ) begin
      COMP_LOOP_COMP_LOOP_and_269_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_6_sva <= 10'b0000000000;
    end
    else if ( mux_2338_nl | (fsm_output[8]) ) begin
      COMP_LOOP_acc_1_cse_6_sva <= nl_COMP_LOOP_acc_1_cse_6_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_6_sva <= 10'b0000000000;
    end
    else if ( mux_2340_nl | (fsm_output[8]) ) begin
      COMP_LOOP_acc_10_cse_10_1_6_sva <= COMP_LOOP_6_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( mux_2341_nl | (fsm_output[8]) ) begin
      COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_7_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_21_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_262 ) begin
      COMP_LOOP_COMP_LOOP_nor_21_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_211_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_262 ) begin
      COMP_LOOP_nor_211_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_212_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_262 ) begin
      COMP_LOOP_nor_212_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[3]) | (COMP_LOOP_6_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_317_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_262 ) begin
      COMP_LOOP_COMP_LOOP_and_317_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_214_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_262 ) begin
      COMP_LOOP_nor_214_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[3]) | (COMP_LOOP_6_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_319_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_262 ) begin
      COMP_LOOP_COMP_LOOP_and_319_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_320_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_262 ) begin
      COMP_LOOP_COMP_LOOP_and_320_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_321_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_262 ) begin
      COMP_LOOP_COMP_LOOP_and_321_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_217_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_262 ) begin
      COMP_LOOP_nor_217_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_323_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_262 ) begin
      COMP_LOOP_COMP_LOOP_and_323_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_324_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_262 ) begin
      COMP_LOOP_COMP_LOOP_and_324_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_325_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_262 ) begin
      COMP_LOOP_COMP_LOOP_and_325_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_326_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_262 ) begin
      COMP_LOOP_COMP_LOOP_and_326_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_327_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_262 ) begin
      COMP_LOOP_COMP_LOOP_and_327_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_328_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_262 ) begin
      COMP_LOOP_COMP_LOOP_and_328_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_329_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_262 ) begin
      COMP_LOOP_COMP_LOOP_and_329_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_14_psp_sva <= 9'b000000000;
    end
    else if ( mux_2346_nl | (fsm_output[8]) ) begin
      COMP_LOOP_acc_14_psp_sva <= nl_COMP_LOOP_acc_14_psp_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_7_sva <= 10'b0000000000;
    end
    else if ( mux_2349_nl | (fsm_output[8]) ) begin
      COMP_LOOP_acc_10_cse_10_1_7_sva <= COMP_LOOP_7_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( mux_2352_nl | (fsm_output[8]) ) begin
      COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm <= readslicef_8_1_7(COMP_LOOP_acc_15_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_25_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_266 ) begin
      COMP_LOOP_COMP_LOOP_nor_25_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_251_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_266 ) begin
      COMP_LOOP_nor_251_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_252_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_266 ) begin
      COMP_LOOP_nor_252_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[3]) | (COMP_LOOP_7_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_377_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_266 ) begin
      COMP_LOOP_COMP_LOOP_and_377_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_254_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_266 ) begin
      COMP_LOOP_nor_254_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[3]) | (COMP_LOOP_7_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_379_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_266 ) begin
      COMP_LOOP_COMP_LOOP_and_379_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_380_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_266 ) begin
      COMP_LOOP_COMP_LOOP_and_380_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_381_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_266 ) begin
      COMP_LOOP_COMP_LOOP_and_381_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_257_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_266 ) begin
      COMP_LOOP_nor_257_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_383_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_266 ) begin
      COMP_LOOP_COMP_LOOP_and_383_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_384_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_266 ) begin
      COMP_LOOP_COMP_LOOP_and_384_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_385_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_266 ) begin
      COMP_LOOP_COMP_LOOP_and_385_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_386_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_266 ) begin
      COMP_LOOP_COMP_LOOP_and_386_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_387_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_266 ) begin
      COMP_LOOP_COMP_LOOP_and_387_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_388_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_266 ) begin
      COMP_LOOP_COMP_LOOP_and_388_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_389_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_266 ) begin
      COMP_LOOP_COMP_LOOP_and_389_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_8_sva <= 10'b0000000000;
    end
    else if ( mux_2354_nl | (fsm_output[8]) ) begin
      COMP_LOOP_acc_1_cse_8_sva <= nl_COMP_LOOP_acc_1_cse_8_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_8_sva <= 10'b0000000000;
    end
    else if ( mux_2355_nl | (fsm_output[8]) ) begin
      COMP_LOOP_acc_10_cse_10_1_8_sva <= COMP_LOOP_8_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( mux_2356_nl | (fsm_output[8]) ) begin
      COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_9_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_29_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_270 ) begin
      COMP_LOOP_COMP_LOOP_nor_29_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_291_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_270 ) begin
      COMP_LOOP_nor_291_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_292_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_270 ) begin
      COMP_LOOP_nor_292_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[3]) | (COMP_LOOP_8_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_437_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_270 ) begin
      COMP_LOOP_COMP_LOOP_and_437_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_294_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_270 ) begin
      COMP_LOOP_nor_294_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[3]) | (COMP_LOOP_8_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_439_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_270 ) begin
      COMP_LOOP_COMP_LOOP_and_439_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_440_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_270 ) begin
      COMP_LOOP_COMP_LOOP_and_440_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_441_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_270 ) begin
      COMP_LOOP_COMP_LOOP_and_441_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_297_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_270 ) begin
      COMP_LOOP_nor_297_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_443_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_270 ) begin
      COMP_LOOP_COMP_LOOP_and_443_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_444_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_270 ) begin
      COMP_LOOP_COMP_LOOP_and_444_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_445_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_270 ) begin
      COMP_LOOP_COMP_LOOP_and_445_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_446_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_270 ) begin
      COMP_LOOP_COMP_LOOP_and_446_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_447_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_270 ) begin
      COMP_LOOP_COMP_LOOP_and_447_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_448_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_270 ) begin
      COMP_LOOP_COMP_LOOP_and_448_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_449_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_270 ) begin
      COMP_LOOP_COMP_LOOP_and_449_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_16_psp_sva <= 7'b0000000;
    end
    else if ( MUX_s_1_2_2(mux_2364_nl, (fsm_output[8]), fsm_output[5]) ) begin
      COMP_LOOP_acc_16_psp_sva <= nl_COMP_LOOP_acc_16_psp_sva[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_9_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_2368_nl, (fsm_output[8]), fsm_output[5]) ) begin
      COMP_LOOP_acc_10_cse_10_1_9_sva <= COMP_LOOP_9_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_2372_nl, (fsm_output[8]), fsm_output[5]) ) begin
      COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_10_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_33_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_271 ) begin
      COMP_LOOP_COMP_LOOP_nor_33_itm <= ~((COMP_LOOP_9_acc_10_itm_10_1_1[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_331_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_271 ) begin
      COMP_LOOP_nor_331_itm <= ~((COMP_LOOP_9_acc_10_itm_10_1_1[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_332_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_271 ) begin
      COMP_LOOP_nor_332_itm <= ~((COMP_LOOP_9_acc_10_itm_10_1_1[3]) | (COMP_LOOP_9_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_9_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_497_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_271 ) begin
      COMP_LOOP_COMP_LOOP_and_497_itm <= (COMP_LOOP_9_acc_10_itm_10_1_1[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_334_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_271 ) begin
      COMP_LOOP_nor_334_itm <= ~((COMP_LOOP_9_acc_10_itm_10_1_1[3]) | (COMP_LOOP_9_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_9_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_499_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_271 ) begin
      COMP_LOOP_COMP_LOOP_and_499_itm <= (COMP_LOOP_9_acc_10_itm_10_1_1[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_500_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_271 ) begin
      COMP_LOOP_COMP_LOOP_and_500_itm <= (COMP_LOOP_9_acc_10_itm_10_1_1[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_501_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_271 ) begin
      COMP_LOOP_COMP_LOOP_and_501_itm <= (COMP_LOOP_9_acc_10_itm_10_1_1[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_337_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_271 ) begin
      COMP_LOOP_nor_337_itm <= ~((COMP_LOOP_9_acc_10_itm_10_1_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_503_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_271 ) begin
      COMP_LOOP_COMP_LOOP_and_503_itm <= (COMP_LOOP_9_acc_10_itm_10_1_1[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_504_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_271 ) begin
      COMP_LOOP_COMP_LOOP_and_504_itm <= (COMP_LOOP_9_acc_10_itm_10_1_1[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_505_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_271 ) begin
      COMP_LOOP_COMP_LOOP_and_505_itm <= (COMP_LOOP_9_acc_10_itm_10_1_1[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_506_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_271 ) begin
      COMP_LOOP_COMP_LOOP_and_506_itm <= (COMP_LOOP_9_acc_10_itm_10_1_1[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_507_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_271 ) begin
      COMP_LOOP_COMP_LOOP_and_507_itm <= (COMP_LOOP_9_acc_10_itm_10_1_1[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_508_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_271 ) begin
      COMP_LOOP_COMP_LOOP_and_508_itm <= (COMP_LOOP_9_acc_10_itm_10_1_1[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_509_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_271 ) begin
      COMP_LOOP_COMP_LOOP_and_509_itm <= (COMP_LOOP_9_acc_10_itm_10_1_1[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_10_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_tmp_2357, mux_2375_nl, fsm_output[5]) ) begin
      COMP_LOOP_acc_1_cse_10_sva <= nl_COMP_LOOP_acc_1_cse_10_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_10_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_tmp_2357, mux_2378_nl, fsm_output[5]) ) begin
      COMP_LOOP_acc_10_cse_10_1_10_sva <= COMP_LOOP_10_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_tmp_2357, and_390_nl, fsm_output[5]) ) begin
      COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_11_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_37_itm <= 1'b0;
      COMP_LOOP_nor_371_itm <= 1'b0;
      COMP_LOOP_nor_372_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_557_itm <= 1'b0;
      COMP_LOOP_nor_374_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_559_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_560_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_561_itm <= 1'b0;
      COMP_LOOP_nor_377_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_563_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_564_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_565_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_566_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_567_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_568_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_569_itm <= 1'b0;
    end
    else if ( mux_2383_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_37_itm <= ~((COMP_LOOP_10_acc_10_itm_10_1_1[3:0]!=4'b0000));
      COMP_LOOP_nor_371_itm <= ~((COMP_LOOP_10_acc_10_itm_10_1_1[3:1]!=3'b000));
      COMP_LOOP_nor_372_itm <= ~((COMP_LOOP_10_acc_10_itm_10_1_1[3]) | (COMP_LOOP_10_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_10_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_557_itm <= (COMP_LOOP_10_acc_10_itm_10_1_1[3:0]==4'b0011);
      COMP_LOOP_nor_374_itm <= ~((COMP_LOOP_10_acc_10_itm_10_1_1[3]) | (COMP_LOOP_10_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_10_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_559_itm <= (COMP_LOOP_10_acc_10_itm_10_1_1[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_560_itm <= (COMP_LOOP_10_acc_10_itm_10_1_1[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_561_itm <= (COMP_LOOP_10_acc_10_itm_10_1_1[3:0]==4'b0111);
      COMP_LOOP_nor_377_itm <= ~((COMP_LOOP_10_acc_10_itm_10_1_1[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_563_itm <= (COMP_LOOP_10_acc_10_itm_10_1_1[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_564_itm <= (COMP_LOOP_10_acc_10_itm_10_1_1[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_565_itm <= (COMP_LOOP_10_acc_10_itm_10_1_1[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_566_itm <= (COMP_LOOP_10_acc_10_itm_10_1_1[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_567_itm <= (COMP_LOOP_10_acc_10_itm_10_1_1[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_568_itm <= (COMP_LOOP_10_acc_10_itm_10_1_1[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_569_itm <= (COMP_LOOP_10_acc_10_itm_10_1_1[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_17_psp_sva <= 9'b000000000;
    end
    else if ( MUX_s_1_2_2(mux_2389_nl, nor_tmp_115, fsm_output[5]) ) begin
      COMP_LOOP_acc_17_psp_sva <= nl_COMP_LOOP_acc_17_psp_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_11_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_2392_nl, nor_tmp_115, fsm_output[5]) ) begin
      COMP_LOOP_acc_10_cse_10_1_11_sva <= COMP_LOOP_11_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_2395_nl, nor_tmp_115, fsm_output[5]) ) begin
      COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm <= readslicef_9_1_8(COMP_LOOP_acc_18_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_41_itm <= 1'b0;
      COMP_LOOP_nor_411_itm <= 1'b0;
      COMP_LOOP_nor_412_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_617_itm <= 1'b0;
      COMP_LOOP_nor_414_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_619_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_620_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_621_itm <= 1'b0;
      COMP_LOOP_nor_417_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_623_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_624_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_625_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_626_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_627_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_628_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_629_itm <= 1'b0;
    end
    else if ( mux_2398_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_41_itm <= ~((COMP_LOOP_11_acc_10_itm_10_1_1[3:0]!=4'b0000));
      COMP_LOOP_nor_411_itm <= ~((COMP_LOOP_11_acc_10_itm_10_1_1[3:1]!=3'b000));
      COMP_LOOP_nor_412_itm <= ~((COMP_LOOP_11_acc_10_itm_10_1_1[3]) | (COMP_LOOP_11_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_11_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_617_itm <= (COMP_LOOP_11_acc_10_itm_10_1_1[3:0]==4'b0011);
      COMP_LOOP_nor_414_itm <= ~((COMP_LOOP_11_acc_10_itm_10_1_1[3]) | (COMP_LOOP_11_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_11_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_619_itm <= (COMP_LOOP_11_acc_10_itm_10_1_1[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_620_itm <= (COMP_LOOP_11_acc_10_itm_10_1_1[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_621_itm <= (COMP_LOOP_11_acc_10_itm_10_1_1[3:0]==4'b0111);
      COMP_LOOP_nor_417_itm <= ~((COMP_LOOP_11_acc_10_itm_10_1_1[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_623_itm <= (COMP_LOOP_11_acc_10_itm_10_1_1[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_624_itm <= (COMP_LOOP_11_acc_10_itm_10_1_1[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_625_itm <= (COMP_LOOP_11_acc_10_itm_10_1_1[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_626_itm <= (COMP_LOOP_11_acc_10_itm_10_1_1[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_627_itm <= (COMP_LOOP_11_acc_10_itm_10_1_1[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_628_itm <= (COMP_LOOP_11_acc_10_itm_10_1_1[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_629_itm <= (COMP_LOOP_11_acc_10_itm_10_1_1[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_12_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_2400_nl, (fsm_output[8]), fsm_output[7]) ) begin
      COMP_LOOP_acc_1_cse_12_sva <= nl_COMP_LOOP_acc_1_cse_12_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_12_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_tmp_2384, mux_2402_nl, fsm_output[5]) ) begin
      COMP_LOOP_acc_10_cse_10_1_12_sva <= COMP_LOOP_12_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_tmp_2384, mux_2405_nl, fsm_output[5]) ) begin
      COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_13_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_45_itm <= 1'b0;
      COMP_LOOP_nor_451_itm <= 1'b0;
      COMP_LOOP_nor_452_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_677_itm <= 1'b0;
      COMP_LOOP_nor_454_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_679_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_680_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_681_itm <= 1'b0;
      COMP_LOOP_nor_457_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_683_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_684_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_685_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_686_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_687_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_688_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_689_itm <= 1'b0;
    end
    else if ( mux_2410_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_45_itm <= ~((COMP_LOOP_12_acc_10_itm_10_1_1[3:0]!=4'b0000));
      COMP_LOOP_nor_451_itm <= ~((COMP_LOOP_12_acc_10_itm_10_1_1[3:1]!=3'b000));
      COMP_LOOP_nor_452_itm <= ~((COMP_LOOP_12_acc_10_itm_10_1_1[3]) | (COMP_LOOP_12_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_12_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_677_itm <= (COMP_LOOP_12_acc_10_itm_10_1_1[3:0]==4'b0011);
      COMP_LOOP_nor_454_itm <= ~((COMP_LOOP_12_acc_10_itm_10_1_1[3]) | (COMP_LOOP_12_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_12_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_679_itm <= (COMP_LOOP_12_acc_10_itm_10_1_1[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_680_itm <= (COMP_LOOP_12_acc_10_itm_10_1_1[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_681_itm <= (COMP_LOOP_12_acc_10_itm_10_1_1[3:0]==4'b0111);
      COMP_LOOP_nor_457_itm <= ~((COMP_LOOP_12_acc_10_itm_10_1_1[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_683_itm <= (COMP_LOOP_12_acc_10_itm_10_1_1[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_684_itm <= (COMP_LOOP_12_acc_10_itm_10_1_1[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_685_itm <= (COMP_LOOP_12_acc_10_itm_10_1_1[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_686_itm <= (COMP_LOOP_12_acc_10_itm_10_1_1[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_687_itm <= (COMP_LOOP_12_acc_10_itm_10_1_1[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_688_itm <= (COMP_LOOP_12_acc_10_itm_10_1_1[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_689_itm <= (COMP_LOOP_12_acc_10_itm_10_1_1[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_19_psp_sva <= 8'b00000000;
    end
    else if ( MUX_s_1_2_2(mux_2415_nl, and_733_cse, fsm_output[5]) ) begin
      COMP_LOOP_acc_19_psp_sva <= nl_COMP_LOOP_acc_19_psp_sva[7:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_13_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_2418_nl, and_733_cse, fsm_output[5]) ) begin
      COMP_LOOP_acc_10_cse_10_1_13_sva <= COMP_LOOP_13_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_2422_nl, and_733_cse, fsm_output[5]) ) begin
      COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_14_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_49_itm <= 1'b0;
      COMP_LOOP_nor_491_itm <= 1'b0;
      COMP_LOOP_nor_492_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_737_itm <= 1'b0;
      COMP_LOOP_nor_494_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_739_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_740_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_741_itm <= 1'b0;
      COMP_LOOP_nor_497_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_743_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_744_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_745_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_746_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_747_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_748_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_749_itm <= 1'b0;
    end
    else if ( mux_2424_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_49_itm <= ~((COMP_LOOP_13_acc_10_itm_10_1_1[3:0]!=4'b0000));
      COMP_LOOP_nor_491_itm <= ~((COMP_LOOP_13_acc_10_itm_10_1_1[3:1]!=3'b000));
      COMP_LOOP_nor_492_itm <= ~((COMP_LOOP_13_acc_10_itm_10_1_1[3]) | (COMP_LOOP_13_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_13_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_737_itm <= (COMP_LOOP_13_acc_10_itm_10_1_1[3:0]==4'b0011);
      COMP_LOOP_nor_494_itm <= ~((COMP_LOOP_13_acc_10_itm_10_1_1[3]) | (COMP_LOOP_13_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_13_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_739_itm <= (COMP_LOOP_13_acc_10_itm_10_1_1[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_740_itm <= (COMP_LOOP_13_acc_10_itm_10_1_1[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_741_itm <= (COMP_LOOP_13_acc_10_itm_10_1_1[3:0]==4'b0111);
      COMP_LOOP_nor_497_itm <= ~((COMP_LOOP_13_acc_10_itm_10_1_1[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_743_itm <= (COMP_LOOP_13_acc_10_itm_10_1_1[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_744_itm <= (COMP_LOOP_13_acc_10_itm_10_1_1[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_745_itm <= (COMP_LOOP_13_acc_10_itm_10_1_1[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_746_itm <= (COMP_LOOP_13_acc_10_itm_10_1_1[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_747_itm <= (COMP_LOOP_13_acc_10_itm_10_1_1[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_748_itm <= (COMP_LOOP_13_acc_10_itm_10_1_1[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_749_itm <= (COMP_LOOP_13_acc_10_itm_10_1_1[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_14_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_2426_nl, and_733_cse, fsm_output[6]) ) begin
      COMP_LOOP_acc_1_cse_14_sva <= nl_COMP_LOOP_acc_1_cse_14_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_14_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_tmp_2410, mux_2428_nl, fsm_output[5]) ) begin
      COMP_LOOP_acc_10_cse_10_1_14_sva <= COMP_LOOP_14_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_tmp_2410, mux_2431_nl, fsm_output[5]) ) begin
      COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_15_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_53_itm <= 1'b0;
      COMP_LOOP_nor_531_itm <= 1'b0;
      COMP_LOOP_nor_532_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_797_itm <= 1'b0;
      COMP_LOOP_nor_534_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_799_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_800_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_801_itm <= 1'b0;
      COMP_LOOP_nor_537_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_803_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_804_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_805_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_806_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_807_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_808_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_809_itm <= 1'b0;
    end
    else if ( mux_2435_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_53_itm <= ~((COMP_LOOP_14_acc_10_itm_10_1_1[3:0]!=4'b0000));
      COMP_LOOP_nor_531_itm <= ~((COMP_LOOP_14_acc_10_itm_10_1_1[3:1]!=3'b000));
      COMP_LOOP_nor_532_itm <= ~((COMP_LOOP_14_acc_10_itm_10_1_1[3]) | (COMP_LOOP_14_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_14_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_797_itm <= (COMP_LOOP_14_acc_10_itm_10_1_1[3:0]==4'b0011);
      COMP_LOOP_nor_534_itm <= ~((COMP_LOOP_14_acc_10_itm_10_1_1[3]) | (COMP_LOOP_14_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_14_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_799_itm <= (COMP_LOOP_14_acc_10_itm_10_1_1[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_800_itm <= (COMP_LOOP_14_acc_10_itm_10_1_1[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_801_itm <= (COMP_LOOP_14_acc_10_itm_10_1_1[3:0]==4'b0111);
      COMP_LOOP_nor_537_itm <= ~((COMP_LOOP_14_acc_10_itm_10_1_1[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_803_itm <= (COMP_LOOP_14_acc_10_itm_10_1_1[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_804_itm <= (COMP_LOOP_14_acc_10_itm_10_1_1[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_805_itm <= (COMP_LOOP_14_acc_10_itm_10_1_1[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_806_itm <= (COMP_LOOP_14_acc_10_itm_10_1_1[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_807_itm <= (COMP_LOOP_14_acc_10_itm_10_1_1[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_808_itm <= (COMP_LOOP_14_acc_10_itm_10_1_1[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_809_itm <= (COMP_LOOP_14_acc_10_itm_10_1_1[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_20_psp_sva <= 9'b000000000;
    end
    else if ( MUX_s_1_2_2(mux_2436_nl, and_dcpl_57, fsm_output[5]) ) begin
      COMP_LOOP_acc_20_psp_sva <= nl_COMP_LOOP_acc_20_psp_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_15_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_2438_nl, and_dcpl_57, fsm_output[5]) ) begin
      COMP_LOOP_acc_10_cse_10_1_15_sva <= COMP_LOOP_15_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( mux_2442_itm ) begin
      COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm <= readslicef_7_1_6(COMP_LOOP_acc_21_nl);
      reg_COMP_LOOP_k_10_4_ftd <= COMP_LOOP_k_10_4_sva_2[5:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_57_itm <= 1'b0;
      COMP_LOOP_nor_571_itm <= 1'b0;
      COMP_LOOP_nor_572_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_857_itm <= 1'b0;
      COMP_LOOP_nor_574_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_859_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_860_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_861_itm <= 1'b0;
      COMP_LOOP_nor_577_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_863_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_864_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_865_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_866_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_867_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_868_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_869_itm <= 1'b0;
    end
    else if ( mux_2444_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_57_itm <= ~((COMP_LOOP_15_acc_10_itm_10_1_1[3:0]!=4'b0000));
      COMP_LOOP_nor_571_itm <= ~((COMP_LOOP_15_acc_10_itm_10_1_1[3:1]!=3'b000));
      COMP_LOOP_nor_572_itm <= ~((COMP_LOOP_15_acc_10_itm_10_1_1[3]) | (COMP_LOOP_15_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_15_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_857_itm <= (COMP_LOOP_15_acc_10_itm_10_1_1[3:0]==4'b0011);
      COMP_LOOP_nor_574_itm <= ~((COMP_LOOP_15_acc_10_itm_10_1_1[3]) | (COMP_LOOP_15_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_15_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_859_itm <= (COMP_LOOP_15_acc_10_itm_10_1_1[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_860_itm <= (COMP_LOOP_15_acc_10_itm_10_1_1[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_861_itm <= (COMP_LOOP_15_acc_10_itm_10_1_1[3:0]==4'b0111);
      COMP_LOOP_nor_577_itm <= ~((COMP_LOOP_15_acc_10_itm_10_1_1[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_863_itm <= (COMP_LOOP_15_acc_10_itm_10_1_1[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_864_itm <= (COMP_LOOP_15_acc_10_itm_10_1_1[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_865_itm <= (COMP_LOOP_15_acc_10_itm_10_1_1[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_866_itm <= (COMP_LOOP_15_acc_10_itm_10_1_1[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_867_itm <= (COMP_LOOP_15_acc_10_itm_10_1_1[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_868_itm <= (COMP_LOOP_15_acc_10_itm_10_1_1[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_869_itm <= (COMP_LOOP_15_acc_10_itm_10_1_1[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_762, and_303_nl, fsm_output[5]) ) begin
      COMP_LOOP_acc_1_cse_sva <= nl_COMP_LOOP_acc_1_cse_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_762, and_363_nl, fsm_output[5]) ) begin
      COMP_LOOP_acc_10_cse_10_1_sva <= COMP_LOOP_16_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(not_tmp_762, and_304_nl, fsm_output[5]) ) begin
      COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_1_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_61_itm <= 1'b0;
      COMP_LOOP_nor_611_itm <= 1'b0;
      COMP_LOOP_nor_612_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_917_itm <= 1'b0;
      COMP_LOOP_nor_614_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_919_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_920_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_921_itm <= 1'b0;
      COMP_LOOP_nor_617_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_923_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_924_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_925_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_926_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_927_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_928_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_929_itm <= 1'b0;
    end
    else if ( mux_2449_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_61_itm <= ~((COMP_LOOP_16_acc_10_itm_10_1_1[3:0]!=4'b0000));
      COMP_LOOP_nor_611_itm <= ~((COMP_LOOP_16_acc_10_itm_10_1_1[3:1]!=3'b000));
      COMP_LOOP_nor_612_itm <= ~((COMP_LOOP_16_acc_10_itm_10_1_1[3]) | (COMP_LOOP_16_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_16_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_917_itm <= (COMP_LOOP_16_acc_10_itm_10_1_1[3:0]==4'b0011);
      COMP_LOOP_nor_614_itm <= ~((COMP_LOOP_16_acc_10_itm_10_1_1[3]) | (COMP_LOOP_16_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_16_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_919_itm <= (COMP_LOOP_16_acc_10_itm_10_1_1[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_920_itm <= (COMP_LOOP_16_acc_10_itm_10_1_1[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_921_itm <= (COMP_LOOP_16_acc_10_itm_10_1_1[3:0]==4'b0111);
      COMP_LOOP_nor_617_itm <= ~((COMP_LOOP_16_acc_10_itm_10_1_1[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_923_itm <= (COMP_LOOP_16_acc_10_itm_10_1_1[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_924_itm <= (COMP_LOOP_16_acc_10_itm_10_1_1[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_925_itm <= (COMP_LOOP_16_acc_10_itm_10_1_1[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_926_itm <= (COMP_LOOP_16_acc_10_itm_10_1_1[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_927_itm <= (COMP_LOOP_16_acc_10_itm_10_1_1[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_928_itm <= (COMP_LOOP_16_acc_10_itm_10_1_1[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_929_itm <= (COMP_LOOP_16_acc_10_itm_10_1_1[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_10_tmp_mul_idiv_sva <= 10'b0000000000;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm <= 1'b0;
      COMP_LOOP_tmp_nor_13_itm <= 1'b0;
      COMP_LOOP_tmp_nor_14_itm <= 1'b0;
      COMP_LOOP_tmp_nor_16_itm <= 1'b0;
      COMP_LOOP_tmp_nor_19_itm <= 1'b0;
    end
    else if ( COMP_LOOP_tmp_or_1_cse ) begin
      COMP_LOOP_10_tmp_mul_idiv_sva <= z_out_3[9:0];
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_23_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_cse,
          {and_dcpl_62 , and_dcpl_189 , COMP_LOOP_or_27_cse});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_24_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_cse,
          {and_dcpl_62 , and_dcpl_189 , COMP_LOOP_or_27_cse});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_25_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_cse,
          {and_dcpl_62 , and_dcpl_189 , COMP_LOOP_or_27_cse});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_26_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse,
          {and_dcpl_62 , and_dcpl_189 , COMP_LOOP_or_27_cse});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_27_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse,
          {and_dcpl_62 , and_dcpl_189 , COMP_LOOP_or_27_cse});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_28_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse,
          {and_dcpl_62 , and_dcpl_189 , COMP_LOOP_or_27_cse});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_29_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse,
          {and_dcpl_62 , and_dcpl_189 , COMP_LOOP_or_27_cse});
      COMP_LOOP_tmp_nor_13_itm <= MUX_s_1_2_2(COMP_LOOP_nor_11_nl, COMP_LOOP_tmp_nor_cse,
          COMP_LOOP_or_23_cse);
      COMP_LOOP_tmp_nor_14_itm <= MUX_s_1_2_2(COMP_LOOP_nor_12_nl, COMP_LOOP_tmp_nor_1_cse,
          COMP_LOOP_or_23_cse);
      COMP_LOOP_tmp_nor_16_itm <= MUX_s_1_2_2(COMP_LOOP_nor_14_nl, COMP_LOOP_tmp_nor_3_cse,
          COMP_LOOP_or_23_cse);
      COMP_LOOP_tmp_nor_19_itm <= MUX_s_1_2_2(COMP_LOOP_nor_17_nl, COMP_LOOP_tmp_nor_6_cse,
          COMP_LOOP_or_23_cse);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm <= 1'b0;
    end
    else if ( COMP_LOOP_tmp_or_2_cse ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_17_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_17_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_cse,
          {and_dcpl_62 , and_dcpl_65 , COMP_LOOP_or_27_cse});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_19_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_19_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_cse,
          {and_dcpl_62 , and_dcpl_65 , COMP_LOOP_or_27_cse});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_20_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_20_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_cse,
          {and_dcpl_62 , and_dcpl_65 , COMP_LOOP_or_27_cse});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_21_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_21_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_cse,
          {and_dcpl_62 , and_dcpl_65 , COMP_LOOP_or_27_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm <= 1'b0;
    end
    else if ( and_dcpl_62 | and_dcpl_189 | and_dcpl_195 | and_dcpl_197 | and_dcpl_198
        ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_nor_1_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_17_cse,
          {and_dcpl_62 , and_dcpl_189 , COMP_LOOP_or_31_cse});
    end
  end
  always @(posedge clk) begin
    if ( ~(or_dcpl_183 | or_dcpl_207) ) begin
      COMP_LOOP_3_tmp_lshift_ncse_sva <= z_out_1[8:0];
    end
  end
  always @(posedge clk) begin
    if ( mux_2565_nl & (fsm_output[6:5]==2'b00) & nor_1630_cse ) begin
      tmp_33_sva_1 <= MUX1HOT_v_64_4_2(twiddle_rsc_0_1_i_q_d, twiddle_rsc_0_6_i_q_d,
          twiddle_rsc_0_12_i_q_d, COMP_LOOP_tmp_mux1h_4_itm_mx0w3, {and_dcpl_175
          , and_dcpl_180 , and_dcpl_277 , and_311_nl});
    end
  end
  always @(posedge clk) begin
    if ( (COMP_LOOP_tmp_nor_1_itm | COMP_LOOP_tmp_nor_14_itm) & (COMP_LOOP_10_tmp_mul_idiv_sva[1])
        ) begin
      tmp_33_sva_2 <= twiddle_rsc_0_2_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm ) begin
      tmp_33_sva_3 <= twiddle_rsc_0_3_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( (COMP_LOOP_tmp_nor_3_itm | COMP_LOOP_tmp_nor_16_itm) & (COMP_LOOP_10_tmp_mul_idiv_sva[2])
        ) begin
      tmp_33_sva_4 <= twiddle_rsc_0_4_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_5 | COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_itm ) begin
      tmp_33_sva_5 <= twiddle_rsc_0_5_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm ) begin
      tmp_33_sva_7 <= twiddle_rsc_0_7_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm ) begin
      tmp_33_sva_9 <= twiddle_rsc_0_9_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_5 | COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm ) begin
      tmp_33_sva_10 <= twiddle_rsc_0_10_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm ) begin
      tmp_33_sva_15 <= twiddle_rsc_0_15_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_itm <= 1'b0;
    end
    else if ( and_dcpl_65 | and_dcpl_181 | and_dcpl_190 | and_dcpl_183 | and_dcpl_191
        | and_dcpl_184 | and_dcpl_192 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_nor_6_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_nor_cse, COMP_LOOP_or_27_cse);
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_2463_nl, and_dcpl_57, fsm_output[5]) ) begin
      COMP_LOOP_tmp_mux1h_12_itm <= MUX1HOT_v_64_6_2(twiddle_rsc_0_0_i_q_d, tmp_33_sva_13,
          tmp_33_sva_1, tmp_33_sva_10, tmp_33_sva_11, tmp_33_sva_12, {COMP_LOOP_tmp_or_33_nl
          , COMP_LOOP_tmp_and_55_nl , COMP_LOOP_tmp_and_56_nl , COMP_LOOP_tmp_and_57_nl
          , COMP_LOOP_tmp_and_58_nl , COMP_LOOP_tmp_and_59_nl});
    end
  end
  always @(posedge clk) begin
    if ( and_dcpl_65 | and_dcpl_189 | COMP_LOOP_10_acc_8_itm_mx0c2 | COMP_LOOP_10_acc_8_itm_mx0c3
        | and_dcpl_70 | and_dcpl_220 | COMP_LOOP_10_acc_8_itm_mx0c6 | and_dcpl_74
        | and_dcpl_222 | COMP_LOOP_10_acc_8_itm_mx0c9 | and_dcpl_81 | and_dcpl_223
        | COMP_LOOP_10_acc_8_itm_mx0c12 | and_dcpl_86 | and_dcpl_225 | COMP_LOOP_10_acc_8_itm_mx0c15
        | and_dcpl_93 | and_dcpl_226 | COMP_LOOP_10_acc_8_itm_mx0c18 | and_dcpl_95
        | and_dcpl_227 | COMP_LOOP_10_acc_8_itm_mx0c21 | and_dcpl_100 | and_dcpl_228
        | COMP_LOOP_10_acc_8_itm_mx0c24 | and_dcpl_102 | and_dcpl_229 | COMP_LOOP_10_acc_8_itm_mx0c27
        | and_dcpl_108 | and_dcpl_230 | COMP_LOOP_10_acc_8_itm_mx0c30 | and_dcpl_110
        | and_dcpl_231 | COMP_LOOP_10_acc_8_itm_mx0c33 | and_dcpl_116 | and_dcpl_232
        | COMP_LOOP_10_acc_8_itm_mx0c36 | and_dcpl_119 | and_dcpl_233 | COMP_LOOP_10_acc_8_itm_mx0c39
        | and_dcpl_125 | and_dcpl_234 | COMP_LOOP_10_acc_8_itm_mx0c42 | and_dcpl_127
        | and_dcpl_235 | and_dcpl_130 | and_dcpl_236 | COMP_LOOP_10_acc_8_itm_mx0c47
        ) begin
      COMP_LOOP_10_acc_8_itm <= MUX1HOT_v_64_19_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d,
          vec_rsc_0_2_i_q_d, vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d,
          vec_rsc_0_6_i_q_d, vec_rsc_0_7_i_q_d, vec_rsc_0_8_i_q_d, vec_rsc_0_9_i_q_d,
          vec_rsc_0_10_i_q_d, vec_rsc_0_11_i_q_d, vec_rsc_0_12_i_q_d, vec_rsc_0_13_i_q_d,
          vec_rsc_0_14_i_q_d, vec_rsc_0_15_i_q_d, COMP_LOOP_acc_23_nl, z_out_3, COMP_LOOP_1_modulo_cmp_return_rsc_z,
          {COMP_LOOP_or_nl , COMP_LOOP_or_1_nl , COMP_LOOP_or_2_nl , COMP_LOOP_or_3_nl
          , COMP_LOOP_or_4_nl , COMP_LOOP_or_5_nl , COMP_LOOP_or_6_nl , COMP_LOOP_or_7_nl
          , COMP_LOOP_or_8_nl , COMP_LOOP_or_9_nl , COMP_LOOP_or_10_nl , COMP_LOOP_or_11_nl
          , COMP_LOOP_or_12_nl , COMP_LOOP_or_13_nl , COMP_LOOP_or_14_nl , COMP_LOOP_or_15_nl
          , COMP_LOOP_or_21_nl , COMP_LOOP_or_22_nl , COMP_LOOP_10_acc_8_itm_mx0c3});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_11_tmp_mul_idiv_sva <= 9'b000000000;
    end
    else if ( COMP_LOOP_tmp_or_19_cse ) begin
      COMP_LOOP_11_tmp_mul_idiv_sva <= z_out_3[8:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ and_332_tmp ) begin
      COMP_LOOP_tmp_mux1h_itm <= MUX1HOT_v_64_16_2(twiddle_rsc_0_0_i_q_d, tmp_33_sva_1,
          tmp_33_sva_2, tmp_33_sva_3, tmp_33_sva_4, tmp_33_sva_5, tmp_33_sva_6, tmp_33_sva_7,
          tmp_33_sva_8, tmp_33_sva_9, tmp_33_sva_10, tmp_33_sva_11, tmp_33_sva_12,
          tmp_33_sva_13, tmp_33_sva_14, tmp_33_sva_15, {COMP_LOOP_tmp_and_42_nl ,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_1_nl
          , COMP_LOOP_tmp_and_43_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl , COMP_LOOP_tmp_and_44_nl
          , COMP_LOOP_tmp_and_45_nl , COMP_LOOP_tmp_and_46_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_7_nl
          , COMP_LOOP_tmp_and_47_nl , COMP_LOOP_tmp_and_48_nl , COMP_LOOP_tmp_and_49_nl
          , COMP_LOOP_tmp_and_50_nl , COMP_LOOP_tmp_and_51_nl , COMP_LOOP_tmp_and_52_nl
          , COMP_LOOP_tmp_and_53_nl});
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_2504_nl, (fsm_output[8]), or_2589_cse) ) begin
      COMP_LOOP_tmp_mux_itm <= MUX1HOT_v_64_3_2(tmp_33_sva_13_mx0w1, twiddle_rsc_0_8_i_q_d,
          twiddle_rsc_0_0_i_q_d, {and_336_nl , and_dcpl_183 , and_340_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_13_tmp_mul_idiv_sva <= 8'b00000000;
    end
    else if ( and_dcpl_189 | and_dcpl_202 ) begin
      COMP_LOOP_13_tmp_mul_idiv_sva <= MUX_v_8_2_2((z_out_1[7:0]), (z_out_3[7:0]),
          and_dcpl_202);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_12_itm <= 1'b0;
    end
    else if ( COMP_LOOP_tmp_or_21_cse ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_19_cse, COMP_LOOP_or_31_cse);
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_20_cse, COMP_LOOP_or_31_cse);
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_21_cse, COMP_LOOP_or_31_cse);
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_12_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_nor_cse,
          COMP_LOOP_tmp_nor_6_cse, COMP_LOOP_or_31_cse);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_5_tmp_mul_idiv_sva <= 8'b00000000;
    end
    else if ( ~(or_dcpl_182 | (fsm_output[2:1]!=2'b10) | or_dcpl_207) ) begin
      COMP_LOOP_5_tmp_mul_idiv_sva <= z_out_3[7:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ and_341_tmp ) begin
      COMP_LOOP_tmp_mux1h_1_itm <= MUX1HOT_v_64_6_2(twiddle_rsc_0_0_i_q_d, COMP_LOOP_tmp_mux_itm,
          tmp_33_sva_1, tmp_33_sva_10, tmp_33_sva_11, tmp_33_sva_12, {COMP_LOOP_tmp_and_36_nl
          , COMP_LOOP_tmp_and_37_nl , COMP_LOOP_tmp_and_38_nl , COMP_LOOP_tmp_and_39_nl
          , COMP_LOOP_tmp_and_40_nl , COMP_LOOP_tmp_and_41_nl});
    end
  end
  always @(posedge clk) begin
    if ( ~ and_342_tmp ) begin
      COMP_LOOP_tmp_mux1h_2_itm <= MUX1HOT_v_64_16_2(twiddle_rsc_0_0_i_q_d, tmp_33_sva_1,
          tmp_33_sva_2, tmp_33_sva_3, tmp_33_sva_4, tmp_33_sva_5, tmp_33_sva_6, tmp_33_sva_7,
          tmp_33_sva_8, tmp_33_sva_9, tmp_33_sva_10, tmp_33_sva_11, tmp_33_sva_12,
          tmp_33_sva_13, tmp_33_sva_14, tmp_33_sva_15, {COMP_LOOP_tmp_and_20_nl ,
          COMP_LOOP_tmp_and_21_nl , COMP_LOOP_tmp_and_22_nl , COMP_LOOP_tmp_and_23_nl
          , COMP_LOOP_tmp_and_24_nl , COMP_LOOP_tmp_and_25_nl , COMP_LOOP_tmp_and_26_nl
          , COMP_LOOP_tmp_and_27_nl , COMP_LOOP_tmp_and_28_nl , COMP_LOOP_tmp_and_29_nl
          , COMP_LOOP_tmp_and_30_nl , COMP_LOOP_tmp_and_31_nl , COMP_LOOP_tmp_and_32_nl
          , COMP_LOOP_tmp_and_33_nl , COMP_LOOP_tmp_and_34_nl , COMP_LOOP_tmp_and_35_nl});
    end
  end
  always @(posedge clk) begin
    if ( (COMP_LOOP_tmp_COMP_LOOP_tmp_nor_14_cse | ((COMP_LOOP_13_tmp_mul_idiv_sva[1:0]==2'b10))
        | ((COMP_LOOP_13_tmp_mul_idiv_sva[1:0]==2'b11)) | and_dcpl_277) & mux_2518_nl
        ) begin
      tmp_36_sva_1 <= MUX1HOT_v_64_4_2(twiddle_rsc_0_4_i_q_d, twiddle_rsc_0_0_i_q_d,
          tmp_36_sva_2, tmp_33_sva_1, {and_dcpl_277 , COMP_LOOP_tmp_and_nl , COMP_LOOP_tmp_and_17_nl
          , COMP_LOOP_tmp_and_18_nl});
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_2520_nl, and_357_nl, fsm_output[5]) ) begin
      tmp_36_sva_2 <= MUX_v_64_2_2(twiddle_rsc_0_8_i_q_d, COMP_LOOP_tmp_mux1h_4_itm_mx0w3,
          and_dcpl_192);
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_nor_16_rgt | COMP_LOOP_tmp_and_14_rgt | COMP_LOOP_tmp_and_15_rgt
        | COMP_LOOP_tmp_and_16_rgt ) begin
      COMP_LOOP_tmp_mux1h_3_itm <= MUX1HOT_v_64_4_2(twiddle_rsc_0_0_i_q_d, tmp_36_sva_1,
          tmp_36_sva_2, tmp_33_sva_1, {COMP_LOOP_tmp_COMP_LOOP_tmp_nor_16_rgt , COMP_LOOP_tmp_and_14_rgt
          , COMP_LOOP_tmp_and_15_rgt , COMP_LOOP_tmp_and_16_rgt});
    end
  end
  always @(posedge clk) begin
    if ( mux_2532_nl | (fsm_output[8]) ) begin
      COMP_LOOP_tmp_mux1h_4_itm <= COMP_LOOP_tmp_mux1h_4_itm_mx0w3;
    end
  end
  always @(posedge clk) begin
    if ( ~ nor_1796_tmp ) begin
      COMP_LOOP_tmp_mux1h_5_itm <= MUX1HOT_v_64_6_2(twiddle_rsc_0_0_i_q_d, COMP_LOOP_tmp_mux_itm,
          tmp_33_sva_1, tmp_33_sva_10, tmp_33_sva_11, tmp_33_sva_12, {COMP_LOOP_tmp_and_7_nl
          , COMP_LOOP_tmp_and_8_nl , COMP_LOOP_tmp_and_9_nl , COMP_LOOP_tmp_and_10_nl
          , COMP_LOOP_tmp_and_11_nl , COMP_LOOP_tmp_and_12_nl});
    end
  end
  always @(posedge clk) begin
    if ( mux_2542_nl | (fsm_output[8]) ) begin
      COMP_LOOP_tmp_mux1h_6_itm <= COMP_LOOP_tmp_mux1h_4_itm_mx0w3;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_2546_nl, and_352_nl, fsm_output[5]) ) begin
      COMP_LOOP_tmp_mux1h_7_itm <= COMP_LOOP_tmp_mux1h_4_itm_mx0w3;
    end
  end
  always @(posedge clk) begin
    if ( ((~(COMP_LOOP_tmp_COMP_LOOP_tmp_and_155 | COMP_LOOP_tmp_COMP_LOOP_tmp_and_157
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_159)) | COMP_LOOP_tmp_COMP_LOOP_tmp_nor_12_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm
        | and_dcpl_191) & mux_2553_nl ) begin
      COMP_LOOP_tmp_mux1h_8_itm <= MUX1HOT_v_64_6_2(tmp_33_sva_13_mx0w1, twiddle_rsc_0_0_i_q_d,
          tmp_33_sva_1, tmp_33_sva_10, tmp_33_sva_11, tmp_33_sva_12, {and_dcpl_191
          , COMP_LOOP_tmp_and_2_nl , COMP_LOOP_tmp_and_3_nl , COMP_LOOP_tmp_and_4_nl
          , COMP_LOOP_tmp_and_5_nl , COMP_LOOP_tmp_and_6_nl});
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_2556_nl, mux_2554_nl, fsm_output[5]) ) begin
      COMP_LOOP_tmp_mux1h_9_itm <= COMP_LOOP_tmp_mux1h_4_itm_mx0w3;
    end
  end
  assign nor_1871_nl = ~((fsm_output[4]) | (fsm_output[0]) | (fsm_output[3]) | (fsm_output[2])
      | (fsm_output[1]) | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[8]));
  assign and_1183_nl = (fsm_output[4]) & mux_tmp_1062;
  assign VEC_LOOP_j_not_1_nl = ~ VEC_LOOP_j_10_0_sva_9_0_mx0c0;
  assign nor_1870_nl = ~((fsm_output[4]) | (fsm_output[3]) | (fsm_output[2]) | (fsm_output[1])
      | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[8]));
  assign and_nl = (fsm_output[4]) & nor_tmp_339;
  assign nor_1622_nl = ~((fsm_output[4]) | (fsm_output[1]) | (fsm_output[6]) | (fsm_output[7])
      | (fsm_output[8]));
  assign and_568_nl = (fsm_output[4]) & (fsm_output[1]) & (fsm_output[6]) & (fsm_output[7])
      & (fsm_output[8]);
  assign mux_1074_nl = MUX_s_1_2_2(nor_1622_nl, and_568_nl, fsm_output[5]);
  assign nand_nl = ~(mux_1074_nl & nor_1624_cse & (fsm_output[0]));
  assign or_nl = (fsm_output[8:6]!=3'b000) | (~((fsm_output[3:1]!=3'b000)));
  assign mux_2558_nl = MUX_s_1_2_2(or_nl, nand_324_cse, fsm_output[5]);
  assign nand_325_nl = ~((fsm_output[8:6]==3'b111) & or_2259_cse_1);
  assign nand_323_nl = ~((fsm_output[8:6]==3'b111) & (~(and_1189_cse | (fsm_output[3:2]!=2'b00))));
  assign mux_nl = MUX_s_1_2_2(nand_325_nl, nand_323_nl, fsm_output[5]);
  assign nl_COMP_LOOP_acc_psp_sva  = (VEC_LOOP_j_10_0_sva_9_0[9:4]) + COMP_LOOP_k_10_4_sva_5_0;
  assign mux_2308_nl = MUX_s_1_2_2(mux_tmp_2288, nor_tmp_489, fsm_output[4]);
  assign mux_2309_nl = MUX_s_1_2_2(mux_2308_nl, (fsm_output[7]), fsm_output[5]);
  assign and_270_nl = (fsm_output[4]) & mux_tmp_2291;
  assign mux_2312_nl = MUX_s_1_2_2(not_tmp_703, and_270_nl, fsm_output[5]);
  assign nand_320_nl = ~((fsm_output[4:0]==5'b11111));
  assign mux_2314_nl = MUX_s_1_2_2(or_tmp_2300, nand_320_nl, fsm_output[5]);
  assign nand_111_nl = ~((fsm_output[4:1]==4'b1111));
  assign mux_2315_nl = MUX_s_1_2_2(or_tmp_2300, nand_111_nl, fsm_output[5]);
  assign nl_COMP_LOOP_3_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_4_sva_5_0 , 4'b0010}) + 11'b00000000001;
  assign COMP_LOOP_3_acc_nl = nl_COMP_LOOP_3_acc_nl[10:0];
  assign nl_COMP_LOOP_acc_11_psp_sva  = (VEC_LOOP_j_10_0_sva_9_0[9:1]) + ({COMP_LOOP_k_10_4_sva_5_0
      , 3'b001});
  assign mux_2316_nl = MUX_s_1_2_2((~ mux_tmp_2292), nor_tmp_10, fsm_output[4]);
  assign mux_2317_nl = MUX_s_1_2_2(mux_2316_nl, (fsm_output[6]), fsm_output[5]);
  assign mux_2318_nl = MUX_s_1_2_2((~ mux_tmp_2292), mux_tmp_2291, fsm_output[4]);
  assign mux_2319_nl = MUX_s_1_2_2(mux_2318_nl, (fsm_output[6]), fsm_output[5]);
  assign nl_COMP_LOOP_acc_12_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:3]))})
      + conv_u2u_8_9({COMP_LOOP_k_10_4_sva_5_0 , 2'b00}) + 9'b000000001;
  assign COMP_LOOP_acc_12_nl = nl_COMP_LOOP_acc_12_nl[8:0];
  assign nand_110_nl = ~((fsm_output[0]) & (fsm_output[3]) & (fsm_output[2]) & (fsm_output[1])
      & (fsm_output[6]));
  assign mux_2320_nl = MUX_s_1_2_2(mux_tmp_2292, nand_110_nl, fsm_output[4]);
  assign mux_2321_nl = MUX_s_1_2_2(mux_2320_nl, (~ (fsm_output[6])), fsm_output[5]);
  assign and_823_nl = (fsm_output[2]) & (fsm_output[3]) & (fsm_output[4]) & (fsm_output[6]);
  assign mux_2326_nl = MUX_s_1_2_2(not_tmp_703, and_823_nl, fsm_output[5]);
  assign nl_COMP_LOOP_5_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_4_sva_5_0 , 4'b0100}) + 11'b00000000001;
  assign COMP_LOOP_5_acc_nl = nl_COMP_LOOP_5_acc_nl[10:0];
  assign and_412_nl = (fsm_output[4]) & (fsm_output[3]) & (fsm_output[2]) & (fsm_output[1])
      & (fsm_output[6]);
  assign mux_2327_nl = MUX_s_1_2_2(not_tmp_703, and_412_nl, fsm_output[5]);
  assign mux_2331_nl = MUX_s_1_2_2(mux_tmp_2288, mux_tmp_2311, fsm_output[4]);
  assign mux_2332_nl = MUX_s_1_2_2(mux_2331_nl, (fsm_output[7]), fsm_output[5]);
  assign nl_COMP_LOOP_6_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_4_sva_5_0 , 4'b0101}) + 11'b00000000001;
  assign COMP_LOOP_6_acc_nl = nl_COMP_LOOP_6_acc_nl[10:0];
  assign and_408_nl = (and_831_cse | (fsm_output[6])) & (fsm_output[7]);
  assign mux_2333_nl = MUX_s_1_2_2(and_408_nl, nor_tmp_489, fsm_output[0]);
  assign mux_2334_nl = MUX_s_1_2_2(mux_tmp_2288, mux_2333_nl, fsm_output[4]);
  assign mux_2335_nl = MUX_s_1_2_2(mux_2334_nl, (fsm_output[7]), fsm_output[5]);
  assign nl_COMP_LOOP_acc_1_cse_6_sva  = VEC_LOOP_j_10_0_sva_9_0 + ({COMP_LOOP_k_10_4_sva_5_0
      , 4'b0101});
  assign mux_2336_nl = MUX_s_1_2_2(nor_tmp_47, mux_tmp_2311, fsm_output[4]);
  assign mux_2338_nl = MUX_s_1_2_2(mux_tmp_2318, mux_2336_nl, fsm_output[5]);
  assign mux_2339_nl = MUX_s_1_2_2(nor_tmp_47, nor_tmp_499, and_407_cse);
  assign mux_2340_nl = MUX_s_1_2_2(mux_tmp_2318, mux_2339_nl, fsm_output[5]);
  assign nl_COMP_LOOP_7_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_4_sva_5_0 , 4'b0110}) + 11'b00000000001;
  assign COMP_LOOP_7_acc_nl = nl_COMP_LOOP_7_acc_nl[10:0];
  assign and_405_nl = (((fsm_output[4:2]==3'b111)) | (fsm_output[6])) & (fsm_output[7]);
  assign mux_2341_nl = MUX_s_1_2_2(mux_tmp_2318, and_405_nl, fsm_output[5]);
  assign nl_COMP_LOOP_acc_14_psp_sva  = (VEC_LOOP_j_10_0_sva_9_0[9:1]) + ({COMP_LOOP_k_10_4_sva_5_0
      , 3'b011});
  assign mux_2345_nl = MUX_s_1_2_2((~ mux_tmp_2325), and_tmp_28, fsm_output[4]);
  assign mux_2346_nl = MUX_s_1_2_2(mux_2345_nl, nor_tmp_47, fsm_output[5]);
  assign mux_2348_nl = MUX_s_1_2_2((~ mux_tmp_2325), mux_tmp_2328, fsm_output[4]);
  assign mux_2349_nl = MUX_s_1_2_2(mux_2348_nl, nor_tmp_47, fsm_output[5]);
  assign nl_COMP_LOOP_acc_15_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:4]))})
      + conv_u2u_7_8({COMP_LOOP_k_10_4_sva_5_0 , 1'b0}) + 8'b00000001;
  assign COMP_LOOP_acc_15_nl = nl_COMP_LOOP_acc_15_nl[7:0];
  assign mux_2350_nl = MUX_s_1_2_2(nor_tmp_509, and_tmp_28, fsm_output[0]);
  assign mux_2351_nl = MUX_s_1_2_2((~ mux_tmp_2325), mux_2350_nl, fsm_output[4]);
  assign mux_2352_nl = MUX_s_1_2_2(mux_2351_nl, nor_tmp_47, fsm_output[5]);
  assign nl_COMP_LOOP_acc_1_cse_8_sva  = VEC_LOOP_j_10_0_sva_9_0 + ({COMP_LOOP_k_10_4_sva_5_0
      , 4'b0111});
  assign and_296_nl = (fsm_output[4]) & mux_tmp_2328;
  assign mux_2354_nl = MUX_s_1_2_2(not_tmp_727, and_296_nl, fsm_output[5]);
  assign and_397_nl = (fsm_output[4]) & (fsm_output[3]) & (fsm_output[6]) & (fsm_output[7]);
  assign mux_2355_nl = MUX_s_1_2_2(not_tmp_727, and_397_nl, fsm_output[5]);
  assign nl_COMP_LOOP_9_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_4_sva_5_0 , 4'b1000}) + 11'b00000000001;
  assign COMP_LOOP_9_acc_nl = nl_COMP_LOOP_9_acc_nl[10:0];
  assign and_299_nl = (fsm_output[4:3]==2'b11) & nor_tmp_507;
  assign mux_2356_nl = MUX_s_1_2_2(not_tmp_727, and_299_nl, fsm_output[5]);
  assign nl_COMP_LOOP_acc_16_psp_sva  = (VEC_LOOP_j_10_0_sva_9_0[9:3]) + ({COMP_LOOP_k_10_4_sva_5_0
      , 1'b1});
  assign mux_2364_nl = MUX_s_1_2_2(mux_tmp_2344, nor_tmp_515, fsm_output[4]);
  assign mux_2368_nl = MUX_s_1_2_2(mux_tmp_2344, mux_tmp_2348, fsm_output[4]);
  assign nl_COMP_LOOP_10_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_4_sva_5_0 , 4'b1001}) + 11'b00000000001;
  assign COMP_LOOP_10_acc_nl = nl_COMP_LOOP_10_acc_nl[10:0];
  assign mux_2371_nl = MUX_s_1_2_2(mux_tmp_2351, nor_tmp_515, fsm_output[0]);
  assign mux_2372_nl = MUX_s_1_2_2(mux_tmp_2344, mux_2371_nl, fsm_output[4]);
  assign nl_COMP_LOOP_acc_1_cse_10_sva  = VEC_LOOP_j_10_0_sva_9_0 + ({COMP_LOOP_k_10_4_sva_5_0
      , 4'b1001});
  assign mux_2375_nl = MUX_s_1_2_2(nor_tmp_115, mux_tmp_2348, fsm_output[4]);
  assign mux_2378_nl = MUX_s_1_2_2(nor_tmp_115, mux_tmp_2347, fsm_output[4]);
  assign nl_COMP_LOOP_11_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_4_sva_5_0 , 4'b1010}) + 11'b00000000001;
  assign COMP_LOOP_11_acc_nl = nl_COMP_LOOP_11_acc_nl[10:0];
  assign and_390_nl = (and_407_cse | (fsm_output[7:6]!=2'b00)) & (fsm_output[8]);
  assign nl_COMP_LOOP_acc_17_psp_sva  = (VEC_LOOP_j_10_0_sva_9_0[9:1]) + ({COMP_LOOP_k_10_4_sva_5_0
      , 3'b101});
  assign mux_2389_nl = MUX_s_1_2_2(mux_tmp_2369, mux_tmp_2365, fsm_output[4]);
  assign mux_2391_nl = MUX_s_1_2_2(mux_tmp_2365, nor_tmp_528, fsm_output[0]);
  assign mux_2392_nl = MUX_s_1_2_2(mux_tmp_2369, mux_2391_nl, fsm_output[4]);
  assign nl_COMP_LOOP_acc_18_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:3]))})
      + conv_u2u_8_9({COMP_LOOP_k_10_4_sva_5_0 , 2'b10}) + 9'b000000001;
  assign COMP_LOOP_acc_18_nl = nl_COMP_LOOP_acc_18_nl[8:0];
  assign mux_2394_nl = MUX_s_1_2_2(nor_tmp_530, mux_tmp_2365, fsm_output[0]);
  assign mux_2395_nl = MUX_s_1_2_2(mux_tmp_2369, mux_2394_nl, fsm_output[4]);
  assign nl_COMP_LOOP_acc_1_cse_12_sva  = VEC_LOOP_j_10_0_sva_9_0 + ({COMP_LOOP_k_10_4_sva_5_0
      , 4'b1011});
  assign nor_581_nl = ~(and_1189_cse | (fsm_output[4]) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[8]));
  assign and_379_nl = ((fsm_output[1:0]!=2'b00)) & (fsm_output[4]) & (fsm_output[5])
      & (fsm_output[6]) & (fsm_output[8]);
  assign mux_2399_nl = MUX_s_1_2_2(nor_581_nl, and_379_nl, fsm_output[2]);
  assign and_380_nl = (fsm_output[4]) & (fsm_output[5]) & (fsm_output[6]) & (fsm_output[8]);
  assign mux_2400_nl = MUX_s_1_2_2(mux_2399_nl, and_380_nl, fsm_output[3]);
  assign mux_2402_nl = MUX_s_1_2_2(and_733_cse, nor_tmp_528, fsm_output[4]);
  assign nl_COMP_LOOP_13_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_4_sva_5_0 , 4'b1100}) + 11'b00000000001;
  assign COMP_LOOP_13_acc_nl = nl_COMP_LOOP_13_acc_nl[10:0];
  assign mux_2405_nl = MUX_s_1_2_2(and_733_cse, mux_tmp_2365, fsm_output[4]);
  assign nl_COMP_LOOP_acc_19_psp_sva  = (VEC_LOOP_j_10_0_sva_9_0[9:2]) + ({COMP_LOOP_k_10_4_sva_5_0
      , 2'b11});
  assign mux_2415_nl = MUX_s_1_2_2(mux_tmp_2395, nor_tmp_537, fsm_output[4]);
  assign mux_2417_nl = MUX_s_1_2_2(nor_tmp_537, nor_tmp_538, fsm_output[0]);
  assign mux_2418_nl = MUX_s_1_2_2(mux_tmp_2395, mux_2417_nl, fsm_output[4]);
  assign nl_COMP_LOOP_14_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_4_sva_5_0 , 4'b1101}) + 11'b00000000001;
  assign COMP_LOOP_14_acc_nl = nl_COMP_LOOP_14_acc_nl[10:0];
  assign mux_2421_nl = MUX_s_1_2_2(mux_tmp_2401, nor_tmp_537, fsm_output[0]);
  assign mux_2422_nl = MUX_s_1_2_2(mux_tmp_2395, mux_2421_nl, fsm_output[4]);
  assign nl_COMP_LOOP_acc_1_cse_14_sva  = VEC_LOOP_j_10_0_sva_9_0 + ({COMP_LOOP_k_10_4_sva_5_0
      , 4'b1101});
  assign nor_580_nl = ~((fsm_output[4]) | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[8]));
  assign mux_2425_nl = MUX_s_1_2_2(nor_580_nl, nor_tmp_544, and_1189_cse);
  assign mux_2426_nl = MUX_s_1_2_2(mux_2425_nl, nor_tmp_544, or_2259_cse_1);
  assign mux_2428_nl = MUX_s_1_2_2(and_dcpl_57, nor_tmp_538, fsm_output[4]);
  assign nl_COMP_LOOP_15_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_4_sva_5_0 , 4'b1110}) + 11'b00000000001;
  assign COMP_LOOP_15_acc_nl = nl_COMP_LOOP_15_acc_nl[10:0];
  assign mux_2431_nl = MUX_s_1_2_2(and_dcpl_57, nor_tmp_537, fsm_output[4]);
  assign nl_COMP_LOOP_acc_20_psp_sva  = (VEC_LOOP_j_10_0_sva_9_0[9:1]) + ({COMP_LOOP_k_10_4_sva_5_0
      , 3'b111});
  assign mux_2436_nl = MUX_s_1_2_2((~ mux_tmp_2282), nor_tmp_547, fsm_output[4]);
  assign mux_2438_nl = MUX_s_1_2_2((~ mux_tmp_2282), nor_tmp_548, fsm_output[4]);
  assign nl_COMP_LOOP_acc_21_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:5]))})
      + conv_u2u_6_7(COMP_LOOP_k_10_4_sva_5_0) + 7'b0000001;
  assign COMP_LOOP_acc_21_nl = nl_COMP_LOOP_acc_21_nl[6:0];
  assign nl_COMP_LOOP_acc_1_cse_sva  = VEC_LOOP_j_10_0_sva_9_0 + ({COMP_LOOP_k_10_4_sva_5_0
      , 4'b1111});
  assign and_303_nl = (fsm_output[4]) & nor_tmp_548;
  assign and_363_nl = (fsm_output[4]) & (fsm_output[6]) & (fsm_output[7]) & (fsm_output[8]);
  assign nl_COMP_LOOP_1_acc_nl = ({COMP_LOOP_k_10_4_sva_2 , 4'b0000}) + ({1'b1 ,
      (~ (STAGE_LOOP_lshift_psp_sva[10:1]))}) + 11'b00000000001;
  assign COMP_LOOP_1_acc_nl = nl_COMP_LOOP_1_acc_nl[10:0];
  assign and_304_nl = (fsm_output[4]) & nor_tmp_547;
  assign COMP_LOOP_COMP_LOOP_and_23_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[3:0]==4'b1001);
  assign COMP_LOOP_COMP_LOOP_and_24_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[3:0]==4'b1010);
  assign COMP_LOOP_COMP_LOOP_and_25_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[3:0]==4'b1011);
  assign COMP_LOOP_COMP_LOOP_and_26_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[3:0]==4'b1100);
  assign COMP_LOOP_COMP_LOOP_and_27_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[3:0]==4'b1101);
  assign COMP_LOOP_COMP_LOOP_and_28_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[3:0]==4'b1110);
  assign COMP_LOOP_COMP_LOOP_and_29_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[3:0]==4'b1111);
  assign COMP_LOOP_nor_11_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:1]!=3'b000));
  assign COMP_LOOP_nor_12_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3]) | (COMP_LOOP_1_acc_10_itm_10_1_1[2])
      | (COMP_LOOP_1_acc_10_itm_10_1_1[0]));
  assign COMP_LOOP_nor_14_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3]) | (COMP_LOOP_1_acc_10_itm_10_1_1[1])
      | (COMP_LOOP_1_acc_10_itm_10_1_1[0]));
  assign COMP_LOOP_nor_17_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[2:0]!=3'b000));
  assign COMP_LOOP_COMP_LOOP_and_17_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[3:0]==4'b0011);
  assign COMP_LOOP_COMP_LOOP_and_19_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[3:0]==4'b0101);
  assign COMP_LOOP_COMP_LOOP_and_20_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[3:0]==4'b0110);
  assign COMP_LOOP_COMP_LOOP_and_21_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[3:0]==4'b0111);
  assign COMP_LOOP_COMP_LOOP_nor_1_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b0000));
  assign and_311_nl = and_dcpl_61 & and_dcpl_123;
  assign or_2758_nl = (fsm_output[0]) | (fsm_output[2]);
  assign mux_2564_nl = MUX_s_1_2_2(or_2259_cse_1, or_2758_nl, fsm_output[1]);
  assign or_2756_nl = (~ (COMP_LOOP_10_tmp_mul_idiv_sva[3])) | (~ COMP_LOOP_tmp_nor_19_itm)
      | (fsm_output[3]) | (fsm_output[0]) | (fsm_output[2]);
  assign mux_2560_nl = MUX_s_1_2_2(or_2756_nl, or_tmp_2410, and_1190_cse);
  assign mux_2561_nl = MUX_s_1_2_2(mux_2560_nl, or_tmp_2410, and_1191_cse);
  assign or_2754_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm
      | COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm
      | COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm
      | COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm
      | COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm
      | COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm;
  assign mux_2562_nl = MUX_s_1_2_2(mux_2561_nl, or_tmp_2410, or_2754_nl);
  assign mux_2563_nl = MUX_s_1_2_2(or_2259_cse_1, mux_2562_nl, fsm_output[1]);
  assign mux_2565_nl = MUX_s_1_2_2(mux_2564_nl, (~ mux_2563_nl), fsm_output[4]);
  assign COMP_LOOP_tmp_or_33_nl = and_dcpl_65 | (COMP_LOOP_tmp_COMP_LOOP_tmp_nor_12_itm
      & and_314_m1c);
  assign COMP_LOOP_tmp_and_55_nl = COMP_LOOP_tmp_or_29_cse & and_314_m1c;
  assign COMP_LOOP_tmp_and_56_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm & and_314_m1c;
  assign COMP_LOOP_tmp_and_57_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm & and_314_m1c;
  assign COMP_LOOP_tmp_and_58_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm & and_314_m1c;
  assign COMP_LOOP_tmp_and_59_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm & and_314_m1c;
  assign mux_2461_nl = MUX_s_1_2_2(and_dcpl_5, and_dcpl_57, or_2259_cse_1);
  assign mux_2459_nl = MUX_s_1_2_2(and_dcpl_5, mux_tmp_2392, fsm_output[1]);
  assign mux_2460_nl = MUX_s_1_2_2(mux_2459_nl, and_dcpl_57, or_2259_cse_1);
  assign mux_2462_nl = MUX_s_1_2_2(mux_2461_nl, mux_2460_nl, fsm_output[0]);
  assign or_2563_nl = (fsm_output[3:0]!=4'b0001);
  assign mux_2458_nl = MUX_s_1_2_2(mux_tmp_2392, and_dcpl_57, or_2563_nl);
  assign mux_2463_nl = MUX_s_1_2_2(mux_2462_nl, mux_2458_nl, fsm_output[4]);
  assign COMP_LOOP_COMP_LOOP_mux_9_nl = MUX_v_64_2_2(COMP_LOOP_10_acc_8_itm, z_out_7,
      COMP_LOOP_or_18_itm);
  assign nl_COMP_LOOP_acc_23_nl = COMP_LOOP_mux_361_cse + COMP_LOOP_COMP_LOOP_mux_9_nl;
  assign COMP_LOOP_acc_23_nl = nl_COMP_LOOP_acc_23_nl[63:0];
  assign COMP_LOOP_or_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm & and_dcpl_65)
      | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_70) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_74) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_81) | (COMP_LOOP_COMP_LOOP_and_72_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_93) | (COMP_LOOP_COMP_LOOP_and_70_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_69_itm & and_dcpl_100) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_dcpl_102) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_108) | (COMP_LOOP_COMP_LOOP_and_66_itm
      & and_dcpl_110) | (COMP_LOOP_COMP_LOOP_and_65_itm & and_dcpl_116) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_dcpl_119) | (COMP_LOOP_COMP_LOOP_and_185_itm & and_dcpl_125) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_127) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_130);
  assign COMP_LOOP_or_1_nl = ((COMP_LOOP_acc_10_cse_10_1_1_sva[0]) & COMP_LOOP_tmp_nor_13_itm
      & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_70) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_74) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_81) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_72_itm & and_dcpl_93) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_70_itm & and_dcpl_100) | (COMP_LOOP_COMP_LOOP_and_69_itm
      & and_dcpl_102) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_108) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_110) | (COMP_LOOP_COMP_LOOP_and_66_itm & and_dcpl_116) | (COMP_LOOP_COMP_LOOP_and_65_itm
      & and_dcpl_119) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_125) | (COMP_LOOP_COMP_LOOP_and_185_itm
      & and_dcpl_127) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_130);
  assign COMP_LOOP_or_2_nl = ((COMP_LOOP_acc_10_cse_10_1_1_sva[1]) & COMP_LOOP_tmp_nor_14_itm
      & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_70) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_74) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_81) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_93) | (COMP_LOOP_COMP_LOOP_and_72_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_100) | (COMP_LOOP_COMP_LOOP_and_70_itm
      & and_dcpl_102) | (COMP_LOOP_COMP_LOOP_and_69_itm & and_dcpl_108) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_dcpl_110) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_116) | (COMP_LOOP_COMP_LOOP_and_66_itm
      & and_dcpl_119) | (COMP_LOOP_COMP_LOOP_and_65_itm & and_dcpl_125) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_dcpl_127) | (COMP_LOOP_COMP_LOOP_and_185_itm & and_dcpl_130);
  assign COMP_LOOP_or_3_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm & and_dcpl_65)
      | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_70) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_dcpl_74) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_81) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_93) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_72_itm & and_dcpl_100) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_102) | (COMP_LOOP_COMP_LOOP_and_70_itm & and_dcpl_108) | (COMP_LOOP_COMP_LOOP_and_69_itm
      & and_dcpl_110) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_116) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_119) | (COMP_LOOP_COMP_LOOP_and_66_itm & and_dcpl_125) | (COMP_LOOP_COMP_LOOP_and_65_itm
      & and_dcpl_127) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_130);
  assign COMP_LOOP_or_4_nl = ((COMP_LOOP_acc_10_cse_10_1_1_sva[2]) & COMP_LOOP_tmp_nor_16_itm
      & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_185_itm & and_dcpl_70) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_74) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_81) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_93) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_100) | (COMP_LOOP_COMP_LOOP_and_72_itm
      & and_dcpl_102) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_108) | (COMP_LOOP_COMP_LOOP_and_70_itm
      & and_dcpl_110) | (COMP_LOOP_COMP_LOOP_and_69_itm & and_dcpl_116) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_dcpl_119) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_125) | (COMP_LOOP_COMP_LOOP_and_66_itm
      & and_dcpl_127) | (COMP_LOOP_COMP_LOOP_and_65_itm & and_dcpl_130);
  assign COMP_LOOP_or_5_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm & and_dcpl_65)
      | (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_70) | (COMP_LOOP_COMP_LOOP_and_185_itm
      & and_dcpl_74) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_81) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_93) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_100) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_102) | (COMP_LOOP_COMP_LOOP_and_72_itm & and_dcpl_108) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_110) | (COMP_LOOP_COMP_LOOP_and_70_itm & and_dcpl_116) | (COMP_LOOP_COMP_LOOP_and_69_itm
      & and_dcpl_119) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_125) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_127) | (COMP_LOOP_COMP_LOOP_and_66_itm & and_dcpl_130);
  assign COMP_LOOP_or_6_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm & and_dcpl_65)
      | (COMP_LOOP_COMP_LOOP_and_65_itm & and_dcpl_70) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_dcpl_74) | (COMP_LOOP_COMP_LOOP_and_185_itm & and_dcpl_81) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_93) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_100) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_102) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_108) | (COMP_LOOP_COMP_LOOP_and_72_itm
      & and_dcpl_110) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_116) | (COMP_LOOP_COMP_LOOP_and_70_itm
      & and_dcpl_119) | (COMP_LOOP_COMP_LOOP_and_69_itm & and_dcpl_125) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_dcpl_127) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_130);
  assign COMP_LOOP_or_7_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm & and_dcpl_65)
      | (COMP_LOOP_COMP_LOOP_and_66_itm & and_dcpl_70) | (COMP_LOOP_COMP_LOOP_and_65_itm
      & and_dcpl_74) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_81) | (COMP_LOOP_COMP_LOOP_and_185_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_93) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_100) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_102) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_108) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_110) | (COMP_LOOP_COMP_LOOP_and_72_itm & and_dcpl_116) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_119) | (COMP_LOOP_COMP_LOOP_and_70_itm & and_dcpl_125) | (COMP_LOOP_COMP_LOOP_and_69_itm
      & and_dcpl_127) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_130);
  assign COMP_LOOP_or_8_nl = ((COMP_LOOP_acc_10_cse_10_1_1_sva[3]) & COMP_LOOP_tmp_nor_19_itm
      & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_70) | (COMP_LOOP_COMP_LOOP_and_66_itm
      & and_dcpl_74) | (COMP_LOOP_COMP_LOOP_and_65_itm & and_dcpl_81) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_185_itm & and_dcpl_93) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_100) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_102) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_108) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_110) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_116) | (COMP_LOOP_COMP_LOOP_and_72_itm
      & and_dcpl_119) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_125) | (COMP_LOOP_COMP_LOOP_and_70_itm
      & and_dcpl_127) | (COMP_LOOP_COMP_LOOP_and_69_itm & and_dcpl_130);
  assign COMP_LOOP_or_9_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm & and_dcpl_65)
      | (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_70) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_74) | (COMP_LOOP_COMP_LOOP_and_66_itm & and_dcpl_81) | (COMP_LOOP_COMP_LOOP_and_65_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_93) | (COMP_LOOP_COMP_LOOP_and_185_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_100) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_dcpl_102) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_108) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_110) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_116) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_119) | (COMP_LOOP_COMP_LOOP_and_72_itm & and_dcpl_125) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_127) | (COMP_LOOP_COMP_LOOP_and_70_itm & and_dcpl_130);
  assign COMP_LOOP_or_10_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm & and_dcpl_65)
      | (COMP_LOOP_COMP_LOOP_and_69_itm & and_dcpl_70) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_dcpl_74) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_81) | (COMP_LOOP_COMP_LOOP_and_66_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_65_itm & and_dcpl_93) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_185_itm & and_dcpl_100) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_102) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_108) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_110) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_116) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_119) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_125) | (COMP_LOOP_COMP_LOOP_and_72_itm
      & and_dcpl_127) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_130);
  assign COMP_LOOP_or_11_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm & and_dcpl_65)
      | (COMP_LOOP_COMP_LOOP_and_70_itm & and_dcpl_70) | (COMP_LOOP_COMP_LOOP_and_69_itm
      & and_dcpl_74) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_81) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_66_itm & and_dcpl_93) | (COMP_LOOP_COMP_LOOP_and_65_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_100) | (COMP_LOOP_COMP_LOOP_and_185_itm
      & and_dcpl_102) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_108) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_dcpl_110) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_116) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_119) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_125) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_127) | (COMP_LOOP_COMP_LOOP_and_72_itm & and_dcpl_130);
  assign COMP_LOOP_or_12_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm & and_dcpl_65)
      | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_70) | (COMP_LOOP_COMP_LOOP_and_70_itm
      & and_dcpl_74) | (COMP_LOOP_COMP_LOOP_and_69_itm & and_dcpl_81) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_93) | (COMP_LOOP_COMP_LOOP_and_66_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_65_itm & and_dcpl_100) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_dcpl_102) | (COMP_LOOP_COMP_LOOP_and_185_itm & and_dcpl_108) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_110) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_116) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_119) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_125) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_127) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_130);
  assign COMP_LOOP_or_13_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm & and_dcpl_65)
      | (COMP_LOOP_COMP_LOOP_and_72_itm & and_dcpl_70) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_74) | (COMP_LOOP_COMP_LOOP_and_70_itm & and_dcpl_81) | (COMP_LOOP_COMP_LOOP_and_69_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_93) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_66_itm & and_dcpl_100) | (COMP_LOOP_COMP_LOOP_and_65_itm
      & and_dcpl_102) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_108) | (COMP_LOOP_COMP_LOOP_and_185_itm
      & and_dcpl_110) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_116) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_dcpl_119) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_125) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_127) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_130);
  assign COMP_LOOP_or_14_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm & and_dcpl_65)
      | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_70) | (COMP_LOOP_COMP_LOOP_and_72_itm
      & and_dcpl_74) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_81) | (COMP_LOOP_COMP_LOOP_and_70_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_69_itm & and_dcpl_93) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_100) | (COMP_LOOP_COMP_LOOP_and_66_itm
      & and_dcpl_102) | (COMP_LOOP_COMP_LOOP_and_65_itm & and_dcpl_108) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_dcpl_110) | (COMP_LOOP_COMP_LOOP_and_185_itm & and_dcpl_116) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_119) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_125) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_127) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_130);
  assign COMP_LOOP_or_15_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm & and_dcpl_65)
      | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_70) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_74) | (COMP_LOOP_COMP_LOOP_and_72_itm & and_dcpl_81) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_70_itm & and_dcpl_93) | (COMP_LOOP_COMP_LOOP_and_69_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_100) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_102) | (COMP_LOOP_COMP_LOOP_and_66_itm & and_dcpl_108) | (COMP_LOOP_COMP_LOOP_and_65_itm
      & and_dcpl_110) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_116) | (COMP_LOOP_COMP_LOOP_and_185_itm
      & and_dcpl_119) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_125) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_dcpl_127) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_130);
  assign COMP_LOOP_or_21_nl = and_dcpl_189 | and_dcpl_220 | and_dcpl_222 | and_dcpl_223
      | and_dcpl_225 | and_dcpl_226 | and_dcpl_227 | and_dcpl_228 | and_dcpl_229
      | and_dcpl_230 | and_dcpl_231 | and_dcpl_232 | and_dcpl_233 | and_dcpl_234
      | and_dcpl_235 | and_dcpl_236;
  assign COMP_LOOP_or_22_nl = COMP_LOOP_10_acc_8_itm_mx0c2 | COMP_LOOP_10_acc_8_itm_mx0c6
      | COMP_LOOP_10_acc_8_itm_mx0c9 | COMP_LOOP_10_acc_8_itm_mx0c12 | COMP_LOOP_10_acc_8_itm_mx0c15
      | COMP_LOOP_10_acc_8_itm_mx0c18 | COMP_LOOP_10_acc_8_itm_mx0c21 | COMP_LOOP_10_acc_8_itm_mx0c24
      | COMP_LOOP_10_acc_8_itm_mx0c27 | COMP_LOOP_10_acc_8_itm_mx0c30 | COMP_LOOP_10_acc_8_itm_mx0c33
      | COMP_LOOP_10_acc_8_itm_mx0c36 | COMP_LOOP_10_acc_8_itm_mx0c39 | COMP_LOOP_10_acc_8_itm_mx0c42
      | COMP_LOOP_10_acc_8_itm_mx0c47;
  assign COMP_LOOP_tmp_and_42_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_nor_itm & (~ and_332_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_nl = (COMP_LOOP_10_tmp_mul_idiv_sva[0])
      & COMP_LOOP_tmp_nor_itm & (~ and_332_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_1_nl = (COMP_LOOP_10_tmp_mul_idiv_sva[1])
      & COMP_LOOP_tmp_nor_1_itm & (~ and_332_tmp);
  assign COMP_LOOP_tmp_and_43_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_itm & (~ and_332_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl = (COMP_LOOP_10_tmp_mul_idiv_sva[2])
      & COMP_LOOP_tmp_nor_3_itm & (~ and_332_tmp);
  assign COMP_LOOP_tmp_and_44_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_itm & (~ and_332_tmp);
  assign COMP_LOOP_tmp_and_45_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_itm & (~ and_332_tmp);
  assign COMP_LOOP_tmp_and_46_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_itm & (~ and_332_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_7_nl = (COMP_LOOP_10_tmp_mul_idiv_sva[3])
      & COMP_LOOP_tmp_nor_6_itm & (~ and_332_tmp);
  assign COMP_LOOP_tmp_and_47_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_itm & (~ and_332_tmp);
  assign COMP_LOOP_tmp_and_48_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_itm & (~ and_332_tmp);
  assign COMP_LOOP_tmp_and_49_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_itm & (~ and_332_tmp);
  assign COMP_LOOP_tmp_and_50_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_itm & (~ and_332_tmp);
  assign COMP_LOOP_tmp_and_51_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_itm & (~ and_332_tmp);
  assign COMP_LOOP_tmp_and_52_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_itm & (~ and_332_tmp);
  assign COMP_LOOP_tmp_and_53_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_itm & (~ and_332_tmp);
  assign and_336_nl = and_dcpl_5 & ((fsm_output[2]) ^ (fsm_output[3])) & (fsm_output[1:0]==2'b00)
      & and_dcpl_45;
  assign and_340_nl = and_dcpl_61 & (~ (COMP_LOOP_9_tmp_lshift_itm[0])) & (fsm_output[3])
      & (fsm_output[0]) & and_dcpl_45;
  assign or_2595_nl = nor_572_cse | (fsm_output[8]);
  assign mux_2501_nl = MUX_s_1_2_2(mux_tmp_439, or_2595_nl, fsm_output[1]);
  assign mux_2502_nl = MUX_s_1_2_2(mux_2501_nl, (fsm_output[8]), fsm_output[2]);
  assign mux_2503_nl = MUX_s_1_2_2(mux_tmp_439, mux_2502_nl, fsm_output[3]);
  assign or_2593_nl = (~((fsm_output[2]) | (fsm_output[6]) | (fsm_output[7]))) |
      (fsm_output[8]);
  assign or_2591_nl = (~((fsm_output[2]) | (fsm_output[1]) | (fsm_output[6]) | (fsm_output[7])))
      | (fsm_output[8]);
  assign mux_2499_nl = MUX_s_1_2_2(or_2593_nl, or_2591_nl, COMP_LOOP_9_tmp_lshift_itm[0]);
  assign mux_2500_nl = MUX_s_1_2_2(mux_tmp_439, mux_2499_nl, fsm_output[3]);
  assign mux_2504_nl = MUX_s_1_2_2(mux_2503_nl, mux_2500_nl, fsm_output[0]);
  assign COMP_LOOP_tmp_and_36_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_itm & (~ and_341_tmp);
  assign COMP_LOOP_tmp_and_37_nl = COMP_LOOP_tmp_or_29_cse & (~ and_341_tmp);
  assign COMP_LOOP_tmp_and_38_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm & (~ and_341_tmp);
  assign COMP_LOOP_tmp_and_39_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm & (~ and_341_tmp);
  assign COMP_LOOP_tmp_and_40_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm & (~ and_341_tmp);
  assign COMP_LOOP_tmp_and_41_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm & (~ and_341_tmp);
  assign COMP_LOOP_tmp_and_20_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_nor_12_itm & (~ and_342_tmp);
  assign COMP_LOOP_tmp_and_21_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_167 & (~ and_342_tmp);
  assign COMP_LOOP_tmp_and_22_nl = and_1191_cse & (~ and_342_tmp);
  assign COMP_LOOP_tmp_and_23_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm & (~ and_342_tmp);
  assign COMP_LOOP_tmp_and_24_nl = and_1190_cse & (~ and_342_tmp);
  assign COMP_LOOP_tmp_and_25_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm & (~ and_342_tmp);
  assign COMP_LOOP_tmp_and_26_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm & (~ and_342_tmp);
  assign COMP_LOOP_tmp_and_27_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm & (~ and_342_tmp);
  assign COMP_LOOP_tmp_and_28_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_161 & (~ and_342_tmp);
  assign COMP_LOOP_tmp_and_29_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm & (~ and_342_tmp);
  assign COMP_LOOP_tmp_and_30_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm & (~ and_342_tmp);
  assign COMP_LOOP_tmp_and_31_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm & (~ and_342_tmp);
  assign COMP_LOOP_tmp_and_32_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm & (~ and_342_tmp);
  assign COMP_LOOP_tmp_and_33_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm & (~ and_342_tmp);
  assign COMP_LOOP_tmp_and_34_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm & (~ and_342_tmp);
  assign COMP_LOOP_tmp_and_35_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm & (~ and_342_tmp);
  assign COMP_LOOP_tmp_and_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_nor_14_cse & and_dcpl_198;
  assign COMP_LOOP_tmp_and_17_nl = (COMP_LOOP_13_tmp_mul_idiv_sva[1:0]==2'b10) &
      and_dcpl_198;
  assign COMP_LOOP_tmp_and_18_nl = (COMP_LOOP_13_tmp_mul_idiv_sva[1:0]==2'b11) &
      and_dcpl_198;
  assign mux_2515_nl = MUX_s_1_2_2(mux_tmp_2392, mux_559_cse, and_674_cse);
  assign mux_2516_nl = MUX_s_1_2_2(mux_2515_nl, mux_559_cse, fsm_output[3]);
  assign mux_2514_nl = MUX_s_1_2_2(mux_tmp_2392, mux_559_cse, or_2259_cse_1);
  assign mux_2517_nl = MUX_s_1_2_2(mux_2516_nl, mux_2514_nl, fsm_output[0]);
  assign mux_2518_nl = MUX_s_1_2_2(mux_2517_nl, and_733_cse, or_2589_cse);
  assign mux_2519_nl = MUX_s_1_2_2(mux_tmp_2392, and_dcpl_57, or_2612_cse);
  assign mux_2520_nl = MUX_s_1_2_2(mux_tmp_2392, mux_2519_nl, fsm_output[4]);
  assign and_357_nl = ((fsm_output[4]) | (fsm_output[3]) | (fsm_output[2]) | (fsm_output[6]))
      & (fsm_output[8:7]==2'b11);
  assign mux_2528_nl = MUX_s_1_2_2(mux_228_cse, nor_tmp_47, or_432_cse);
  assign mux_2529_nl = MUX_s_1_2_2(mux_228_cse, mux_2528_nl, fsm_output[3]);
  assign mux_2527_nl = MUX_s_1_2_2(mux_228_cse, nor_tmp_47, fsm_output[3]);
  assign mux_2530_nl = MUX_s_1_2_2(mux_2529_nl, mux_2527_nl, fsm_output[0]);
  assign mux_2531_nl = MUX_s_1_2_2(mux_2530_nl, nor_tmp_47, fsm_output[4]);
  assign mux_2526_nl = MUX_s_1_2_2(nor_tmp_489, (fsm_output[7]), fsm_output[4]);
  assign mux_2532_nl = MUX_s_1_2_2(mux_2531_nl, mux_2526_nl, fsm_output[5]);
  assign COMP_LOOP_tmp_and_7_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_nor_12_itm & (~ nor_1796_tmp);
  assign COMP_LOOP_tmp_and_8_nl = COMP_LOOP_tmp_or_29_cse & (~ nor_1796_tmp);
  assign COMP_LOOP_tmp_and_9_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm & (~ nor_1796_tmp);
  assign COMP_LOOP_tmp_and_10_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm & (~ nor_1796_tmp);
  assign COMP_LOOP_tmp_and_11_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm & (~ nor_1796_tmp);
  assign COMP_LOOP_tmp_and_12_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm & (~ nor_1796_tmp);
  assign mux_2540_nl = MUX_s_1_2_2(or_2732_cse, or_2729_cse, fsm_output[3]);
  assign mux_2541_nl = MUX_s_1_2_2(or_2621_cse, mux_2540_nl, fsm_output[0]);
  assign nor_568_nl = ~((fsm_output[4]) | mux_2541_nl);
  assign mux_2539_nl = MUX_s_1_2_2(and_tmp_28, nor_tmp_47, fsm_output[4]);
  assign mux_2542_nl = MUX_s_1_2_2(nor_568_nl, mux_2539_nl, fsm_output[5]);
  assign mux_2544_nl = MUX_s_1_2_2(mux_tmp_439, nor_tmp_115, and_831_cse);
  assign mux_2543_nl = MUX_s_1_2_2(mux_tmp_439, nor_tmp_115, and_570_cse);
  assign mux_2545_nl = MUX_s_1_2_2(mux_2544_nl, mux_2543_nl, fsm_output[0]);
  assign mux_2546_nl = MUX_s_1_2_2(mux_2545_nl, nor_tmp_115, fsm_output[4]);
  assign and_352_nl = ((fsm_output[4]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[7]))
      & (fsm_output[8]);
  assign COMP_LOOP_tmp_and_2_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_nor_12_itm & and_dcpl_202;
  assign COMP_LOOP_tmp_and_3_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm & and_dcpl_202;
  assign COMP_LOOP_tmp_and_4_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm & and_dcpl_202;
  assign COMP_LOOP_tmp_and_5_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm & and_dcpl_202;
  assign COMP_LOOP_tmp_and_6_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm & and_dcpl_202;
  assign mux_2551_nl = MUX_s_1_2_2(mux_559_cse, mux_tmp_538, fsm_output[3]);
  assign mux_560_nl = MUX_s_1_2_2(mux_559_cse, mux_tmp_439, and_674_cse);
  assign mux_561_nl = MUX_s_1_2_2(mux_560_nl, mux_tmp_538, fsm_output[3]);
  assign mux_2552_nl = MUX_s_1_2_2(mux_2551_nl, mux_561_nl, fsm_output[0]);
  assign mux_2553_nl = MUX_s_1_2_2(mux_2552_nl, nor_tmp_115, or_2589_cse);
  assign mux_2555_nl = MUX_s_1_2_2(mux_464_cse, and_733_cse, or_2626_cse);
  assign mux_2556_nl = MUX_s_1_2_2(mux_2555_nl, and_733_cse, fsm_output[4]);
  assign or_2625_nl = (fsm_output[4:3]!=2'b00);
  assign mux_2554_nl = MUX_s_1_2_2(and_655_cse, nor_tmp_115, or_2625_nl);
  assign COMP_LOOP_mux_358_nl = MUX_v_11_2_2(({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))}),
      STAGE_LOOP_lshift_psp_sva, and_dcpl_356);
  assign COMP_LOOP_COMP_LOOP_nand_1_nl = ~(and_dcpl_356 & (~((fsm_output[8:6]==3'b000)
      & nor_1624_cse & (fsm_output[1:0]==2'b10) & and_dcpl_45)));
  assign COMP_LOOP_mux_359_nl = MUX_v_10_2_2(({COMP_LOOP_k_10_4_sva_5_0 , 4'b0001}),
      VEC_LOOP_j_10_0_sva_9_0, and_dcpl_356);
  assign nl_acc_nl = ({COMP_LOOP_mux_358_nl , COMP_LOOP_COMP_LOOP_nand_1_nl}) + conv_u2u_11_12({COMP_LOOP_mux_359_nl
      , 1'b1});
  assign acc_nl = nl_acc_nl[11:0];
  assign z_out_2 = readslicef_12_11_1(acc_nl);
  assign COMP_LOOP_mux1h_710_nl = MUX1HOT_v_54_15_2((COMP_LOOP_tmp_mux1h_12_itm[63:10]),
      (COMP_LOOP_tmp_mux1h_itm[63:10]), (COMP_LOOP_tmp_mux1h_1_itm[63:10]), (COMP_LOOP_tmp_mux1h_2_itm[63:10]),
      (COMP_LOOP_tmp_mux1h_3_itm[63:10]), (COMP_LOOP_tmp_mux1h_4_itm[63:10]), (COMP_LOOP_tmp_mux1h_5_itm[63:10]),
      (COMP_LOOP_tmp_mux1h_6_itm[63:10]), (COMP_LOOP_tmp_mux_itm[63:10]), (COMP_LOOP_tmp_mux1h_7_itm[63:10]),
      (COMP_LOOP_tmp_mux1h_8_itm[63:10]), (COMP_LOOP_tmp_mux1h_9_itm[63:10]), (tmp_36_sva_1[63:10]),
      (tmp_36_sva_2[63:10]), (tmp_33_sva_1[63:10]), {and_dcpl_360 , and_dcpl_367
      , and_dcpl_374 , and_dcpl_378 , and_dcpl_384 , and_dcpl_386 , and_dcpl_390
      , and_dcpl_391 , and_dcpl_395 , and_dcpl_396 , and_dcpl_400 , and_dcpl_401
      , and_dcpl_405 , and_dcpl_406 , and_dcpl_409});
  assign COMP_LOOP_and_260_nl = MUX_v_54_2_2(54'b000000000000000000000000000000000000000000000000000000,
      COMP_LOOP_mux1h_710_nl, COMP_LOOP_nor_itm);
  assign COMP_LOOP_mux1h_711_nl = MUX1HOT_s_1_17_2((COMP_LOOP_tmp_mux1h_12_itm[9]),
      (COMP_LOOP_tmp_mux1h_itm[9]), (COMP_LOOP_tmp_mux1h_1_itm[9]), (COMP_LOOP_tmp_mux1h_2_itm[9]),
      (COMP_LOOP_tmp_mux1h_3_itm[9]), (COMP_LOOP_tmp_mux1h_4_itm[9]), (COMP_LOOP_tmp_mux1h_5_itm[9]),
      (COMP_LOOP_tmp_mux1h_6_itm[9]), (COMP_LOOP_tmp_mux_itm[9]), (COMP_LOOP_tmp_mux1h_7_itm[9]),
      (COMP_LOOP_tmp_mux1h_8_itm[9]), (COMP_LOOP_tmp_mux1h_9_itm[9]), (tmp_36_sva_1[9]),
      (tmp_36_sva_2[9]), (tmp_33_sva_1[9]), (z_out_1[9]), (COMP_LOOP_2_tmp_lshift_ncse_sva[9]),
      {and_dcpl_360 , and_dcpl_367 , and_dcpl_374 , and_dcpl_378 , and_dcpl_384 ,
      and_dcpl_386 , and_dcpl_390 , and_dcpl_391 , and_dcpl_395 , and_dcpl_396 ,
      and_dcpl_400 , and_dcpl_401 , and_dcpl_405 , and_dcpl_406 , and_dcpl_409 ,
      and_dcpl_411 , COMP_LOOP_or_40_itm});
  assign COMP_LOOP_and_261_nl = COMP_LOOP_mux1h_711_nl & COMP_LOOP_nor_621_itm;
  assign COMP_LOOP_mux1h_712_nl = MUX1HOT_s_1_18_2((COMP_LOOP_tmp_mux1h_12_itm[8]),
      (COMP_LOOP_tmp_mux1h_itm[8]), (COMP_LOOP_tmp_mux1h_1_itm[8]), (COMP_LOOP_tmp_mux1h_2_itm[8]),
      (COMP_LOOP_tmp_mux1h_3_itm[8]), (COMP_LOOP_tmp_mux1h_4_itm[8]), (COMP_LOOP_tmp_mux1h_5_itm[8]),
      (COMP_LOOP_tmp_mux1h_6_itm[8]), (COMP_LOOP_tmp_mux_itm[8]), (COMP_LOOP_tmp_mux1h_7_itm[8]),
      (COMP_LOOP_tmp_mux1h_8_itm[8]), (COMP_LOOP_tmp_mux1h_9_itm[8]), (tmp_36_sva_1[8]),
      (tmp_36_sva_2[8]), (tmp_33_sva_1[8]), (z_out_1[8]), (COMP_LOOP_2_tmp_lshift_ncse_sva[8]),
      (COMP_LOOP_3_tmp_lshift_ncse_sva[8]), {and_dcpl_360 , and_dcpl_367 , and_dcpl_374
      , and_dcpl_378 , and_dcpl_384 , and_dcpl_386 , and_dcpl_390 , and_dcpl_391
      , and_dcpl_395 , and_dcpl_396 , and_dcpl_400 , and_dcpl_401 , and_dcpl_405
      , and_dcpl_406 , and_dcpl_409 , COMP_LOOP_or_41_itm , COMP_LOOP_or_40_itm ,
      COMP_LOOP_or_43_itm});
  assign COMP_LOOP_and_262_nl = COMP_LOOP_mux1h_712_nl & COMP_LOOP_nor_622_itm;
  assign COMP_LOOP_mux1h_713_nl = MUX1HOT_v_8_20_2((COMP_LOOP_tmp_mux1h_12_itm[7:0]),
      (COMP_LOOP_tmp_mux1h_itm[7:0]), (COMP_LOOP_tmp_mux1h_1_itm[7:0]), (COMP_LOOP_tmp_mux1h_2_itm[7:0]),
      (COMP_LOOP_tmp_mux1h_3_itm[7:0]), (COMP_LOOP_tmp_mux1h_4_itm[7:0]), (COMP_LOOP_tmp_mux1h_5_itm[7:0]),
      (COMP_LOOP_tmp_mux1h_6_itm[7:0]), (COMP_LOOP_tmp_mux_itm[7:0]), (COMP_LOOP_tmp_mux1h_7_itm[7:0]),
      (COMP_LOOP_tmp_mux1h_8_itm[7:0]), (COMP_LOOP_tmp_mux1h_9_itm[7:0]), (tmp_36_sva_1[7:0]),
      (tmp_36_sva_2[7:0]), (tmp_33_sva_1[7:0]), (z_out_1[7:0]), ({1'b0 , COMP_LOOP_9_tmp_lshift_itm}),
      (COMP_LOOP_2_tmp_lshift_ncse_sva[7:0]), (COMP_LOOP_3_tmp_lshift_ncse_sva[7:0]),
      COMP_LOOP_13_tmp_mul_idiv_sva, {and_dcpl_360 , and_dcpl_367 , and_dcpl_374
      , and_dcpl_378 , and_dcpl_384 , and_dcpl_386 , and_dcpl_390 , and_dcpl_391
      , and_dcpl_395 , and_dcpl_396 , and_dcpl_400 , and_dcpl_401 , and_dcpl_405
      , and_dcpl_406 , and_dcpl_409 , COMP_LOOP_or_41_itm , and_dcpl_413 , COMP_LOOP_or_40_itm
      , COMP_LOOP_or_43_itm , COMP_LOOP_or_47_itm});
  assign COMP_LOOP_COMP_LOOP_and_983_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[63])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_984_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[62])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_985_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[61])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_986_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[60])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_987_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[59])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_988_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[58])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_989_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[57])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_990_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[56])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_991_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[55])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_992_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[54])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_993_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[53])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_994_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[52])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_995_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[51])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_996_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[50])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_997_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[49])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_998_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[48])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_999_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[47])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1000_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[46])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1001_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[45])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1002_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[44])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1003_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[43])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1004_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[42])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1005_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[41])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1006_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[40])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1007_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[39])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1008_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[38])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1009_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[37])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1010_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[36])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1011_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[35])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1012_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[34])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1013_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[33])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1014_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[32])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1015_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[31])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1016_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[30])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1017_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[29])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1018_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[28])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1019_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[27])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1020_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[26])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1021_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[25])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1022_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[24])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1023_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[23])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1024_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[22])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1025_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[21])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1026_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[20])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1027_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[19])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1028_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[18])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1029_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[17])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1030_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[16])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1031_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[15])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1032_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[14])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1033_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[13])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1034_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[12])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1035_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[11])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_and_1036_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[10])
      & COMP_LOOP_nor_itm;
  assign COMP_LOOP_COMP_LOOP_mux_8_nl = MUX_s_1_2_2((COMP_LOOP_1_modulo_cmp_return_rsc_z[9]),
      (COMP_LOOP_k_10_4_sva_5_0[5]), COMP_LOOP_or_52_itm);
  assign COMP_LOOP_and_263_nl = COMP_LOOP_COMP_LOOP_mux_8_nl & COMP_LOOP_nor_621_itm;
  assign COMP_LOOP_mux1h_714_nl = MUX1HOT_s_1_3_2((COMP_LOOP_1_modulo_cmp_return_rsc_z[8]),
      (COMP_LOOP_k_10_4_sva_5_0[4]), (COMP_LOOP_k_10_4_sva_5_0[5]), {COMP_LOOP_or_17_ssc
      , COMP_LOOP_or_52_itm , COMP_LOOP_or_54_itm});
  assign COMP_LOOP_and_264_nl = COMP_LOOP_mux1h_714_nl & COMP_LOOP_nor_622_itm;
  assign COMP_LOOP_mux1h_715_nl = MUX1HOT_v_4_5_2((COMP_LOOP_1_modulo_cmp_return_rsc_z[7:4]),
      (COMP_LOOP_k_10_4_sva_5_0[3:0]), ({1'b0 , (COMP_LOOP_k_10_4_sva_5_0[5:3])}),
      (COMP_LOOP_k_10_4_sva_5_0[4:1]), (COMP_LOOP_k_10_4_sva_5_0[5:2]), {COMP_LOOP_or_17_ssc
      , COMP_LOOP_or_52_itm , and_dcpl_413 , COMP_LOOP_or_54_itm , COMP_LOOP_or_47_itm});
  assign COMP_LOOP_mux1h_716_nl = MUX1HOT_s_1_4_2((COMP_LOOP_1_modulo_cmp_return_rsc_z[3]),
      (COMP_LOOP_k_10_4_sva_5_0[2]), (COMP_LOOP_k_10_4_sva_5_0[0]), (COMP_LOOP_k_10_4_sva_5_0[1]),
      {COMP_LOOP_or_17_ssc , and_dcpl_413 , COMP_LOOP_or_54_itm , COMP_LOOP_or_47_itm});
  assign COMP_LOOP_or_61_nl = (COMP_LOOP_mux1h_716_nl & (~(and_dcpl_411 | and_dcpl_416
      | and_dcpl_417 | and_dcpl_418))) | and_dcpl_419 | and_dcpl_421 | and_dcpl_422
      | and_dcpl_425;
  assign COMP_LOOP_mux1h_717_nl = MUX1HOT_s_1_3_2((COMP_LOOP_1_modulo_cmp_return_rsc_z[2]),
      (COMP_LOOP_k_10_4_sva_5_0[1]), (COMP_LOOP_k_10_4_sva_5_0[0]), {COMP_LOOP_or_17_ssc
      , and_dcpl_413 , COMP_LOOP_or_47_itm});
  assign COMP_LOOP_or_62_nl = (COMP_LOOP_mux1h_717_nl & (~(and_dcpl_411 | and_dcpl_416
      | and_dcpl_419 | and_dcpl_421 | and_dcpl_426 | and_dcpl_427))) | and_dcpl_417
      | and_dcpl_418 | and_dcpl_422 | and_dcpl_425 | and_dcpl_428 | and_dcpl_429;
  assign COMP_LOOP_mux_360_nl = MUX_s_1_2_2((COMP_LOOP_1_modulo_cmp_return_rsc_z[1]),
      (COMP_LOOP_k_10_4_sva_5_0[0]), and_dcpl_413);
  assign COMP_LOOP_COMP_LOOP_or_2_nl = (COMP_LOOP_mux_360_nl & (~(and_dcpl_411 |
      and_dcpl_417 | and_dcpl_419 | and_dcpl_422 | and_dcpl_426 | and_dcpl_428 |
      and_dcpl_431))) | and_dcpl_416 | and_dcpl_418 | and_dcpl_421 | and_dcpl_425
      | and_dcpl_427 | and_dcpl_429 | and_dcpl_430;
  assign COMP_LOOP_COMP_LOOP_or_3_nl = (COMP_LOOP_1_modulo_cmp_return_rsc_z[0]) |
      and_dcpl_411 | and_dcpl_416 | and_dcpl_417 | and_dcpl_418 | and_dcpl_419 |
      and_dcpl_421 | and_dcpl_422 | and_dcpl_425 | and_dcpl_426 | and_dcpl_427 |
      and_dcpl_428 | and_dcpl_429 | and_dcpl_430 | and_dcpl_431 | and_dcpl_413;
  assign nl_z_out_3 = ({COMP_LOOP_and_260_nl , COMP_LOOP_and_261_nl , COMP_LOOP_and_262_nl
      , COMP_LOOP_mux1h_713_nl}) * ({COMP_LOOP_COMP_LOOP_and_983_nl , COMP_LOOP_COMP_LOOP_and_984_nl
      , COMP_LOOP_COMP_LOOP_and_985_nl , COMP_LOOP_COMP_LOOP_and_986_nl , COMP_LOOP_COMP_LOOP_and_987_nl
      , COMP_LOOP_COMP_LOOP_and_988_nl , COMP_LOOP_COMP_LOOP_and_989_nl , COMP_LOOP_COMP_LOOP_and_990_nl
      , COMP_LOOP_COMP_LOOP_and_991_nl , COMP_LOOP_COMP_LOOP_and_992_nl , COMP_LOOP_COMP_LOOP_and_993_nl
      , COMP_LOOP_COMP_LOOP_and_994_nl , COMP_LOOP_COMP_LOOP_and_995_nl , COMP_LOOP_COMP_LOOP_and_996_nl
      , COMP_LOOP_COMP_LOOP_and_997_nl , COMP_LOOP_COMP_LOOP_and_998_nl , COMP_LOOP_COMP_LOOP_and_999_nl
      , COMP_LOOP_COMP_LOOP_and_1000_nl , COMP_LOOP_COMP_LOOP_and_1001_nl , COMP_LOOP_COMP_LOOP_and_1002_nl
      , COMP_LOOP_COMP_LOOP_and_1003_nl , COMP_LOOP_COMP_LOOP_and_1004_nl , COMP_LOOP_COMP_LOOP_and_1005_nl
      , COMP_LOOP_COMP_LOOP_and_1006_nl , COMP_LOOP_COMP_LOOP_and_1007_nl , COMP_LOOP_COMP_LOOP_and_1008_nl
      , COMP_LOOP_COMP_LOOP_and_1009_nl , COMP_LOOP_COMP_LOOP_and_1010_nl , COMP_LOOP_COMP_LOOP_and_1011_nl
      , COMP_LOOP_COMP_LOOP_and_1012_nl , COMP_LOOP_COMP_LOOP_and_1013_nl , COMP_LOOP_COMP_LOOP_and_1014_nl
      , COMP_LOOP_COMP_LOOP_and_1015_nl , COMP_LOOP_COMP_LOOP_and_1016_nl , COMP_LOOP_COMP_LOOP_and_1017_nl
      , COMP_LOOP_COMP_LOOP_and_1018_nl , COMP_LOOP_COMP_LOOP_and_1019_nl , COMP_LOOP_COMP_LOOP_and_1020_nl
      , COMP_LOOP_COMP_LOOP_and_1021_nl , COMP_LOOP_COMP_LOOP_and_1022_nl , COMP_LOOP_COMP_LOOP_and_1023_nl
      , COMP_LOOP_COMP_LOOP_and_1024_nl , COMP_LOOP_COMP_LOOP_and_1025_nl , COMP_LOOP_COMP_LOOP_and_1026_nl
      , COMP_LOOP_COMP_LOOP_and_1027_nl , COMP_LOOP_COMP_LOOP_and_1028_nl , COMP_LOOP_COMP_LOOP_and_1029_nl
      , COMP_LOOP_COMP_LOOP_and_1030_nl , COMP_LOOP_COMP_LOOP_and_1031_nl , COMP_LOOP_COMP_LOOP_and_1032_nl
      , COMP_LOOP_COMP_LOOP_and_1033_nl , COMP_LOOP_COMP_LOOP_and_1034_nl , COMP_LOOP_COMP_LOOP_and_1035_nl
      , COMP_LOOP_COMP_LOOP_and_1036_nl , COMP_LOOP_and_263_nl , COMP_LOOP_and_264_nl
      , COMP_LOOP_mux1h_715_nl , COMP_LOOP_or_61_nl , COMP_LOOP_or_62_nl , COMP_LOOP_COMP_LOOP_or_2_nl
      , COMP_LOOP_COMP_LOOP_or_3_nl});
  assign z_out_3 = nl_z_out_3[63:0];
  assign STAGE_LOOP_mux_4_nl = MUX_v_4_2_2(STAGE_LOOP_i_3_0_sva, (~ STAGE_LOOP_i_3_0_sva),
      and_dcpl_447);
  assign nl_z_out_4 = STAGE_LOOP_mux_4_nl + ({1'b1 , (~ and_dcpl_447) , 2'b11});
  assign z_out_4 = nl_z_out_4[3:0];
  assign COMP_LOOP_mux_361_cse = MUX_v_64_2_2(z_out_7, COMP_LOOP_10_acc_8_itm, COMP_LOOP_or_18_itm);
  assign COMP_LOOP_mux1h_718_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_nor_itm, COMP_LOOP_COMP_LOOP_nor_5_itm,
      COMP_LOOP_COMP_LOOP_nor_9_itm, COMP_LOOP_COMP_LOOP_nor_13_itm, COMP_LOOP_COMP_LOOP_nor_17_itm,
      COMP_LOOP_COMP_LOOP_nor_21_itm, COMP_LOOP_COMP_LOOP_nor_25_itm, COMP_LOOP_COMP_LOOP_nor_29_itm,
      COMP_LOOP_COMP_LOOP_nor_33_itm, COMP_LOOP_COMP_LOOP_nor_37_itm, COMP_LOOP_COMP_LOOP_nor_41_itm,
      COMP_LOOP_COMP_LOOP_nor_45_itm, COMP_LOOP_COMP_LOOP_nor_49_itm, COMP_LOOP_COMP_LOOP_nor_53_itm,
      COMP_LOOP_COMP_LOOP_nor_57_itm, COMP_LOOP_COMP_LOOP_nor_61_itm, {and_dcpl_571
      , and_dcpl_577 , and_1025_cse , and_1028_cse , and_dcpl_589 , and_1037_cse
      , and_1040_cse , and_1044_cse , and_1046_cse , and_1051_cse , and_1052_cse
      , and_1055_cse , and_1056_cse , and_1060_cse , and_1061_cse , and_1064_cse});
  assign COMP_LOOP_COMP_LOOP_and_1037_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[0]) &
      COMP_LOOP_nor_51_itm;
  assign COMP_LOOP_COMP_LOOP_and_1038_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[0]) &
      COMP_LOOP_nor_91_itm;
  assign COMP_LOOP_COMP_LOOP_and_1039_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[0]) &
      COMP_LOOP_nor_131_itm;
  assign COMP_LOOP_COMP_LOOP_and_1040_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[0]) &
      COMP_LOOP_nor_171_itm;
  assign COMP_LOOP_COMP_LOOP_and_1041_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[0]) &
      COMP_LOOP_nor_211_itm;
  assign COMP_LOOP_COMP_LOOP_and_1042_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) &
      COMP_LOOP_nor_251_itm;
  assign COMP_LOOP_COMP_LOOP_and_1043_nl = (COMP_LOOP_acc_10_cse_10_1_8_sva[0]) &
      COMP_LOOP_nor_291_itm;
  assign COMP_LOOP_COMP_LOOP_and_1044_nl = (COMP_LOOP_acc_10_cse_10_1_9_sva[0]) &
      COMP_LOOP_nor_331_itm;
  assign COMP_LOOP_COMP_LOOP_and_1045_nl = (COMP_LOOP_acc_10_cse_10_1_10_sva[0])
      & COMP_LOOP_nor_371_itm;
  assign COMP_LOOP_COMP_LOOP_and_1046_nl = (COMP_LOOP_acc_10_cse_10_1_11_sva[0])
      & COMP_LOOP_nor_411_itm;
  assign COMP_LOOP_COMP_LOOP_and_1047_nl = (COMP_LOOP_acc_10_cse_10_1_12_sva[0])
      & COMP_LOOP_nor_451_itm;
  assign COMP_LOOP_COMP_LOOP_and_1048_nl = (COMP_LOOP_acc_10_cse_10_1_13_sva[0])
      & COMP_LOOP_nor_491_itm;
  assign COMP_LOOP_COMP_LOOP_and_1049_nl = (COMP_LOOP_acc_10_cse_10_1_14_sva[0])
      & COMP_LOOP_nor_531_itm;
  assign COMP_LOOP_COMP_LOOP_and_1050_nl = (COMP_LOOP_acc_10_cse_10_1_15_sva[0])
      & COMP_LOOP_nor_571_itm;
  assign COMP_LOOP_COMP_LOOP_and_1051_nl = (COMP_LOOP_acc_10_cse_10_1_sva[0]) & COMP_LOOP_nor_611_itm;
  assign COMP_LOOP_mux1h_719_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_244_itm,
      COMP_LOOP_COMP_LOOP_and_1037_nl, COMP_LOOP_COMP_LOOP_and_1038_nl, COMP_LOOP_COMP_LOOP_and_1039_nl,
      COMP_LOOP_COMP_LOOP_and_1040_nl, COMP_LOOP_COMP_LOOP_and_1041_nl, COMP_LOOP_COMP_LOOP_and_1042_nl,
      COMP_LOOP_COMP_LOOP_and_1043_nl, COMP_LOOP_COMP_LOOP_and_1044_nl, COMP_LOOP_COMP_LOOP_and_1045_nl,
      COMP_LOOP_COMP_LOOP_and_1046_nl, COMP_LOOP_COMP_LOOP_and_1047_nl, COMP_LOOP_COMP_LOOP_and_1048_nl,
      COMP_LOOP_COMP_LOOP_and_1049_nl, COMP_LOOP_COMP_LOOP_and_1050_nl, COMP_LOOP_COMP_LOOP_and_1051_nl,
      {and_dcpl_571 , and_dcpl_577 , and_1025_cse , and_1028_cse , and_dcpl_589 ,
      and_1037_cse , and_1040_cse , and_1044_cse , and_1046_cse , and_1051_cse ,
      and_1052_cse , and_1055_cse , and_1056_cse , and_1060_cse , and_1061_cse ,
      and_1064_cse});
  assign COMP_LOOP_COMP_LOOP_and_1052_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[1]) &
      COMP_LOOP_nor_52_itm;
  assign COMP_LOOP_COMP_LOOP_and_1053_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[1]) &
      COMP_LOOP_nor_92_itm;
  assign COMP_LOOP_COMP_LOOP_and_1054_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[1]) &
      COMP_LOOP_nor_132_itm;
  assign COMP_LOOP_COMP_LOOP_and_1055_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[1]) &
      COMP_LOOP_nor_172_itm;
  assign COMP_LOOP_COMP_LOOP_and_1056_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[1]) &
      COMP_LOOP_nor_212_itm;
  assign COMP_LOOP_COMP_LOOP_and_1057_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[1]) &
      COMP_LOOP_nor_252_itm;
  assign COMP_LOOP_COMP_LOOP_and_1058_nl = (COMP_LOOP_acc_10_cse_10_1_8_sva[1]) &
      COMP_LOOP_nor_292_itm;
  assign COMP_LOOP_COMP_LOOP_and_1059_nl = (COMP_LOOP_acc_10_cse_10_1_9_sva[1]) &
      COMP_LOOP_nor_332_itm;
  assign COMP_LOOP_COMP_LOOP_and_1060_nl = (COMP_LOOP_acc_10_cse_10_1_10_sva[1])
      & COMP_LOOP_nor_372_itm;
  assign COMP_LOOP_COMP_LOOP_and_1061_nl = (COMP_LOOP_acc_10_cse_10_1_11_sva[1])
      & COMP_LOOP_nor_412_itm;
  assign COMP_LOOP_COMP_LOOP_and_1062_nl = (COMP_LOOP_acc_10_cse_10_1_12_sva[1])
      & COMP_LOOP_nor_452_itm;
  assign COMP_LOOP_COMP_LOOP_and_1063_nl = (COMP_LOOP_acc_10_cse_10_1_13_sva[1])
      & COMP_LOOP_nor_492_itm;
  assign COMP_LOOP_COMP_LOOP_and_1064_nl = (COMP_LOOP_acc_10_cse_10_1_14_sva[1])
      & COMP_LOOP_nor_532_itm;
  assign COMP_LOOP_COMP_LOOP_and_1065_nl = (COMP_LOOP_acc_10_cse_10_1_15_sva[1])
      & COMP_LOOP_nor_572_itm;
  assign COMP_LOOP_COMP_LOOP_and_1066_nl = (COMP_LOOP_acc_10_cse_10_1_sva[1]) & COMP_LOOP_nor_612_itm;
  assign COMP_LOOP_mux1h_720_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_62_itm,
      COMP_LOOP_COMP_LOOP_and_1052_nl, COMP_LOOP_COMP_LOOP_and_1053_nl, COMP_LOOP_COMP_LOOP_and_1054_nl,
      COMP_LOOP_COMP_LOOP_and_1055_nl, COMP_LOOP_COMP_LOOP_and_1056_nl, COMP_LOOP_COMP_LOOP_and_1057_nl,
      COMP_LOOP_COMP_LOOP_and_1058_nl, COMP_LOOP_COMP_LOOP_and_1059_nl, COMP_LOOP_COMP_LOOP_and_1060_nl,
      COMP_LOOP_COMP_LOOP_and_1061_nl, COMP_LOOP_COMP_LOOP_and_1062_nl, COMP_LOOP_COMP_LOOP_and_1063_nl,
      COMP_LOOP_COMP_LOOP_and_1064_nl, COMP_LOOP_COMP_LOOP_and_1065_nl, COMP_LOOP_COMP_LOOP_and_1066_nl,
      {and_dcpl_571 , and_dcpl_577 , and_1025_cse , and_1028_cse , and_dcpl_589 ,
      and_1037_cse , and_1040_cse , and_1044_cse , and_1046_cse , and_1051_cse ,
      and_1052_cse , and_1055_cse , and_1056_cse , and_1060_cse , and_1061_cse ,
      and_1064_cse});
  assign COMP_LOOP_mux1h_721_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_185_itm,
      COMP_LOOP_COMP_LOOP_and_77_itm, COMP_LOOP_COMP_LOOP_and_137_itm, COMP_LOOP_COMP_LOOP_and_197_itm,
      COMP_LOOP_COMP_LOOP_and_257_itm, COMP_LOOP_COMP_LOOP_and_317_itm, COMP_LOOP_COMP_LOOP_and_377_itm,
      COMP_LOOP_COMP_LOOP_and_437_itm, COMP_LOOP_COMP_LOOP_and_497_itm, COMP_LOOP_COMP_LOOP_and_557_itm,
      COMP_LOOP_COMP_LOOP_and_617_itm, COMP_LOOP_COMP_LOOP_and_677_itm, COMP_LOOP_COMP_LOOP_and_737_itm,
      COMP_LOOP_COMP_LOOP_and_797_itm, COMP_LOOP_COMP_LOOP_and_857_itm, COMP_LOOP_COMP_LOOP_and_917_itm,
      {and_dcpl_571 , and_dcpl_577 , and_1025_cse , and_1028_cse , and_dcpl_589 ,
      and_1037_cse , and_1040_cse , and_1044_cse , and_1046_cse , and_1051_cse ,
      and_1052_cse , and_1055_cse , and_1056_cse , and_1060_cse , and_1061_cse ,
      and_1064_cse});
  assign COMP_LOOP_COMP_LOOP_and_1067_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[2]) &
      COMP_LOOP_nor_54_itm;
  assign COMP_LOOP_COMP_LOOP_and_1068_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[2]) &
      COMP_LOOP_nor_94_itm;
  assign COMP_LOOP_COMP_LOOP_and_1069_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[2]) &
      COMP_LOOP_nor_134_itm;
  assign COMP_LOOP_COMP_LOOP_and_1070_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[2]) &
      COMP_LOOP_nor_174_itm;
  assign COMP_LOOP_COMP_LOOP_and_1071_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[2]) &
      COMP_LOOP_nor_214_itm;
  assign COMP_LOOP_COMP_LOOP_and_1072_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[2]) &
      COMP_LOOP_nor_254_itm;
  assign COMP_LOOP_COMP_LOOP_and_1073_nl = (COMP_LOOP_acc_10_cse_10_1_8_sva[2]) &
      COMP_LOOP_nor_294_itm;
  assign COMP_LOOP_COMP_LOOP_and_1074_nl = (COMP_LOOP_acc_10_cse_10_1_9_sva[2]) &
      COMP_LOOP_nor_334_itm;
  assign COMP_LOOP_COMP_LOOP_and_1075_nl = (COMP_LOOP_acc_10_cse_10_1_10_sva[2])
      & COMP_LOOP_nor_374_itm;
  assign COMP_LOOP_COMP_LOOP_and_1076_nl = (COMP_LOOP_acc_10_cse_10_1_11_sva[2])
      & COMP_LOOP_nor_414_itm;
  assign COMP_LOOP_COMP_LOOP_and_1077_nl = (COMP_LOOP_acc_10_cse_10_1_12_sva[2])
      & COMP_LOOP_nor_454_itm;
  assign COMP_LOOP_COMP_LOOP_and_1078_nl = (COMP_LOOP_acc_10_cse_10_1_13_sva[2])
      & COMP_LOOP_nor_494_itm;
  assign COMP_LOOP_COMP_LOOP_and_1079_nl = (COMP_LOOP_acc_10_cse_10_1_14_sva[2])
      & COMP_LOOP_nor_534_itm;
  assign COMP_LOOP_COMP_LOOP_and_1080_nl = (COMP_LOOP_acc_10_cse_10_1_15_sva[2])
      & COMP_LOOP_nor_574_itm;
  assign COMP_LOOP_COMP_LOOP_and_1081_nl = (COMP_LOOP_acc_10_cse_10_1_sva[2]) & COMP_LOOP_nor_614_itm;
  assign COMP_LOOP_mux1h_722_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_64_itm,
      COMP_LOOP_COMP_LOOP_and_1067_nl, COMP_LOOP_COMP_LOOP_and_1068_nl, COMP_LOOP_COMP_LOOP_and_1069_nl,
      COMP_LOOP_COMP_LOOP_and_1070_nl, COMP_LOOP_COMP_LOOP_and_1071_nl, COMP_LOOP_COMP_LOOP_and_1072_nl,
      COMP_LOOP_COMP_LOOP_and_1073_nl, COMP_LOOP_COMP_LOOP_and_1074_nl, COMP_LOOP_COMP_LOOP_and_1075_nl,
      COMP_LOOP_COMP_LOOP_and_1076_nl, COMP_LOOP_COMP_LOOP_and_1077_nl, COMP_LOOP_COMP_LOOP_and_1078_nl,
      COMP_LOOP_COMP_LOOP_and_1079_nl, COMP_LOOP_COMP_LOOP_and_1080_nl, COMP_LOOP_COMP_LOOP_and_1081_nl,
      {and_dcpl_571 , and_dcpl_577 , and_1025_cse , and_1028_cse , and_dcpl_589 ,
      and_1037_cse , and_1040_cse , and_1044_cse , and_1046_cse , and_1051_cse ,
      and_1052_cse , and_1055_cse , and_1056_cse , and_1060_cse , and_1061_cse ,
      and_1064_cse});
  assign COMP_LOOP_mux1h_723_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_65_itm,
      COMP_LOOP_COMP_LOOP_and_79_itm, COMP_LOOP_COMP_LOOP_and_139_itm, COMP_LOOP_COMP_LOOP_and_199_itm,
      COMP_LOOP_COMP_LOOP_and_259_itm, COMP_LOOP_COMP_LOOP_and_319_itm, COMP_LOOP_COMP_LOOP_and_379_itm,
      COMP_LOOP_COMP_LOOP_and_439_itm, COMP_LOOP_COMP_LOOP_and_499_itm, COMP_LOOP_COMP_LOOP_and_559_itm,
      COMP_LOOP_COMP_LOOP_and_619_itm, COMP_LOOP_COMP_LOOP_and_679_itm, COMP_LOOP_COMP_LOOP_and_739_itm,
      COMP_LOOP_COMP_LOOP_and_799_itm, COMP_LOOP_COMP_LOOP_and_859_itm, COMP_LOOP_COMP_LOOP_and_919_itm,
      {and_dcpl_571 , and_dcpl_577 , and_1025_cse , and_1028_cse , and_dcpl_589 ,
      and_1037_cse , and_1040_cse , and_1044_cse , and_1046_cse , and_1051_cse ,
      and_1052_cse , and_1055_cse , and_1056_cse , and_1060_cse , and_1061_cse ,
      and_1064_cse});
  assign COMP_LOOP_mux1h_724_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_66_itm,
      COMP_LOOP_COMP_LOOP_and_80_itm, COMP_LOOP_COMP_LOOP_and_140_itm, COMP_LOOP_COMP_LOOP_and_200_itm,
      COMP_LOOP_COMP_LOOP_and_260_itm, COMP_LOOP_COMP_LOOP_and_320_itm, COMP_LOOP_COMP_LOOP_and_380_itm,
      COMP_LOOP_COMP_LOOP_and_440_itm, COMP_LOOP_COMP_LOOP_and_500_itm, COMP_LOOP_COMP_LOOP_and_560_itm,
      COMP_LOOP_COMP_LOOP_and_620_itm, COMP_LOOP_COMP_LOOP_and_680_itm, COMP_LOOP_COMP_LOOP_and_740_itm,
      COMP_LOOP_COMP_LOOP_and_800_itm, COMP_LOOP_COMP_LOOP_and_860_itm, COMP_LOOP_COMP_LOOP_and_920_itm,
      {and_dcpl_571 , and_dcpl_577 , and_1025_cse , and_1028_cse , and_dcpl_589 ,
      and_1037_cse , and_1040_cse , and_1044_cse , and_1046_cse , and_1051_cse ,
      and_1052_cse , and_1055_cse , and_1056_cse , and_1060_cse , and_1061_cse ,
      and_1064_cse});
  assign COMP_LOOP_mux1h_725_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_6_itm,
      COMP_LOOP_COMP_LOOP_and_81_itm, COMP_LOOP_COMP_LOOP_and_141_itm, COMP_LOOP_COMP_LOOP_and_201_itm,
      COMP_LOOP_COMP_LOOP_and_261_itm, COMP_LOOP_COMP_LOOP_and_321_itm, COMP_LOOP_COMP_LOOP_and_381_itm,
      COMP_LOOP_COMP_LOOP_and_441_itm, COMP_LOOP_COMP_LOOP_and_501_itm, COMP_LOOP_COMP_LOOP_and_561_itm,
      COMP_LOOP_COMP_LOOP_and_621_itm, COMP_LOOP_COMP_LOOP_and_681_itm, COMP_LOOP_COMP_LOOP_and_741_itm,
      COMP_LOOP_COMP_LOOP_and_801_itm, COMP_LOOP_COMP_LOOP_and_861_itm, COMP_LOOP_COMP_LOOP_and_921_itm,
      {and_dcpl_571 , and_dcpl_577 , and_1025_cse , and_1028_cse , and_dcpl_589 ,
      and_1037_cse , and_1040_cse , and_1044_cse , and_1046_cse , and_1051_cse ,
      and_1052_cse , and_1055_cse , and_1056_cse , and_1060_cse , and_1061_cse ,
      and_1064_cse});
  assign COMP_LOOP_COMP_LOOP_and_1082_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[3]) &
      COMP_LOOP_nor_57_itm;
  assign COMP_LOOP_COMP_LOOP_and_1083_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[3]) &
      COMP_LOOP_nor_97_itm;
  assign COMP_LOOP_COMP_LOOP_and_1084_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[3]) &
      COMP_LOOP_nor_137_itm;
  assign COMP_LOOP_COMP_LOOP_and_1085_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[3]) &
      COMP_LOOP_nor_177_itm;
  assign COMP_LOOP_COMP_LOOP_and_1086_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3]) &
      COMP_LOOP_nor_217_itm;
  assign COMP_LOOP_COMP_LOOP_and_1087_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3]) &
      COMP_LOOP_nor_257_itm;
  assign COMP_LOOP_COMP_LOOP_and_1088_nl = (COMP_LOOP_acc_10_cse_10_1_8_sva[3]) &
      COMP_LOOP_nor_297_itm;
  assign COMP_LOOP_COMP_LOOP_and_1089_nl = (COMP_LOOP_acc_10_cse_10_1_9_sva[3]) &
      COMP_LOOP_nor_337_itm;
  assign COMP_LOOP_COMP_LOOP_and_1090_nl = (COMP_LOOP_acc_10_cse_10_1_10_sva[3])
      & COMP_LOOP_nor_377_itm;
  assign COMP_LOOP_COMP_LOOP_and_1091_nl = (COMP_LOOP_acc_10_cse_10_1_11_sva[3])
      & COMP_LOOP_nor_417_itm;
  assign COMP_LOOP_COMP_LOOP_and_1092_nl = (COMP_LOOP_acc_10_cse_10_1_12_sva[3])
      & COMP_LOOP_nor_457_itm;
  assign COMP_LOOP_COMP_LOOP_and_1093_nl = (COMP_LOOP_acc_10_cse_10_1_13_sva[3])
      & COMP_LOOP_nor_497_itm;
  assign COMP_LOOP_COMP_LOOP_and_1094_nl = (COMP_LOOP_acc_10_cse_10_1_14_sva[3])
      & COMP_LOOP_nor_537_itm;
  assign COMP_LOOP_COMP_LOOP_and_1095_nl = (COMP_LOOP_acc_10_cse_10_1_15_sva[3])
      & COMP_LOOP_nor_577_itm;
  assign COMP_LOOP_COMP_LOOP_and_1096_nl = (COMP_LOOP_acc_10_cse_10_1_sva[3]) & COMP_LOOP_nor_617_itm;
  assign COMP_LOOP_mux1h_726_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_68_itm,
      COMP_LOOP_COMP_LOOP_and_1082_nl, COMP_LOOP_COMP_LOOP_and_1083_nl, COMP_LOOP_COMP_LOOP_and_1084_nl,
      COMP_LOOP_COMP_LOOP_and_1085_nl, COMP_LOOP_COMP_LOOP_and_1086_nl, COMP_LOOP_COMP_LOOP_and_1087_nl,
      COMP_LOOP_COMP_LOOP_and_1088_nl, COMP_LOOP_COMP_LOOP_and_1089_nl, COMP_LOOP_COMP_LOOP_and_1090_nl,
      COMP_LOOP_COMP_LOOP_and_1091_nl, COMP_LOOP_COMP_LOOP_and_1092_nl, COMP_LOOP_COMP_LOOP_and_1093_nl,
      COMP_LOOP_COMP_LOOP_and_1094_nl, COMP_LOOP_COMP_LOOP_and_1095_nl, COMP_LOOP_COMP_LOOP_and_1096_nl,
      {and_dcpl_571 , and_dcpl_577 , and_1025_cse , and_1028_cse , and_dcpl_589 ,
      and_1037_cse , and_1040_cse , and_1044_cse , and_1046_cse , and_1051_cse ,
      and_1052_cse , and_1055_cse , and_1056_cse , and_1060_cse , and_1061_cse ,
      and_1064_cse});
  assign COMP_LOOP_mux1h_727_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_69_itm,
      COMP_LOOP_COMP_LOOP_and_83_itm, COMP_LOOP_COMP_LOOP_and_143_itm, COMP_LOOP_COMP_LOOP_and_203_itm,
      COMP_LOOP_COMP_LOOP_and_263_itm, COMP_LOOP_COMP_LOOP_and_323_itm, COMP_LOOP_COMP_LOOP_and_383_itm,
      COMP_LOOP_COMP_LOOP_and_443_itm, COMP_LOOP_COMP_LOOP_and_503_itm, COMP_LOOP_COMP_LOOP_and_563_itm,
      COMP_LOOP_COMP_LOOP_and_623_itm, COMP_LOOP_COMP_LOOP_and_683_itm, COMP_LOOP_COMP_LOOP_and_743_itm,
      COMP_LOOP_COMP_LOOP_and_803_itm, COMP_LOOP_COMP_LOOP_and_863_itm, COMP_LOOP_COMP_LOOP_and_923_itm,
      {and_dcpl_571 , and_dcpl_577 , and_1025_cse , and_1028_cse , and_dcpl_589 ,
      and_1037_cse , and_1040_cse , and_1044_cse , and_1046_cse , and_1051_cse ,
      and_1052_cse , and_1055_cse , and_1056_cse , and_1060_cse , and_1061_cse ,
      and_1064_cse});
  assign COMP_LOOP_mux1h_728_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_70_itm,
      COMP_LOOP_COMP_LOOP_and_84_itm, COMP_LOOP_COMP_LOOP_and_144_itm, COMP_LOOP_COMP_LOOP_and_204_itm,
      COMP_LOOP_COMP_LOOP_and_264_itm, COMP_LOOP_COMP_LOOP_and_324_itm, COMP_LOOP_COMP_LOOP_and_384_itm,
      COMP_LOOP_COMP_LOOP_and_444_itm, COMP_LOOP_COMP_LOOP_and_504_itm, COMP_LOOP_COMP_LOOP_and_564_itm,
      COMP_LOOP_COMP_LOOP_and_624_itm, COMP_LOOP_COMP_LOOP_and_684_itm, COMP_LOOP_COMP_LOOP_and_744_itm,
      COMP_LOOP_COMP_LOOP_and_804_itm, COMP_LOOP_COMP_LOOP_and_864_itm, COMP_LOOP_COMP_LOOP_and_924_itm,
      {and_dcpl_571 , and_dcpl_577 , and_1025_cse , and_1028_cse , and_dcpl_589 ,
      and_1037_cse , and_1040_cse , and_1044_cse , and_1046_cse , and_1051_cse ,
      and_1052_cse , and_1055_cse , and_1056_cse , and_1060_cse , and_1061_cse ,
      and_1064_cse});
  assign COMP_LOOP_mux1h_729_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_10_itm,
      COMP_LOOP_COMP_LOOP_and_85_itm, COMP_LOOP_COMP_LOOP_and_145_itm, COMP_LOOP_COMP_LOOP_and_205_itm,
      COMP_LOOP_COMP_LOOP_and_265_itm, COMP_LOOP_COMP_LOOP_and_325_itm, COMP_LOOP_COMP_LOOP_and_385_itm,
      COMP_LOOP_COMP_LOOP_and_445_itm, COMP_LOOP_COMP_LOOP_and_505_itm, COMP_LOOP_COMP_LOOP_and_565_itm,
      COMP_LOOP_COMP_LOOP_and_625_itm, COMP_LOOP_COMP_LOOP_and_685_itm, COMP_LOOP_COMP_LOOP_and_745_itm,
      COMP_LOOP_COMP_LOOP_and_805_itm, COMP_LOOP_COMP_LOOP_and_865_itm, COMP_LOOP_COMP_LOOP_and_925_itm,
      {and_dcpl_571 , and_dcpl_577 , and_1025_cse , and_1028_cse , and_dcpl_589 ,
      and_1037_cse , and_1040_cse , and_1044_cse , and_1046_cse , and_1051_cse ,
      and_1052_cse , and_1055_cse , and_1056_cse , and_1060_cse , and_1061_cse ,
      and_1064_cse});
  assign COMP_LOOP_mux1h_730_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_72_itm,
      COMP_LOOP_COMP_LOOP_and_86_itm, COMP_LOOP_COMP_LOOP_and_146_itm, COMP_LOOP_COMP_LOOP_and_206_itm,
      COMP_LOOP_COMP_LOOP_and_266_itm, COMP_LOOP_COMP_LOOP_and_326_itm, COMP_LOOP_COMP_LOOP_and_386_itm,
      COMP_LOOP_COMP_LOOP_and_446_itm, COMP_LOOP_COMP_LOOP_and_506_itm, COMP_LOOP_COMP_LOOP_and_566_itm,
      COMP_LOOP_COMP_LOOP_and_626_itm, COMP_LOOP_COMP_LOOP_and_686_itm, COMP_LOOP_COMP_LOOP_and_746_itm,
      COMP_LOOP_COMP_LOOP_and_806_itm, COMP_LOOP_COMP_LOOP_and_866_itm, COMP_LOOP_COMP_LOOP_and_926_itm,
      {and_dcpl_571 , and_dcpl_577 , and_1025_cse , and_1028_cse , and_dcpl_589 ,
      and_1037_cse , and_1040_cse , and_1044_cse , and_1046_cse , and_1051_cse ,
      and_1052_cse , and_1055_cse , and_1056_cse , and_1060_cse , and_1061_cse ,
      and_1064_cse});
  assign COMP_LOOP_mux1h_731_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_12_itm,
      COMP_LOOP_COMP_LOOP_and_87_itm, COMP_LOOP_COMP_LOOP_and_147_itm, COMP_LOOP_COMP_LOOP_and_207_itm,
      COMP_LOOP_COMP_LOOP_and_267_itm, COMP_LOOP_COMP_LOOP_and_327_itm, COMP_LOOP_COMP_LOOP_and_387_itm,
      COMP_LOOP_COMP_LOOP_and_447_itm, COMP_LOOP_COMP_LOOP_and_507_itm, COMP_LOOP_COMP_LOOP_and_567_itm,
      COMP_LOOP_COMP_LOOP_and_627_itm, COMP_LOOP_COMP_LOOP_and_687_itm, COMP_LOOP_COMP_LOOP_and_747_itm,
      COMP_LOOP_COMP_LOOP_and_807_itm, COMP_LOOP_COMP_LOOP_and_867_itm, COMP_LOOP_COMP_LOOP_and_927_itm,
      {and_dcpl_571 , and_dcpl_577 , and_1025_cse , and_1028_cse , and_dcpl_589 ,
      and_1037_cse , and_1040_cse , and_1044_cse , and_1046_cse , and_1051_cse ,
      and_1052_cse , and_1055_cse , and_1056_cse , and_1060_cse , and_1061_cse ,
      and_1064_cse});
  assign COMP_LOOP_mux1h_732_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_13_itm,
      COMP_LOOP_COMP_LOOP_and_88_itm, COMP_LOOP_COMP_LOOP_and_148_itm, COMP_LOOP_COMP_LOOP_and_208_itm,
      COMP_LOOP_COMP_LOOP_and_268_itm, COMP_LOOP_COMP_LOOP_and_328_itm, COMP_LOOP_COMP_LOOP_and_388_itm,
      COMP_LOOP_COMP_LOOP_and_448_itm, COMP_LOOP_COMP_LOOP_and_508_itm, COMP_LOOP_COMP_LOOP_and_568_itm,
      COMP_LOOP_COMP_LOOP_and_628_itm, COMP_LOOP_COMP_LOOP_and_688_itm, COMP_LOOP_COMP_LOOP_and_748_itm,
      COMP_LOOP_COMP_LOOP_and_808_itm, COMP_LOOP_COMP_LOOP_and_868_itm, COMP_LOOP_COMP_LOOP_and_928_itm,
      {and_dcpl_571 , and_dcpl_577 , and_1025_cse , and_1028_cse , and_dcpl_589 ,
      and_1037_cse , and_1040_cse , and_1044_cse , and_1046_cse , and_1051_cse ,
      and_1052_cse , and_1055_cse , and_1056_cse , and_1060_cse , and_1061_cse ,
      and_1064_cse});
  assign COMP_LOOP_mux1h_733_nl = MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_14_itm,
      COMP_LOOP_COMP_LOOP_and_89_itm, COMP_LOOP_COMP_LOOP_and_149_itm, COMP_LOOP_COMP_LOOP_and_209_itm,
      COMP_LOOP_COMP_LOOP_and_269_itm, COMP_LOOP_COMP_LOOP_and_329_itm, COMP_LOOP_COMP_LOOP_and_389_itm,
      COMP_LOOP_COMP_LOOP_and_449_itm, COMP_LOOP_COMP_LOOP_and_509_itm, COMP_LOOP_COMP_LOOP_and_569_itm,
      COMP_LOOP_COMP_LOOP_and_629_itm, COMP_LOOP_COMP_LOOP_and_689_itm, COMP_LOOP_COMP_LOOP_and_749_itm,
      COMP_LOOP_COMP_LOOP_and_809_itm, COMP_LOOP_COMP_LOOP_and_869_itm, COMP_LOOP_COMP_LOOP_and_929_itm,
      {and_dcpl_571 , and_dcpl_577 , and_1025_cse , and_1028_cse , and_dcpl_589 ,
      and_1037_cse , and_1040_cse , and_1044_cse , and_1046_cse , and_1051_cse ,
      and_1052_cse , and_1055_cse , and_1056_cse , and_1060_cse , and_1061_cse ,
      and_1064_cse});
  assign z_out_7 = MUX1HOT_v_64_16_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d, vec_rsc_0_2_i_q_d,
      vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d, vec_rsc_0_6_i_q_d,
      vec_rsc_0_7_i_q_d, vec_rsc_0_8_i_q_d, vec_rsc_0_9_i_q_d, vec_rsc_0_10_i_q_d,
      vec_rsc_0_11_i_q_d, vec_rsc_0_12_i_q_d, vec_rsc_0_13_i_q_d, vec_rsc_0_14_i_q_d,
      vec_rsc_0_15_i_q_d, {COMP_LOOP_mux1h_718_nl , COMP_LOOP_mux1h_719_nl , COMP_LOOP_mux1h_720_nl
      , COMP_LOOP_mux1h_721_nl , COMP_LOOP_mux1h_722_nl , COMP_LOOP_mux1h_723_nl
      , COMP_LOOP_mux1h_724_nl , COMP_LOOP_mux1h_725_nl , COMP_LOOP_mux1h_726_nl
      , COMP_LOOP_mux1h_727_nl , COMP_LOOP_mux1h_728_nl , COMP_LOOP_mux1h_729_nl
      , COMP_LOOP_mux1h_730_nl , COMP_LOOP_mux1h_731_nl , COMP_LOOP_mux1h_732_nl
      , COMP_LOOP_mux1h_733_nl});

  function automatic [0:0] MUX1HOT_s_1_16_2;
    input [0:0] input_15;
    input [0:0] input_14;
    input [0:0] input_13;
    input [0:0] input_12;
    input [0:0] input_11;
    input [0:0] input_10;
    input [0:0] input_9;
    input [0:0] input_8;
    input [0:0] input_7;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [15:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    result = result | ( input_7 & {1{sel[7]}});
    result = result | ( input_8 & {1{sel[8]}});
    result = result | ( input_9 & {1{sel[9]}});
    result = result | ( input_10 & {1{sel[10]}});
    result = result | ( input_11 & {1{sel[11]}});
    result = result | ( input_12 & {1{sel[12]}});
    result = result | ( input_13 & {1{sel[13]}});
    result = result | ( input_14 & {1{sel[14]}});
    result = result | ( input_15 & {1{sel[15]}});
    MUX1HOT_s_1_16_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_17_2;
    input [0:0] input_16;
    input [0:0] input_15;
    input [0:0] input_14;
    input [0:0] input_13;
    input [0:0] input_12;
    input [0:0] input_11;
    input [0:0] input_10;
    input [0:0] input_9;
    input [0:0] input_8;
    input [0:0] input_7;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [16:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    result = result | ( input_7 & {1{sel[7]}});
    result = result | ( input_8 & {1{sel[8]}});
    result = result | ( input_9 & {1{sel[9]}});
    result = result | ( input_10 & {1{sel[10]}});
    result = result | ( input_11 & {1{sel[11]}});
    result = result | ( input_12 & {1{sel[12]}});
    result = result | ( input_13 & {1{sel[13]}});
    result = result | ( input_14 & {1{sel[14]}});
    result = result | ( input_15 & {1{sel[15]}});
    result = result | ( input_16 & {1{sel[16]}});
    MUX1HOT_s_1_17_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_18_2;
    input [0:0] input_17;
    input [0:0] input_16;
    input [0:0] input_15;
    input [0:0] input_14;
    input [0:0] input_13;
    input [0:0] input_12;
    input [0:0] input_11;
    input [0:0] input_10;
    input [0:0] input_9;
    input [0:0] input_8;
    input [0:0] input_7;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [17:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    result = result | ( input_7 & {1{sel[7]}});
    result = result | ( input_8 & {1{sel[8]}});
    result = result | ( input_9 & {1{sel[9]}});
    result = result | ( input_10 & {1{sel[10]}});
    result = result | ( input_11 & {1{sel[11]}});
    result = result | ( input_12 & {1{sel[12]}});
    result = result | ( input_13 & {1{sel[13]}});
    result = result | ( input_14 & {1{sel[14]}});
    result = result | ( input_15 & {1{sel[15]}});
    result = result | ( input_16 & {1{sel[16]}});
    result = result | ( input_17 & {1{sel[17]}});
    MUX1HOT_s_1_18_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_5_2;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [4:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    MUX1HOT_v_4_5_2 = result;
  end
  endfunction


  function automatic [53:0] MUX1HOT_v_54_15_2;
    input [53:0] input_14;
    input [53:0] input_13;
    input [53:0] input_12;
    input [53:0] input_11;
    input [53:0] input_10;
    input [53:0] input_9;
    input [53:0] input_8;
    input [53:0] input_7;
    input [53:0] input_6;
    input [53:0] input_5;
    input [53:0] input_4;
    input [53:0] input_3;
    input [53:0] input_2;
    input [53:0] input_1;
    input [53:0] input_0;
    input [14:0] sel;
    reg [53:0] result;
  begin
    result = input_0 & {54{sel[0]}};
    result = result | ( input_1 & {54{sel[1]}});
    result = result | ( input_2 & {54{sel[2]}});
    result = result | ( input_3 & {54{sel[3]}});
    result = result | ( input_4 & {54{sel[4]}});
    result = result | ( input_5 & {54{sel[5]}});
    result = result | ( input_6 & {54{sel[6]}});
    result = result | ( input_7 & {54{sel[7]}});
    result = result | ( input_8 & {54{sel[8]}});
    result = result | ( input_9 & {54{sel[9]}});
    result = result | ( input_10 & {54{sel[10]}});
    result = result | ( input_11 & {54{sel[11]}});
    result = result | ( input_12 & {54{sel[12]}});
    result = result | ( input_13 & {54{sel[13]}});
    result = result | ( input_14 & {54{sel[14]}});
    MUX1HOT_v_54_15_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_16_2;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [15:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    MUX1HOT_v_64_16_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_19_2;
    input [63:0] input_18;
    input [63:0] input_17;
    input [63:0] input_16;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [18:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    result = result | ( input_16 & {64{sel[16]}});
    result = result | ( input_17 & {64{sel[17]}});
    result = result | ( input_18 & {64{sel[18]}});
    MUX1HOT_v_64_19_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_4_2;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [3:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    MUX1HOT_v_64_4_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_6_2;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [5:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    MUX1HOT_v_64_6_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_32_2;
    input [5:0] input_31;
    input [5:0] input_30;
    input [5:0] input_29;
    input [5:0] input_28;
    input [5:0] input_27;
    input [5:0] input_26;
    input [5:0] input_25;
    input [5:0] input_24;
    input [5:0] input_23;
    input [5:0] input_22;
    input [5:0] input_21;
    input [5:0] input_20;
    input [5:0] input_19;
    input [5:0] input_18;
    input [5:0] input_17;
    input [5:0] input_16;
    input [5:0] input_15;
    input [5:0] input_14;
    input [5:0] input_13;
    input [5:0] input_12;
    input [5:0] input_11;
    input [5:0] input_10;
    input [5:0] input_9;
    input [5:0] input_8;
    input [5:0] input_7;
    input [5:0] input_6;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [31:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    result = result | ( input_3 & {6{sel[3]}});
    result = result | ( input_4 & {6{sel[4]}});
    result = result | ( input_5 & {6{sel[5]}});
    result = result | ( input_6 & {6{sel[6]}});
    result = result | ( input_7 & {6{sel[7]}});
    result = result | ( input_8 & {6{sel[8]}});
    result = result | ( input_9 & {6{sel[9]}});
    result = result | ( input_10 & {6{sel[10]}});
    result = result | ( input_11 & {6{sel[11]}});
    result = result | ( input_12 & {6{sel[12]}});
    result = result | ( input_13 & {6{sel[13]}});
    result = result | ( input_14 & {6{sel[14]}});
    result = result | ( input_15 & {6{sel[15]}});
    result = result | ( input_16 & {6{sel[16]}});
    result = result | ( input_17 & {6{sel[17]}});
    result = result | ( input_18 & {6{sel[18]}});
    result = result | ( input_19 & {6{sel[19]}});
    result = result | ( input_20 & {6{sel[20]}});
    result = result | ( input_21 & {6{sel[21]}});
    result = result | ( input_22 & {6{sel[22]}});
    result = result | ( input_23 & {6{sel[23]}});
    result = result | ( input_24 & {6{sel[24]}});
    result = result | ( input_25 & {6{sel[25]}});
    result = result | ( input_26 & {6{sel[26]}});
    result = result | ( input_27 & {6{sel[27]}});
    result = result | ( input_28 & {6{sel[28]}});
    result = result | ( input_29 & {6{sel[29]}});
    result = result | ( input_30 & {6{sel[30]}});
    result = result | ( input_31 & {6{sel[31]}});
    MUX1HOT_v_6_32_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    result = result | ( input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_6_2;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [5:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    result = result | ( input_3 & {6{sel[3]}});
    result = result | ( input_4 & {6{sel[4]}});
    result = result | ( input_5 & {6{sel[5]}});
    MUX1HOT_v_6_6_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_20_2;
    input [7:0] input_19;
    input [7:0] input_18;
    input [7:0] input_17;
    input [7:0] input_16;
    input [7:0] input_15;
    input [7:0] input_14;
    input [7:0] input_13;
    input [7:0] input_12;
    input [7:0] input_11;
    input [7:0] input_10;
    input [7:0] input_9;
    input [7:0] input_8;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [19:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    result = result | ( input_5 & {8{sel[5]}});
    result = result | ( input_6 & {8{sel[6]}});
    result = result | ( input_7 & {8{sel[7]}});
    result = result | ( input_8 & {8{sel[8]}});
    result = result | ( input_9 & {8{sel[9]}});
    result = result | ( input_10 & {8{sel[10]}});
    result = result | ( input_11 & {8{sel[11]}});
    result = result | ( input_12 & {8{sel[12]}});
    result = result | ( input_13 & {8{sel[13]}});
    result = result | ( input_14 & {8{sel[14]}});
    result = result | ( input_15 & {8{sel[15]}});
    result = result | ( input_16 & {8{sel[16]}});
    result = result | ( input_17 & {8{sel[17]}});
    result = result | ( input_18 & {8{sel[18]}});
    result = result | ( input_19 & {8{sel[19]}});
    MUX1HOT_v_8_20_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [53:0] MUX_v_54_2_2;
    input [53:0] input_0;
    input [53:0] input_1;
    input [0:0] sel;
    reg [53:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_54_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [9:0] readslicef_11_10_1;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_11_10_1 = tmp[9:0];
  end
  endfunction


  function automatic [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function automatic [10:0] readslicef_12_11_1;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_12_11_1 = tmp[10:0];
  end
  endfunction


  function automatic [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function automatic [63:0] readslicef_65_64_1;
    input [64:0] vector;
    reg [64:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_65_64_1 = tmp[63:0];
  end
  endfunction


  function automatic [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_12 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF
// ------------------------------------------------------------------


module inPlaceNTT_DIF (
  clk, rst, vec_rsc_0_0_wadr, vec_rsc_0_0_d, vec_rsc_0_0_we, vec_rsc_0_0_radr, vec_rsc_0_0_q,
      vec_rsc_triosy_0_0_lz, vec_rsc_0_1_wadr, vec_rsc_0_1_d, vec_rsc_0_1_we, vec_rsc_0_1_radr,
      vec_rsc_0_1_q, vec_rsc_triosy_0_1_lz, vec_rsc_0_2_wadr, vec_rsc_0_2_d, vec_rsc_0_2_we,
      vec_rsc_0_2_radr, vec_rsc_0_2_q, vec_rsc_triosy_0_2_lz, vec_rsc_0_3_wadr, vec_rsc_0_3_d,
      vec_rsc_0_3_we, vec_rsc_0_3_radr, vec_rsc_0_3_q, vec_rsc_triosy_0_3_lz, vec_rsc_0_4_wadr,
      vec_rsc_0_4_d, vec_rsc_0_4_we, vec_rsc_0_4_radr, vec_rsc_0_4_q, vec_rsc_triosy_0_4_lz,
      vec_rsc_0_5_wadr, vec_rsc_0_5_d, vec_rsc_0_5_we, vec_rsc_0_5_radr, vec_rsc_0_5_q,
      vec_rsc_triosy_0_5_lz, vec_rsc_0_6_wadr, vec_rsc_0_6_d, vec_rsc_0_6_we, vec_rsc_0_6_radr,
      vec_rsc_0_6_q, vec_rsc_triosy_0_6_lz, vec_rsc_0_7_wadr, vec_rsc_0_7_d, vec_rsc_0_7_we,
      vec_rsc_0_7_radr, vec_rsc_0_7_q, vec_rsc_triosy_0_7_lz, vec_rsc_0_8_wadr, vec_rsc_0_8_d,
      vec_rsc_0_8_we, vec_rsc_0_8_radr, vec_rsc_0_8_q, vec_rsc_triosy_0_8_lz, vec_rsc_0_9_wadr,
      vec_rsc_0_9_d, vec_rsc_0_9_we, vec_rsc_0_9_radr, vec_rsc_0_9_q, vec_rsc_triosy_0_9_lz,
      vec_rsc_0_10_wadr, vec_rsc_0_10_d, vec_rsc_0_10_we, vec_rsc_0_10_radr, vec_rsc_0_10_q,
      vec_rsc_triosy_0_10_lz, vec_rsc_0_11_wadr, vec_rsc_0_11_d, vec_rsc_0_11_we,
      vec_rsc_0_11_radr, vec_rsc_0_11_q, vec_rsc_triosy_0_11_lz, vec_rsc_0_12_wadr,
      vec_rsc_0_12_d, vec_rsc_0_12_we, vec_rsc_0_12_radr, vec_rsc_0_12_q, vec_rsc_triosy_0_12_lz,
      vec_rsc_0_13_wadr, vec_rsc_0_13_d, vec_rsc_0_13_we, vec_rsc_0_13_radr, vec_rsc_0_13_q,
      vec_rsc_triosy_0_13_lz, vec_rsc_0_14_wadr, vec_rsc_0_14_d, vec_rsc_0_14_we,
      vec_rsc_0_14_radr, vec_rsc_0_14_q, vec_rsc_triosy_0_14_lz, vec_rsc_0_15_wadr,
      vec_rsc_0_15_d, vec_rsc_0_15_we, vec_rsc_0_15_radr, vec_rsc_0_15_q, vec_rsc_triosy_0_15_lz,
      p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz, twiddle_rsc_0_0_radr,
      twiddle_rsc_0_0_q, twiddle_rsc_triosy_0_0_lz, twiddle_rsc_0_1_radr, twiddle_rsc_0_1_q,
      twiddle_rsc_triosy_0_1_lz, twiddle_rsc_0_2_radr, twiddle_rsc_0_2_q, twiddle_rsc_triosy_0_2_lz,
      twiddle_rsc_0_3_radr, twiddle_rsc_0_3_q, twiddle_rsc_triosy_0_3_lz, twiddle_rsc_0_4_radr,
      twiddle_rsc_0_4_q, twiddle_rsc_triosy_0_4_lz, twiddle_rsc_0_5_radr, twiddle_rsc_0_5_q,
      twiddle_rsc_triosy_0_5_lz, twiddle_rsc_0_6_radr, twiddle_rsc_0_6_q, twiddle_rsc_triosy_0_6_lz,
      twiddle_rsc_0_7_radr, twiddle_rsc_0_7_q, twiddle_rsc_triosy_0_7_lz, twiddle_rsc_0_8_radr,
      twiddle_rsc_0_8_q, twiddle_rsc_triosy_0_8_lz, twiddle_rsc_0_9_radr, twiddle_rsc_0_9_q,
      twiddle_rsc_triosy_0_9_lz, twiddle_rsc_0_10_radr, twiddle_rsc_0_10_q, twiddle_rsc_triosy_0_10_lz,
      twiddle_rsc_0_11_radr, twiddle_rsc_0_11_q, twiddle_rsc_triosy_0_11_lz, twiddle_rsc_0_12_radr,
      twiddle_rsc_0_12_q, twiddle_rsc_triosy_0_12_lz, twiddle_rsc_0_13_radr, twiddle_rsc_0_13_q,
      twiddle_rsc_triosy_0_13_lz, twiddle_rsc_0_14_radr, twiddle_rsc_0_14_q, twiddle_rsc_triosy_0_14_lz,
      twiddle_rsc_0_15_radr, twiddle_rsc_0_15_q, twiddle_rsc_triosy_0_15_lz
);
  input clk;
  input rst;
  output [5:0] vec_rsc_0_0_wadr;
  output [63:0] vec_rsc_0_0_d;
  output vec_rsc_0_0_we;
  output [5:0] vec_rsc_0_0_radr;
  input [63:0] vec_rsc_0_0_q;
  output vec_rsc_triosy_0_0_lz;
  output [5:0] vec_rsc_0_1_wadr;
  output [63:0] vec_rsc_0_1_d;
  output vec_rsc_0_1_we;
  output [5:0] vec_rsc_0_1_radr;
  input [63:0] vec_rsc_0_1_q;
  output vec_rsc_triosy_0_1_lz;
  output [5:0] vec_rsc_0_2_wadr;
  output [63:0] vec_rsc_0_2_d;
  output vec_rsc_0_2_we;
  output [5:0] vec_rsc_0_2_radr;
  input [63:0] vec_rsc_0_2_q;
  output vec_rsc_triosy_0_2_lz;
  output [5:0] vec_rsc_0_3_wadr;
  output [63:0] vec_rsc_0_3_d;
  output vec_rsc_0_3_we;
  output [5:0] vec_rsc_0_3_radr;
  input [63:0] vec_rsc_0_3_q;
  output vec_rsc_triosy_0_3_lz;
  output [5:0] vec_rsc_0_4_wadr;
  output [63:0] vec_rsc_0_4_d;
  output vec_rsc_0_4_we;
  output [5:0] vec_rsc_0_4_radr;
  input [63:0] vec_rsc_0_4_q;
  output vec_rsc_triosy_0_4_lz;
  output [5:0] vec_rsc_0_5_wadr;
  output [63:0] vec_rsc_0_5_d;
  output vec_rsc_0_5_we;
  output [5:0] vec_rsc_0_5_radr;
  input [63:0] vec_rsc_0_5_q;
  output vec_rsc_triosy_0_5_lz;
  output [5:0] vec_rsc_0_6_wadr;
  output [63:0] vec_rsc_0_6_d;
  output vec_rsc_0_6_we;
  output [5:0] vec_rsc_0_6_radr;
  input [63:0] vec_rsc_0_6_q;
  output vec_rsc_triosy_0_6_lz;
  output [5:0] vec_rsc_0_7_wadr;
  output [63:0] vec_rsc_0_7_d;
  output vec_rsc_0_7_we;
  output [5:0] vec_rsc_0_7_radr;
  input [63:0] vec_rsc_0_7_q;
  output vec_rsc_triosy_0_7_lz;
  output [5:0] vec_rsc_0_8_wadr;
  output [63:0] vec_rsc_0_8_d;
  output vec_rsc_0_8_we;
  output [5:0] vec_rsc_0_8_radr;
  input [63:0] vec_rsc_0_8_q;
  output vec_rsc_triosy_0_8_lz;
  output [5:0] vec_rsc_0_9_wadr;
  output [63:0] vec_rsc_0_9_d;
  output vec_rsc_0_9_we;
  output [5:0] vec_rsc_0_9_radr;
  input [63:0] vec_rsc_0_9_q;
  output vec_rsc_triosy_0_9_lz;
  output [5:0] vec_rsc_0_10_wadr;
  output [63:0] vec_rsc_0_10_d;
  output vec_rsc_0_10_we;
  output [5:0] vec_rsc_0_10_radr;
  input [63:0] vec_rsc_0_10_q;
  output vec_rsc_triosy_0_10_lz;
  output [5:0] vec_rsc_0_11_wadr;
  output [63:0] vec_rsc_0_11_d;
  output vec_rsc_0_11_we;
  output [5:0] vec_rsc_0_11_radr;
  input [63:0] vec_rsc_0_11_q;
  output vec_rsc_triosy_0_11_lz;
  output [5:0] vec_rsc_0_12_wadr;
  output [63:0] vec_rsc_0_12_d;
  output vec_rsc_0_12_we;
  output [5:0] vec_rsc_0_12_radr;
  input [63:0] vec_rsc_0_12_q;
  output vec_rsc_triosy_0_12_lz;
  output [5:0] vec_rsc_0_13_wadr;
  output [63:0] vec_rsc_0_13_d;
  output vec_rsc_0_13_we;
  output [5:0] vec_rsc_0_13_radr;
  input [63:0] vec_rsc_0_13_q;
  output vec_rsc_triosy_0_13_lz;
  output [5:0] vec_rsc_0_14_wadr;
  output [63:0] vec_rsc_0_14_d;
  output vec_rsc_0_14_we;
  output [5:0] vec_rsc_0_14_radr;
  input [63:0] vec_rsc_0_14_q;
  output vec_rsc_triosy_0_14_lz;
  output [5:0] vec_rsc_0_15_wadr;
  output [63:0] vec_rsc_0_15_d;
  output vec_rsc_0_15_we;
  output [5:0] vec_rsc_0_15_radr;
  input [63:0] vec_rsc_0_15_q;
  output vec_rsc_triosy_0_15_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  output [5:0] twiddle_rsc_0_0_radr;
  input [63:0] twiddle_rsc_0_0_q;
  output twiddle_rsc_triosy_0_0_lz;
  output [5:0] twiddle_rsc_0_1_radr;
  input [63:0] twiddle_rsc_0_1_q;
  output twiddle_rsc_triosy_0_1_lz;
  output [5:0] twiddle_rsc_0_2_radr;
  input [63:0] twiddle_rsc_0_2_q;
  output twiddle_rsc_triosy_0_2_lz;
  output [5:0] twiddle_rsc_0_3_radr;
  input [63:0] twiddle_rsc_0_3_q;
  output twiddle_rsc_triosy_0_3_lz;
  output [5:0] twiddle_rsc_0_4_radr;
  input [63:0] twiddle_rsc_0_4_q;
  output twiddle_rsc_triosy_0_4_lz;
  output [5:0] twiddle_rsc_0_5_radr;
  input [63:0] twiddle_rsc_0_5_q;
  output twiddle_rsc_triosy_0_5_lz;
  output [5:0] twiddle_rsc_0_6_radr;
  input [63:0] twiddle_rsc_0_6_q;
  output twiddle_rsc_triosy_0_6_lz;
  output [5:0] twiddle_rsc_0_7_radr;
  input [63:0] twiddle_rsc_0_7_q;
  output twiddle_rsc_triosy_0_7_lz;
  output [5:0] twiddle_rsc_0_8_radr;
  input [63:0] twiddle_rsc_0_8_q;
  output twiddle_rsc_triosy_0_8_lz;
  output [5:0] twiddle_rsc_0_9_radr;
  input [63:0] twiddle_rsc_0_9_q;
  output twiddle_rsc_triosy_0_9_lz;
  output [5:0] twiddle_rsc_0_10_radr;
  input [63:0] twiddle_rsc_0_10_q;
  output twiddle_rsc_triosy_0_10_lz;
  output [5:0] twiddle_rsc_0_11_radr;
  input [63:0] twiddle_rsc_0_11_q;
  output twiddle_rsc_triosy_0_11_lz;
  output [5:0] twiddle_rsc_0_12_radr;
  input [63:0] twiddle_rsc_0_12_q;
  output twiddle_rsc_triosy_0_12_lz;
  output [5:0] twiddle_rsc_0_13_radr;
  input [63:0] twiddle_rsc_0_13_q;
  output twiddle_rsc_triosy_0_13_lz;
  output [5:0] twiddle_rsc_0_14_radr;
  input [63:0] twiddle_rsc_0_14_q;
  output twiddle_rsc_triosy_0_14_lz;
  output [5:0] twiddle_rsc_0_15_radr;
  input [63:0] twiddle_rsc_0_15_q;
  output twiddle_rsc_triosy_0_15_lz;


  // Interconnect Declarations
  wire [63:0] vec_rsc_0_0_i_q_d;
  wire vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_1_i_q_d;
  wire vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_2_i_q_d;
  wire vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_3_i_q_d;
  wire vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_4_i_q_d;
  wire vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_5_i_q_d;
  wire vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_6_i_q_d;
  wire vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_7_i_q_d;
  wire vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_8_i_q_d;
  wire vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_9_i_q_d;
  wire vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_10_i_q_d;
  wire vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_11_i_q_d;
  wire vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_12_i_q_d;
  wire vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_13_i_q_d;
  wire vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_14_i_q_d;
  wire vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_15_i_q_d;
  wire vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_0_i_q_d;
  wire [5:0] twiddle_rsc_0_0_i_radr_d;
  wire twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_1_i_q_d;
  wire twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_2_i_q_d;
  wire twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_3_i_q_d;
  wire twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_4_i_q_d;
  wire twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_5_i_q_d;
  wire twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_6_i_q_d;
  wire twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_7_i_q_d;
  wire twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_8_i_q_d;
  wire [5:0] twiddle_rsc_0_8_i_radr_d;
  wire twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_9_i_q_d;
  wire twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_10_i_q_d;
  wire twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_11_i_q_d;
  wire twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_12_i_q_d;
  wire twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_13_i_q_d;
  wire twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_14_i_q_d;
  wire twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_15_i_q_d;
  wire twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_0_i_d_d_iff;
  wire [5:0] vec_rsc_0_0_i_radr_d_iff;
  wire [5:0] vec_rsc_0_0_i_wadr_d_iff;
  wire vec_rsc_0_0_i_we_d_iff;
  wire vec_rsc_0_1_i_we_d_iff;
  wire vec_rsc_0_2_i_we_d_iff;
  wire vec_rsc_0_3_i_we_d_iff;
  wire vec_rsc_0_4_i_we_d_iff;
  wire vec_rsc_0_5_i_we_d_iff;
  wire vec_rsc_0_6_i_we_d_iff;
  wire vec_rsc_0_7_i_we_d_iff;
  wire vec_rsc_0_8_i_we_d_iff;
  wire vec_rsc_0_9_i_we_d_iff;
  wire vec_rsc_0_10_i_we_d_iff;
  wire vec_rsc_0_11_i_we_d_iff;
  wire vec_rsc_0_12_i_we_d_iff;
  wire vec_rsc_0_13_i_we_d_iff;
  wire vec_rsc_0_14_i_we_d_iff;
  wire vec_rsc_0_15_i_we_d_iff;
  wire [5:0] twiddle_rsc_0_1_i_radr_d_iff;
  wire [5:0] twiddle_rsc_0_2_i_radr_d_iff;
  wire [5:0] twiddle_rsc_0_4_i_radr_d_iff;


  // Interconnect Declarations for Component Instantiations 
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen vec_rsc_0_0_i
      (
      .q(vec_rsc_0_0_q),
      .radr(vec_rsc_0_0_radr),
      .we(vec_rsc_0_0_we),
      .d(vec_rsc_0_0_d),
      .wadr(vec_rsc_0_0_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_0_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen vec_rsc_0_1_i
      (
      .q(vec_rsc_0_1_q),
      .radr(vec_rsc_0_1_radr),
      .we(vec_rsc_0_1_we),
      .d(vec_rsc_0_1_d),
      .wadr(vec_rsc_0_1_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_1_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_1_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_1_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen vec_rsc_0_2_i
      (
      .q(vec_rsc_0_2_q),
      .radr(vec_rsc_0_2_radr),
      .we(vec_rsc_0_2_we),
      .d(vec_rsc_0_2_d),
      .wadr(vec_rsc_0_2_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_2_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_2_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_2_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen vec_rsc_0_3_i
      (
      .q(vec_rsc_0_3_q),
      .radr(vec_rsc_0_3_radr),
      .we(vec_rsc_0_3_we),
      .d(vec_rsc_0_3_d),
      .wadr(vec_rsc_0_3_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_3_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_3_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_3_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen vec_rsc_0_4_i
      (
      .q(vec_rsc_0_4_q),
      .radr(vec_rsc_0_4_radr),
      .we(vec_rsc_0_4_we),
      .d(vec_rsc_0_4_d),
      .wadr(vec_rsc_0_4_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_4_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_4_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_4_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen vec_rsc_0_5_i
      (
      .q(vec_rsc_0_5_q),
      .radr(vec_rsc_0_5_radr),
      .we(vec_rsc_0_5_we),
      .d(vec_rsc_0_5_d),
      .wadr(vec_rsc_0_5_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_5_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_5_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_5_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen vec_rsc_0_6_i
      (
      .q(vec_rsc_0_6_q),
      .radr(vec_rsc_0_6_radr),
      .we(vec_rsc_0_6_we),
      .d(vec_rsc_0_6_d),
      .wadr(vec_rsc_0_6_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_6_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_6_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_6_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen vec_rsc_0_7_i
      (
      .q(vec_rsc_0_7_q),
      .radr(vec_rsc_0_7_radr),
      .we(vec_rsc_0_7_we),
      .d(vec_rsc_0_7_d),
      .wadr(vec_rsc_0_7_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_7_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_7_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_7_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen vec_rsc_0_8_i
      (
      .q(vec_rsc_0_8_q),
      .radr(vec_rsc_0_8_radr),
      .we(vec_rsc_0_8_we),
      .d(vec_rsc_0_8_d),
      .wadr(vec_rsc_0_8_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_8_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_8_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_8_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen vec_rsc_0_9_i
      (
      .q(vec_rsc_0_9_q),
      .radr(vec_rsc_0_9_radr),
      .we(vec_rsc_0_9_we),
      .d(vec_rsc_0_9_d),
      .wadr(vec_rsc_0_9_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_9_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_9_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_9_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen vec_rsc_0_10_i
      (
      .q(vec_rsc_0_10_q),
      .radr(vec_rsc_0_10_radr),
      .we(vec_rsc_0_10_we),
      .d(vec_rsc_0_10_d),
      .wadr(vec_rsc_0_10_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_10_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_10_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_10_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen vec_rsc_0_11_i
      (
      .q(vec_rsc_0_11_q),
      .radr(vec_rsc_0_11_radr),
      .we(vec_rsc_0_11_we),
      .d(vec_rsc_0_11_d),
      .wadr(vec_rsc_0_11_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_11_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_11_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_11_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen vec_rsc_0_12_i
      (
      .q(vec_rsc_0_12_q),
      .radr(vec_rsc_0_12_radr),
      .we(vec_rsc_0_12_we),
      .d(vec_rsc_0_12_d),
      .wadr(vec_rsc_0_12_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_12_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_12_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_12_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen vec_rsc_0_13_i
      (
      .q(vec_rsc_0_13_q),
      .radr(vec_rsc_0_13_radr),
      .we(vec_rsc_0_13_we),
      .d(vec_rsc_0_13_d),
      .wadr(vec_rsc_0_13_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_13_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_13_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_13_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen vec_rsc_0_14_i
      (
      .q(vec_rsc_0_14_q),
      .radr(vec_rsc_0_14_radr),
      .we(vec_rsc_0_14_we),
      .d(vec_rsc_0_14_d),
      .wadr(vec_rsc_0_14_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_14_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_14_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_14_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_6_64_64_64_64_1_gen vec_rsc_0_15_i
      (
      .q(vec_rsc_0_15_q),
      .radr(vec_rsc_0_15_radr),
      .we(vec_rsc_0_15_we),
      .d(vec_rsc_0_15_d),
      .wadr(vec_rsc_0_15_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_15_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_15_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_15_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_25_6_64_64_64_64_1_gen twiddle_rsc_0_0_i
      (
      .q(twiddle_rsc_0_0_q),
      .radr(twiddle_rsc_0_0_radr),
      .q_d(twiddle_rsc_0_0_i_q_d),
      .radr_d(twiddle_rsc_0_0_i_radr_d),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_26_6_64_64_64_64_1_gen twiddle_rsc_0_1_i
      (
      .q(twiddle_rsc_0_1_q),
      .radr(twiddle_rsc_0_1_radr),
      .q_d(twiddle_rsc_0_1_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_27_6_64_64_64_64_1_gen twiddle_rsc_0_2_i
      (
      .q(twiddle_rsc_0_2_q),
      .radr(twiddle_rsc_0_2_radr),
      .q_d(twiddle_rsc_0_2_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_28_6_64_64_64_64_1_gen twiddle_rsc_0_3_i
      (
      .q(twiddle_rsc_0_3_q),
      .radr(twiddle_rsc_0_3_radr),
      .q_d(twiddle_rsc_0_3_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_29_6_64_64_64_64_1_gen twiddle_rsc_0_4_i
      (
      .q(twiddle_rsc_0_4_q),
      .radr(twiddle_rsc_0_4_radr),
      .q_d(twiddle_rsc_0_4_i_q_d),
      .radr_d(twiddle_rsc_0_4_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_30_6_64_64_64_64_1_gen twiddle_rsc_0_5_i
      (
      .q(twiddle_rsc_0_5_q),
      .radr(twiddle_rsc_0_5_radr),
      .q_d(twiddle_rsc_0_5_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_31_6_64_64_64_64_1_gen twiddle_rsc_0_6_i
      (
      .q(twiddle_rsc_0_6_q),
      .radr(twiddle_rsc_0_6_radr),
      .q_d(twiddle_rsc_0_6_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_32_6_64_64_64_64_1_gen twiddle_rsc_0_7_i
      (
      .q(twiddle_rsc_0_7_q),
      .radr(twiddle_rsc_0_7_radr),
      .q_d(twiddle_rsc_0_7_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_33_6_64_64_64_64_1_gen twiddle_rsc_0_8_i
      (
      .q(twiddle_rsc_0_8_q),
      .radr(twiddle_rsc_0_8_radr),
      .q_d(twiddle_rsc_0_8_i_q_d),
      .radr_d(twiddle_rsc_0_8_i_radr_d),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_34_6_64_64_64_64_1_gen twiddle_rsc_0_9_i
      (
      .q(twiddle_rsc_0_9_q),
      .radr(twiddle_rsc_0_9_radr),
      .q_d(twiddle_rsc_0_9_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_35_6_64_64_64_64_1_gen twiddle_rsc_0_10_i
      (
      .q(twiddle_rsc_0_10_q),
      .radr(twiddle_rsc_0_10_radr),
      .q_d(twiddle_rsc_0_10_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_36_6_64_64_64_64_1_gen twiddle_rsc_0_11_i
      (
      .q(twiddle_rsc_0_11_q),
      .radr(twiddle_rsc_0_11_radr),
      .q_d(twiddle_rsc_0_11_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_37_6_64_64_64_64_1_gen twiddle_rsc_0_12_i
      (
      .q(twiddle_rsc_0_12_q),
      .radr(twiddle_rsc_0_12_radr),
      .q_d(twiddle_rsc_0_12_i_q_d),
      .radr_d(twiddle_rsc_0_4_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_38_6_64_64_64_64_1_gen twiddle_rsc_0_13_i
      (
      .q(twiddle_rsc_0_13_q),
      .radr(twiddle_rsc_0_13_radr),
      .q_d(twiddle_rsc_0_13_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_39_6_64_64_64_64_1_gen twiddle_rsc_0_14_i
      (
      .q(twiddle_rsc_0_14_q),
      .radr(twiddle_rsc_0_14_radr),
      .q_d(twiddle_rsc_0_14_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_40_6_64_64_64_64_1_gen twiddle_rsc_0_15_i
      (
      .q(twiddle_rsc_0_15_q),
      .radr(twiddle_rsc_0_15_radr),
      .q_d(twiddle_rsc_0_15_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_core inPlaceNTT_DIF_core_inst (
      .clk(clk),
      .rst(rst),
      .vec_rsc_triosy_0_0_lz(vec_rsc_triosy_0_0_lz),
      .vec_rsc_triosy_0_1_lz(vec_rsc_triosy_0_1_lz),
      .vec_rsc_triosy_0_2_lz(vec_rsc_triosy_0_2_lz),
      .vec_rsc_triosy_0_3_lz(vec_rsc_triosy_0_3_lz),
      .vec_rsc_triosy_0_4_lz(vec_rsc_triosy_0_4_lz),
      .vec_rsc_triosy_0_5_lz(vec_rsc_triosy_0_5_lz),
      .vec_rsc_triosy_0_6_lz(vec_rsc_triosy_0_6_lz),
      .vec_rsc_triosy_0_7_lz(vec_rsc_triosy_0_7_lz),
      .vec_rsc_triosy_0_8_lz(vec_rsc_triosy_0_8_lz),
      .vec_rsc_triosy_0_9_lz(vec_rsc_triosy_0_9_lz),
      .vec_rsc_triosy_0_10_lz(vec_rsc_triosy_0_10_lz),
      .vec_rsc_triosy_0_11_lz(vec_rsc_triosy_0_11_lz),
      .vec_rsc_triosy_0_12_lz(vec_rsc_triosy_0_12_lz),
      .vec_rsc_triosy_0_13_lz(vec_rsc_triosy_0_13_lz),
      .vec_rsc_triosy_0_14_lz(vec_rsc_triosy_0_14_lz),
      .vec_rsc_triosy_0_15_lz(vec_rsc_triosy_0_15_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .twiddle_rsc_triosy_0_0_lz(twiddle_rsc_triosy_0_0_lz),
      .twiddle_rsc_triosy_0_1_lz(twiddle_rsc_triosy_0_1_lz),
      .twiddle_rsc_triosy_0_2_lz(twiddle_rsc_triosy_0_2_lz),
      .twiddle_rsc_triosy_0_3_lz(twiddle_rsc_triosy_0_3_lz),
      .twiddle_rsc_triosy_0_4_lz(twiddle_rsc_triosy_0_4_lz),
      .twiddle_rsc_triosy_0_5_lz(twiddle_rsc_triosy_0_5_lz),
      .twiddle_rsc_triosy_0_6_lz(twiddle_rsc_triosy_0_6_lz),
      .twiddle_rsc_triosy_0_7_lz(twiddle_rsc_triosy_0_7_lz),
      .twiddle_rsc_triosy_0_8_lz(twiddle_rsc_triosy_0_8_lz),
      .twiddle_rsc_triosy_0_9_lz(twiddle_rsc_triosy_0_9_lz),
      .twiddle_rsc_triosy_0_10_lz(twiddle_rsc_triosy_0_10_lz),
      .twiddle_rsc_triosy_0_11_lz(twiddle_rsc_triosy_0_11_lz),
      .twiddle_rsc_triosy_0_12_lz(twiddle_rsc_triosy_0_12_lz),
      .twiddle_rsc_triosy_0_13_lz(twiddle_rsc_triosy_0_13_lz),
      .twiddle_rsc_triosy_0_14_lz(twiddle_rsc_triosy_0_14_lz),
      .twiddle_rsc_triosy_0_15_lz(twiddle_rsc_triosy_0_15_lz),
      .vec_rsc_0_0_i_q_d(vec_rsc_0_0_i_q_d),
      .vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_1_i_q_d(vec_rsc_0_1_i_q_d),
      .vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_2_i_q_d(vec_rsc_0_2_i_q_d),
      .vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_3_i_q_d(vec_rsc_0_3_i_q_d),
      .vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_4_i_q_d(vec_rsc_0_4_i_q_d),
      .vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_5_i_q_d(vec_rsc_0_5_i_q_d),
      .vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_6_i_q_d(vec_rsc_0_6_i_q_d),
      .vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_7_i_q_d(vec_rsc_0_7_i_q_d),
      .vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_8_i_q_d(vec_rsc_0_8_i_q_d),
      .vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_9_i_q_d(vec_rsc_0_9_i_q_d),
      .vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_10_i_q_d(vec_rsc_0_10_i_q_d),
      .vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_11_i_q_d(vec_rsc_0_11_i_q_d),
      .vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_12_i_q_d(vec_rsc_0_12_i_q_d),
      .vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_13_i_q_d(vec_rsc_0_13_i_q_d),
      .vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_14_i_q_d(vec_rsc_0_14_i_q_d),
      .vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_15_i_q_d(vec_rsc_0_15_i_q_d),
      .vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_0_i_q_d(twiddle_rsc_0_0_i_q_d),
      .twiddle_rsc_0_0_i_radr_d(twiddle_rsc_0_0_i_radr_d),
      .twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_1_i_q_d(twiddle_rsc_0_1_i_q_d),
      .twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_2_i_q_d(twiddle_rsc_0_2_i_q_d),
      .twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_3_i_q_d(twiddle_rsc_0_3_i_q_d),
      .twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_4_i_q_d(twiddle_rsc_0_4_i_q_d),
      .twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_5_i_q_d(twiddle_rsc_0_5_i_q_d),
      .twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_6_i_q_d(twiddle_rsc_0_6_i_q_d),
      .twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_7_i_q_d(twiddle_rsc_0_7_i_q_d),
      .twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_8_i_q_d(twiddle_rsc_0_8_i_q_d),
      .twiddle_rsc_0_8_i_radr_d(twiddle_rsc_0_8_i_radr_d),
      .twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_9_i_q_d(twiddle_rsc_0_9_i_q_d),
      .twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_10_i_q_d(twiddle_rsc_0_10_i_q_d),
      .twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_11_i_q_d(twiddle_rsc_0_11_i_q_d),
      .twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_12_i_q_d(twiddle_rsc_0_12_i_q_d),
      .twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_13_i_q_d(twiddle_rsc_0_13_i_q_d),
      .twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_14_i_q_d(twiddle_rsc_0_14_i_q_d),
      .twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_15_i_q_d(twiddle_rsc_0_15_i_q_d),
      .twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_0_i_d_d_pff(vec_rsc_0_0_i_d_d_iff),
      .vec_rsc_0_0_i_radr_d_pff(vec_rsc_0_0_i_radr_d_iff),
      .vec_rsc_0_0_i_wadr_d_pff(vec_rsc_0_0_i_wadr_d_iff),
      .vec_rsc_0_0_i_we_d_pff(vec_rsc_0_0_i_we_d_iff),
      .vec_rsc_0_1_i_we_d_pff(vec_rsc_0_1_i_we_d_iff),
      .vec_rsc_0_2_i_we_d_pff(vec_rsc_0_2_i_we_d_iff),
      .vec_rsc_0_3_i_we_d_pff(vec_rsc_0_3_i_we_d_iff),
      .vec_rsc_0_4_i_we_d_pff(vec_rsc_0_4_i_we_d_iff),
      .vec_rsc_0_5_i_we_d_pff(vec_rsc_0_5_i_we_d_iff),
      .vec_rsc_0_6_i_we_d_pff(vec_rsc_0_6_i_we_d_iff),
      .vec_rsc_0_7_i_we_d_pff(vec_rsc_0_7_i_we_d_iff),
      .vec_rsc_0_8_i_we_d_pff(vec_rsc_0_8_i_we_d_iff),
      .vec_rsc_0_9_i_we_d_pff(vec_rsc_0_9_i_we_d_iff),
      .vec_rsc_0_10_i_we_d_pff(vec_rsc_0_10_i_we_d_iff),
      .vec_rsc_0_11_i_we_d_pff(vec_rsc_0_11_i_we_d_iff),
      .vec_rsc_0_12_i_we_d_pff(vec_rsc_0_12_i_we_d_iff),
      .vec_rsc_0_13_i_we_d_pff(vec_rsc_0_13_i_we_d_iff),
      .vec_rsc_0_14_i_we_d_pff(vec_rsc_0_14_i_we_d_iff),
      .vec_rsc_0_15_i_we_d_pff(vec_rsc_0_15_i_we_d_iff),
      .twiddle_rsc_0_1_i_radr_d_pff(twiddle_rsc_0_1_i_radr_d_iff),
      .twiddle_rsc_0_2_i_radr_d_pff(twiddle_rsc_0_2_i_radr_d_iff),
      .twiddle_rsc_0_4_i_radr_d_pff(twiddle_rsc_0_4_i_radr_d_iff)
    );
endmodule



