// check_properties -prop -list spec.prop_ovf_spec_wrapper_ln65_1 ; # ( ovf ) (l1=1, l2=0)
module GOTH_58 ( M1TU__P_18_14 , M1TU__P_36_15 , M1TU__clk , M1TU__asm_sym_data_21
 , M1TU__asm_sym_data_17 , M1TU__OOB_X_1 , M1TU__asm_sym_data_16 , M1TU__OOB_X_2
 , M1TU__asm_sym_data_11 , M1TU__asm_sym_data_8 , M1TU__asm_sym_data_9 , M1TU__asm_sym_data_10
 , M1TU__OOB_X_3 , M1TU__asm_sym_data_3 , M1TU__asm_sym_data_0 , M1TU__asm_sym_data_1
 , M1TU__asm_sym_data_2 , M1TU__OOB_X_4 , M1TU__P_56 , M1TU__OOB_X_6 , M1TU__asm_sym_data_20
 , M1TU__OOB_X_7 , M1TU__OOB_X_8 , M1TU__OOB_X_9 ) ;
 input wire  M1TU__clk ; 
 input wire  [31:0]  M1TU__asm_sym_data_21 ; 
 input wire  [31:0]  M1TU__asm_sym_data_17 ; 
 input wire  [31:0]  M1TU__OOB_X_1 ; 
 input wire  [31:0]  M1TU__asm_sym_data_16 ; 
 input wire  [31:0]  M1TU__OOB_X_2 ; 
 input wire  [31:0]  M1TU__asm_sym_data_11 ; 
 input wire  [31:0]  M1TU__asm_sym_data_8 ; 
 input wire  [31:0]  M1TU__asm_sym_data_9 ; 
 input wire  [31:0]  M1TU__asm_sym_data_10 ; 
 input wire  [31:0]  M1TU__OOB_X_3 ; 
 input wire  [31:0]  M1TU__asm_sym_data_3 ; 
 input wire  [31:0]  M1TU__asm_sym_data_0 ; 
 input wire  [31:0]  M1TU__asm_sym_data_1 ; 
 input wire  [31:0]  M1TU__asm_sym_data_2 ; 
 input wire  [31:0]  M1TU__OOB_X_4 ; 
 input wire  [31:0]  M1TU__P_56 ; 
 input wire  [31:0]  M1TU__OOB_X_6 ; 
 input wire  [31:0]  M1TU__asm_sym_data_20 ; 
 input wire  [31:0]  M1TU__OOB_X_7 ; 
 input wire  [31:0]  M1TU__OOB_X_8 ; 
 input wire  [31:0]  M1TU__OOB_X_9 ; 
 output wire  M1TU__P_18_14 ; 
 output wire  [0:0]  M1TU__P_36_15 ; 
 wire  [0:0] E_48092 ; 
assign M1TU__P_36_15 = E_48092 ;
 wire  [0:0] E_48220 ; 
assign M1TU__P_18_14 = E_48220 ;
 wire  [0:0] E_47863 ; 
 wire  [0:0] E_47862 ; 
 wire  [0:0] E_47861 ; 
 wire  [32:0] E_48018 ; 
 wire  [31:0] E_48055 ; 
 wire  [0:0] E_48412 ; 
 wire  [19:0] E_51353 ; 
 wire  [19:0] E_48053 ; 
 wire  [18:0] E_48052 ; 
 wire  [19:0] E_48016 ; 
 wire  [0:0] E_48170 ; 
 wire  [0:0] E_48169 ; 
 wire  [0:0] E_48168 ; 
 wire  [19:0] E_48167 ; 
 wire  [19:0] E_48068 ; 
 wire  [0:0] E_48165 ; 
 wire  [0:0] E_48164 ; 
 wire  [2:0] E_48189 ; 
 wire  [2:0] E_48205 ; 
 wire  [0:0] E_48203 ; 
 wire  [0:0] E_48202 ; 
 wire  [0:0] E_48201 ; 
 wire  [0:0] E_48200 ; 
 wire  [0:0] E_48199 ; 
 wire  [19:0] E_48198 ; 
 wire  [19:0] E_48197 ; 
 wire  [0:0] E_48196 ; 
 wire  [0:0] E_48195 ; 
 wire  [0:0] E_48194 ; 
 wire  [19:0] E_48193 ; 
 wire  [19:0] E_47976 ; 
 wire  [0:0] E_48191 ; 
 wire  [0:0] E_48190 ; 
 wire  [2:0] E_48188 ; 
 wire  [0:0] E_48187 ; 
 wire  [0:0] E_48186 ; 
 wire  [0:0] E_48185 ; 
 wire  [0:0] E_48184 ; 
 wire  [19:0] E_48183 ; 
 wire  signed  [20:0] E_48036 ; 
 wire  [19:0] E_48182 ; 
 wire  [0:0] E_48181 ; 
 wire  [0:0] E_48115 ; 
 wire  [19:0] E_48179 ; 
 wire  [19:0] E_48206 ; 
 wire  [19:0] E_48141 ; 
 wire  [0:0] E_48175 ; 
 wire  [0:0] E_48174 ; 
 wire  [0:0] E_48173 ; 
 wire  [19:0] E_48172 ; 
 wire  [9:0] E_48075 ; 
 wire  [0:0] E_48156 ; 
 wire  [0:0] E_48155 ; 
 wire  [1:0] E_47804 ; 
 wire  [19:0] E_48142 ; 
 wire  signed  [20:0] E_47957 ; 
 wire  [1:0] E_47806 ; 
 wire clk ; 
assign clk = M1TU__clk ;
 wire  [19:0] E_48253 ; 
 wire  [19:0] E_48178_68655 ; 
 wire  [3:0] E_48178 ; 
 wire  [2:0] E_48176 ; 
 wire  [0:0] E_48152 ; 
 wire  [19:0] E_48151 ; 
 wire  [19:0] E_48209 ; 
 wire  [0:0] E_48150 ; 
 wire  [0:0] E_48149 ; 
 wire  [2:0] E_48148 ; 
 wire  [19:0] E_48256 ; 
 wire  [19:0] E_48092_68651 ; 
 wire  [19:0] E_48147 ; 
 wire  [19:0] E_48210 ; 
 wire  [0:0] E_48146 ; 
 wire  [0:0] E_48145 ; 
 wire  [19:0] E_48257 ; 
 wire  [0:0] E_48144 ; 
 wire  [0:0] E_48143 ; 
 wire  [0:0] E_48140 ; 
 wire  [0:0] E_48139 ; 
 wire  [2:0] E_47813 ; 
 wire  [2:0] E_47812 ; 
 wire  [2:0] E_47811 ; 
 wire  [2:0] E_47810 ; 
 wire  [0:0] E_48159 ; 
 wire  [0:0] E_48158 ; 
 wire  [2:0] E_47809 ; 
 wire  [0:0] E_48136 ; 
 wire  [2:0] E_48115_68642 ; 
 wire  [2:0] E_47807 ; 
 wire  [2:0] E_47806_68640 ; 
 wire  [2:0] E_47805 ; 
 wire  [2:0] E_47804_68639 ; 
 wire  [2:0] E_47803 ; 
 wire  [2:0] E_48163 ; 
 wire  [2:0] E_47802 ; 
 wire  [2:0] E_47801 ; 
 wire  [2:0] E_47800 ; 
 wire  [2:0] E_60005 ; 
 wire  [19:0] E_48162 ; 
 wire  [19:0] E_48207 ; 
 wire  [19:0] E_48254 ; 
 wire  [19:0] E_48157 ; 
 wire  [19:0] E_48208 ; 
 wire  [19:0] E_48255 ; 
 wire  [9:0] E_51065 ; 
 wire  [31:0] E_48055_clone_48407 ; 
 wire  [31:0] asm_sym_data_21 ; 
assign asm_sym_data_21 = M1TU__asm_sym_data_21 ;
 wire  [31:0] E_49059 ; 
 wire  [0:0] E_49046 ; 
 wire  [20:0] E_48076 ; 
 wire  [31:0] E_49057 ; 
 wire  [0:0] E_51058 ; 
 wire  [31:0] E_48073 ; 
 wire  [0:0] E_48072 ; 
 wire  [31:0] E_48071 ; 
 wire  [31:0] E_48120 ; 
 wire  [0:0] E_48347 ; 
 wire  [19:0] E_51359 ; 
 wire  [19:0] E_48117 ; 
 wire  [18:0] E_48116 ; 
 wire  [31:0] E_48120_clone_48342 ; 
assign E_48120_clone_48342 = M1TU__asm_sym_data_17 ;
 wire  [31:0] OOB_X_1 ; 
assign OOB_X_1 = M1TU__OOB_X_1 ;
 wire  [31:0] E_48114 ; 
 wire  [0:0] E_48113 ; 
 wire  [31:0] E_48112 ; 
 wire  [31:0] E_48110 ; 
 wire  [31:0] E_48108 ; 
 wire  [31:0] E_48108_clone_48355 ; 
assign E_48108_clone_48355 = M1TU__asm_sym_data_16 ;
 wire  [31:0] OOB_X_2 ; 
assign OOB_X_2 = M1TU__OOB_X_2 ;
 wire  [31:0] E_48106 ; 
 wire  [0:0] E_48373 ; 
 wire  [19:0] E_51357 ; 
 wire  [19:0] E_48102 ; 
 wire  [19:0] E_48101 ; 
 wire  [19:0] E_48040 ; 
 wire  [19:0] E_48039 ; 
 wire  signed  [31:0] E_48038 ; 
 wire  [0:0] E_48037 ; 
 wire  [5:0] E_48096 ; 
 wire  signed  [31:0] E_48035_68647 ; 
 wire  [31:0] E_48035 ; 
 wire  signed  [0:0] E_48093 ; 
 wire  signed  [31:0] E_48092_68644 ; 
 wire  [19:0] E_48258 ; 
 wire  [19:0] E_48100 ; 
 wire  [0:0] E_48098 ; 
 wire  signed  [20:0] E_48097 ; 
 wire  [19:0] E_48095 ; 
 wire  [31:0] E_48106_clone_48368 ; 
 wire  [0:0] E_51002 ; 
 wire  [19:0] E_51351 ; 
 wire  [31:0] E_50825 ; 
 wire  [0:0] E_51018 ; 
 wire  [19:0] E_51345 ; 
 wire  [19:0] E_48001 ; 
 wire  [19:0] E_48000 ; 
 wire  [19:0] E_47961 ; 
 wire  [19:0] E_47960 ; 
 wire  signed  [31:0] E_47959 ; 
 wire  [0:0] E_47958 ; 
 wire  signed  [31:0] E_47956_68643 ; 
 wire  [31:0] E_47956 ; 
 wire  [19:0] E_48260 ; 
 wire  [19:0] E_47999 ; 
 wire  signed  [31:0] E_47998 ; 
 wire  [0:0] E_47997 ; 
 wire  signed  [20:0] E_47996 ; 
 wire  signed  [31:0] E_47995_68645 ; 
 wire  [31:0] E_47995 ; 
 wire  [31:0] E_50829 ; 
 wire  [0:0] E_51038 ; 
 wire  [19:0] E_51339 ; 
 wire  [31:0] asm_sym_data_11 ; 
assign asm_sym_data_11 = M1TU__asm_sym_data_11 ;
 wire  [31:0] asm_sym_data_8 ; 
assign asm_sym_data_8 = M1TU__asm_sym_data_8 ;
 wire  [31:0] E_50905 ; 
 wire  [0:0] E_51014 ; 
 wire  [31:0] asm_sym_data_9 ; 
assign asm_sym_data_9 = M1TU__asm_sym_data_9 ;
 wire  [31:0] E_50865 ; 
 wire  [0:0] E_50994 ; 
 wire  [31:0] E_50869 ; 
 wire  [0:0] E_50998 ; 
 wire  [31:0] asm_sym_data_10 ; 
assign asm_sym_data_10 = M1TU__asm_sym_data_10 ;
 wire  [31:0] OOB_X_3 ; 
assign OOB_X_3 = M1TU__OOB_X_3 ;
 wire  [31:0] E_48091 ; 
 wire  [31:0] E_48089 ; 
 wire  [51:0] E_48087 ; 
 wire  [31:0] E_48086 ; 
 wire  [31:0] E_48086_clone_48381 ; 
 wire  [31:0] E_51037 ; 
 wire  [31:0] E_51041 ; 
 wire  [31:0] asm_sym_data_3 ; 
assign asm_sym_data_3 = M1TU__asm_sym_data_3 ;
 wire  [31:0] E_47949_clone_48524 ; 
assign E_47949_clone_48524 = M1TU__asm_sym_data_0 ;
 wire  [31:0] E_51053 ; 
 wire  [31:0] asm_sym_data_1 ; 
assign asm_sym_data_1 = M1TU__asm_sym_data_1 ;
 wire  [31:0] E_48028_clone_48446 ; 
 wire  [31:0] E_51049 ; 
 wire  [31:0] asm_sym_data_2 ; 
assign asm_sym_data_2 = M1TU__asm_sym_data_2 ;
 wire  [31:0] OOB_X_4 ; 
assign OOB_X_4 = M1TU__OOB_X_4 ;
 wire  [4:0] E_48084 ; 
 wire  [31:0] E_48083 ; 
 wire  [31:0] E_48082 ; 
 wire  [31:0] E_48259 ; 
 wire  [31:0] E_48081 ; 
assign E_48081 = M1TU__P_56 ;
 wire  [31:0] E_48080 ; 
 wire  signed  [32:0] E_48079 ; 
 wire  [31:0] E_48069 ; 
 wire  [31:0] E_48124 ; 
 wire  [0:0] E_48123 ; 
 wire  signed  [31:0] E_48122 ; 
 wire  [31:0] E_48122_68652 ; 
 wire  [31:0] E_48077 ; 
 wire  [31:0] OOB_X_6 ; 
assign OOB_X_6 = M1TU__OOB_X_6 ;
 wire  [31:0] E_48051 ; 
 wire  [0:0] E_48050 ; 
 wire  [31:0] E_48049 ; 
 wire  signed  [32:0] E_48048 ; 
 wire  [31:0] E_48047 ; 
 wire  [63:0] E_48046 ; 
 wire  [31:0] E_48045 ; 
 wire  [31:0] E_48045_clone_48420 ; 
 wire  [31:0] asm_sym_data_20 ; 
assign asm_sym_data_20 = M1TU__asm_sym_data_20 ;
 wire  [31:0] E_49053 ; 
 wire  [0:0] E_49037 ; 
 wire  [31:0] E_49051 ; 
 wire  [0:0] E_51057 ; 
 wire  [31:0] OOB_X_7 ; 
assign OOB_X_7 = M1TU__OOB_X_7 ;
 wire  [31:0] E_48043 ; 
 wire  [0:0] E_48438 ; 
 wire  [31:0] E_48043_clone_48433 ; 
 wire  [31:0] E_50681 ; 
 wire  [31:0] E_47964_clone_48511 ; 
 wire  [31:0] E_50781 ; 
 wire  [31:0] E_48004_clone_48472 ; 
 wire  [31:0] E_50733 ; 
 wire  [31:0] OOB_X_8 ; 
assign OOB_X_8 = M1TU__OOB_X_8 ;
 wire  [31:0] E_48033 ; 
 wire  [63:0] E_48032 ; 
 wire  [31:0] E_48031 ; 
 wire  [43:0] E_48030 ; 
 wire  [63:0] E_48029 ; 
 wire  [31:0] E_48028 ; 
 wire  [31:0] OOB_X_9 ; 
assign OOB_X_9 = M1TU__OOB_X_9 ;
 wire  [31:0] E_48027 ; 
 wire  signed  [32:0] E_48026 ; 
 wire  [31:0] E_47937 ; 
 wire  [0:0] E_47860 ; 
      assign E_48092 = 1'h0;
    CPL_MUX_2  I_47710 ( .o ( E_48220 )  , .s ( E_47863 )  , .d0 ( E_47860 )  , .d1 ( E_48115 )  );
    CPL_LAND  I_47709 ( .o ( E_47863 )  , .l ( E_47862 )  , .r ( E_48156 )  );
    CPL_NOT  I_47708 ( .o ( E_47862 )  , .l ( E_47861 )  );
    CPL_LE  I_47707 ( .o ( E_47861 )  , .l ( E_48018 )  , .r ( E_47937 )  );
    CPL_ADD  I_47863 ( .o ( E_48018 )  , .l ( E_48055 )  , .r ( E_48051 )  );
    CPL_MUX_2  I_48200 ( .o ( E_48055 )  , .s ( E_48412 )  , .d0 ( E_48055_clone_48407 )  , 
		.d1 ( OOB_X_6 )  );
    CPL_GT  I_48205 ( .o ( E_48412 )  , .l ( E_51353 )  , .r ( E_51065 )  );
    CPL_ADD  I_47889 ( .o ( E_51353 )  , .l ( E_48053 )  , .r ( E_48115 )  );
    CPL_LASFT  I_47898 ( .o ( E_48053 )  , .d ( E_48052 )  , .s ( E_48115 )  );
    CPL_TYPE  I_51609 ( .o ( E_48052 )  , .l ( E_48016 )  );
    CPL_MUX_2  I_48005 ( .o ( E_48016 )  , .s ( E_48170 )  , .d0 ( E_48157 )  , .d1 ( E_48092_68651 )  );
    CPL_LAND  I_48004 ( .o ( E_48170 )  , .l ( E_48169 )  , .r ( E_48159 )  );
    CPL_NOT  I_48003 ( .o ( E_48169 )  , .l ( E_48168 )  );
    CPL_LT  I_48002 ( .o ( E_48168 )  , .l ( E_48167 )  , .r ( E_48075 )  );
    CPL_ADD  I_48001 ( .o ( E_48167 )  , .l ( E_48068 )  , .r ( E_48115 )  );
    CPL_MUX_2  I_48000 ( .o ( E_48068 )  , .s ( E_48165 )  , .d0 ( E_48162 )  , .d1 ( E_48092_68651 )  );
    CPL_LOR  I_47999 ( .o ( E_48165 )  , .l ( E_48164 )  , .r ( E_48181 )  );
    CPL_EQ  I_47998 ( .o ( E_48164 )  , .l ( E_48189 )  , .r ( E_48163 )  );
    CPL_FF#3  I_48047_reg ( .q ( E_48189 )  , .qbar (  )  , .d ( E_48205 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_60005 )  );
    CPL_MUX_2  I_47653 ( .o ( E_48205 )  , .s ( E_48203 )  , .d0 ( E_47813 )  , .d1 ( E_48115_68642 )  );
    CPL_LOR  I_48035 ( .o ( E_48203 )  , .l ( E_48202 )  , .r ( E_48140 )  );
    CPL_MUX_2  I_48034 ( .o ( E_48202 )  , .s ( E_48201 )  , .d0 ( E_48092 )  , .d1 ( E_48144 )  );
    CPL_LAND  I_48033 ( .o ( E_48201 )  , .l ( E_48200 )  , .r ( E_48146 )  );
    CPL_NOT  I_48032 ( .o ( E_48200 )  , .l ( E_48199 )  );
    CPL_LT  I_48031 ( .o ( E_48199 )  , .l ( E_48198 )  , .r ( E_48075 )  );
    CPL_ADD  I_48030 ( .o ( E_48198 )  , .l ( E_48197 )  , .r ( E_48115 )  );
    CPL_MUX_2  I_48029 ( .o ( E_48197 )  , .s ( E_48196 )  , .d0 ( E_48147 )  , .d1 ( E_48092_68651 )  );
    CPL_LAND  I_48028 ( .o ( E_48196 )  , .l ( E_48195 )  , .r ( E_48150 )  );
    CPL_NOT  I_48027 ( .o ( E_48195 )  , .l ( E_48194 )  );
    CPL_LT  I_48026 ( .o ( E_48194 )  , .l ( E_48193 )  , .r ( E_48075 )  );
    CPL_ADD  I_48025 ( .o ( E_48193 )  , .l ( E_47976 )  , .r ( E_48115 )  );
    CPL_MUX_2  I_48024 ( .o ( E_47976 )  , .s ( E_48191 )  , .d0 ( E_48151 )  , .d1 ( E_48092_68651 )  );
    CPL_LOR  I_48023 ( .o ( E_48191 )  , .l ( E_48190 )  , .r ( E_48187 )  );
    CPL_EQ  I_48022 ( .o ( E_48190 )  , .l ( E_48189 )  , .r ( E_48188 )  );
      assign E_48188 = 3'h7;
    CPL_MUX_2  I_48020 ( .o ( E_48187 )  , .s ( E_48186 )  , .d0 ( E_48092 )  , .d1 ( E_48152 )  );
    CPL_LAND  I_48019 ( .o ( E_48186 )  , .l ( E_48185 )  , .r ( E_48175 )  );
    CPL_NOT  I_48018 ( .o ( E_48185 )  , .l ( E_48184 )  );
    CPL_GE  I_48017 ( .o ( E_48184 )  , .l ( E_48183 )  , .r ( E_48176 )  );
    CPL_TYPE  I_51614 ( .o ( E_48183 )  , .l ( E_48036 )  );
    CPL_SUB  I_47881 ( .o ( E_48036 )  , .l ( E_48182 )  , .r ( E_47806 )  );
    CPL_MUX_2  I_48015 ( .o ( E_48182 )  , .s ( E_48181 )  , .d0 ( E_48179 )  , .d1 ( E_48178_68655 )  );
    CPL_EQ  I_48014 ( .o ( E_48181 )  , .l ( E_48189 )  , .r ( E_48115 )  );
      assign E_48115 = 1'h1;
    CPL_FF#20  I_48049_reg ( .q ( E_48179 )  , .qbar (  )  , .d ( E_48206 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48253 )  );
    CPL_MUX_2  I_47654 ( .o ( E_48206 )  , .s ( E_48201 )  , .d0 ( E_48141 )  , .d1 ( E_48142 )  );
    CPL_MUX_2  I_47979 ( .o ( E_48141 )  , .s ( E_48175 )  , .d0 ( E_48182 )  , .d1 ( E_48183 )  );
    CPL_LAND  I_48009 ( .o ( E_48175 )  , .l ( E_48174 )  , .r ( E_48156 )  );
    CPL_NOT  I_48008 ( .o ( E_48174 )  , .l ( E_48173 )  );
    CPL_LT  I_48007 ( .o ( E_48173 )  , .l ( E_48172 )  , .r ( E_48075 )  );
    CPL_ADD  I_48006 ( .o ( E_48172 )  , .l ( E_48016 )  , .r ( E_48115 )  );
      assign E_48075 = 10'h200;
    CPL_LOR  I_47992 ( .o ( E_48156 )  , .l ( E_48155 )  , .r ( E_48170 )  );
    CPL_EQ  I_47991 ( .o ( E_48155 )  , .l ( E_48189 )  , .r ( E_47804 )  );
      assign E_47804 = 2'h3;
    CPL_TYPE  I_51597 ( .o ( E_48142 )  , .l ( E_47957 )  );
    CPL_SUB  I_47803 ( .o ( E_47957 )  , .l ( E_48141 )  , .r ( E_47806 )  );
      assign E_47806 = 2'h2;
      assign E_48253 = 20'hX; /*CDBImplicitXNone*/
    CPL_TYPE  I_69221 ( .o ( E_48178_68655 )  , .l ( E_48178 )  );
      assign E_48178 = 4'ha;
      assign E_48176 = 3'h6;
    CPL_GE  I_47988 ( .o ( E_48152 )  , .l ( E_48183 )  , .r ( E_47806 )  );
    CPL_FF#20  I_48054_reg ( .q ( E_48151 )  , .qbar (  )  , .d ( E_48209 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48256 )  );
    CPL_MUX_2  I_47657 ( .o ( E_48209 )  , .s ( E_48150 )  , .d0 ( E_47976 )  , .d1 ( E_48193 )  );
    CPL_LOR  I_47987 ( .o ( E_48150 )  , .l ( E_48149 )  , .r ( E_48191 )  );
    CPL_EQ  I_47986 ( .o ( E_48149 )  , .l ( E_48189 )  , .r ( E_48148 )  );
      assign E_48148 = 3'h5;
      assign E_48256 = 20'hX; /*CDBImplicitXNone*/
    CPL_TYPE  I_69217 ( .o ( E_48092_68651 )  , .l ( E_48092 )  );
    CPL_FF#20  I_48056_reg ( .q ( E_48147 )  , .qbar (  )  , .d ( E_48210 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48257 )  );
    CPL_MUX_2  I_47658 ( .o ( E_48210 )  , .s ( E_48146 )  , .d0 ( E_48197 )  , .d1 ( E_48198 )  );
    CPL_LOR  I_47984 ( .o ( E_48146 )  , .l ( E_48145 )  , .r ( E_48196 )  );
    CPL_EQ  I_47983 ( .o ( E_48145 )  , .l ( E_48189 )  , .r ( E_48176 )  );
      assign E_48257 = 20'hX; /*CDBImplicitXNone*/
    CPL_NOT  I_47982 ( .o ( E_48144 )  , .l ( E_48143 )  );
    CPL_GE  I_47981 ( .o ( E_48143 )  , .l ( E_48142 )  , .r ( E_47806 )  );
    CPL_MUX_2  I_47978 ( .o ( E_48140 )  , .s ( E_48186 )  , .d0 ( E_48092 )  , .d1 ( E_48139 )  );
    CPL_NOT  I_47977 ( .o ( E_48139 )  , .l ( E_48152 )  );
    CPL_MUX_2  I_47652 ( .o ( E_47813 )  , .s ( E_48146 )  , .d0 ( E_47812 )  , .d1 ( E_47801 )  );
    CPL_MUX_2  I_47651 ( .o ( E_47812 )  , .s ( E_48150 )  , .d0 ( E_47811 )  , .d1 ( E_47802 )  );
    CPL_MUX_2  I_47650 ( .o ( E_47811 )  , .s ( E_48156 )  , .d0 ( E_47810 )  , .d1 ( E_47805 )  );
    CPL_MUX_2  I_47649 ( .o ( E_47810 )  , .s ( E_48159 )  , .d0 ( E_47809 )  , .d1 ( E_47807 )  );
    CPL_LOR  I_47994 ( .o ( E_48159 )  , .l ( E_48158 )  , .r ( E_48165 )  );
    CPL_EQ  I_47993 ( .o ( E_48158 )  , .l ( E_48189 )  , .r ( E_47806 )  );
    CPL_MUX_2  I_47648 ( .o ( E_47809 )  , .s ( E_48136 )  , .d0 ( E_48189 )  , .d1 ( E_48115_68642 )  );
    CPL_EQ  I_47974 ( .o ( E_48136 )  , .l ( E_48189 )  , .r ( E_48092 )  );
    CPL_TYPE  I_69208 ( .o ( E_48115_68642 )  , .l ( E_48115 )  );
    CPL_MUX_2  I_47646 ( .o ( E_47807 )  , .s ( E_48169 )  , .d0 ( E_47806_68640 )  , .d1 ( E_47809 )  );
    CPL_TYPE  I_69206 ( .o ( E_47806_68640 )  , .l ( E_47806 )  );
    CPL_MUX_2  I_47644 ( .o ( E_47805 )  , .s ( E_48174 )  , .d0 ( E_47804_68639 )  , .d1 ( E_47803 )  );
    CPL_TYPE  I_69205 ( .o ( E_47804_68639 )  , .l ( E_47804 )  );
    CPL_MUX_2  I_47642 ( .o ( E_47803 )  , .s ( E_48185 )  , .d0 ( E_48163 )  , .d1 ( E_47810 )  );
      assign E_48163 = 3'h4;
    CPL_MUX_2  I_47641 ( .o ( E_47802 )  , .s ( E_48195 )  , .d0 ( E_48148 )  , .d1 ( E_47811 )  );
    CPL_MUX_2  I_47640 ( .o ( E_47801 )  , .s ( E_48200 )  , .d0 ( E_48176 )  , .d1 ( E_47800 )  );
    CPL_MUX_2  I_47639 ( .o ( E_47800 )  , .s ( E_48144 )  , .d0 ( E_48188 )  , .d1 ( E_47812 )  );
      assign E_60005 = 3'h1;
    CPL_FF#20  I_48050_reg ( .q ( E_48162 )  , .qbar (  )  , .d ( E_48207 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48254 )  );
    CPL_MUX_2  I_47655 ( .o ( E_48207 )  , .s ( E_48159 )  , .d0 ( E_48068 )  , .d1 ( E_48167 )  );
      assign E_48254 = 20'hX; /*CDBImplicitXNone*/
    CPL_FF#20  I_48052_reg ( .q ( E_48157 )  , .qbar (  )  , .d ( E_48208 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48255 )  );
    CPL_MUX_2  I_47656 ( .o ( E_48208 )  , .s ( E_48156 )  , .d0 ( E_48016 )  , .d1 ( E_48172 )  );
      assign E_48255 = 20'hX; /*CDBImplicitXNone*/
      assign E_51065 = 10'h3ff;
    CPL_MUX_2  I_48957 ( .o ( E_48055_clone_48407 )  , .s ( E_48159 )  , .d0 ( asm_sym_data_21 )  , 
		.d1 ( E_49059 )  );
    CPL_MUX_2  I_48956 ( .o ( E_49059 )  , .s ( E_49046 )  , .d0 ( E_49057 )  , .d1 ( E_48124 )  );
    CPL_EQ  I_48941 ( .o ( E_49046 )  , .l ( E_48076 )  , .r ( E_48053 )  );
    CPL_ADD  I_47921 ( .o ( E_48076 )  , .l ( E_48068 )  , .r ( E_48075 )  );
    CPL_MUX_2  I_48954 ( .o ( E_49057 )  , .s ( E_51058 )  , .d0 ( asm_sym_data_21 )  , 
		.d1 ( E_48073 )  );
    CPL_EQ  I_48938 ( .o ( E_51058 )  , .l ( E_48068 )  , .r ( E_48053 )  );
    CPL_MUX_2  I_47918 ( .o ( E_48073 )  , .s ( E_48072 )  , .d0 ( E_48071 )  , .d1 ( E_48069 )  );
    CPL_GT  I_47917 ( .o ( E_48072 )  , .l ( E_48071 )  , .r ( E_48083 )  );
    CPL_ADD  I_47915 ( .o ( E_48071 )  , .l ( E_48120 )  , .r ( E_48114 )  );
    CPL_MUX_2  I_48135 ( .o ( E_48120 )  , .s ( E_48347 )  , .d0 ( E_48120_clone_48342 )  , 
		.d1 ( OOB_X_1 )  );
    CPL_GT  I_48140 ( .o ( E_48347 )  , .l ( E_51359 )  , .r ( E_51065 )  );
    CPL_ADD  I_47947 ( .o ( E_51359 )  , .l ( E_48117 )  , .r ( E_48115 )  );
    CPL_LASFT  I_47957 ( .o ( E_48117 )  , .d ( E_48116 )  , .s ( E_48115 )  );
    CPL_TYPE  I_51620 ( .o ( E_48116 )  , .l ( E_48068 )  );
    CPL_MUX_2  I_47954 ( .o ( E_48114 )  , .s ( E_48113 )  , .d0 ( E_48112 )  , .d1 ( E_48080 )  );
    CPL_GE  I_47953 ( .o ( E_48113 )  , .l ( E_48112 )  , .r ( E_48083 )  );
    CPL_SUB  I_47951 ( .o ( E_48112 )  , .l ( E_48110 )  , .r ( E_48091 )  );
    CPL_MULT  I_47949 ( .o ( E_48110 )  , .l ( E_48108 )  , .r ( E_48106 )  );
    CPL_MUX_2  I_48148 ( .o ( E_48108 )  , .s ( E_48347 )  , .d0 ( E_48108_clone_48355 )  , 
		.d1 ( OOB_X_2 )  );
    CPL_MUX_2  I_48161 ( .o ( E_48106 )  , .s ( E_48373 )  , .d0 ( E_48106_clone_48368 )  , 
		.d1 ( OOB_X_3 )  );
    CPL_GT  I_48166 ( .o ( E_48373 )  , .l ( E_51357 )  , .r ( E_51065 )  );
    CPL_AND  I_47944 ( .o ( E_51357 )  , .l ( E_48102 )  , .r ( E_48068 )  );
    CPL_MUX_2  I_47943 ( .o ( E_48102 )  , .s ( E_48165 )  , .d0 ( E_48101 )  , .d1 ( E_48100 )  );
    CPL_FF#20  I_48058_reg ( .q ( E_48101 )  , .qbar (  )  , .d ( E_48040 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48258 )  );
    CPL_MUX_2  I_47885 ( .o ( E_48040 )  , .s ( E_48170 )  , .d0 ( E_48102 )  , .d1 ( E_48039 )  );
    CPL_TYPE  I_51615 ( .o ( E_48039 )  , .l ( E_48038 )  );
    CPL_MUX_2  I_47883 ( .o ( E_48038 )  , .s ( E_48037 )  , .d0 ( E_48035_68647 )  , .d1 ( E_48092_68644 )  );
    CPL_GT  I_47882 ( .o ( E_48037 )  , .l ( E_48036 )  , .r ( E_48096 )  );
      assign E_48096 = 6'h20;
    CPL_TYPE  I_69213 ( .o ( E_48035_68647 )  , .l ( E_48035 )  );
    CPL_LASFT  I_47879 ( .o ( E_48035 )  , .d ( E_48093 )  , .s ( E_48036 )  );
      assign E_48093 = 1'sh1;
    CPL_TYPE  I_69210 ( .o ( E_48092_68644 )  , .l ( E_48092 )  );
      assign E_48258 = 20'hX; /*CDBImplicitXNone*/
    CPL_MUX_2  I_47941 ( .o ( E_48100 )  , .s ( E_48098 )  , .d0 ( E_48095 )  , .d1 ( E_48092_68651 )  );
    CPL_GT  I_47940 ( .o ( E_48098 )  , .l ( E_48097 )  , .r ( E_48096 )  );
    CPL_SUB  I_47939 ( .o ( E_48097 )  , .l ( E_48182 )  , .r ( E_48115 )  );
    CPL_LASFT  I_47936 ( .o ( E_48095 )  , .d ( E_48093 )  , .s ( E_48097 )  );
    CPL_MUX_2  I_51145 ( .o ( E_48106_clone_48368 )  , .s ( E_51002 )  , .d0 ( E_50825 )  , 
		.d1 ( E_50865 )  );
    CPL_EQ  I_51372 ( .o ( E_51002 )  , .l ( E_51351 )  , .r ( E_51357 )  );
    CPL_AND  I_47886 ( .o ( E_51351 )  , .l ( E_48040 )  , .r ( E_48016 )  );
    CPL_MUX_2  I_51150 ( .o ( E_50825 )  , .s ( E_51018 )  , .d0 ( E_50829 )  , .d1 ( E_50905 )  );
    CPL_EQ  I_51392 ( .o ( E_51018 )  , .l ( E_51345 )  , .r ( E_51357 )  );
    CPL_AND  I_47847 ( .o ( E_51345 )  , .l ( E_48001 )  , .r ( E_47976 )  );
    CPL_MUX_2  I_47846 ( .o ( E_48001 )  , .s ( E_48191 )  , .d0 ( E_48000 )  , .d1 ( E_47999 )  );
    CPL_FF#20  I_48062_reg ( .q ( E_48000 )  , .qbar (  )  , .d ( E_47961 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48260 )  );
    CPL_MUX_2  I_47807 ( .o ( E_47961 )  , .s ( E_48196 )  , .d0 ( E_48001 )  , .d1 ( E_47960 )  );
    CPL_TYPE  I_51598 ( .o ( E_47960 )  , .l ( E_47959 )  );
    CPL_MUX_2  I_47805 ( .o ( E_47959 )  , .s ( E_47958 )  , .d0 ( E_47956_68643 )  , .d1 ( E_48092_68644 )  );
    CPL_GT  I_47804 ( .o ( E_47958 )  , .l ( E_47957 )  , .r ( E_48096 )  );
    CPL_TYPE  I_69209 ( .o ( E_47956_68643 )  , .l ( E_47956 )  );
    CPL_LASFT  I_47801 ( .o ( E_47956 )  , .d ( E_48093 )  , .s ( E_47957 )  );
      assign E_48260 = 20'hX; /*CDBImplicitXNone*/
    CPL_TYPE  I_51606 ( .o ( E_47999 )  , .l ( E_47998 )  );
    CPL_MUX_2  I_47844 ( .o ( E_47998 )  , .s ( E_47997 )  , .d0 ( E_47995_68645 )  , .d1 ( E_48092_68644 )  );
    CPL_GT  I_47843 ( .o ( E_47997 )  , .l ( E_47996 )  , .r ( E_48096 )  );
    CPL_SUB  I_47842 ( .o ( E_47996 )  , .l ( E_48141 )  , .r ( E_48115 )  );
    CPL_TYPE  I_69211 ( .o ( E_47995_68645 )  , .l ( E_47995 )  );
    CPL_LASFT  I_47840 ( .o ( E_47995 )  , .d ( E_48093 )  , .s ( E_47996 )  );
    CPL_MUX_2  I_51155 ( .o ( E_50829 )  , .s ( E_51038 )  , .d0 ( asm_sym_data_11 )  , 
		.d1 ( asm_sym_data_8 )  );
    CPL_EQ  I_51417 ( .o ( E_51038 )  , .l ( E_51357 )  , .r ( E_51339 )  );
    CPL_AND  I_47808 ( .o ( E_51339 )  , .l ( E_47961 )  , .r ( E_48197 )  );
    CPL_MUX_2  I_51250 ( .o ( E_50905 )  , .s ( E_51014 )  , .d0 ( asm_sym_data_9 )  , 
		.d1 ( asm_sym_data_8 )  );
    CPL_EQ  I_51387 ( .o ( E_51014 )  , .l ( E_51345 )  , .r ( E_51339 )  );
    CPL_MUX_2  I_51200 ( .o ( E_50865 )  , .s ( E_50994 )  , .d0 ( E_50869 )  , .d1 ( E_50905 )  );
    CPL_EQ  I_51362 ( .o ( E_50994 )  , .l ( E_51351 )  , .r ( E_51345 )  );
    CPL_MUX_2  I_51205 ( .o ( E_50869 )  , .s ( E_50998 )  , .d0 ( asm_sym_data_10 )  , 
		.d1 ( asm_sym_data_8 )  );
    CPL_EQ  I_51367 ( .o ( E_50998 )  , .l ( E_51351 )  , .r ( E_51339 )  );
    CPL_MULT  I_47932 ( .o ( E_48091 )  , .l ( E_48089 )  , .r ( E_48083 )  );
    CPL_RASFT  I_47930 ( .o ( E_48089 )  , .d ( E_48087 )  , .s ( E_48084 )  );
    CPL_MULT  I_47929 ( .o ( E_48087 )  , .l ( E_48108 )  , .r ( E_48086 )  );
    CPL_MUX_2  I_48174 ( .o ( E_48086 )  , .s ( E_48373 )  , .d0 ( E_48086_clone_48381 )  , 
		.d1 ( OOB_X_4 )  );
    CPL_MUX_2  I_51410 ( .o ( E_48086_clone_48381 )  , .s ( E_51002 )  , .d0 ( E_51037 )  , 
		.d1 ( E_48028_clone_48446 )  );
    CPL_MUX_2  I_51415 ( .o ( E_51037 )  , .s ( E_51018 )  , .d0 ( E_51041 )  , .d1 ( E_51053 )  );
    CPL_MUX_2  I_51420 ( .o ( E_51041 )  , .s ( E_51038 )  , .d0 ( asm_sym_data_3 )  , 
		.d1 ( E_47949_clone_48524 )  );
    CPL_MUX_2  I_51435 ( .o ( E_51053 )  , .s ( E_51014 )  , .d0 ( asm_sym_data_1 )  , 
		.d1 ( E_47949_clone_48524 )  );
    CPL_MUX_2  I_51425 ( .o ( E_48028_clone_48446 )  , .s ( E_50994 )  , .d0 ( E_51049 )  , 
		.d1 ( E_51053 )  );
    CPL_MUX_2  I_51430 ( .o ( E_51049 )  , .s ( E_50998 )  , .d0 ( asm_sym_data_2 )  , 
		.d1 ( E_47949_clone_48524 )  );
      assign E_48084 = 5'h14;
    CPL_MUX_2  I_47926 ( .o ( E_48083 )  , .s ( E_48181 )  , .d0 ( E_48082 )  , .d1 ( E_48081 )  );
    CPL_FF#32  I_48060_reg ( .q ( E_48082 )  , .qbar (  )  , .d ( E_48083 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48259 )  );
      assign E_48259 = 32'hX; /*CDBImplicitXNone*/
    CPL_TYPE  I_51621 ( .o ( E_48080 )  , .l ( E_48079 )  );
    CPL_SUB  I_47924 ( .o ( E_48079 )  , .l ( E_48112 )  , .r ( E_48083 )  );
    CPL_SUB  I_47914 ( .o ( E_48069 )  , .l ( E_48071 )  , .r ( E_48083 )  );
    CPL_MUX_2  I_47963 ( .o ( E_48124 )  , .s ( E_48123 )  , .d0 ( E_48122_68652 )  , .d1 ( E_48077 )  );
    CPL_LT  I_47962 ( .o ( E_48123 )  , .l ( E_48122 )  , .r ( E_48092 )  );
    CPL_SUB  I_47960 ( .o ( E_48122 )  , .l ( E_48120 )  , .r ( E_48114 )  );
    CPL_TYPE  I_69218 ( .o ( E_48122_68652 )  , .l ( E_48122 )  );
    CPL_ADD  I_47922 ( .o ( E_48077 )  , .l ( E_48122 )  , .r ( E_48083 )  );
    CPL_MUX_2  I_47896 ( .o ( E_48051 )  , .s ( E_48050 )  , .d0 ( E_48049 )  , .d1 ( E_48027 )  );
    CPL_GE  I_47895 ( .o ( E_48050 )  , .l ( E_48049 )  , .r ( E_48083 )  );
    CPL_TYPE  I_51617 ( .o ( E_48049 )  , .l ( E_48048 )  );
    CPL_SUB  I_47893 ( .o ( E_48048 )  , .l ( E_48047 )  , .r ( E_48033 )  );
    CPL_TYPE  I_51616 ( .o ( E_48047 )  , .l ( E_48046 )  );
    CPL_MULT  I_47891 ( .o ( E_48046 )  , .l ( E_48045 )  , .r ( E_48043 )  );
    CPL_MUX_2  I_48213 ( .o ( E_48045 )  , .s ( E_48412 )  , .d0 ( E_48045_clone_48420 )  , 
		.d1 ( OOB_X_7 )  );
    CPL_MUX_2  I_48950 ( .o ( E_48045_clone_48420 )  , .s ( E_48159 )  , .d0 ( asm_sym_data_20 )  , 
		.d1 ( E_49053 )  );
    CPL_MUX_2  I_48949 ( .o ( E_49053 )  , .s ( E_49037 )  , .d0 ( E_49051 )  , .d1 ( E_48124 )  );
    CPL_EQ  I_48931 ( .o ( E_49037 )  , .l ( E_48076 )  , .r ( E_51353 )  );
    CPL_MUX_2  I_48947 ( .o ( E_49051 )  , .s ( E_51057 )  , .d0 ( asm_sym_data_20 )  , 
		.d1 ( E_48073 )  );
    CPL_EQ  I_48928 ( .o ( E_51057 )  , .l ( E_48068 )  , .r ( E_51353 )  );
    CPL_MUX_2  I_48226 ( .o ( E_48043 )  , .s ( E_48438 )  , .d0 ( E_48043_clone_48433 )  , 
		.d1 ( OOB_X_8 )  );
    CPL_GT  I_48231 ( .o ( E_48438 )  , .l ( E_51351 )  , .r ( E_51065 )  );
    CPL_MUX_2  I_50965 ( .o ( E_48043_clone_48433 )  , .s ( E_50994 )  , .d0 ( E_50681 )  , 
		.d1 ( E_48004_clone_48472 )  );
    CPL_MUX_2  I_50970 ( .o ( E_50681 )  , .s ( E_50998 )  , .d0 ( E_50865 )  , .d1 ( E_47964_clone_48511 )  );
    CPL_MUX_2  I_51090 ( .o ( E_47964_clone_48511 )  , .s ( E_51038 )  , .d0 ( E_50781 )  , 
		.d1 ( E_48106_clone_48368 )  );
    CPL_MUX_2  I_51095 ( .o ( E_50781 )  , .s ( E_50998 )  , .d0 ( asm_sym_data_8 )  , 
		.d1 ( E_50865 )  );
    CPL_MUX_2  I_51030 ( .o ( E_48004_clone_48472 )  , .s ( E_51014 )  , .d0 ( E_50733 )  , 
		.d1 ( E_47964_clone_48511 )  );
    CPL_MUX_2  I_51035 ( .o ( E_50733 )  , .s ( E_51018 )  , .d0 ( E_50905 )  , .d1 ( E_48106_clone_48368 )  );
    CPL_TYPE  I_51613 ( .o ( E_48033 )  , .l ( E_48032 )  );
    CPL_MULT  I_47877 ( .o ( E_48032 )  , .l ( E_48031 )  , .r ( E_48083 )  );
    CPL_TYPE  I_51612 ( .o ( E_48031 )  , .l ( E_48030 )  );
    CPL_RASFT  I_47875 ( .o ( E_48030 )  , .d ( E_48029 )  , .s ( E_48084 )  );
    CPL_MULT  I_47874 ( .o ( E_48029 )  , .l ( E_48045 )  , .r ( E_48028 )  );
    CPL_MUX_2  I_48239 ( .o ( E_48028 )  , .s ( E_48438 )  , .d0 ( E_48028_clone_48446 )  , 
		.d1 ( OOB_X_9 )  );
    CPL_TYPE  I_51611 ( .o ( E_48027 )  , .l ( E_48026 )  );
    CPL_SUB  I_47871 ( .o ( E_48026 )  , .l ( E_48049 )  , .r ( E_48083 )  );
      assign E_47937 = 32'hffffffff;
    CPL_FF  I_48081_reg ( .q ( E_47860 )  , .qbar (  )  , .d ( E_48220 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48092 )  );
endmodule

