
--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_pkg_v1 IS

COMPONENT ccs_in_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    dat    : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_in_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    dat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_in_v1;

ARCHITECTURE beh OF ccs_in_v1 IS
BEGIN

  idat <= dat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/src/funcs.vhd 

-- a package of attributes that give verification tools a hint about
-- the function being implemented
PACKAGE attributes IS
  ATTRIBUTE CALYPTO_FUNC : string;
  ATTRIBUTE CALYPTO_DATA_ORDER : string;
end attributes;

-----------------------------------------------------------------------
-- Package that declares synthesizable functions needed for RTL output
-----------------------------------------------------------------------

LIBRARY ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

PACKAGE funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

   FUNCTION maximum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION minimum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2 : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;
   
-----------------------------------------------------------------
-- logic functions
-----------------------------------------------------------------

   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION or_v (inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- mux functions
-----------------------------------------------------------------

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC_VECTOR;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- latch functions
-----------------------------------------------------------------
   FUNCTION lat_s(dinput: STD_LOGIC       ; clk: STD_LOGIC; doutput: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- tristate functions
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC       ; control: STD_LOGIC) RETURN STD_LOGIC;
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: SIGNED  ) RETURN STD_LOGIC;

   -- RETURN 2 bits (left => lt, right => eq)
   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED;
 
   FUNCTION fabs(arg1: SIGNED  ) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "**" (l, r: UNSIGNED) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "**" (l, r: SIGNED  ) RETURN SIGNED  ;

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-- *_stdar functions use shift functions from std_logic_arith
-----------------------------------------------------------------

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;

   -----------------------------------------------------------------
   -- *_stdar functions use shift functions from std_logic_arith
   -----------------------------------------------------------------
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC;
   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE;
   --FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR ;

   FUNCTION ceil_log2(size : NATURAL) return NATURAL;
   FUNCTION bits(size : NATURAL) return NATURAL;    

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   
END funcs;


--------------------------- B O D Y ----------------------------


PACKAGE BODY funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC IS
     BEGIN IF arg1 THEN RETURN '1'; ELSE RETURN '0'; END IF; END;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
--     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;

   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
     VARIABLE result: STD_LOGIC_VECTOR(0 DOWNTO 0);
   BEGIN
     result := (0 => arg1);
     RETURN result;
   END;

   FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 > arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION minimum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 < arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;

   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := input1'LENGTH;
     ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
     ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     --synopsys translate_off
     FOR i IN len-1 DOWNTO 0 LOOP
       result(i) := resolved(input1a(i) & input2a(i));
     END LOOP;
     --synopsys translate_on
     RETURN result;
   END;

   FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED) RETURN UNSIGNED IS
   BEGIN RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

   FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED) RETURN SIGNED IS
   BEGIN RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

-----------------------------------------------------------------
-- Logic Functions
-----------------------------------------------------------------

   FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;
   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(and_v(inputs, 1)); END;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(or_v(inputs, 1)); END;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(xor_v(inputs, 1)); END;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result AND inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

   FUNCTION or_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     -- this if is added as a quick fix for a bug in catapult evaluating the loop even if inputs'LENGTH==1
     -- see dts0100971279
     IF icnt2 > 1 THEN
       FOR i IN icnt2-1 DOWNTO 1 LOOP
         inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
         result := result OR inputsx(olenM1 DOWNTO 0);
       END LOOP;
     END IF;
     RETURN result;
   END;

   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result XOR inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

-----------------------------------------------------------------
-- Muxes
-----------------------------------------------------------------
   
   FUNCTION mux_sel2_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(1 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 4;
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector( size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "01" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "10" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "11" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel3_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(2 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 8;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "001" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "010" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "011" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN "100" =>
       result := inputs0(5*size-1 DOWNTO 4*size);
     WHEN "101" =>
       result := inputs0(6*size-1 DOWNTO 5*size);
     WHEN "110" =>
       result := inputs0(7*size-1 DOWNTO 6*size);
     WHEN "111" =>
       result := inputs0(8*size-1 DOWNTO 7*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel4_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(3 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 16;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "0000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "0001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "0010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "0011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "0100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "0101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "0110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "0111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "1000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "1001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "1010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "1011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "1100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "1101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "1110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "1111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel5_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(4 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 32;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0 );
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "00001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "00010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "00011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "00100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "00101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "00110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "00111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "01000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "01001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "01010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "01011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "01100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "01101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "01110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "01111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "10000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "10001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "10010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "10011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "10100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "10101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "10110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "10111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "11000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "11001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "11010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "11011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "11100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "11101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "11110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "11111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel6_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(5 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 64;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "000001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "000010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "000011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "000100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "000101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "000110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "000111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "001000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "001001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "001010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "001011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "001100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "001101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "001110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "001111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "010000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "010001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "010010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "010011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "010100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "010101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "010110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "010111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "011000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "011001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "011010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "011011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "011100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "011101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "011110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "011111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN "100000" =>
       result := inputs0( 33*size-1 DOWNTO 32*size);
     WHEN "100001" =>
       result := inputs0( 34*size-1 DOWNTO 33*size);
     WHEN "100010" =>
       result := inputs0( 35*size-1 DOWNTO 34*size);
     WHEN "100011" =>
       result := inputs0( 36*size-1 DOWNTO 35*size);
     WHEN "100100" =>
       result := inputs0( 37*size-1 DOWNTO 36*size);
     WHEN "100101" =>
       result := inputs0( 38*size-1 DOWNTO 37*size);
     WHEN "100110" =>
       result := inputs0( 39*size-1 DOWNTO 38*size);
     WHEN "100111" =>
       result := inputs0( 40*size-1 DOWNTO 39*size);
     WHEN "101000" =>
       result := inputs0( 41*size-1 DOWNTO 40*size);
     WHEN "101001" =>
       result := inputs0( 42*size-1 DOWNTO 41*size);
     WHEN "101010" =>
       result := inputs0( 43*size-1 DOWNTO 42*size);
     WHEN "101011" =>
       result := inputs0( 44*size-1 DOWNTO 43*size);
     WHEN "101100" =>
       result := inputs0( 45*size-1 DOWNTO 44*size);
     WHEN "101101" =>
       result := inputs0( 46*size-1 DOWNTO 45*size);
     WHEN "101110" =>
       result := inputs0( 47*size-1 DOWNTO 46*size);
     WHEN "101111" =>
       result := inputs0( 48*size-1 DOWNTO 47*size);
     WHEN "110000" =>
       result := inputs0( 49*size-1 DOWNTO 48*size);
     WHEN "110001" =>
       result := inputs0( 50*size-1 DOWNTO 49*size);
     WHEN "110010" =>
       result := inputs0( 51*size-1 DOWNTO 50*size);
     WHEN "110011" =>
       result := inputs0( 52*size-1 DOWNTO 51*size);
     WHEN "110100" =>
       result := inputs0( 53*size-1 DOWNTO 52*size);
     WHEN "110101" =>
       result := inputs0( 54*size-1 DOWNTO 53*size);
     WHEN "110110" =>
       result := inputs0( 55*size-1 DOWNTO 54*size);
     WHEN "110111" =>
       result := inputs0( 56*size-1 DOWNTO 55*size);
     WHEN "111000" =>
       result := inputs0( 57*size-1 DOWNTO 56*size);
     WHEN "111001" =>
       result := inputs0( 58*size-1 DOWNTO 57*size);
     WHEN "111010" =>
       result := inputs0( 59*size-1 DOWNTO 58*size);
     WHEN "111011" =>
       result := inputs0( 60*size-1 DOWNTO 59*size);
     WHEN "111100" =>
       result := inputs0( 61*size-1 DOWNTO 60*size);
     WHEN "111101" =>
       result := inputs0( 62*size-1 DOWNTO 61*size);
     WHEN "111110" =>
       result := inputs0( 63*size-1 DOWNTO 62*size);
     WHEN "111111" =>
       result := inputs0( 64*size-1 DOWNTO 63*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS  --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2 SEVERITY FAILURE;
     --synopsys translate_on
       CASE sel IS
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0( size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1  DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0(size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
       RETURN result;
   END;
--   BEGIN RETURN mux_v(inputs, TO_STDLOGICVECTOR(sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     ALIAS    sel0   : STD_LOGIC_VECTOR( sel'LENGTH-1 DOWNTO 0 ) IS sel;

     VARIABLE sellen : INTEGER RANGE 2-sel'LENGTH TO sel'LENGTH;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2**sel'LENGTH;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
     TYPE inputs_array_type is array(natural range <>) of std_logic_vector( olen - 1 DOWNTO 0);
     VARIABLE inputs_array : inputs_array_type( 2**sel'LENGTH - 1 DOWNTO 0);
   BEGIN
     sellen := sel'LENGTH;
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2**sellen SEVERITY FAILURE;
     sellen := 2-sellen;
     --synopsys translate_on
     CASE sellen IS
     WHEN 1 =>
       CASE sel0(0) IS

       WHEN '1' 
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0(  size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1 DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0( size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
     WHEN 2 =>
       result := mux_sel2_v(inputs, not sel);
     WHEN 3 =>
       result := mux_sel3_v(inputs, not sel);
     WHEN 4 =>
       result := mux_sel4_v(inputs, not sel);
     WHEN 5 =>
       result := mux_sel5_v(inputs, not sel);
     WHEN 6 =>
       result := mux_sel6_v(inputs, not sel);
     WHEN others =>
       -- synopsys translate_off
       IF(Is_X(sel0)) THEN
         result := (others => 'X');
       ELSE
       -- synopsys translate_on
         FOR i in 0 to 2**sel'LENGTH - 1 LOOP
           inputs_array(i) := inputs0( ((i + 1) * olen) - 1  DOWNTO i*olen);
         END LOOP;
         result := inputs_array(CONV_INTEGER( (UNSIGNED(NOT sel0)) ));
       -- synopsys translate_off
       END IF;
       -- synopsys translate_on
     END CASE;
     RETURN result;
   END;

 
-----------------------------------------------------------------
-- Latches
-----------------------------------------------------------------

   FUNCTION lat_s(dinput: STD_LOGIC; clk: STD_LOGIC; doutput: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN mux_s(STD_LOGIC_VECTOR'(doutput & dinput), clk); END;

   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR ; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR ) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     --synopsys translate_off
     ASSERT dinput'LENGTH = doutput'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN mux_v(doutput & dinput, clk);
   END;

-----------------------------------------------------------------
-- Tri-States
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC; control: STD_LOGIC) RETURN STD_LOGIC IS
--   BEGIN RETURN TO_STDLOGIC(tri_v(TO_STDLOGICVECTOR(dinput), control)); END;
--
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR ; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
--     VARIABLE result: STD_LOGIC_VECTOR(dinput'range);
--   BEGIN
--     CASE control IS
--     WHEN '0' | 'L' =>
--       result := (others => 'Z');
--     WHEN '1' | 'H' =>
--       FOR i IN dinput'range LOOP
--         result(i) := to_UX01(dinput(i));
--       END LOOP;
--     WHEN others =>
--       -- synopsys translate_off
--       result := (others => 'X');
--       -- synopsys translate_on
--     END CASE;
--     RETURN result;
--   END;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;

   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     VARIABLE diff: UNSIGNED(l'LENGTH DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     diff := ('0'&l) - ('0'&r);
     RETURN diff(l'LENGTH);
   END;
   FUNCTION "<"(l, r: SIGNED  ) RETURN STD_LOGIC IS
   BEGIN
     RETURN (UNSIGNED(l) < UNSIGNED(r)) xor (l(l'LEFT) xor r(r'LEFT));
   END;

   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION "<=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">"(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;
   FUNCTION ">=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;

   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN not or_s(l xor r);
   END;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   --some functions to placate spyglass
   FUNCTION mult_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a*b;
   END mult_natural;

   FUNCTION div_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a/b;
   END div_natural;

   FUNCTION mod_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a mod b;
   END mod_natural;

   FUNCTION add_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a+b;
   END add_unsigned;

   FUNCTION sub_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a-b;
   END sub_unsigned;

   FUNCTION sub_int(a,b : INTEGER) RETURN INTEGER IS
   BEGIN
     return a-b;
   END sub_int;

   FUNCTION concat_0(b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return '0' & b;
   END concat_0;

   FUNCTION concat_uns(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a&b;
   END concat_uns;

   FUNCTION concat_vect(a,b : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     return a&b;
   END concat_vect;





   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED IS
     CONSTANT ninps : NATURAL := arg'LENGTH / width;
     ALIAS    arg0  : UNSIGNED(arg'LENGTH-1 DOWNTO 0) IS arg;
     VARIABLE result: UNSIGNED(width-1 DOWNTO 0);
     VARIABLE from  : INTEGER;
     VARIABLE dto   : INTEGER;
   BEGIN
     --synopsys translate_off
     ASSERT arg'LENGTH = width * ninps SEVERITY FAILURE;
     --synopsys translate_on
     result := (OTHERS => '0');
     FOR i IN ninps-1 DOWNTO 0 LOOP
       --result := result + arg0((i+1)*width-1 DOWNTO i*width);
       from := mult_natural((i+1), width)-1; --2.1.6.3
       dto  := mult_natural(i,width); --2.1.6.3
       result := add_unsigned(result , arg0(from DOWNTO dto) );
     END LOOP;
     RETURN result;
   END faccu;

   FUNCTION  fabs (arg1: SIGNED) RETURN UNSIGNED IS
   BEGIN
     CASE arg1(arg1'LEFT) IS
     WHEN '1'
     --synopsys translate_off
          | 'H'
     --synopsys translate_on
       =>
       RETURN UNSIGNED'("0") - UNSIGNED(arg1);
     WHEN '0'
     --synopsys translate_off
          | 'L'
     --synopsys translate_on
       =>
       RETURN UNSIGNED(arg1);
     WHEN others =>
       RETURN resolve_unsigned(UNSIGNED(arg1), UNSIGNED'("0") - UNSIGNED(arg1));
     END CASE;
   END;

   PROCEDURE divmod(l, r: UNSIGNED; rdiv, rmod: OUT UNSIGNED) IS
     CONSTANT llen: INTEGER := l'LENGTH;
     CONSTANT rlen: INTEGER := r'LENGTH;
     CONSTANT llen_plus_rlen: INTEGER := llen + rlen;
     VARIABLE lbuf: UNSIGNED(llen+rlen-1 DOWNTO 0);
     VARIABLE diff: UNSIGNED(rlen DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT rdiv'LENGTH = llen AND rmod'LENGTH = rlen SEVERITY FAILURE;
     --synopsys translate_on
     lbuf := (others => '0');
     lbuf(llen-1 DOWNTO 0) := l;
     FOR i IN rdiv'range LOOP
       diff := sub_unsigned(lbuf(llen_plus_rlen-1 DOWNTO llen-1) ,(concat_0(r)));
       rdiv(i) := not diff(rlen);
       IF diff(rlen) = '0' THEN
         lbuf(llen_plus_rlen-1 DOWNTO llen-1) := diff;
       END IF;
       lbuf(llen_plus_rlen-1 DOWNTO 1) := lbuf(llen_plus_rlen-2 DOWNTO 0);
     END LOOP;
     rmod := lbuf(llen_plus_rlen-1 DOWNTO llen);
   END divmod;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rdiv;
   END "/";

   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rmod;
   END;

   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN l MOD r; END;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rdiv := UNSIGNED'("0") - rdiv;
     END IF;
     RETURN SIGNED(rdiv); -- overflow problem "1000" / "11"
   END "/";

   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
     CONSTANT rnul: UNSIGNED(r'LENGTH-1 DOWNTO 0) := (others => '0');
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     IF rmod /= rnul AND to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rmod := UNSIGNED(r) + rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "MOD";

   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "REM";

   FUNCTION mult_unsigned(l,r : UNSIGNED) return UNSIGNED is
   BEGIN
     return l*r; 
   END mult_unsigned;

   FUNCTION "**" (l, r : UNSIGNED) RETURN UNSIGNED IS
     CONSTANT llen  : NATURAL := l'LENGTH;
     VARIABLE result: UNSIGNED(llen-1 DOWNTO 0);
     VARIABLE fak   : UNSIGNED(llen-1 DOWNTO 0);
   BEGIN
     fak := l;
     result := (others => '0'); result(0) := '1';
     FOR i IN r'reverse_range LOOP
       --was:result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(result & (result*fak)), r(i)));
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR( concat_uns(result , mult_unsigned(result,fak) )), r(i)));

       fak := mult_unsigned(fak , fak);
     END LOOP;
     RETURN result;
   END "**";

   FUNCTION "**" (l, r : SIGNED) RETURN SIGNED IS
     CONSTANT rlen  : NATURAL := r'LENGTH;
     ALIAS    r0    : SIGNED(0 TO r'LENGTH-1) IS r;
     VARIABLE result: SIGNED(l'range);
   BEGIN
     CASE r(r'LEFT) IS
     WHEN '0'
   --synopsys translate_off
          | 'L'
   --synopsys translate_on
     =>
       result := SIGNED(UNSIGNED(l) ** UNSIGNED(r0(1 TO r'LENGTH-1)));
     WHEN '1'
   --synopsys translate_off
          | 'H'
   --synopsys translate_on
     =>
       result := (others => '0');
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END "**";

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-----------------------------------------------------------------

   FUNCTION add_nat(arg1 : NATURAL; arg2 : NATURAL ) RETURN NATURAL IS
   BEGIN
     return (arg1 + arg2);
   END;
   
--   FUNCTION UNSIGNED_2_BIT_VECTOR(arg1 : NATURAL; arg2 : NATURAL ) RETURN BIT_VECTOR IS
--   BEGIN
--     return (arg1 + arg2);
--   END;
   
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(SIGNED(result), arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
        =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
        =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;


   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     --SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: NATURAL range 1 TO len;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => '0');
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         --was:temp(i2+sw) := result(i2);
         temp_idx := add_nat(i2,sw);
         temp(temp_idx) := result(i2);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: sw_range;
     VARIABLE result_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => sbit);
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         -- was: temp(i2) := result(i2+sw);
         result_idx := add_nat(i2,sw);
         temp(i2) := result(result_idx);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;


   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := arg1'LENGTH;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     VARIABLE temp: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     SUBTYPE sw_range IS NATURAL range 0 TO len-1;
     VARIABLE sw: sw_range;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     result := (others=>'0');
     result := arg1;
     sw := sdir MOD len;
     FOR i IN arg2'reverse_range LOOP
       EXIT WHEN sw = 0;
       IF signd2 AND i = arg2'LEFT THEN 
         sw := sub_int(len,sw); 
       END IF;
       -- temp := result(len-sw-1 DOWNTO 0) & result(len-1 DOWNTO len-sw)
       FOR i2 IN len-1 DOWNTO 0 LOOP
         --was: temp((i2+sw) MOD len) := result(i2);
         temp_idx := add_nat(i2,sw) MOD len;
         temp(temp_idx) := result(i2);
       END LOOP;
       result := mux_v(STD_LOGIC_VECTOR(concat_vect(result,temp)), arg2(i));
       sw := mod_natural(mult_natural(sw,2), len);
     END LOOP;
     RETURN result;
   END frot;

   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, -1); END;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, -1); END;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC IS
     CONSTANT len : INTEGER := vec'LENGTH;
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
   BEGIN
     IF index >= len OR index < 0 THEN
       RETURN 'X';
     END IF;
     RETURN vec0(index);
   END;

   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     CONSTANT indexPwidthM1 : INTEGER := index+width-1; --2.1.6.3
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
     CONSTANT xxx : STD_LOGIC_VECTOR(width-1 DOWNTO 0) := (others => 'X');
   BEGIN
     IF index+width > len OR index < 0 THEN
       RETURN xxx;
     END IF;
     RETURN vec0(indexPwidthM1 DOWNTO index);
   END;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     VARIABLE vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     CONSTANT xxx : STD_LOGIC_VECTOR(len-1 DOWNTO 0) := (others => 'X');
   BEGIN
     vec0 := vec;
     IF index >= len OR index < 0 THEN
       RETURN xxx;
     END IF;
     vec0(index) := dinput;
     RETURN vec0;
   END;

   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE IS
     VARIABLE n_b : POSITIVE;
     VARIABLE p_v : NATURAL;
   BEGIN
     p_v := p;
     FOR i IN 1 TO 32 LOOP
       p_v := div_natural(p_v,2);
       n_b := i;
       EXIT WHEN (p_v = 0);
     END LOOP;
     RETURN n_b;
   END;


--   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
--
--     CONSTANT vlen: INTEGER := vec'LENGTH;
--     CONSTANT ilen: INTEGER := dinput'LENGTH;
--     CONSTANT max_shift: INTEGER := vlen-ilen;
--     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
--     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
--     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
--     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
--     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
--     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
--   BEGIN
--     inp := (others => '0');
--     mask := (others => '0');
--
--     IF index > max_shift OR index < 0 THEN
--       RETURN xxx;
--     END IF;
--
--     shift := CONV_UNSIGNED(index, shift'LENGTH);
--     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
--     mask(ilen-1 DOWNTO 0) := ones;
--     inp := fshl(inp, shift, vlen);
--     mask := fshl(mask, shift, vlen);
--     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
--     RETURN vec0;
--   END;

   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR IS

     type enable_matrix is array (0 to enable'LENGTH-1 ) of std_logic_vector(byte_width-1 downto 0);
     CONSTANT vlen: INTEGER := vec'LENGTH;
     CONSTANT ilen: INTEGER := dinput'LENGTH;
     CONSTANT max_shift: INTEGER := vlen-ilen;
     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask2: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE enables: enable_matrix;
     VARIABLE cat_enables: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0 );
     VARIABLE lsbi : INTEGER;
     VARIABLE msbi : INTEGER;

   BEGIN
     cat_enables := (others => '0');
     lsbi := 0;
     msbi := byte_width-1;
     inp := (others => '0');
     mask := (others => '0');

     IF index > max_shift OR index < 0 THEN
       RETURN xxx;
     END IF;

     --initialize enables
     for i in 0 TO (enable'LENGTH-1) loop
       enables(i)  := (others => enable(i));
       cat_enables(msbi downto lsbi) := enables(i) ;
       lsbi := msbi+1;
       msbi := msbi+byte_width;
     end loop;


     shift := CONV_UNSIGNED(index, shift'LENGTH);
     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
     mask(ilen-1 DOWNTO 0) := UNSIGNED((STD_LOGIC_VECTOR(ones) AND cat_enables));
     inp := fshl(inp, shift, vlen);
     mask := fshl(mask, shift, vlen);
     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
     RETURN vec0;
   END;


   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;
   
   FUNCTION bits(size : NATURAL) return NATURAL is
   begin
     return ceil_log2(size);
   END;

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH) xor conv_std_logic_vector(c, s'LENGTH);
     cout := ( (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH)) or (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) or (conv_std_logic_vector(b, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) );
   END PROCEDURE csa;

   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH);
     cout := (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH));
   END PROCEDURE csha;

END funcs;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_comps.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_comps IS
 
FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
FUNCTION ceil_log2(size : NATURAL) return NATURAL;
 

COMPONENT mgc_not
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_and
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nand
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_or
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xnor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux
  GENERIC (
    width  :  NATURAL;
    ctrlw  :  NATURAL;
    p2ctrlw : NATURAL := 0
  );
  PORT (
    a: in  std_logic_vector(width*(2**ctrlw) - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw            - 1 DOWNTO 0);
    z: out std_logic_vector(width            - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux1hot
  GENERIC (
    width  : NATURAL;
    ctrlw  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ctrlw - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw       - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_reg_pos
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;  -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL  -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_reg_neg
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;   -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_generic_reg
  GENERIC(
   width: natural := 8;
   ph_clk: integer range 0 to 1 := 1; -- clock polarity, 1=rising_edge
   ph_en: integer range 0 to 1 := 1;
   ph_a_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   ph_s_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   a_rst_used: integer range 0 to 1 := 1;
   s_rst_used: integer range 0 to 1 := 0;
   en_used: integer range 0 to 1 := 1
  );
  PORT(
   d: std_logic_vector(width-1 downto 0);
   clk: in std_logic;
   en: in std_logic;
   a_rst: in std_logic;
   s_rst: in std_logic;
   q: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_equal
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a : in  std_logic_vector(width-1 DOWNTO 0);
    b : in  std_logic_vector(width-1 DOWNTO 0);
    eq: out std_logic;
    ne: out std_logic
  );
END COMPONENT;

COMPONENT mgc_shift_l
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rot
  GENERIC (
    width  : NATURAL;
    width_s: NATURAL;
    signd_s: NATURAL;      -- 0:unsigned 1:signed
    sleft  : NATURAL;      -- 0:right 1:left;
    log2w  : NATURAL := 0; -- LOG2(width)
    l2wp2  : NATURAL := 0  --2**LOG2(width)
  );
  PORT (
    a : in  std_logic_vector(width  -1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width  -1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_sub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_ci
  GENERIC (
    width_a : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width_a, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width_a, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width_a,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width_a,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_addc
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add3
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_c : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_c : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(ifeqsel(width_c,0,width,width_c)-1 DOWNTO 0);
    d: in  std_logic_vector(0 DOWNTO 0);
    e: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_sub_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addc_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     c: in std_logic_vector(0 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addsub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    add: in  std_logic;
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_accu
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_abs
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_fast
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_pipe
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2  : NATURAL;
    add_d2  : NATURAL
  );
  PORT (
    a   : in  std_logic_vector(width_a-1 DOWNTO 0);
    b   : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2  : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c   : in  std_logic_vector(width_c-1 DOWNTO 0);
    d   : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2  : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst : in  std_logic_vector(width_e-1 DOWNTO 0);
    z   : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1_pipe
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2   : NATURAL;
    add_d2   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2     : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2     : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_e-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL
  );
  PORT (
    a:   in  std_logic_vector(width_a-1 DOWNTO 0);
    b:   in  std_logic_vector(width_b-1 DOWNTO 0);
    c:   in  std_logic_vector(width_c-1 DOWNTO 0);
    cst: in  std_logic_vector(width_cst-1 DOWNTO 0);
    d:   in  std_logic_vector(width_d-1 DOWNTO 0);
    z:   out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1_pipe
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_cst-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mulacc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2acc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    add_cxd : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    d         : in  std_logic_vector(width_d-1 DOWNTO 0);
    e         : in  std_logic_vector(width_e-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_div
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mod
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rem
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_csa
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     c: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_csha
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_rom
    GENERIC (
      rom_id : natural := 1;
      size : natural := 33;
      width : natural := 32
      );
    PORT (
      data_in : std_logic_vector((size*width)-1 downto 0);
      addr : std_logic_vector(ceil_log2(size)-1 downto 0);
      data_out : out std_logic_vector(width-1 downto 0)
    );
END COMPONENT;

END mgc_comps;

PACKAGE BODY mgc_comps IS
 
   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;
 
END mgc_comps;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_rem IS
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END mgc_rem;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

USE work.funcs.all;

ARCHITECTURE beh OF mgc_rem IS
BEGIN
  z <= std_logic_vector(unsigned(a) rem unsigned(b)) WHEN signd = 0 ELSE
       std_logic_vector(  signed(a) rem   signed(b));
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_div IS
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END mgc_div;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

USE work.funcs.all;

ARCHITECTURE beh OF mgc_div IS
BEGIN
  z <= std_logic_vector(unsigned(a) / unsigned(b)) WHEN signd = 0 ELSE
       std_logic_vector(  signed(a) /   signed(b));
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_comps_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_shift_comps_v5 IS

COMPONENT mgc_shift_l_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_shift_comps_v5;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_shift_l_v5 IS
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_shift_l_v5;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_shift_l_v5 IS

  FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1 > arg2) THEN
      RETURN(arg1) ;
    ELSE
      RETURN(arg2) ;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(SIGNED(result), arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE)
  RETURN UNSIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, '0', olen);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE)
  RETURN SIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen);
  END;

BEGIN
UNSGNED:  IF signd_a = 0 GENERATE
    z <= std_logic_vector(fshl_stdar(unsigned(a), unsigned(s), width_z));
  END GENERATE;
SGNED:  IF signd_a /= 0 GENERATE
    z <= std_logic_vector(fshl_stdar(  signed(a), unsigned(s), width_z));
  END GENERATE;
END beh;

--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Wed Jun 30 21:42:10 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_9_64_512_512_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_9_64_512_512_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_9_64_512_512_64_1_gen;

ARCHITECTURE v40 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_9_64_512_512_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v40;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_9_64_512_512_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_9_64_512_512_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_9_64_512_512_64_1_gen;

ARCHITECTURE v40 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_9_64_512_512_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v40;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_9_64_512_512_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_9_64_512_512_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_9_64_512_512_64_1_gen;

ARCHITECTURE v40 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_9_64_512_512_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v40;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_9_64_512_512_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_9_64_512_512_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_9_64_512_512_64_1_gen;

ARCHITECTURE v40 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_9_64_512_512_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v40;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_9_64_512_512_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_9_64_512_512_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_9_64_512_512_64_1_gen;

ARCHITECTURE v40 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_9_64_512_512_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v40;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_9_64_512_512_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_9_64_512_512_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_9_64_512_512_64_1_gen;

ARCHITECTURE v40 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_9_64_512_512_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v40;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_9_64_512_512_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_9_64_512_512_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_9_64_512_512_64_1_gen;

ARCHITECTURE v40 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_9_64_512_512_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v40;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_9_64_512_512_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_9_64_512_512_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_9_64_512_512_64_1_gen;

ARCHITECTURE v40 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_9_64_512_512_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v40;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    STAGE_LOOP_C_8_tr0 : IN STD_LOGIC;
    modExp_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_1_tr0 : IN STD_LOGIC;
    COMP_LOOP_1_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_62_tr0 : IN STD_LOGIC;
    COMP_LOOP_2_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_124_tr0 : IN STD_LOGIC;
    COMP_LOOP_3_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_186_tr0 : IN STD_LOGIC;
    COMP_LOOP_4_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_248_tr0 : IN STD_LOGIC;
    COMP_LOOP_5_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_310_tr0 : IN STD_LOGIC;
    COMP_LOOP_6_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_372_tr0 : IN STD_LOGIC;
    COMP_LOOP_7_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_434_tr0 : IN STD_LOGIC;
    COMP_LOOP_8_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_496_tr0 : IN STD_LOGIC;
    VEC_LOOP_C_0_tr0 : IN STD_LOGIC;
    STAGE_LOOP_C_9_tr0 : IN STD_LOGIC
  );
END inPlaceNTT_DIT_core_core_fsm;

ARCHITECTURE v40 OF inPlaceNTT_DIT_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for inPlaceNTT_DIT_core_core_fsm_1
  TYPE inPlaceNTT_DIT_core_core_fsm_1_ST IS (main_C_0, STAGE_LOOP_C_0, STAGE_LOOP_C_1,
      STAGE_LOOP_C_2, STAGE_LOOP_C_3, STAGE_LOOP_C_4, STAGE_LOOP_C_5, STAGE_LOOP_C_6,
      STAGE_LOOP_C_7, STAGE_LOOP_C_8, modExp_while_C_0, modExp_while_C_1, modExp_while_C_2,
      modExp_while_C_3, modExp_while_C_4, modExp_while_C_5, modExp_while_C_6, modExp_while_C_7,
      modExp_while_C_8, modExp_while_C_9, modExp_while_C_10, modExp_while_C_11, modExp_while_C_12,
      modExp_while_C_13, modExp_while_C_14, modExp_while_C_15, modExp_while_C_16,
      modExp_while_C_17, modExp_while_C_18, modExp_while_C_19, modExp_while_C_20,
      modExp_while_C_21, modExp_while_C_22, modExp_while_C_23, modExp_while_C_24,
      modExp_while_C_25, modExp_while_C_26, modExp_while_C_27, modExp_while_C_28,
      modExp_while_C_29, modExp_while_C_30, modExp_while_C_31, modExp_while_C_32,
      modExp_while_C_33, modExp_while_C_34, modExp_while_C_35, modExp_while_C_36,
      modExp_while_C_37, modExp_while_C_38, COMP_LOOP_C_0, COMP_LOOP_C_1, COMP_LOOP_1_modExp_1_while_C_0,
      COMP_LOOP_1_modExp_1_while_C_1, COMP_LOOP_1_modExp_1_while_C_2, COMP_LOOP_1_modExp_1_while_C_3,
      COMP_LOOP_1_modExp_1_while_C_4, COMP_LOOP_1_modExp_1_while_C_5, COMP_LOOP_1_modExp_1_while_C_6,
      COMP_LOOP_1_modExp_1_while_C_7, COMP_LOOP_1_modExp_1_while_C_8, COMP_LOOP_1_modExp_1_while_C_9,
      COMP_LOOP_1_modExp_1_while_C_10, COMP_LOOP_1_modExp_1_while_C_11, COMP_LOOP_1_modExp_1_while_C_12,
      COMP_LOOP_1_modExp_1_while_C_13, COMP_LOOP_1_modExp_1_while_C_14, COMP_LOOP_1_modExp_1_while_C_15,
      COMP_LOOP_1_modExp_1_while_C_16, COMP_LOOP_1_modExp_1_while_C_17, COMP_LOOP_1_modExp_1_while_C_18,
      COMP_LOOP_1_modExp_1_while_C_19, COMP_LOOP_1_modExp_1_while_C_20, COMP_LOOP_1_modExp_1_while_C_21,
      COMP_LOOP_1_modExp_1_while_C_22, COMP_LOOP_1_modExp_1_while_C_23, COMP_LOOP_1_modExp_1_while_C_24,
      COMP_LOOP_1_modExp_1_while_C_25, COMP_LOOP_1_modExp_1_while_C_26, COMP_LOOP_1_modExp_1_while_C_27,
      COMP_LOOP_1_modExp_1_while_C_28, COMP_LOOP_1_modExp_1_while_C_29, COMP_LOOP_1_modExp_1_while_C_30,
      COMP_LOOP_1_modExp_1_while_C_31, COMP_LOOP_1_modExp_1_while_C_32, COMP_LOOP_1_modExp_1_while_C_33,
      COMP_LOOP_1_modExp_1_while_C_34, COMP_LOOP_1_modExp_1_while_C_35, COMP_LOOP_1_modExp_1_while_C_36,
      COMP_LOOP_1_modExp_1_while_C_37, COMP_LOOP_1_modExp_1_while_C_38, COMP_LOOP_C_2,
      COMP_LOOP_C_3, COMP_LOOP_C_4, COMP_LOOP_C_5, COMP_LOOP_C_6, COMP_LOOP_C_7,
      COMP_LOOP_C_8, COMP_LOOP_C_9, COMP_LOOP_C_10, COMP_LOOP_C_11, COMP_LOOP_C_12,
      COMP_LOOP_C_13, COMP_LOOP_C_14, COMP_LOOP_C_15, COMP_LOOP_C_16, COMP_LOOP_C_17,
      COMP_LOOP_C_18, COMP_LOOP_C_19, COMP_LOOP_C_20, COMP_LOOP_C_21, COMP_LOOP_C_22,
      COMP_LOOP_C_23, COMP_LOOP_C_24, COMP_LOOP_C_25, COMP_LOOP_C_26, COMP_LOOP_C_27,
      COMP_LOOP_C_28, COMP_LOOP_C_29, COMP_LOOP_C_30, COMP_LOOP_C_31, COMP_LOOP_C_32,
      COMP_LOOP_C_33, COMP_LOOP_C_34, COMP_LOOP_C_35, COMP_LOOP_C_36, COMP_LOOP_C_37,
      COMP_LOOP_C_38, COMP_LOOP_C_39, COMP_LOOP_C_40, COMP_LOOP_C_41, COMP_LOOP_C_42,
      COMP_LOOP_C_43, COMP_LOOP_C_44, COMP_LOOP_C_45, COMP_LOOP_C_46, COMP_LOOP_C_47,
      COMP_LOOP_C_48, COMP_LOOP_C_49, COMP_LOOP_C_50, COMP_LOOP_C_51, COMP_LOOP_C_52,
      COMP_LOOP_C_53, COMP_LOOP_C_54, COMP_LOOP_C_55, COMP_LOOP_C_56, COMP_LOOP_C_57,
      COMP_LOOP_C_58, COMP_LOOP_C_59, COMP_LOOP_C_60, COMP_LOOP_C_61, COMP_LOOP_C_62,
      COMP_LOOP_C_63, COMP_LOOP_2_modExp_1_while_C_0, COMP_LOOP_2_modExp_1_while_C_1,
      COMP_LOOP_2_modExp_1_while_C_2, COMP_LOOP_2_modExp_1_while_C_3, COMP_LOOP_2_modExp_1_while_C_4,
      COMP_LOOP_2_modExp_1_while_C_5, COMP_LOOP_2_modExp_1_while_C_6, COMP_LOOP_2_modExp_1_while_C_7,
      COMP_LOOP_2_modExp_1_while_C_8, COMP_LOOP_2_modExp_1_while_C_9, COMP_LOOP_2_modExp_1_while_C_10,
      COMP_LOOP_2_modExp_1_while_C_11, COMP_LOOP_2_modExp_1_while_C_12, COMP_LOOP_2_modExp_1_while_C_13,
      COMP_LOOP_2_modExp_1_while_C_14, COMP_LOOP_2_modExp_1_while_C_15, COMP_LOOP_2_modExp_1_while_C_16,
      COMP_LOOP_2_modExp_1_while_C_17, COMP_LOOP_2_modExp_1_while_C_18, COMP_LOOP_2_modExp_1_while_C_19,
      COMP_LOOP_2_modExp_1_while_C_20, COMP_LOOP_2_modExp_1_while_C_21, COMP_LOOP_2_modExp_1_while_C_22,
      COMP_LOOP_2_modExp_1_while_C_23, COMP_LOOP_2_modExp_1_while_C_24, COMP_LOOP_2_modExp_1_while_C_25,
      COMP_LOOP_2_modExp_1_while_C_26, COMP_LOOP_2_modExp_1_while_C_27, COMP_LOOP_2_modExp_1_while_C_28,
      COMP_LOOP_2_modExp_1_while_C_29, COMP_LOOP_2_modExp_1_while_C_30, COMP_LOOP_2_modExp_1_while_C_31,
      COMP_LOOP_2_modExp_1_while_C_32, COMP_LOOP_2_modExp_1_while_C_33, COMP_LOOP_2_modExp_1_while_C_34,
      COMP_LOOP_2_modExp_1_while_C_35, COMP_LOOP_2_modExp_1_while_C_36, COMP_LOOP_2_modExp_1_while_C_37,
      COMP_LOOP_2_modExp_1_while_C_38, COMP_LOOP_C_64, COMP_LOOP_C_65, COMP_LOOP_C_66,
      COMP_LOOP_C_67, COMP_LOOP_C_68, COMP_LOOP_C_69, COMP_LOOP_C_70, COMP_LOOP_C_71,
      COMP_LOOP_C_72, COMP_LOOP_C_73, COMP_LOOP_C_74, COMP_LOOP_C_75, COMP_LOOP_C_76,
      COMP_LOOP_C_77, COMP_LOOP_C_78, COMP_LOOP_C_79, COMP_LOOP_C_80, COMP_LOOP_C_81,
      COMP_LOOP_C_82, COMP_LOOP_C_83, COMP_LOOP_C_84, COMP_LOOP_C_85, COMP_LOOP_C_86,
      COMP_LOOP_C_87, COMP_LOOP_C_88, COMP_LOOP_C_89, COMP_LOOP_C_90, COMP_LOOP_C_91,
      COMP_LOOP_C_92, COMP_LOOP_C_93, COMP_LOOP_C_94, COMP_LOOP_C_95, COMP_LOOP_C_96,
      COMP_LOOP_C_97, COMP_LOOP_C_98, COMP_LOOP_C_99, COMP_LOOP_C_100, COMP_LOOP_C_101,
      COMP_LOOP_C_102, COMP_LOOP_C_103, COMP_LOOP_C_104, COMP_LOOP_C_105, COMP_LOOP_C_106,
      COMP_LOOP_C_107, COMP_LOOP_C_108, COMP_LOOP_C_109, COMP_LOOP_C_110, COMP_LOOP_C_111,
      COMP_LOOP_C_112, COMP_LOOP_C_113, COMP_LOOP_C_114, COMP_LOOP_C_115, COMP_LOOP_C_116,
      COMP_LOOP_C_117, COMP_LOOP_C_118, COMP_LOOP_C_119, COMP_LOOP_C_120, COMP_LOOP_C_121,
      COMP_LOOP_C_122, COMP_LOOP_C_123, COMP_LOOP_C_124, COMP_LOOP_C_125, COMP_LOOP_3_modExp_1_while_C_0,
      COMP_LOOP_3_modExp_1_while_C_1, COMP_LOOP_3_modExp_1_while_C_2, COMP_LOOP_3_modExp_1_while_C_3,
      COMP_LOOP_3_modExp_1_while_C_4, COMP_LOOP_3_modExp_1_while_C_5, COMP_LOOP_3_modExp_1_while_C_6,
      COMP_LOOP_3_modExp_1_while_C_7, COMP_LOOP_3_modExp_1_while_C_8, COMP_LOOP_3_modExp_1_while_C_9,
      COMP_LOOP_3_modExp_1_while_C_10, COMP_LOOP_3_modExp_1_while_C_11, COMP_LOOP_3_modExp_1_while_C_12,
      COMP_LOOP_3_modExp_1_while_C_13, COMP_LOOP_3_modExp_1_while_C_14, COMP_LOOP_3_modExp_1_while_C_15,
      COMP_LOOP_3_modExp_1_while_C_16, COMP_LOOP_3_modExp_1_while_C_17, COMP_LOOP_3_modExp_1_while_C_18,
      COMP_LOOP_3_modExp_1_while_C_19, COMP_LOOP_3_modExp_1_while_C_20, COMP_LOOP_3_modExp_1_while_C_21,
      COMP_LOOP_3_modExp_1_while_C_22, COMP_LOOP_3_modExp_1_while_C_23, COMP_LOOP_3_modExp_1_while_C_24,
      COMP_LOOP_3_modExp_1_while_C_25, COMP_LOOP_3_modExp_1_while_C_26, COMP_LOOP_3_modExp_1_while_C_27,
      COMP_LOOP_3_modExp_1_while_C_28, COMP_LOOP_3_modExp_1_while_C_29, COMP_LOOP_3_modExp_1_while_C_30,
      COMP_LOOP_3_modExp_1_while_C_31, COMP_LOOP_3_modExp_1_while_C_32, COMP_LOOP_3_modExp_1_while_C_33,
      COMP_LOOP_3_modExp_1_while_C_34, COMP_LOOP_3_modExp_1_while_C_35, COMP_LOOP_3_modExp_1_while_C_36,
      COMP_LOOP_3_modExp_1_while_C_37, COMP_LOOP_3_modExp_1_while_C_38, COMP_LOOP_C_126,
      COMP_LOOP_C_127, COMP_LOOP_C_128, COMP_LOOP_C_129, COMP_LOOP_C_130, COMP_LOOP_C_131,
      COMP_LOOP_C_132, COMP_LOOP_C_133, COMP_LOOP_C_134, COMP_LOOP_C_135, COMP_LOOP_C_136,
      COMP_LOOP_C_137, COMP_LOOP_C_138, COMP_LOOP_C_139, COMP_LOOP_C_140, COMP_LOOP_C_141,
      COMP_LOOP_C_142, COMP_LOOP_C_143, COMP_LOOP_C_144, COMP_LOOP_C_145, COMP_LOOP_C_146,
      COMP_LOOP_C_147, COMP_LOOP_C_148, COMP_LOOP_C_149, COMP_LOOP_C_150, COMP_LOOP_C_151,
      COMP_LOOP_C_152, COMP_LOOP_C_153, COMP_LOOP_C_154, COMP_LOOP_C_155, COMP_LOOP_C_156,
      COMP_LOOP_C_157, COMP_LOOP_C_158, COMP_LOOP_C_159, COMP_LOOP_C_160, COMP_LOOP_C_161,
      COMP_LOOP_C_162, COMP_LOOP_C_163, COMP_LOOP_C_164, COMP_LOOP_C_165, COMP_LOOP_C_166,
      COMP_LOOP_C_167, COMP_LOOP_C_168, COMP_LOOP_C_169, COMP_LOOP_C_170, COMP_LOOP_C_171,
      COMP_LOOP_C_172, COMP_LOOP_C_173, COMP_LOOP_C_174, COMP_LOOP_C_175, COMP_LOOP_C_176,
      COMP_LOOP_C_177, COMP_LOOP_C_178, COMP_LOOP_C_179, COMP_LOOP_C_180, COMP_LOOP_C_181,
      COMP_LOOP_C_182, COMP_LOOP_C_183, COMP_LOOP_C_184, COMP_LOOP_C_185, COMP_LOOP_C_186,
      COMP_LOOP_C_187, COMP_LOOP_4_modExp_1_while_C_0, COMP_LOOP_4_modExp_1_while_C_1,
      COMP_LOOP_4_modExp_1_while_C_2, COMP_LOOP_4_modExp_1_while_C_3, COMP_LOOP_4_modExp_1_while_C_4,
      COMP_LOOP_4_modExp_1_while_C_5, COMP_LOOP_4_modExp_1_while_C_6, COMP_LOOP_4_modExp_1_while_C_7,
      COMP_LOOP_4_modExp_1_while_C_8, COMP_LOOP_4_modExp_1_while_C_9, COMP_LOOP_4_modExp_1_while_C_10,
      COMP_LOOP_4_modExp_1_while_C_11, COMP_LOOP_4_modExp_1_while_C_12, COMP_LOOP_4_modExp_1_while_C_13,
      COMP_LOOP_4_modExp_1_while_C_14, COMP_LOOP_4_modExp_1_while_C_15, COMP_LOOP_4_modExp_1_while_C_16,
      COMP_LOOP_4_modExp_1_while_C_17, COMP_LOOP_4_modExp_1_while_C_18, COMP_LOOP_4_modExp_1_while_C_19,
      COMP_LOOP_4_modExp_1_while_C_20, COMP_LOOP_4_modExp_1_while_C_21, COMP_LOOP_4_modExp_1_while_C_22,
      COMP_LOOP_4_modExp_1_while_C_23, COMP_LOOP_4_modExp_1_while_C_24, COMP_LOOP_4_modExp_1_while_C_25,
      COMP_LOOP_4_modExp_1_while_C_26, COMP_LOOP_4_modExp_1_while_C_27, COMP_LOOP_4_modExp_1_while_C_28,
      COMP_LOOP_4_modExp_1_while_C_29, COMP_LOOP_4_modExp_1_while_C_30, COMP_LOOP_4_modExp_1_while_C_31,
      COMP_LOOP_4_modExp_1_while_C_32, COMP_LOOP_4_modExp_1_while_C_33, COMP_LOOP_4_modExp_1_while_C_34,
      COMP_LOOP_4_modExp_1_while_C_35, COMP_LOOP_4_modExp_1_while_C_36, COMP_LOOP_4_modExp_1_while_C_37,
      COMP_LOOP_4_modExp_1_while_C_38, COMP_LOOP_C_188, COMP_LOOP_C_189, COMP_LOOP_C_190,
      COMP_LOOP_C_191, COMP_LOOP_C_192, COMP_LOOP_C_193, COMP_LOOP_C_194, COMP_LOOP_C_195,
      COMP_LOOP_C_196, COMP_LOOP_C_197, COMP_LOOP_C_198, COMP_LOOP_C_199, COMP_LOOP_C_200,
      COMP_LOOP_C_201, COMP_LOOP_C_202, COMP_LOOP_C_203, COMP_LOOP_C_204, COMP_LOOP_C_205,
      COMP_LOOP_C_206, COMP_LOOP_C_207, COMP_LOOP_C_208, COMP_LOOP_C_209, COMP_LOOP_C_210,
      COMP_LOOP_C_211, COMP_LOOP_C_212, COMP_LOOP_C_213, COMP_LOOP_C_214, COMP_LOOP_C_215,
      COMP_LOOP_C_216, COMP_LOOP_C_217, COMP_LOOP_C_218, COMP_LOOP_C_219, COMP_LOOP_C_220,
      COMP_LOOP_C_221, COMP_LOOP_C_222, COMP_LOOP_C_223, COMP_LOOP_C_224, COMP_LOOP_C_225,
      COMP_LOOP_C_226, COMP_LOOP_C_227, COMP_LOOP_C_228, COMP_LOOP_C_229, COMP_LOOP_C_230,
      COMP_LOOP_C_231, COMP_LOOP_C_232, COMP_LOOP_C_233, COMP_LOOP_C_234, COMP_LOOP_C_235,
      COMP_LOOP_C_236, COMP_LOOP_C_237, COMP_LOOP_C_238, COMP_LOOP_C_239, COMP_LOOP_C_240,
      COMP_LOOP_C_241, COMP_LOOP_C_242, COMP_LOOP_C_243, COMP_LOOP_C_244, COMP_LOOP_C_245,
      COMP_LOOP_C_246, COMP_LOOP_C_247, COMP_LOOP_C_248, COMP_LOOP_C_249, COMP_LOOP_5_modExp_1_while_C_0,
      COMP_LOOP_5_modExp_1_while_C_1, COMP_LOOP_5_modExp_1_while_C_2, COMP_LOOP_5_modExp_1_while_C_3,
      COMP_LOOP_5_modExp_1_while_C_4, COMP_LOOP_5_modExp_1_while_C_5, COMP_LOOP_5_modExp_1_while_C_6,
      COMP_LOOP_5_modExp_1_while_C_7, COMP_LOOP_5_modExp_1_while_C_8, COMP_LOOP_5_modExp_1_while_C_9,
      COMP_LOOP_5_modExp_1_while_C_10, COMP_LOOP_5_modExp_1_while_C_11, COMP_LOOP_5_modExp_1_while_C_12,
      COMP_LOOP_5_modExp_1_while_C_13, COMP_LOOP_5_modExp_1_while_C_14, COMP_LOOP_5_modExp_1_while_C_15,
      COMP_LOOP_5_modExp_1_while_C_16, COMP_LOOP_5_modExp_1_while_C_17, COMP_LOOP_5_modExp_1_while_C_18,
      COMP_LOOP_5_modExp_1_while_C_19, COMP_LOOP_5_modExp_1_while_C_20, COMP_LOOP_5_modExp_1_while_C_21,
      COMP_LOOP_5_modExp_1_while_C_22, COMP_LOOP_5_modExp_1_while_C_23, COMP_LOOP_5_modExp_1_while_C_24,
      COMP_LOOP_5_modExp_1_while_C_25, COMP_LOOP_5_modExp_1_while_C_26, COMP_LOOP_5_modExp_1_while_C_27,
      COMP_LOOP_5_modExp_1_while_C_28, COMP_LOOP_5_modExp_1_while_C_29, COMP_LOOP_5_modExp_1_while_C_30,
      COMP_LOOP_5_modExp_1_while_C_31, COMP_LOOP_5_modExp_1_while_C_32, COMP_LOOP_5_modExp_1_while_C_33,
      COMP_LOOP_5_modExp_1_while_C_34, COMP_LOOP_5_modExp_1_while_C_35, COMP_LOOP_5_modExp_1_while_C_36,
      COMP_LOOP_5_modExp_1_while_C_37, COMP_LOOP_5_modExp_1_while_C_38, COMP_LOOP_C_250,
      COMP_LOOP_C_251, COMP_LOOP_C_252, COMP_LOOP_C_253, COMP_LOOP_C_254, COMP_LOOP_C_255,
      COMP_LOOP_C_256, COMP_LOOP_C_257, COMP_LOOP_C_258, COMP_LOOP_C_259, COMP_LOOP_C_260,
      COMP_LOOP_C_261, COMP_LOOP_C_262, COMP_LOOP_C_263, COMP_LOOP_C_264, COMP_LOOP_C_265,
      COMP_LOOP_C_266, COMP_LOOP_C_267, COMP_LOOP_C_268, COMP_LOOP_C_269, COMP_LOOP_C_270,
      COMP_LOOP_C_271, COMP_LOOP_C_272, COMP_LOOP_C_273, COMP_LOOP_C_274, COMP_LOOP_C_275,
      COMP_LOOP_C_276, COMP_LOOP_C_277, COMP_LOOP_C_278, COMP_LOOP_C_279, COMP_LOOP_C_280,
      COMP_LOOP_C_281, COMP_LOOP_C_282, COMP_LOOP_C_283, COMP_LOOP_C_284, COMP_LOOP_C_285,
      COMP_LOOP_C_286, COMP_LOOP_C_287, COMP_LOOP_C_288, COMP_LOOP_C_289, COMP_LOOP_C_290,
      COMP_LOOP_C_291, COMP_LOOP_C_292, COMP_LOOP_C_293, COMP_LOOP_C_294, COMP_LOOP_C_295,
      COMP_LOOP_C_296, COMP_LOOP_C_297, COMP_LOOP_C_298, COMP_LOOP_C_299, COMP_LOOP_C_300,
      COMP_LOOP_C_301, COMP_LOOP_C_302, COMP_LOOP_C_303, COMP_LOOP_C_304, COMP_LOOP_C_305,
      COMP_LOOP_C_306, COMP_LOOP_C_307, COMP_LOOP_C_308, COMP_LOOP_C_309, COMP_LOOP_C_310,
      COMP_LOOP_C_311, COMP_LOOP_6_modExp_1_while_C_0, COMP_LOOP_6_modExp_1_while_C_1,
      COMP_LOOP_6_modExp_1_while_C_2, COMP_LOOP_6_modExp_1_while_C_3, COMP_LOOP_6_modExp_1_while_C_4,
      COMP_LOOP_6_modExp_1_while_C_5, COMP_LOOP_6_modExp_1_while_C_6, COMP_LOOP_6_modExp_1_while_C_7,
      COMP_LOOP_6_modExp_1_while_C_8, COMP_LOOP_6_modExp_1_while_C_9, COMP_LOOP_6_modExp_1_while_C_10,
      COMP_LOOP_6_modExp_1_while_C_11, COMP_LOOP_6_modExp_1_while_C_12, COMP_LOOP_6_modExp_1_while_C_13,
      COMP_LOOP_6_modExp_1_while_C_14, COMP_LOOP_6_modExp_1_while_C_15, COMP_LOOP_6_modExp_1_while_C_16,
      COMP_LOOP_6_modExp_1_while_C_17, COMP_LOOP_6_modExp_1_while_C_18, COMP_LOOP_6_modExp_1_while_C_19,
      COMP_LOOP_6_modExp_1_while_C_20, COMP_LOOP_6_modExp_1_while_C_21, COMP_LOOP_6_modExp_1_while_C_22,
      COMP_LOOP_6_modExp_1_while_C_23, COMP_LOOP_6_modExp_1_while_C_24, COMP_LOOP_6_modExp_1_while_C_25,
      COMP_LOOP_6_modExp_1_while_C_26, COMP_LOOP_6_modExp_1_while_C_27, COMP_LOOP_6_modExp_1_while_C_28,
      COMP_LOOP_6_modExp_1_while_C_29, COMP_LOOP_6_modExp_1_while_C_30, COMP_LOOP_6_modExp_1_while_C_31,
      COMP_LOOP_6_modExp_1_while_C_32, COMP_LOOP_6_modExp_1_while_C_33, COMP_LOOP_6_modExp_1_while_C_34,
      COMP_LOOP_6_modExp_1_while_C_35, COMP_LOOP_6_modExp_1_while_C_36, COMP_LOOP_6_modExp_1_while_C_37,
      COMP_LOOP_6_modExp_1_while_C_38, COMP_LOOP_C_312, COMP_LOOP_C_313, COMP_LOOP_C_314,
      COMP_LOOP_C_315, COMP_LOOP_C_316, COMP_LOOP_C_317, COMP_LOOP_C_318, COMP_LOOP_C_319,
      COMP_LOOP_C_320, COMP_LOOP_C_321, COMP_LOOP_C_322, COMP_LOOP_C_323, COMP_LOOP_C_324,
      COMP_LOOP_C_325, COMP_LOOP_C_326, COMP_LOOP_C_327, COMP_LOOP_C_328, COMP_LOOP_C_329,
      COMP_LOOP_C_330, COMP_LOOP_C_331, COMP_LOOP_C_332, COMP_LOOP_C_333, COMP_LOOP_C_334,
      COMP_LOOP_C_335, COMP_LOOP_C_336, COMP_LOOP_C_337, COMP_LOOP_C_338, COMP_LOOP_C_339,
      COMP_LOOP_C_340, COMP_LOOP_C_341, COMP_LOOP_C_342, COMP_LOOP_C_343, COMP_LOOP_C_344,
      COMP_LOOP_C_345, COMP_LOOP_C_346, COMP_LOOP_C_347, COMP_LOOP_C_348, COMP_LOOP_C_349,
      COMP_LOOP_C_350, COMP_LOOP_C_351, COMP_LOOP_C_352, COMP_LOOP_C_353, COMP_LOOP_C_354,
      COMP_LOOP_C_355, COMP_LOOP_C_356, COMP_LOOP_C_357, COMP_LOOP_C_358, COMP_LOOP_C_359,
      COMP_LOOP_C_360, COMP_LOOP_C_361, COMP_LOOP_C_362, COMP_LOOP_C_363, COMP_LOOP_C_364,
      COMP_LOOP_C_365, COMP_LOOP_C_366, COMP_LOOP_C_367, COMP_LOOP_C_368, COMP_LOOP_C_369,
      COMP_LOOP_C_370, COMP_LOOP_C_371, COMP_LOOP_C_372, COMP_LOOP_C_373, COMP_LOOP_7_modExp_1_while_C_0,
      COMP_LOOP_7_modExp_1_while_C_1, COMP_LOOP_7_modExp_1_while_C_2, COMP_LOOP_7_modExp_1_while_C_3,
      COMP_LOOP_7_modExp_1_while_C_4, COMP_LOOP_7_modExp_1_while_C_5, COMP_LOOP_7_modExp_1_while_C_6,
      COMP_LOOP_7_modExp_1_while_C_7, COMP_LOOP_7_modExp_1_while_C_8, COMP_LOOP_7_modExp_1_while_C_9,
      COMP_LOOP_7_modExp_1_while_C_10, COMP_LOOP_7_modExp_1_while_C_11, COMP_LOOP_7_modExp_1_while_C_12,
      COMP_LOOP_7_modExp_1_while_C_13, COMP_LOOP_7_modExp_1_while_C_14, COMP_LOOP_7_modExp_1_while_C_15,
      COMP_LOOP_7_modExp_1_while_C_16, COMP_LOOP_7_modExp_1_while_C_17, COMP_LOOP_7_modExp_1_while_C_18,
      COMP_LOOP_7_modExp_1_while_C_19, COMP_LOOP_7_modExp_1_while_C_20, COMP_LOOP_7_modExp_1_while_C_21,
      COMP_LOOP_7_modExp_1_while_C_22, COMP_LOOP_7_modExp_1_while_C_23, COMP_LOOP_7_modExp_1_while_C_24,
      COMP_LOOP_7_modExp_1_while_C_25, COMP_LOOP_7_modExp_1_while_C_26, COMP_LOOP_7_modExp_1_while_C_27,
      COMP_LOOP_7_modExp_1_while_C_28, COMP_LOOP_7_modExp_1_while_C_29, COMP_LOOP_7_modExp_1_while_C_30,
      COMP_LOOP_7_modExp_1_while_C_31, COMP_LOOP_7_modExp_1_while_C_32, COMP_LOOP_7_modExp_1_while_C_33,
      COMP_LOOP_7_modExp_1_while_C_34, COMP_LOOP_7_modExp_1_while_C_35, COMP_LOOP_7_modExp_1_while_C_36,
      COMP_LOOP_7_modExp_1_while_C_37, COMP_LOOP_7_modExp_1_while_C_38, COMP_LOOP_C_374,
      COMP_LOOP_C_375, COMP_LOOP_C_376, COMP_LOOP_C_377, COMP_LOOP_C_378, COMP_LOOP_C_379,
      COMP_LOOP_C_380, COMP_LOOP_C_381, COMP_LOOP_C_382, COMP_LOOP_C_383, COMP_LOOP_C_384,
      COMP_LOOP_C_385, COMP_LOOP_C_386, COMP_LOOP_C_387, COMP_LOOP_C_388, COMP_LOOP_C_389,
      COMP_LOOP_C_390, COMP_LOOP_C_391, COMP_LOOP_C_392, COMP_LOOP_C_393, COMP_LOOP_C_394,
      COMP_LOOP_C_395, COMP_LOOP_C_396, COMP_LOOP_C_397, COMP_LOOP_C_398, COMP_LOOP_C_399,
      COMP_LOOP_C_400, COMP_LOOP_C_401, COMP_LOOP_C_402, COMP_LOOP_C_403, COMP_LOOP_C_404,
      COMP_LOOP_C_405, COMP_LOOP_C_406, COMP_LOOP_C_407, COMP_LOOP_C_408, COMP_LOOP_C_409,
      COMP_LOOP_C_410, COMP_LOOP_C_411, COMP_LOOP_C_412, COMP_LOOP_C_413, COMP_LOOP_C_414,
      COMP_LOOP_C_415, COMP_LOOP_C_416, COMP_LOOP_C_417, COMP_LOOP_C_418, COMP_LOOP_C_419,
      COMP_LOOP_C_420, COMP_LOOP_C_421, COMP_LOOP_C_422, COMP_LOOP_C_423, COMP_LOOP_C_424,
      COMP_LOOP_C_425, COMP_LOOP_C_426, COMP_LOOP_C_427, COMP_LOOP_C_428, COMP_LOOP_C_429,
      COMP_LOOP_C_430, COMP_LOOP_C_431, COMP_LOOP_C_432, COMP_LOOP_C_433, COMP_LOOP_C_434,
      COMP_LOOP_C_435, COMP_LOOP_8_modExp_1_while_C_0, COMP_LOOP_8_modExp_1_while_C_1,
      COMP_LOOP_8_modExp_1_while_C_2, COMP_LOOP_8_modExp_1_while_C_3, COMP_LOOP_8_modExp_1_while_C_4,
      COMP_LOOP_8_modExp_1_while_C_5, COMP_LOOP_8_modExp_1_while_C_6, COMP_LOOP_8_modExp_1_while_C_7,
      COMP_LOOP_8_modExp_1_while_C_8, COMP_LOOP_8_modExp_1_while_C_9, COMP_LOOP_8_modExp_1_while_C_10,
      COMP_LOOP_8_modExp_1_while_C_11, COMP_LOOP_8_modExp_1_while_C_12, COMP_LOOP_8_modExp_1_while_C_13,
      COMP_LOOP_8_modExp_1_while_C_14, COMP_LOOP_8_modExp_1_while_C_15, COMP_LOOP_8_modExp_1_while_C_16,
      COMP_LOOP_8_modExp_1_while_C_17, COMP_LOOP_8_modExp_1_while_C_18, COMP_LOOP_8_modExp_1_while_C_19,
      COMP_LOOP_8_modExp_1_while_C_20, COMP_LOOP_8_modExp_1_while_C_21, COMP_LOOP_8_modExp_1_while_C_22,
      COMP_LOOP_8_modExp_1_while_C_23, COMP_LOOP_8_modExp_1_while_C_24, COMP_LOOP_8_modExp_1_while_C_25,
      COMP_LOOP_8_modExp_1_while_C_26, COMP_LOOP_8_modExp_1_while_C_27, COMP_LOOP_8_modExp_1_while_C_28,
      COMP_LOOP_8_modExp_1_while_C_29, COMP_LOOP_8_modExp_1_while_C_30, COMP_LOOP_8_modExp_1_while_C_31,
      COMP_LOOP_8_modExp_1_while_C_32, COMP_LOOP_8_modExp_1_while_C_33, COMP_LOOP_8_modExp_1_while_C_34,
      COMP_LOOP_8_modExp_1_while_C_35, COMP_LOOP_8_modExp_1_while_C_36, COMP_LOOP_8_modExp_1_while_C_37,
      COMP_LOOP_8_modExp_1_while_C_38, COMP_LOOP_C_436, COMP_LOOP_C_437, COMP_LOOP_C_438,
      COMP_LOOP_C_439, COMP_LOOP_C_440, COMP_LOOP_C_441, COMP_LOOP_C_442, COMP_LOOP_C_443,
      COMP_LOOP_C_444, COMP_LOOP_C_445, COMP_LOOP_C_446, COMP_LOOP_C_447, COMP_LOOP_C_448,
      COMP_LOOP_C_449, COMP_LOOP_C_450, COMP_LOOP_C_451, COMP_LOOP_C_452, COMP_LOOP_C_453,
      COMP_LOOP_C_454, COMP_LOOP_C_455, COMP_LOOP_C_456, COMP_LOOP_C_457, COMP_LOOP_C_458,
      COMP_LOOP_C_459, COMP_LOOP_C_460, COMP_LOOP_C_461, COMP_LOOP_C_462, COMP_LOOP_C_463,
      COMP_LOOP_C_464, COMP_LOOP_C_465, COMP_LOOP_C_466, COMP_LOOP_C_467, COMP_LOOP_C_468,
      COMP_LOOP_C_469, COMP_LOOP_C_470, COMP_LOOP_C_471, COMP_LOOP_C_472, COMP_LOOP_C_473,
      COMP_LOOP_C_474, COMP_LOOP_C_475, COMP_LOOP_C_476, COMP_LOOP_C_477, COMP_LOOP_C_478,
      COMP_LOOP_C_479, COMP_LOOP_C_480, COMP_LOOP_C_481, COMP_LOOP_C_482, COMP_LOOP_C_483,
      COMP_LOOP_C_484, COMP_LOOP_C_485, COMP_LOOP_C_486, COMP_LOOP_C_487, COMP_LOOP_C_488,
      COMP_LOOP_C_489, COMP_LOOP_C_490, COMP_LOOP_C_491, COMP_LOOP_C_492, COMP_LOOP_C_493,
      COMP_LOOP_C_494, COMP_LOOP_C_495, COMP_LOOP_C_496, VEC_LOOP_C_0, STAGE_LOOP_C_9,
      main_C_1);

  SIGNAL state_var : inPlaceNTT_DIT_core_core_fsm_1_ST;
  SIGNAL state_var_NS : inPlaceNTT_DIT_core_core_fsm_1_ST;

BEGIN
  inPlaceNTT_DIT_core_core_fsm_1 : PROCESS (STAGE_LOOP_C_8_tr0, modExp_while_C_38_tr0,
      COMP_LOOP_C_1_tr0, COMP_LOOP_1_modExp_1_while_C_38_tr0, COMP_LOOP_C_62_tr0,
      COMP_LOOP_2_modExp_1_while_C_38_tr0, COMP_LOOP_C_124_tr0, COMP_LOOP_3_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_186_tr0, COMP_LOOP_4_modExp_1_while_C_38_tr0, COMP_LOOP_C_248_tr0,
      COMP_LOOP_5_modExp_1_while_C_38_tr0, COMP_LOOP_C_310_tr0, COMP_LOOP_6_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_372_tr0, COMP_LOOP_7_modExp_1_while_C_38_tr0, COMP_LOOP_C_434_tr0,
      COMP_LOOP_8_modExp_1_while_C_38_tr0, COMP_LOOP_C_496_tr0, VEC_LOOP_C_0_tr0,
      STAGE_LOOP_C_9_tr0, state_var)
  BEGIN
    CASE state_var IS
      WHEN STAGE_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000001");
        state_var_NS <= STAGE_LOOP_C_1;
      WHEN STAGE_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000010");
        state_var_NS <= STAGE_LOOP_C_2;
      WHEN STAGE_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000011");
        state_var_NS <= STAGE_LOOP_C_3;
      WHEN STAGE_LOOP_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000100");
        state_var_NS <= STAGE_LOOP_C_4;
      WHEN STAGE_LOOP_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000101");
        state_var_NS <= STAGE_LOOP_C_5;
      WHEN STAGE_LOOP_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000110");
        state_var_NS <= STAGE_LOOP_C_6;
      WHEN STAGE_LOOP_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000111");
        state_var_NS <= STAGE_LOOP_C_7;
      WHEN STAGE_LOOP_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001000");
        state_var_NS <= STAGE_LOOP_C_8;
      WHEN STAGE_LOOP_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001001");
        IF ( STAGE_LOOP_C_8_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_0;
        ELSE
          state_var_NS <= modExp_while_C_0;
        END IF;
      WHEN modExp_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001010");
        state_var_NS <= modExp_while_C_1;
      WHEN modExp_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001011");
        state_var_NS <= modExp_while_C_2;
      WHEN modExp_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001100");
        state_var_NS <= modExp_while_C_3;
      WHEN modExp_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001101");
        state_var_NS <= modExp_while_C_4;
      WHEN modExp_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001110");
        state_var_NS <= modExp_while_C_5;
      WHEN modExp_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001111");
        state_var_NS <= modExp_while_C_6;
      WHEN modExp_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010000");
        state_var_NS <= modExp_while_C_7;
      WHEN modExp_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010001");
        state_var_NS <= modExp_while_C_8;
      WHEN modExp_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010010");
        state_var_NS <= modExp_while_C_9;
      WHEN modExp_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010011");
        state_var_NS <= modExp_while_C_10;
      WHEN modExp_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010100");
        state_var_NS <= modExp_while_C_11;
      WHEN modExp_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010101");
        state_var_NS <= modExp_while_C_12;
      WHEN modExp_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010110");
        state_var_NS <= modExp_while_C_13;
      WHEN modExp_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010111");
        state_var_NS <= modExp_while_C_14;
      WHEN modExp_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011000");
        state_var_NS <= modExp_while_C_15;
      WHEN modExp_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011001");
        state_var_NS <= modExp_while_C_16;
      WHEN modExp_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011010");
        state_var_NS <= modExp_while_C_17;
      WHEN modExp_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011011");
        state_var_NS <= modExp_while_C_18;
      WHEN modExp_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011100");
        state_var_NS <= modExp_while_C_19;
      WHEN modExp_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011101");
        state_var_NS <= modExp_while_C_20;
      WHEN modExp_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011110");
        state_var_NS <= modExp_while_C_21;
      WHEN modExp_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011111");
        state_var_NS <= modExp_while_C_22;
      WHEN modExp_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100000");
        state_var_NS <= modExp_while_C_23;
      WHEN modExp_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100001");
        state_var_NS <= modExp_while_C_24;
      WHEN modExp_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100010");
        state_var_NS <= modExp_while_C_25;
      WHEN modExp_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100011");
        state_var_NS <= modExp_while_C_26;
      WHEN modExp_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100100");
        state_var_NS <= modExp_while_C_27;
      WHEN modExp_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100101");
        state_var_NS <= modExp_while_C_28;
      WHEN modExp_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100110");
        state_var_NS <= modExp_while_C_29;
      WHEN modExp_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100111");
        state_var_NS <= modExp_while_C_30;
      WHEN modExp_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101000");
        state_var_NS <= modExp_while_C_31;
      WHEN modExp_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101001");
        state_var_NS <= modExp_while_C_32;
      WHEN modExp_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101010");
        state_var_NS <= modExp_while_C_33;
      WHEN modExp_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101011");
        state_var_NS <= modExp_while_C_34;
      WHEN modExp_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101100");
        state_var_NS <= modExp_while_C_35;
      WHEN modExp_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101101");
        state_var_NS <= modExp_while_C_36;
      WHEN modExp_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101110");
        state_var_NS <= modExp_while_C_37;
      WHEN modExp_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101111");
        state_var_NS <= modExp_while_C_38;
      WHEN modExp_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110000");
        IF ( modExp_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_0;
        ELSE
          state_var_NS <= modExp_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110001");
        state_var_NS <= COMP_LOOP_C_1;
      WHEN COMP_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110010");
        IF ( COMP_LOOP_C_1_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_2;
        ELSE
          state_var_NS <= COMP_LOOP_1_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_1_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110011");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_1;
      WHEN COMP_LOOP_1_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110100");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_2;
      WHEN COMP_LOOP_1_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110101");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_3;
      WHEN COMP_LOOP_1_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110110");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_4;
      WHEN COMP_LOOP_1_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110111");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_5;
      WHEN COMP_LOOP_1_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111000");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_6;
      WHEN COMP_LOOP_1_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111001");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_7;
      WHEN COMP_LOOP_1_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111010");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_8;
      WHEN COMP_LOOP_1_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111011");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_9;
      WHEN COMP_LOOP_1_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111100");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_10;
      WHEN COMP_LOOP_1_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111101");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_11;
      WHEN COMP_LOOP_1_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111110");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_12;
      WHEN COMP_LOOP_1_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111111");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_13;
      WHEN COMP_LOOP_1_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000000");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_14;
      WHEN COMP_LOOP_1_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000001");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_15;
      WHEN COMP_LOOP_1_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000010");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_16;
      WHEN COMP_LOOP_1_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000011");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_17;
      WHEN COMP_LOOP_1_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000100");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_18;
      WHEN COMP_LOOP_1_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000101");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_19;
      WHEN COMP_LOOP_1_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000110");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_20;
      WHEN COMP_LOOP_1_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000111");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_21;
      WHEN COMP_LOOP_1_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001000");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_22;
      WHEN COMP_LOOP_1_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001001");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_23;
      WHEN COMP_LOOP_1_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001010");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_24;
      WHEN COMP_LOOP_1_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001011");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_25;
      WHEN COMP_LOOP_1_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001100");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_26;
      WHEN COMP_LOOP_1_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001101");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_27;
      WHEN COMP_LOOP_1_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001110");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_28;
      WHEN COMP_LOOP_1_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001111");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_29;
      WHEN COMP_LOOP_1_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010000");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_30;
      WHEN COMP_LOOP_1_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010001");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_31;
      WHEN COMP_LOOP_1_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010010");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_32;
      WHEN COMP_LOOP_1_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010011");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_33;
      WHEN COMP_LOOP_1_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010100");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_34;
      WHEN COMP_LOOP_1_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010101");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_35;
      WHEN COMP_LOOP_1_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010110");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_36;
      WHEN COMP_LOOP_1_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010111");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_37;
      WHEN COMP_LOOP_1_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011000");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_38;
      WHEN COMP_LOOP_1_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011001");
        IF ( COMP_LOOP_1_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_2;
        ELSE
          state_var_NS <= COMP_LOOP_1_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011010");
        state_var_NS <= COMP_LOOP_C_3;
      WHEN COMP_LOOP_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011011");
        state_var_NS <= COMP_LOOP_C_4;
      WHEN COMP_LOOP_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011100");
        state_var_NS <= COMP_LOOP_C_5;
      WHEN COMP_LOOP_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011101");
        state_var_NS <= COMP_LOOP_C_6;
      WHEN COMP_LOOP_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011110");
        state_var_NS <= COMP_LOOP_C_7;
      WHEN COMP_LOOP_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011111");
        state_var_NS <= COMP_LOOP_C_8;
      WHEN COMP_LOOP_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100000");
        state_var_NS <= COMP_LOOP_C_9;
      WHEN COMP_LOOP_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100001");
        state_var_NS <= COMP_LOOP_C_10;
      WHEN COMP_LOOP_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100010");
        state_var_NS <= COMP_LOOP_C_11;
      WHEN COMP_LOOP_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100011");
        state_var_NS <= COMP_LOOP_C_12;
      WHEN COMP_LOOP_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100100");
        state_var_NS <= COMP_LOOP_C_13;
      WHEN COMP_LOOP_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100101");
        state_var_NS <= COMP_LOOP_C_14;
      WHEN COMP_LOOP_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100110");
        state_var_NS <= COMP_LOOP_C_15;
      WHEN COMP_LOOP_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100111");
        state_var_NS <= COMP_LOOP_C_16;
      WHEN COMP_LOOP_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101000");
        state_var_NS <= COMP_LOOP_C_17;
      WHEN COMP_LOOP_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101001");
        state_var_NS <= COMP_LOOP_C_18;
      WHEN COMP_LOOP_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101010");
        state_var_NS <= COMP_LOOP_C_19;
      WHEN COMP_LOOP_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101011");
        state_var_NS <= COMP_LOOP_C_20;
      WHEN COMP_LOOP_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101100");
        state_var_NS <= COMP_LOOP_C_21;
      WHEN COMP_LOOP_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101101");
        state_var_NS <= COMP_LOOP_C_22;
      WHEN COMP_LOOP_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101110");
        state_var_NS <= COMP_LOOP_C_23;
      WHEN COMP_LOOP_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101111");
        state_var_NS <= COMP_LOOP_C_24;
      WHEN COMP_LOOP_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110000");
        state_var_NS <= COMP_LOOP_C_25;
      WHEN COMP_LOOP_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110001");
        state_var_NS <= COMP_LOOP_C_26;
      WHEN COMP_LOOP_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110010");
        state_var_NS <= COMP_LOOP_C_27;
      WHEN COMP_LOOP_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110011");
        state_var_NS <= COMP_LOOP_C_28;
      WHEN COMP_LOOP_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110100");
        state_var_NS <= COMP_LOOP_C_29;
      WHEN COMP_LOOP_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110101");
        state_var_NS <= COMP_LOOP_C_30;
      WHEN COMP_LOOP_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110110");
        state_var_NS <= COMP_LOOP_C_31;
      WHEN COMP_LOOP_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110111");
        state_var_NS <= COMP_LOOP_C_32;
      WHEN COMP_LOOP_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111000");
        state_var_NS <= COMP_LOOP_C_33;
      WHEN COMP_LOOP_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111001");
        state_var_NS <= COMP_LOOP_C_34;
      WHEN COMP_LOOP_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111010");
        state_var_NS <= COMP_LOOP_C_35;
      WHEN COMP_LOOP_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111011");
        state_var_NS <= COMP_LOOP_C_36;
      WHEN COMP_LOOP_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111100");
        state_var_NS <= COMP_LOOP_C_37;
      WHEN COMP_LOOP_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111101");
        state_var_NS <= COMP_LOOP_C_38;
      WHEN COMP_LOOP_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111110");
        state_var_NS <= COMP_LOOP_C_39;
      WHEN COMP_LOOP_C_39 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111111");
        state_var_NS <= COMP_LOOP_C_40;
      WHEN COMP_LOOP_C_40 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000000");
        state_var_NS <= COMP_LOOP_C_41;
      WHEN COMP_LOOP_C_41 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000001");
        state_var_NS <= COMP_LOOP_C_42;
      WHEN COMP_LOOP_C_42 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000010");
        state_var_NS <= COMP_LOOP_C_43;
      WHEN COMP_LOOP_C_43 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000011");
        state_var_NS <= COMP_LOOP_C_44;
      WHEN COMP_LOOP_C_44 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000100");
        state_var_NS <= COMP_LOOP_C_45;
      WHEN COMP_LOOP_C_45 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000101");
        state_var_NS <= COMP_LOOP_C_46;
      WHEN COMP_LOOP_C_46 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000110");
        state_var_NS <= COMP_LOOP_C_47;
      WHEN COMP_LOOP_C_47 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000111");
        state_var_NS <= COMP_LOOP_C_48;
      WHEN COMP_LOOP_C_48 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001000");
        state_var_NS <= COMP_LOOP_C_49;
      WHEN COMP_LOOP_C_49 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001001");
        state_var_NS <= COMP_LOOP_C_50;
      WHEN COMP_LOOP_C_50 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001010");
        state_var_NS <= COMP_LOOP_C_51;
      WHEN COMP_LOOP_C_51 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001011");
        state_var_NS <= COMP_LOOP_C_52;
      WHEN COMP_LOOP_C_52 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001100");
        state_var_NS <= COMP_LOOP_C_53;
      WHEN COMP_LOOP_C_53 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001101");
        state_var_NS <= COMP_LOOP_C_54;
      WHEN COMP_LOOP_C_54 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001110");
        state_var_NS <= COMP_LOOP_C_55;
      WHEN COMP_LOOP_C_55 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001111");
        state_var_NS <= COMP_LOOP_C_56;
      WHEN COMP_LOOP_C_56 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010000");
        state_var_NS <= COMP_LOOP_C_57;
      WHEN COMP_LOOP_C_57 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010001");
        state_var_NS <= COMP_LOOP_C_58;
      WHEN COMP_LOOP_C_58 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010010");
        state_var_NS <= COMP_LOOP_C_59;
      WHEN COMP_LOOP_C_59 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010011");
        state_var_NS <= COMP_LOOP_C_60;
      WHEN COMP_LOOP_C_60 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010100");
        state_var_NS <= COMP_LOOP_C_61;
      WHEN COMP_LOOP_C_61 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010101");
        state_var_NS <= COMP_LOOP_C_62;
      WHEN COMP_LOOP_C_62 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010110");
        IF ( COMP_LOOP_C_62_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_63;
        END IF;
      WHEN COMP_LOOP_C_63 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010111");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_0;
      WHEN COMP_LOOP_2_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011000");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_1;
      WHEN COMP_LOOP_2_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011001");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_2;
      WHEN COMP_LOOP_2_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011010");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_3;
      WHEN COMP_LOOP_2_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011011");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_4;
      WHEN COMP_LOOP_2_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011100");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_5;
      WHEN COMP_LOOP_2_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011101");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_6;
      WHEN COMP_LOOP_2_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011110");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_7;
      WHEN COMP_LOOP_2_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011111");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_8;
      WHEN COMP_LOOP_2_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100000");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_9;
      WHEN COMP_LOOP_2_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100001");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_10;
      WHEN COMP_LOOP_2_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100010");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_11;
      WHEN COMP_LOOP_2_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100011");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_12;
      WHEN COMP_LOOP_2_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100100");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_13;
      WHEN COMP_LOOP_2_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100101");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_14;
      WHEN COMP_LOOP_2_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100110");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_15;
      WHEN COMP_LOOP_2_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100111");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_16;
      WHEN COMP_LOOP_2_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101000");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_17;
      WHEN COMP_LOOP_2_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101001");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_18;
      WHEN COMP_LOOP_2_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101010");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_19;
      WHEN COMP_LOOP_2_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101011");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_20;
      WHEN COMP_LOOP_2_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101100");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_21;
      WHEN COMP_LOOP_2_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101101");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_22;
      WHEN COMP_LOOP_2_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101110");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_23;
      WHEN COMP_LOOP_2_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101111");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_24;
      WHEN COMP_LOOP_2_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110000");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_25;
      WHEN COMP_LOOP_2_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110001");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_26;
      WHEN COMP_LOOP_2_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110010");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_27;
      WHEN COMP_LOOP_2_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110011");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_28;
      WHEN COMP_LOOP_2_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110100");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_29;
      WHEN COMP_LOOP_2_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110101");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_30;
      WHEN COMP_LOOP_2_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110110");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_31;
      WHEN COMP_LOOP_2_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110111");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_32;
      WHEN COMP_LOOP_2_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111000");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_33;
      WHEN COMP_LOOP_2_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111001");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_34;
      WHEN COMP_LOOP_2_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111010");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_35;
      WHEN COMP_LOOP_2_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111011");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_36;
      WHEN COMP_LOOP_2_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111100");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_37;
      WHEN COMP_LOOP_2_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111101");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_38;
      WHEN COMP_LOOP_2_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111110");
        IF ( COMP_LOOP_2_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_64;
        ELSE
          state_var_NS <= COMP_LOOP_2_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_64 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111111");
        state_var_NS <= COMP_LOOP_C_65;
      WHEN COMP_LOOP_C_65 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000000");
        state_var_NS <= COMP_LOOP_C_66;
      WHEN COMP_LOOP_C_66 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000001");
        state_var_NS <= COMP_LOOP_C_67;
      WHEN COMP_LOOP_C_67 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000010");
        state_var_NS <= COMP_LOOP_C_68;
      WHEN COMP_LOOP_C_68 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000011");
        state_var_NS <= COMP_LOOP_C_69;
      WHEN COMP_LOOP_C_69 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000100");
        state_var_NS <= COMP_LOOP_C_70;
      WHEN COMP_LOOP_C_70 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000101");
        state_var_NS <= COMP_LOOP_C_71;
      WHEN COMP_LOOP_C_71 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000110");
        state_var_NS <= COMP_LOOP_C_72;
      WHEN COMP_LOOP_C_72 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000111");
        state_var_NS <= COMP_LOOP_C_73;
      WHEN COMP_LOOP_C_73 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001000");
        state_var_NS <= COMP_LOOP_C_74;
      WHEN COMP_LOOP_C_74 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001001");
        state_var_NS <= COMP_LOOP_C_75;
      WHEN COMP_LOOP_C_75 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001010");
        state_var_NS <= COMP_LOOP_C_76;
      WHEN COMP_LOOP_C_76 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001011");
        state_var_NS <= COMP_LOOP_C_77;
      WHEN COMP_LOOP_C_77 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001100");
        state_var_NS <= COMP_LOOP_C_78;
      WHEN COMP_LOOP_C_78 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001101");
        state_var_NS <= COMP_LOOP_C_79;
      WHEN COMP_LOOP_C_79 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001110");
        state_var_NS <= COMP_LOOP_C_80;
      WHEN COMP_LOOP_C_80 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001111");
        state_var_NS <= COMP_LOOP_C_81;
      WHEN COMP_LOOP_C_81 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010000");
        state_var_NS <= COMP_LOOP_C_82;
      WHEN COMP_LOOP_C_82 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010001");
        state_var_NS <= COMP_LOOP_C_83;
      WHEN COMP_LOOP_C_83 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010010");
        state_var_NS <= COMP_LOOP_C_84;
      WHEN COMP_LOOP_C_84 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010011");
        state_var_NS <= COMP_LOOP_C_85;
      WHEN COMP_LOOP_C_85 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010100");
        state_var_NS <= COMP_LOOP_C_86;
      WHEN COMP_LOOP_C_86 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010101");
        state_var_NS <= COMP_LOOP_C_87;
      WHEN COMP_LOOP_C_87 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010110");
        state_var_NS <= COMP_LOOP_C_88;
      WHEN COMP_LOOP_C_88 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010111");
        state_var_NS <= COMP_LOOP_C_89;
      WHEN COMP_LOOP_C_89 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011000");
        state_var_NS <= COMP_LOOP_C_90;
      WHEN COMP_LOOP_C_90 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011001");
        state_var_NS <= COMP_LOOP_C_91;
      WHEN COMP_LOOP_C_91 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011010");
        state_var_NS <= COMP_LOOP_C_92;
      WHEN COMP_LOOP_C_92 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011011");
        state_var_NS <= COMP_LOOP_C_93;
      WHEN COMP_LOOP_C_93 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011100");
        state_var_NS <= COMP_LOOP_C_94;
      WHEN COMP_LOOP_C_94 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011101");
        state_var_NS <= COMP_LOOP_C_95;
      WHEN COMP_LOOP_C_95 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011110");
        state_var_NS <= COMP_LOOP_C_96;
      WHEN COMP_LOOP_C_96 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011111");
        state_var_NS <= COMP_LOOP_C_97;
      WHEN COMP_LOOP_C_97 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100000");
        state_var_NS <= COMP_LOOP_C_98;
      WHEN COMP_LOOP_C_98 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100001");
        state_var_NS <= COMP_LOOP_C_99;
      WHEN COMP_LOOP_C_99 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100010");
        state_var_NS <= COMP_LOOP_C_100;
      WHEN COMP_LOOP_C_100 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100011");
        state_var_NS <= COMP_LOOP_C_101;
      WHEN COMP_LOOP_C_101 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100100");
        state_var_NS <= COMP_LOOP_C_102;
      WHEN COMP_LOOP_C_102 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100101");
        state_var_NS <= COMP_LOOP_C_103;
      WHEN COMP_LOOP_C_103 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100110");
        state_var_NS <= COMP_LOOP_C_104;
      WHEN COMP_LOOP_C_104 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100111");
        state_var_NS <= COMP_LOOP_C_105;
      WHEN COMP_LOOP_C_105 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101000");
        state_var_NS <= COMP_LOOP_C_106;
      WHEN COMP_LOOP_C_106 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101001");
        state_var_NS <= COMP_LOOP_C_107;
      WHEN COMP_LOOP_C_107 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101010");
        state_var_NS <= COMP_LOOP_C_108;
      WHEN COMP_LOOP_C_108 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101011");
        state_var_NS <= COMP_LOOP_C_109;
      WHEN COMP_LOOP_C_109 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101100");
        state_var_NS <= COMP_LOOP_C_110;
      WHEN COMP_LOOP_C_110 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101101");
        state_var_NS <= COMP_LOOP_C_111;
      WHEN COMP_LOOP_C_111 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101110");
        state_var_NS <= COMP_LOOP_C_112;
      WHEN COMP_LOOP_C_112 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101111");
        state_var_NS <= COMP_LOOP_C_113;
      WHEN COMP_LOOP_C_113 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110000");
        state_var_NS <= COMP_LOOP_C_114;
      WHEN COMP_LOOP_C_114 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110001");
        state_var_NS <= COMP_LOOP_C_115;
      WHEN COMP_LOOP_C_115 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110010");
        state_var_NS <= COMP_LOOP_C_116;
      WHEN COMP_LOOP_C_116 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110011");
        state_var_NS <= COMP_LOOP_C_117;
      WHEN COMP_LOOP_C_117 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110100");
        state_var_NS <= COMP_LOOP_C_118;
      WHEN COMP_LOOP_C_118 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110101");
        state_var_NS <= COMP_LOOP_C_119;
      WHEN COMP_LOOP_C_119 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110110");
        state_var_NS <= COMP_LOOP_C_120;
      WHEN COMP_LOOP_C_120 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110111");
        state_var_NS <= COMP_LOOP_C_121;
      WHEN COMP_LOOP_C_121 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111000");
        state_var_NS <= COMP_LOOP_C_122;
      WHEN COMP_LOOP_C_122 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111001");
        state_var_NS <= COMP_LOOP_C_123;
      WHEN COMP_LOOP_C_123 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111010");
        state_var_NS <= COMP_LOOP_C_124;
      WHEN COMP_LOOP_C_124 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111011");
        IF ( COMP_LOOP_C_124_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_125;
        END IF;
      WHEN COMP_LOOP_C_125 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111100");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_0;
      WHEN COMP_LOOP_3_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111101");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_1;
      WHEN COMP_LOOP_3_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111110");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_2;
      WHEN COMP_LOOP_3_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111111");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_3;
      WHEN COMP_LOOP_3_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000000");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_4;
      WHEN COMP_LOOP_3_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000001");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_5;
      WHEN COMP_LOOP_3_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000010");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_6;
      WHEN COMP_LOOP_3_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000011");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_7;
      WHEN COMP_LOOP_3_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000100");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_8;
      WHEN COMP_LOOP_3_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000101");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_9;
      WHEN COMP_LOOP_3_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000110");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_10;
      WHEN COMP_LOOP_3_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000111");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_11;
      WHEN COMP_LOOP_3_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001000");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_12;
      WHEN COMP_LOOP_3_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001001");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_13;
      WHEN COMP_LOOP_3_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001010");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_14;
      WHEN COMP_LOOP_3_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001011");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_15;
      WHEN COMP_LOOP_3_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001100");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_16;
      WHEN COMP_LOOP_3_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001101");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_17;
      WHEN COMP_LOOP_3_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001110");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_18;
      WHEN COMP_LOOP_3_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001111");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_19;
      WHEN COMP_LOOP_3_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010000");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_20;
      WHEN COMP_LOOP_3_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010001");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_21;
      WHEN COMP_LOOP_3_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010010");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_22;
      WHEN COMP_LOOP_3_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010011");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_23;
      WHEN COMP_LOOP_3_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010100");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_24;
      WHEN COMP_LOOP_3_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010101");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_25;
      WHEN COMP_LOOP_3_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010110");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_26;
      WHEN COMP_LOOP_3_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010111");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_27;
      WHEN COMP_LOOP_3_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011000");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_28;
      WHEN COMP_LOOP_3_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011001");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_29;
      WHEN COMP_LOOP_3_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011010");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_30;
      WHEN COMP_LOOP_3_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011011");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_31;
      WHEN COMP_LOOP_3_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011100");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_32;
      WHEN COMP_LOOP_3_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011101");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_33;
      WHEN COMP_LOOP_3_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011110");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_34;
      WHEN COMP_LOOP_3_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011111");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_35;
      WHEN COMP_LOOP_3_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100000");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_36;
      WHEN COMP_LOOP_3_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100001");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_37;
      WHEN COMP_LOOP_3_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100010");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_38;
      WHEN COMP_LOOP_3_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100011");
        IF ( COMP_LOOP_3_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_126;
        ELSE
          state_var_NS <= COMP_LOOP_3_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_126 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100100");
        state_var_NS <= COMP_LOOP_C_127;
      WHEN COMP_LOOP_C_127 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100101");
        state_var_NS <= COMP_LOOP_C_128;
      WHEN COMP_LOOP_C_128 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100110");
        state_var_NS <= COMP_LOOP_C_129;
      WHEN COMP_LOOP_C_129 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100111");
        state_var_NS <= COMP_LOOP_C_130;
      WHEN COMP_LOOP_C_130 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101000");
        state_var_NS <= COMP_LOOP_C_131;
      WHEN COMP_LOOP_C_131 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101001");
        state_var_NS <= COMP_LOOP_C_132;
      WHEN COMP_LOOP_C_132 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101010");
        state_var_NS <= COMP_LOOP_C_133;
      WHEN COMP_LOOP_C_133 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101011");
        state_var_NS <= COMP_LOOP_C_134;
      WHEN COMP_LOOP_C_134 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101100");
        state_var_NS <= COMP_LOOP_C_135;
      WHEN COMP_LOOP_C_135 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101101");
        state_var_NS <= COMP_LOOP_C_136;
      WHEN COMP_LOOP_C_136 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101110");
        state_var_NS <= COMP_LOOP_C_137;
      WHEN COMP_LOOP_C_137 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101111");
        state_var_NS <= COMP_LOOP_C_138;
      WHEN COMP_LOOP_C_138 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110000");
        state_var_NS <= COMP_LOOP_C_139;
      WHEN COMP_LOOP_C_139 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110001");
        state_var_NS <= COMP_LOOP_C_140;
      WHEN COMP_LOOP_C_140 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110010");
        state_var_NS <= COMP_LOOP_C_141;
      WHEN COMP_LOOP_C_141 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110011");
        state_var_NS <= COMP_LOOP_C_142;
      WHEN COMP_LOOP_C_142 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110100");
        state_var_NS <= COMP_LOOP_C_143;
      WHEN COMP_LOOP_C_143 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110101");
        state_var_NS <= COMP_LOOP_C_144;
      WHEN COMP_LOOP_C_144 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110110");
        state_var_NS <= COMP_LOOP_C_145;
      WHEN COMP_LOOP_C_145 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110111");
        state_var_NS <= COMP_LOOP_C_146;
      WHEN COMP_LOOP_C_146 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111000");
        state_var_NS <= COMP_LOOP_C_147;
      WHEN COMP_LOOP_C_147 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111001");
        state_var_NS <= COMP_LOOP_C_148;
      WHEN COMP_LOOP_C_148 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111010");
        state_var_NS <= COMP_LOOP_C_149;
      WHEN COMP_LOOP_C_149 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111011");
        state_var_NS <= COMP_LOOP_C_150;
      WHEN COMP_LOOP_C_150 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111100");
        state_var_NS <= COMP_LOOP_C_151;
      WHEN COMP_LOOP_C_151 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111101");
        state_var_NS <= COMP_LOOP_C_152;
      WHEN COMP_LOOP_C_152 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111110");
        state_var_NS <= COMP_LOOP_C_153;
      WHEN COMP_LOOP_C_153 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111111");
        state_var_NS <= COMP_LOOP_C_154;
      WHEN COMP_LOOP_C_154 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000000");
        state_var_NS <= COMP_LOOP_C_155;
      WHEN COMP_LOOP_C_155 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000001");
        state_var_NS <= COMP_LOOP_C_156;
      WHEN COMP_LOOP_C_156 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000010");
        state_var_NS <= COMP_LOOP_C_157;
      WHEN COMP_LOOP_C_157 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000011");
        state_var_NS <= COMP_LOOP_C_158;
      WHEN COMP_LOOP_C_158 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000100");
        state_var_NS <= COMP_LOOP_C_159;
      WHEN COMP_LOOP_C_159 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000101");
        state_var_NS <= COMP_LOOP_C_160;
      WHEN COMP_LOOP_C_160 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000110");
        state_var_NS <= COMP_LOOP_C_161;
      WHEN COMP_LOOP_C_161 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000111");
        state_var_NS <= COMP_LOOP_C_162;
      WHEN COMP_LOOP_C_162 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001000");
        state_var_NS <= COMP_LOOP_C_163;
      WHEN COMP_LOOP_C_163 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001001");
        state_var_NS <= COMP_LOOP_C_164;
      WHEN COMP_LOOP_C_164 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001010");
        state_var_NS <= COMP_LOOP_C_165;
      WHEN COMP_LOOP_C_165 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001011");
        state_var_NS <= COMP_LOOP_C_166;
      WHEN COMP_LOOP_C_166 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001100");
        state_var_NS <= COMP_LOOP_C_167;
      WHEN COMP_LOOP_C_167 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001101");
        state_var_NS <= COMP_LOOP_C_168;
      WHEN COMP_LOOP_C_168 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001110");
        state_var_NS <= COMP_LOOP_C_169;
      WHEN COMP_LOOP_C_169 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001111");
        state_var_NS <= COMP_LOOP_C_170;
      WHEN COMP_LOOP_C_170 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010000");
        state_var_NS <= COMP_LOOP_C_171;
      WHEN COMP_LOOP_C_171 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010001");
        state_var_NS <= COMP_LOOP_C_172;
      WHEN COMP_LOOP_C_172 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010010");
        state_var_NS <= COMP_LOOP_C_173;
      WHEN COMP_LOOP_C_173 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010011");
        state_var_NS <= COMP_LOOP_C_174;
      WHEN COMP_LOOP_C_174 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010100");
        state_var_NS <= COMP_LOOP_C_175;
      WHEN COMP_LOOP_C_175 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010101");
        state_var_NS <= COMP_LOOP_C_176;
      WHEN COMP_LOOP_C_176 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010110");
        state_var_NS <= COMP_LOOP_C_177;
      WHEN COMP_LOOP_C_177 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010111");
        state_var_NS <= COMP_LOOP_C_178;
      WHEN COMP_LOOP_C_178 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011000");
        state_var_NS <= COMP_LOOP_C_179;
      WHEN COMP_LOOP_C_179 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011001");
        state_var_NS <= COMP_LOOP_C_180;
      WHEN COMP_LOOP_C_180 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011010");
        state_var_NS <= COMP_LOOP_C_181;
      WHEN COMP_LOOP_C_181 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011011");
        state_var_NS <= COMP_LOOP_C_182;
      WHEN COMP_LOOP_C_182 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011100");
        state_var_NS <= COMP_LOOP_C_183;
      WHEN COMP_LOOP_C_183 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011101");
        state_var_NS <= COMP_LOOP_C_184;
      WHEN COMP_LOOP_C_184 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011110");
        state_var_NS <= COMP_LOOP_C_185;
      WHEN COMP_LOOP_C_185 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011111");
        state_var_NS <= COMP_LOOP_C_186;
      WHEN COMP_LOOP_C_186 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100000");
        IF ( COMP_LOOP_C_186_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_187;
        END IF;
      WHEN COMP_LOOP_C_187 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100001");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_0;
      WHEN COMP_LOOP_4_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100010");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_1;
      WHEN COMP_LOOP_4_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100011");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_2;
      WHEN COMP_LOOP_4_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100100");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_3;
      WHEN COMP_LOOP_4_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100101");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_4;
      WHEN COMP_LOOP_4_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100110");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_5;
      WHEN COMP_LOOP_4_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100111");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_6;
      WHEN COMP_LOOP_4_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101000");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_7;
      WHEN COMP_LOOP_4_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101001");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_8;
      WHEN COMP_LOOP_4_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101010");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_9;
      WHEN COMP_LOOP_4_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101011");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_10;
      WHEN COMP_LOOP_4_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101100");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_11;
      WHEN COMP_LOOP_4_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101101");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_12;
      WHEN COMP_LOOP_4_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101110");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_13;
      WHEN COMP_LOOP_4_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101111");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_14;
      WHEN COMP_LOOP_4_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110000");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_15;
      WHEN COMP_LOOP_4_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110001");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_16;
      WHEN COMP_LOOP_4_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110010");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_17;
      WHEN COMP_LOOP_4_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110011");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_18;
      WHEN COMP_LOOP_4_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110100");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_19;
      WHEN COMP_LOOP_4_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110101");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_20;
      WHEN COMP_LOOP_4_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110110");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_21;
      WHEN COMP_LOOP_4_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110111");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_22;
      WHEN COMP_LOOP_4_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111000");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_23;
      WHEN COMP_LOOP_4_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111001");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_24;
      WHEN COMP_LOOP_4_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111010");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_25;
      WHEN COMP_LOOP_4_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111011");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_26;
      WHEN COMP_LOOP_4_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111100");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_27;
      WHEN COMP_LOOP_4_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111101");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_28;
      WHEN COMP_LOOP_4_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111110");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_29;
      WHEN COMP_LOOP_4_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111111");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_30;
      WHEN COMP_LOOP_4_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000000");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_31;
      WHEN COMP_LOOP_4_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000001");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_32;
      WHEN COMP_LOOP_4_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000010");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_33;
      WHEN COMP_LOOP_4_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000011");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_34;
      WHEN COMP_LOOP_4_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000100");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_35;
      WHEN COMP_LOOP_4_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000101");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_36;
      WHEN COMP_LOOP_4_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000110");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_37;
      WHEN COMP_LOOP_4_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000111");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_38;
      WHEN COMP_LOOP_4_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001000");
        IF ( COMP_LOOP_4_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_188;
        ELSE
          state_var_NS <= COMP_LOOP_4_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_188 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001001");
        state_var_NS <= COMP_LOOP_C_189;
      WHEN COMP_LOOP_C_189 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001010");
        state_var_NS <= COMP_LOOP_C_190;
      WHEN COMP_LOOP_C_190 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001011");
        state_var_NS <= COMP_LOOP_C_191;
      WHEN COMP_LOOP_C_191 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001100");
        state_var_NS <= COMP_LOOP_C_192;
      WHEN COMP_LOOP_C_192 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001101");
        state_var_NS <= COMP_LOOP_C_193;
      WHEN COMP_LOOP_C_193 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001110");
        state_var_NS <= COMP_LOOP_C_194;
      WHEN COMP_LOOP_C_194 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001111");
        state_var_NS <= COMP_LOOP_C_195;
      WHEN COMP_LOOP_C_195 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010000");
        state_var_NS <= COMP_LOOP_C_196;
      WHEN COMP_LOOP_C_196 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010001");
        state_var_NS <= COMP_LOOP_C_197;
      WHEN COMP_LOOP_C_197 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010010");
        state_var_NS <= COMP_LOOP_C_198;
      WHEN COMP_LOOP_C_198 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010011");
        state_var_NS <= COMP_LOOP_C_199;
      WHEN COMP_LOOP_C_199 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010100");
        state_var_NS <= COMP_LOOP_C_200;
      WHEN COMP_LOOP_C_200 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010101");
        state_var_NS <= COMP_LOOP_C_201;
      WHEN COMP_LOOP_C_201 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010110");
        state_var_NS <= COMP_LOOP_C_202;
      WHEN COMP_LOOP_C_202 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010111");
        state_var_NS <= COMP_LOOP_C_203;
      WHEN COMP_LOOP_C_203 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011000");
        state_var_NS <= COMP_LOOP_C_204;
      WHEN COMP_LOOP_C_204 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011001");
        state_var_NS <= COMP_LOOP_C_205;
      WHEN COMP_LOOP_C_205 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011010");
        state_var_NS <= COMP_LOOP_C_206;
      WHEN COMP_LOOP_C_206 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011011");
        state_var_NS <= COMP_LOOP_C_207;
      WHEN COMP_LOOP_C_207 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011100");
        state_var_NS <= COMP_LOOP_C_208;
      WHEN COMP_LOOP_C_208 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011101");
        state_var_NS <= COMP_LOOP_C_209;
      WHEN COMP_LOOP_C_209 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011110");
        state_var_NS <= COMP_LOOP_C_210;
      WHEN COMP_LOOP_C_210 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011111");
        state_var_NS <= COMP_LOOP_C_211;
      WHEN COMP_LOOP_C_211 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100000");
        state_var_NS <= COMP_LOOP_C_212;
      WHEN COMP_LOOP_C_212 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100001");
        state_var_NS <= COMP_LOOP_C_213;
      WHEN COMP_LOOP_C_213 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100010");
        state_var_NS <= COMP_LOOP_C_214;
      WHEN COMP_LOOP_C_214 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100011");
        state_var_NS <= COMP_LOOP_C_215;
      WHEN COMP_LOOP_C_215 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100100");
        state_var_NS <= COMP_LOOP_C_216;
      WHEN COMP_LOOP_C_216 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100101");
        state_var_NS <= COMP_LOOP_C_217;
      WHEN COMP_LOOP_C_217 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100110");
        state_var_NS <= COMP_LOOP_C_218;
      WHEN COMP_LOOP_C_218 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100111");
        state_var_NS <= COMP_LOOP_C_219;
      WHEN COMP_LOOP_C_219 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101000");
        state_var_NS <= COMP_LOOP_C_220;
      WHEN COMP_LOOP_C_220 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101001");
        state_var_NS <= COMP_LOOP_C_221;
      WHEN COMP_LOOP_C_221 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101010");
        state_var_NS <= COMP_LOOP_C_222;
      WHEN COMP_LOOP_C_222 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101011");
        state_var_NS <= COMP_LOOP_C_223;
      WHEN COMP_LOOP_C_223 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101100");
        state_var_NS <= COMP_LOOP_C_224;
      WHEN COMP_LOOP_C_224 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101101");
        state_var_NS <= COMP_LOOP_C_225;
      WHEN COMP_LOOP_C_225 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101110");
        state_var_NS <= COMP_LOOP_C_226;
      WHEN COMP_LOOP_C_226 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101111");
        state_var_NS <= COMP_LOOP_C_227;
      WHEN COMP_LOOP_C_227 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110000");
        state_var_NS <= COMP_LOOP_C_228;
      WHEN COMP_LOOP_C_228 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110001");
        state_var_NS <= COMP_LOOP_C_229;
      WHEN COMP_LOOP_C_229 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110010");
        state_var_NS <= COMP_LOOP_C_230;
      WHEN COMP_LOOP_C_230 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110011");
        state_var_NS <= COMP_LOOP_C_231;
      WHEN COMP_LOOP_C_231 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110100");
        state_var_NS <= COMP_LOOP_C_232;
      WHEN COMP_LOOP_C_232 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110101");
        state_var_NS <= COMP_LOOP_C_233;
      WHEN COMP_LOOP_C_233 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110110");
        state_var_NS <= COMP_LOOP_C_234;
      WHEN COMP_LOOP_C_234 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110111");
        state_var_NS <= COMP_LOOP_C_235;
      WHEN COMP_LOOP_C_235 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111000");
        state_var_NS <= COMP_LOOP_C_236;
      WHEN COMP_LOOP_C_236 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111001");
        state_var_NS <= COMP_LOOP_C_237;
      WHEN COMP_LOOP_C_237 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111010");
        state_var_NS <= COMP_LOOP_C_238;
      WHEN COMP_LOOP_C_238 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111011");
        state_var_NS <= COMP_LOOP_C_239;
      WHEN COMP_LOOP_C_239 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111100");
        state_var_NS <= COMP_LOOP_C_240;
      WHEN COMP_LOOP_C_240 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111101");
        state_var_NS <= COMP_LOOP_C_241;
      WHEN COMP_LOOP_C_241 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111110");
        state_var_NS <= COMP_LOOP_C_242;
      WHEN COMP_LOOP_C_242 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111111");
        state_var_NS <= COMP_LOOP_C_243;
      WHEN COMP_LOOP_C_243 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000000");
        state_var_NS <= COMP_LOOP_C_244;
      WHEN COMP_LOOP_C_244 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000001");
        state_var_NS <= COMP_LOOP_C_245;
      WHEN COMP_LOOP_C_245 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000010");
        state_var_NS <= COMP_LOOP_C_246;
      WHEN COMP_LOOP_C_246 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000011");
        state_var_NS <= COMP_LOOP_C_247;
      WHEN COMP_LOOP_C_247 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000100");
        state_var_NS <= COMP_LOOP_C_248;
      WHEN COMP_LOOP_C_248 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000101");
        IF ( COMP_LOOP_C_248_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_249;
        END IF;
      WHEN COMP_LOOP_C_249 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000110");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_0;
      WHEN COMP_LOOP_5_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000111");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_1;
      WHEN COMP_LOOP_5_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001000");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_2;
      WHEN COMP_LOOP_5_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001001");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_3;
      WHEN COMP_LOOP_5_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001010");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_4;
      WHEN COMP_LOOP_5_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001011");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_5;
      WHEN COMP_LOOP_5_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001100");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_6;
      WHEN COMP_LOOP_5_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001101");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_7;
      WHEN COMP_LOOP_5_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001110");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_8;
      WHEN COMP_LOOP_5_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001111");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_9;
      WHEN COMP_LOOP_5_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010000");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_10;
      WHEN COMP_LOOP_5_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010001");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_11;
      WHEN COMP_LOOP_5_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010010");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_12;
      WHEN COMP_LOOP_5_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010011");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_13;
      WHEN COMP_LOOP_5_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010100");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_14;
      WHEN COMP_LOOP_5_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010101");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_15;
      WHEN COMP_LOOP_5_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010110");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_16;
      WHEN COMP_LOOP_5_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010111");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_17;
      WHEN COMP_LOOP_5_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011000");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_18;
      WHEN COMP_LOOP_5_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011001");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_19;
      WHEN COMP_LOOP_5_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011010");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_20;
      WHEN COMP_LOOP_5_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011011");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_21;
      WHEN COMP_LOOP_5_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011100");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_22;
      WHEN COMP_LOOP_5_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011101");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_23;
      WHEN COMP_LOOP_5_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011110");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_24;
      WHEN COMP_LOOP_5_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011111");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_25;
      WHEN COMP_LOOP_5_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100000");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_26;
      WHEN COMP_LOOP_5_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100001");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_27;
      WHEN COMP_LOOP_5_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100010");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_28;
      WHEN COMP_LOOP_5_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100011");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_29;
      WHEN COMP_LOOP_5_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100100");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_30;
      WHEN COMP_LOOP_5_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100101");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_31;
      WHEN COMP_LOOP_5_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100110");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_32;
      WHEN COMP_LOOP_5_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100111");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_33;
      WHEN COMP_LOOP_5_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101000");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_34;
      WHEN COMP_LOOP_5_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101001");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_35;
      WHEN COMP_LOOP_5_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101010");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_36;
      WHEN COMP_LOOP_5_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101011");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_37;
      WHEN COMP_LOOP_5_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101100");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_38;
      WHEN COMP_LOOP_5_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101101");
        IF ( COMP_LOOP_5_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_250;
        ELSE
          state_var_NS <= COMP_LOOP_5_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_250 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101110");
        state_var_NS <= COMP_LOOP_C_251;
      WHEN COMP_LOOP_C_251 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101111");
        state_var_NS <= COMP_LOOP_C_252;
      WHEN COMP_LOOP_C_252 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110000");
        state_var_NS <= COMP_LOOP_C_253;
      WHEN COMP_LOOP_C_253 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110001");
        state_var_NS <= COMP_LOOP_C_254;
      WHEN COMP_LOOP_C_254 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110010");
        state_var_NS <= COMP_LOOP_C_255;
      WHEN COMP_LOOP_C_255 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110011");
        state_var_NS <= COMP_LOOP_C_256;
      WHEN COMP_LOOP_C_256 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110100");
        state_var_NS <= COMP_LOOP_C_257;
      WHEN COMP_LOOP_C_257 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110101");
        state_var_NS <= COMP_LOOP_C_258;
      WHEN COMP_LOOP_C_258 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110110");
        state_var_NS <= COMP_LOOP_C_259;
      WHEN COMP_LOOP_C_259 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110111");
        state_var_NS <= COMP_LOOP_C_260;
      WHEN COMP_LOOP_C_260 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111000");
        state_var_NS <= COMP_LOOP_C_261;
      WHEN COMP_LOOP_C_261 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111001");
        state_var_NS <= COMP_LOOP_C_262;
      WHEN COMP_LOOP_C_262 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111010");
        state_var_NS <= COMP_LOOP_C_263;
      WHEN COMP_LOOP_C_263 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111011");
        state_var_NS <= COMP_LOOP_C_264;
      WHEN COMP_LOOP_C_264 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111100");
        state_var_NS <= COMP_LOOP_C_265;
      WHEN COMP_LOOP_C_265 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111101");
        state_var_NS <= COMP_LOOP_C_266;
      WHEN COMP_LOOP_C_266 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111110");
        state_var_NS <= COMP_LOOP_C_267;
      WHEN COMP_LOOP_C_267 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111111");
        state_var_NS <= COMP_LOOP_C_268;
      WHEN COMP_LOOP_C_268 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000000");
        state_var_NS <= COMP_LOOP_C_269;
      WHEN COMP_LOOP_C_269 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000001");
        state_var_NS <= COMP_LOOP_C_270;
      WHEN COMP_LOOP_C_270 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000010");
        state_var_NS <= COMP_LOOP_C_271;
      WHEN COMP_LOOP_C_271 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000011");
        state_var_NS <= COMP_LOOP_C_272;
      WHEN COMP_LOOP_C_272 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000100");
        state_var_NS <= COMP_LOOP_C_273;
      WHEN COMP_LOOP_C_273 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000101");
        state_var_NS <= COMP_LOOP_C_274;
      WHEN COMP_LOOP_C_274 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000110");
        state_var_NS <= COMP_LOOP_C_275;
      WHEN COMP_LOOP_C_275 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000111");
        state_var_NS <= COMP_LOOP_C_276;
      WHEN COMP_LOOP_C_276 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001000");
        state_var_NS <= COMP_LOOP_C_277;
      WHEN COMP_LOOP_C_277 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001001");
        state_var_NS <= COMP_LOOP_C_278;
      WHEN COMP_LOOP_C_278 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001010");
        state_var_NS <= COMP_LOOP_C_279;
      WHEN COMP_LOOP_C_279 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001011");
        state_var_NS <= COMP_LOOP_C_280;
      WHEN COMP_LOOP_C_280 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001100");
        state_var_NS <= COMP_LOOP_C_281;
      WHEN COMP_LOOP_C_281 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001101");
        state_var_NS <= COMP_LOOP_C_282;
      WHEN COMP_LOOP_C_282 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001110");
        state_var_NS <= COMP_LOOP_C_283;
      WHEN COMP_LOOP_C_283 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001111");
        state_var_NS <= COMP_LOOP_C_284;
      WHEN COMP_LOOP_C_284 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010000");
        state_var_NS <= COMP_LOOP_C_285;
      WHEN COMP_LOOP_C_285 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010001");
        state_var_NS <= COMP_LOOP_C_286;
      WHEN COMP_LOOP_C_286 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010010");
        state_var_NS <= COMP_LOOP_C_287;
      WHEN COMP_LOOP_C_287 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010011");
        state_var_NS <= COMP_LOOP_C_288;
      WHEN COMP_LOOP_C_288 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010100");
        state_var_NS <= COMP_LOOP_C_289;
      WHEN COMP_LOOP_C_289 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010101");
        state_var_NS <= COMP_LOOP_C_290;
      WHEN COMP_LOOP_C_290 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010110");
        state_var_NS <= COMP_LOOP_C_291;
      WHEN COMP_LOOP_C_291 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010111");
        state_var_NS <= COMP_LOOP_C_292;
      WHEN COMP_LOOP_C_292 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011000");
        state_var_NS <= COMP_LOOP_C_293;
      WHEN COMP_LOOP_C_293 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011001");
        state_var_NS <= COMP_LOOP_C_294;
      WHEN COMP_LOOP_C_294 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011010");
        state_var_NS <= COMP_LOOP_C_295;
      WHEN COMP_LOOP_C_295 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011011");
        state_var_NS <= COMP_LOOP_C_296;
      WHEN COMP_LOOP_C_296 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011100");
        state_var_NS <= COMP_LOOP_C_297;
      WHEN COMP_LOOP_C_297 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011101");
        state_var_NS <= COMP_LOOP_C_298;
      WHEN COMP_LOOP_C_298 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011110");
        state_var_NS <= COMP_LOOP_C_299;
      WHEN COMP_LOOP_C_299 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011111");
        state_var_NS <= COMP_LOOP_C_300;
      WHEN COMP_LOOP_C_300 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100000");
        state_var_NS <= COMP_LOOP_C_301;
      WHEN COMP_LOOP_C_301 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100001");
        state_var_NS <= COMP_LOOP_C_302;
      WHEN COMP_LOOP_C_302 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100010");
        state_var_NS <= COMP_LOOP_C_303;
      WHEN COMP_LOOP_C_303 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100011");
        state_var_NS <= COMP_LOOP_C_304;
      WHEN COMP_LOOP_C_304 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100100");
        state_var_NS <= COMP_LOOP_C_305;
      WHEN COMP_LOOP_C_305 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100101");
        state_var_NS <= COMP_LOOP_C_306;
      WHEN COMP_LOOP_C_306 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100110");
        state_var_NS <= COMP_LOOP_C_307;
      WHEN COMP_LOOP_C_307 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100111");
        state_var_NS <= COMP_LOOP_C_308;
      WHEN COMP_LOOP_C_308 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101000");
        state_var_NS <= COMP_LOOP_C_309;
      WHEN COMP_LOOP_C_309 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101001");
        state_var_NS <= COMP_LOOP_C_310;
      WHEN COMP_LOOP_C_310 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101010");
        IF ( COMP_LOOP_C_310_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_311;
        END IF;
      WHEN COMP_LOOP_C_311 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101011");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_0;
      WHEN COMP_LOOP_6_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101100");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_1;
      WHEN COMP_LOOP_6_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101101");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_2;
      WHEN COMP_LOOP_6_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101110");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_3;
      WHEN COMP_LOOP_6_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101111");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_4;
      WHEN COMP_LOOP_6_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110000");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_5;
      WHEN COMP_LOOP_6_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110001");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_6;
      WHEN COMP_LOOP_6_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110010");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_7;
      WHEN COMP_LOOP_6_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110011");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_8;
      WHEN COMP_LOOP_6_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110100");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_9;
      WHEN COMP_LOOP_6_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110101");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_10;
      WHEN COMP_LOOP_6_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110110");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_11;
      WHEN COMP_LOOP_6_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110111");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_12;
      WHEN COMP_LOOP_6_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111000");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_13;
      WHEN COMP_LOOP_6_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111001");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_14;
      WHEN COMP_LOOP_6_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111010");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_15;
      WHEN COMP_LOOP_6_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111011");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_16;
      WHEN COMP_LOOP_6_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111100");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_17;
      WHEN COMP_LOOP_6_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111101");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_18;
      WHEN COMP_LOOP_6_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111110");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_19;
      WHEN COMP_LOOP_6_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111111");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_20;
      WHEN COMP_LOOP_6_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000000");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_21;
      WHEN COMP_LOOP_6_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000001");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_22;
      WHEN COMP_LOOP_6_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000010");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_23;
      WHEN COMP_LOOP_6_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000011");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_24;
      WHEN COMP_LOOP_6_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000100");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_25;
      WHEN COMP_LOOP_6_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000101");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_26;
      WHEN COMP_LOOP_6_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000110");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_27;
      WHEN COMP_LOOP_6_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000111");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_28;
      WHEN COMP_LOOP_6_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001000");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_29;
      WHEN COMP_LOOP_6_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001001");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_30;
      WHEN COMP_LOOP_6_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001010");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_31;
      WHEN COMP_LOOP_6_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001011");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_32;
      WHEN COMP_LOOP_6_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001100");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_33;
      WHEN COMP_LOOP_6_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001101");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_34;
      WHEN COMP_LOOP_6_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001110");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_35;
      WHEN COMP_LOOP_6_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001111");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_36;
      WHEN COMP_LOOP_6_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010000");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_37;
      WHEN COMP_LOOP_6_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010001");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_38;
      WHEN COMP_LOOP_6_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010010");
        IF ( COMP_LOOP_6_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_312;
        ELSE
          state_var_NS <= COMP_LOOP_6_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_312 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010011");
        state_var_NS <= COMP_LOOP_C_313;
      WHEN COMP_LOOP_C_313 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010100");
        state_var_NS <= COMP_LOOP_C_314;
      WHEN COMP_LOOP_C_314 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010101");
        state_var_NS <= COMP_LOOP_C_315;
      WHEN COMP_LOOP_C_315 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010110");
        state_var_NS <= COMP_LOOP_C_316;
      WHEN COMP_LOOP_C_316 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010111");
        state_var_NS <= COMP_LOOP_C_317;
      WHEN COMP_LOOP_C_317 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011000");
        state_var_NS <= COMP_LOOP_C_318;
      WHEN COMP_LOOP_C_318 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011001");
        state_var_NS <= COMP_LOOP_C_319;
      WHEN COMP_LOOP_C_319 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011010");
        state_var_NS <= COMP_LOOP_C_320;
      WHEN COMP_LOOP_C_320 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011011");
        state_var_NS <= COMP_LOOP_C_321;
      WHEN COMP_LOOP_C_321 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011100");
        state_var_NS <= COMP_LOOP_C_322;
      WHEN COMP_LOOP_C_322 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011101");
        state_var_NS <= COMP_LOOP_C_323;
      WHEN COMP_LOOP_C_323 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011110");
        state_var_NS <= COMP_LOOP_C_324;
      WHEN COMP_LOOP_C_324 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011111");
        state_var_NS <= COMP_LOOP_C_325;
      WHEN COMP_LOOP_C_325 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100000");
        state_var_NS <= COMP_LOOP_C_326;
      WHEN COMP_LOOP_C_326 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100001");
        state_var_NS <= COMP_LOOP_C_327;
      WHEN COMP_LOOP_C_327 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100010");
        state_var_NS <= COMP_LOOP_C_328;
      WHEN COMP_LOOP_C_328 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100011");
        state_var_NS <= COMP_LOOP_C_329;
      WHEN COMP_LOOP_C_329 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100100");
        state_var_NS <= COMP_LOOP_C_330;
      WHEN COMP_LOOP_C_330 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100101");
        state_var_NS <= COMP_LOOP_C_331;
      WHEN COMP_LOOP_C_331 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100110");
        state_var_NS <= COMP_LOOP_C_332;
      WHEN COMP_LOOP_C_332 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100111");
        state_var_NS <= COMP_LOOP_C_333;
      WHEN COMP_LOOP_C_333 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101000");
        state_var_NS <= COMP_LOOP_C_334;
      WHEN COMP_LOOP_C_334 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101001");
        state_var_NS <= COMP_LOOP_C_335;
      WHEN COMP_LOOP_C_335 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101010");
        state_var_NS <= COMP_LOOP_C_336;
      WHEN COMP_LOOP_C_336 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101011");
        state_var_NS <= COMP_LOOP_C_337;
      WHEN COMP_LOOP_C_337 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101100");
        state_var_NS <= COMP_LOOP_C_338;
      WHEN COMP_LOOP_C_338 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101101");
        state_var_NS <= COMP_LOOP_C_339;
      WHEN COMP_LOOP_C_339 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101110");
        state_var_NS <= COMP_LOOP_C_340;
      WHEN COMP_LOOP_C_340 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101111");
        state_var_NS <= COMP_LOOP_C_341;
      WHEN COMP_LOOP_C_341 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110000");
        state_var_NS <= COMP_LOOP_C_342;
      WHEN COMP_LOOP_C_342 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110001");
        state_var_NS <= COMP_LOOP_C_343;
      WHEN COMP_LOOP_C_343 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110010");
        state_var_NS <= COMP_LOOP_C_344;
      WHEN COMP_LOOP_C_344 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110011");
        state_var_NS <= COMP_LOOP_C_345;
      WHEN COMP_LOOP_C_345 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110100");
        state_var_NS <= COMP_LOOP_C_346;
      WHEN COMP_LOOP_C_346 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110101");
        state_var_NS <= COMP_LOOP_C_347;
      WHEN COMP_LOOP_C_347 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110110");
        state_var_NS <= COMP_LOOP_C_348;
      WHEN COMP_LOOP_C_348 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110111");
        state_var_NS <= COMP_LOOP_C_349;
      WHEN COMP_LOOP_C_349 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111000");
        state_var_NS <= COMP_LOOP_C_350;
      WHEN COMP_LOOP_C_350 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111001");
        state_var_NS <= COMP_LOOP_C_351;
      WHEN COMP_LOOP_C_351 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111010");
        state_var_NS <= COMP_LOOP_C_352;
      WHEN COMP_LOOP_C_352 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111011");
        state_var_NS <= COMP_LOOP_C_353;
      WHEN COMP_LOOP_C_353 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111100");
        state_var_NS <= COMP_LOOP_C_354;
      WHEN COMP_LOOP_C_354 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111101");
        state_var_NS <= COMP_LOOP_C_355;
      WHEN COMP_LOOP_C_355 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111110");
        state_var_NS <= COMP_LOOP_C_356;
      WHEN COMP_LOOP_C_356 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111111");
        state_var_NS <= COMP_LOOP_C_357;
      WHEN COMP_LOOP_C_357 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000000");
        state_var_NS <= COMP_LOOP_C_358;
      WHEN COMP_LOOP_C_358 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000001");
        state_var_NS <= COMP_LOOP_C_359;
      WHEN COMP_LOOP_C_359 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000010");
        state_var_NS <= COMP_LOOP_C_360;
      WHEN COMP_LOOP_C_360 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000011");
        state_var_NS <= COMP_LOOP_C_361;
      WHEN COMP_LOOP_C_361 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000100");
        state_var_NS <= COMP_LOOP_C_362;
      WHEN COMP_LOOP_C_362 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000101");
        state_var_NS <= COMP_LOOP_C_363;
      WHEN COMP_LOOP_C_363 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000110");
        state_var_NS <= COMP_LOOP_C_364;
      WHEN COMP_LOOP_C_364 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000111");
        state_var_NS <= COMP_LOOP_C_365;
      WHEN COMP_LOOP_C_365 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001000");
        state_var_NS <= COMP_LOOP_C_366;
      WHEN COMP_LOOP_C_366 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001001");
        state_var_NS <= COMP_LOOP_C_367;
      WHEN COMP_LOOP_C_367 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001010");
        state_var_NS <= COMP_LOOP_C_368;
      WHEN COMP_LOOP_C_368 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001011");
        state_var_NS <= COMP_LOOP_C_369;
      WHEN COMP_LOOP_C_369 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001100");
        state_var_NS <= COMP_LOOP_C_370;
      WHEN COMP_LOOP_C_370 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001101");
        state_var_NS <= COMP_LOOP_C_371;
      WHEN COMP_LOOP_C_371 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001110");
        state_var_NS <= COMP_LOOP_C_372;
      WHEN COMP_LOOP_C_372 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001111");
        IF ( COMP_LOOP_C_372_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_373;
        END IF;
      WHEN COMP_LOOP_C_373 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010000");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_0;
      WHEN COMP_LOOP_7_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010001");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_1;
      WHEN COMP_LOOP_7_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010010");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_2;
      WHEN COMP_LOOP_7_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010011");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_3;
      WHEN COMP_LOOP_7_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010100");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_4;
      WHEN COMP_LOOP_7_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010101");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_5;
      WHEN COMP_LOOP_7_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010110");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_6;
      WHEN COMP_LOOP_7_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010111");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_7;
      WHEN COMP_LOOP_7_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011000");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_8;
      WHEN COMP_LOOP_7_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011001");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_9;
      WHEN COMP_LOOP_7_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011010");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_10;
      WHEN COMP_LOOP_7_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011011");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_11;
      WHEN COMP_LOOP_7_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011100");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_12;
      WHEN COMP_LOOP_7_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011101");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_13;
      WHEN COMP_LOOP_7_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011110");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_14;
      WHEN COMP_LOOP_7_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011111");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_15;
      WHEN COMP_LOOP_7_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100000");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_16;
      WHEN COMP_LOOP_7_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100001");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_17;
      WHEN COMP_LOOP_7_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100010");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_18;
      WHEN COMP_LOOP_7_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100011");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_19;
      WHEN COMP_LOOP_7_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100100");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_20;
      WHEN COMP_LOOP_7_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100101");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_21;
      WHEN COMP_LOOP_7_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100110");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_22;
      WHEN COMP_LOOP_7_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100111");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_23;
      WHEN COMP_LOOP_7_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101000");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_24;
      WHEN COMP_LOOP_7_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101001");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_25;
      WHEN COMP_LOOP_7_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101010");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_26;
      WHEN COMP_LOOP_7_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101011");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_27;
      WHEN COMP_LOOP_7_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101100");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_28;
      WHEN COMP_LOOP_7_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101101");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_29;
      WHEN COMP_LOOP_7_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101110");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_30;
      WHEN COMP_LOOP_7_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101111");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_31;
      WHEN COMP_LOOP_7_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110000");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_32;
      WHEN COMP_LOOP_7_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110001");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_33;
      WHEN COMP_LOOP_7_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110010");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_34;
      WHEN COMP_LOOP_7_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110011");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_35;
      WHEN COMP_LOOP_7_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110100");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_36;
      WHEN COMP_LOOP_7_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110101");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_37;
      WHEN COMP_LOOP_7_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110110");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_38;
      WHEN COMP_LOOP_7_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110111");
        IF ( COMP_LOOP_7_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_374;
        ELSE
          state_var_NS <= COMP_LOOP_7_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_374 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111000");
        state_var_NS <= COMP_LOOP_C_375;
      WHEN COMP_LOOP_C_375 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111001");
        state_var_NS <= COMP_LOOP_C_376;
      WHEN COMP_LOOP_C_376 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111010");
        state_var_NS <= COMP_LOOP_C_377;
      WHEN COMP_LOOP_C_377 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111011");
        state_var_NS <= COMP_LOOP_C_378;
      WHEN COMP_LOOP_C_378 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111100");
        state_var_NS <= COMP_LOOP_C_379;
      WHEN COMP_LOOP_C_379 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111101");
        state_var_NS <= COMP_LOOP_C_380;
      WHEN COMP_LOOP_C_380 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111110");
        state_var_NS <= COMP_LOOP_C_381;
      WHEN COMP_LOOP_C_381 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111111");
        state_var_NS <= COMP_LOOP_C_382;
      WHEN COMP_LOOP_C_382 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000000");
        state_var_NS <= COMP_LOOP_C_383;
      WHEN COMP_LOOP_C_383 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000001");
        state_var_NS <= COMP_LOOP_C_384;
      WHEN COMP_LOOP_C_384 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000010");
        state_var_NS <= COMP_LOOP_C_385;
      WHEN COMP_LOOP_C_385 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000011");
        state_var_NS <= COMP_LOOP_C_386;
      WHEN COMP_LOOP_C_386 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000100");
        state_var_NS <= COMP_LOOP_C_387;
      WHEN COMP_LOOP_C_387 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000101");
        state_var_NS <= COMP_LOOP_C_388;
      WHEN COMP_LOOP_C_388 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000110");
        state_var_NS <= COMP_LOOP_C_389;
      WHEN COMP_LOOP_C_389 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000111");
        state_var_NS <= COMP_LOOP_C_390;
      WHEN COMP_LOOP_C_390 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001000");
        state_var_NS <= COMP_LOOP_C_391;
      WHEN COMP_LOOP_C_391 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001001");
        state_var_NS <= COMP_LOOP_C_392;
      WHEN COMP_LOOP_C_392 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001010");
        state_var_NS <= COMP_LOOP_C_393;
      WHEN COMP_LOOP_C_393 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001011");
        state_var_NS <= COMP_LOOP_C_394;
      WHEN COMP_LOOP_C_394 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001100");
        state_var_NS <= COMP_LOOP_C_395;
      WHEN COMP_LOOP_C_395 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001101");
        state_var_NS <= COMP_LOOP_C_396;
      WHEN COMP_LOOP_C_396 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001110");
        state_var_NS <= COMP_LOOP_C_397;
      WHEN COMP_LOOP_C_397 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001111");
        state_var_NS <= COMP_LOOP_C_398;
      WHEN COMP_LOOP_C_398 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010000");
        state_var_NS <= COMP_LOOP_C_399;
      WHEN COMP_LOOP_C_399 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010001");
        state_var_NS <= COMP_LOOP_C_400;
      WHEN COMP_LOOP_C_400 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010010");
        state_var_NS <= COMP_LOOP_C_401;
      WHEN COMP_LOOP_C_401 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010011");
        state_var_NS <= COMP_LOOP_C_402;
      WHEN COMP_LOOP_C_402 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010100");
        state_var_NS <= COMP_LOOP_C_403;
      WHEN COMP_LOOP_C_403 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010101");
        state_var_NS <= COMP_LOOP_C_404;
      WHEN COMP_LOOP_C_404 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010110");
        state_var_NS <= COMP_LOOP_C_405;
      WHEN COMP_LOOP_C_405 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010111");
        state_var_NS <= COMP_LOOP_C_406;
      WHEN COMP_LOOP_C_406 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011000");
        state_var_NS <= COMP_LOOP_C_407;
      WHEN COMP_LOOP_C_407 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011001");
        state_var_NS <= COMP_LOOP_C_408;
      WHEN COMP_LOOP_C_408 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011010");
        state_var_NS <= COMP_LOOP_C_409;
      WHEN COMP_LOOP_C_409 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011011");
        state_var_NS <= COMP_LOOP_C_410;
      WHEN COMP_LOOP_C_410 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011100");
        state_var_NS <= COMP_LOOP_C_411;
      WHEN COMP_LOOP_C_411 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011101");
        state_var_NS <= COMP_LOOP_C_412;
      WHEN COMP_LOOP_C_412 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011110");
        state_var_NS <= COMP_LOOP_C_413;
      WHEN COMP_LOOP_C_413 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011111");
        state_var_NS <= COMP_LOOP_C_414;
      WHEN COMP_LOOP_C_414 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100000");
        state_var_NS <= COMP_LOOP_C_415;
      WHEN COMP_LOOP_C_415 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100001");
        state_var_NS <= COMP_LOOP_C_416;
      WHEN COMP_LOOP_C_416 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100010");
        state_var_NS <= COMP_LOOP_C_417;
      WHEN COMP_LOOP_C_417 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100011");
        state_var_NS <= COMP_LOOP_C_418;
      WHEN COMP_LOOP_C_418 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100100");
        state_var_NS <= COMP_LOOP_C_419;
      WHEN COMP_LOOP_C_419 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100101");
        state_var_NS <= COMP_LOOP_C_420;
      WHEN COMP_LOOP_C_420 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100110");
        state_var_NS <= COMP_LOOP_C_421;
      WHEN COMP_LOOP_C_421 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100111");
        state_var_NS <= COMP_LOOP_C_422;
      WHEN COMP_LOOP_C_422 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101000");
        state_var_NS <= COMP_LOOP_C_423;
      WHEN COMP_LOOP_C_423 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101001");
        state_var_NS <= COMP_LOOP_C_424;
      WHEN COMP_LOOP_C_424 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101010");
        state_var_NS <= COMP_LOOP_C_425;
      WHEN COMP_LOOP_C_425 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101011");
        state_var_NS <= COMP_LOOP_C_426;
      WHEN COMP_LOOP_C_426 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101100");
        state_var_NS <= COMP_LOOP_C_427;
      WHEN COMP_LOOP_C_427 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101101");
        state_var_NS <= COMP_LOOP_C_428;
      WHEN COMP_LOOP_C_428 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101110");
        state_var_NS <= COMP_LOOP_C_429;
      WHEN COMP_LOOP_C_429 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101111");
        state_var_NS <= COMP_LOOP_C_430;
      WHEN COMP_LOOP_C_430 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110000");
        state_var_NS <= COMP_LOOP_C_431;
      WHEN COMP_LOOP_C_431 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110001");
        state_var_NS <= COMP_LOOP_C_432;
      WHEN COMP_LOOP_C_432 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110010");
        state_var_NS <= COMP_LOOP_C_433;
      WHEN COMP_LOOP_C_433 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110011");
        state_var_NS <= COMP_LOOP_C_434;
      WHEN COMP_LOOP_C_434 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110100");
        IF ( COMP_LOOP_C_434_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_435;
        END IF;
      WHEN COMP_LOOP_C_435 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110101");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_0;
      WHEN COMP_LOOP_8_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110110");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_1;
      WHEN COMP_LOOP_8_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110111");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_2;
      WHEN COMP_LOOP_8_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111000");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_3;
      WHEN COMP_LOOP_8_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111001");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_4;
      WHEN COMP_LOOP_8_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111010");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_5;
      WHEN COMP_LOOP_8_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111011");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_6;
      WHEN COMP_LOOP_8_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111100");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_7;
      WHEN COMP_LOOP_8_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111101");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_8;
      WHEN COMP_LOOP_8_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111110");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_9;
      WHEN COMP_LOOP_8_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111111");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_10;
      WHEN COMP_LOOP_8_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000000");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_11;
      WHEN COMP_LOOP_8_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000001");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_12;
      WHEN COMP_LOOP_8_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000010");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_13;
      WHEN COMP_LOOP_8_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000011");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_14;
      WHEN COMP_LOOP_8_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000100");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_15;
      WHEN COMP_LOOP_8_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000101");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_16;
      WHEN COMP_LOOP_8_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000110");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_17;
      WHEN COMP_LOOP_8_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000111");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_18;
      WHEN COMP_LOOP_8_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100001000");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_19;
      WHEN COMP_LOOP_8_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100001001");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_20;
      WHEN COMP_LOOP_8_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100001010");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_21;
      WHEN COMP_LOOP_8_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100001011");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_22;
      WHEN COMP_LOOP_8_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100001100");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_23;
      WHEN COMP_LOOP_8_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100001101");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_24;
      WHEN COMP_LOOP_8_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100001110");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_25;
      WHEN COMP_LOOP_8_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100001111");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_26;
      WHEN COMP_LOOP_8_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100010000");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_27;
      WHEN COMP_LOOP_8_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100010001");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_28;
      WHEN COMP_LOOP_8_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100010010");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_29;
      WHEN COMP_LOOP_8_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100010011");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_30;
      WHEN COMP_LOOP_8_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100010100");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_31;
      WHEN COMP_LOOP_8_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100010101");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_32;
      WHEN COMP_LOOP_8_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100010110");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_33;
      WHEN COMP_LOOP_8_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100010111");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_34;
      WHEN COMP_LOOP_8_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100011000");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_35;
      WHEN COMP_LOOP_8_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100011001");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_36;
      WHEN COMP_LOOP_8_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100011010");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_37;
      WHEN COMP_LOOP_8_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100011011");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_38;
      WHEN COMP_LOOP_8_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100011100");
        IF ( COMP_LOOP_8_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_436;
        ELSE
          state_var_NS <= COMP_LOOP_8_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_436 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100011101");
        state_var_NS <= COMP_LOOP_C_437;
      WHEN COMP_LOOP_C_437 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100011110");
        state_var_NS <= COMP_LOOP_C_438;
      WHEN COMP_LOOP_C_438 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100011111");
        state_var_NS <= COMP_LOOP_C_439;
      WHEN COMP_LOOP_C_439 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100100000");
        state_var_NS <= COMP_LOOP_C_440;
      WHEN COMP_LOOP_C_440 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100100001");
        state_var_NS <= COMP_LOOP_C_441;
      WHEN COMP_LOOP_C_441 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100100010");
        state_var_NS <= COMP_LOOP_C_442;
      WHEN COMP_LOOP_C_442 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100100011");
        state_var_NS <= COMP_LOOP_C_443;
      WHEN COMP_LOOP_C_443 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100100100");
        state_var_NS <= COMP_LOOP_C_444;
      WHEN COMP_LOOP_C_444 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100100101");
        state_var_NS <= COMP_LOOP_C_445;
      WHEN COMP_LOOP_C_445 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100100110");
        state_var_NS <= COMP_LOOP_C_446;
      WHEN COMP_LOOP_C_446 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100100111");
        state_var_NS <= COMP_LOOP_C_447;
      WHEN COMP_LOOP_C_447 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100101000");
        state_var_NS <= COMP_LOOP_C_448;
      WHEN COMP_LOOP_C_448 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100101001");
        state_var_NS <= COMP_LOOP_C_449;
      WHEN COMP_LOOP_C_449 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100101010");
        state_var_NS <= COMP_LOOP_C_450;
      WHEN COMP_LOOP_C_450 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100101011");
        state_var_NS <= COMP_LOOP_C_451;
      WHEN COMP_LOOP_C_451 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100101100");
        state_var_NS <= COMP_LOOP_C_452;
      WHEN COMP_LOOP_C_452 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100101101");
        state_var_NS <= COMP_LOOP_C_453;
      WHEN COMP_LOOP_C_453 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100101110");
        state_var_NS <= COMP_LOOP_C_454;
      WHEN COMP_LOOP_C_454 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100101111");
        state_var_NS <= COMP_LOOP_C_455;
      WHEN COMP_LOOP_C_455 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100110000");
        state_var_NS <= COMP_LOOP_C_456;
      WHEN COMP_LOOP_C_456 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100110001");
        state_var_NS <= COMP_LOOP_C_457;
      WHEN COMP_LOOP_C_457 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100110010");
        state_var_NS <= COMP_LOOP_C_458;
      WHEN COMP_LOOP_C_458 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100110011");
        state_var_NS <= COMP_LOOP_C_459;
      WHEN COMP_LOOP_C_459 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100110100");
        state_var_NS <= COMP_LOOP_C_460;
      WHEN COMP_LOOP_C_460 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100110101");
        state_var_NS <= COMP_LOOP_C_461;
      WHEN COMP_LOOP_C_461 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100110110");
        state_var_NS <= COMP_LOOP_C_462;
      WHEN COMP_LOOP_C_462 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100110111");
        state_var_NS <= COMP_LOOP_C_463;
      WHEN COMP_LOOP_C_463 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100111000");
        state_var_NS <= COMP_LOOP_C_464;
      WHEN COMP_LOOP_C_464 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100111001");
        state_var_NS <= COMP_LOOP_C_465;
      WHEN COMP_LOOP_C_465 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100111010");
        state_var_NS <= COMP_LOOP_C_466;
      WHEN COMP_LOOP_C_466 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100111011");
        state_var_NS <= COMP_LOOP_C_467;
      WHEN COMP_LOOP_C_467 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100111100");
        state_var_NS <= COMP_LOOP_C_468;
      WHEN COMP_LOOP_C_468 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100111101");
        state_var_NS <= COMP_LOOP_C_469;
      WHEN COMP_LOOP_C_469 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100111110");
        state_var_NS <= COMP_LOOP_C_470;
      WHEN COMP_LOOP_C_470 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100111111");
        state_var_NS <= COMP_LOOP_C_471;
      WHEN COMP_LOOP_C_471 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101000000");
        state_var_NS <= COMP_LOOP_C_472;
      WHEN COMP_LOOP_C_472 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101000001");
        state_var_NS <= COMP_LOOP_C_473;
      WHEN COMP_LOOP_C_473 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101000010");
        state_var_NS <= COMP_LOOP_C_474;
      WHEN COMP_LOOP_C_474 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101000011");
        state_var_NS <= COMP_LOOP_C_475;
      WHEN COMP_LOOP_C_475 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101000100");
        state_var_NS <= COMP_LOOP_C_476;
      WHEN COMP_LOOP_C_476 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101000101");
        state_var_NS <= COMP_LOOP_C_477;
      WHEN COMP_LOOP_C_477 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101000110");
        state_var_NS <= COMP_LOOP_C_478;
      WHEN COMP_LOOP_C_478 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101000111");
        state_var_NS <= COMP_LOOP_C_479;
      WHEN COMP_LOOP_C_479 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101001000");
        state_var_NS <= COMP_LOOP_C_480;
      WHEN COMP_LOOP_C_480 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101001001");
        state_var_NS <= COMP_LOOP_C_481;
      WHEN COMP_LOOP_C_481 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101001010");
        state_var_NS <= COMP_LOOP_C_482;
      WHEN COMP_LOOP_C_482 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101001011");
        state_var_NS <= COMP_LOOP_C_483;
      WHEN COMP_LOOP_C_483 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101001100");
        state_var_NS <= COMP_LOOP_C_484;
      WHEN COMP_LOOP_C_484 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101001101");
        state_var_NS <= COMP_LOOP_C_485;
      WHEN COMP_LOOP_C_485 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101001110");
        state_var_NS <= COMP_LOOP_C_486;
      WHEN COMP_LOOP_C_486 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101001111");
        state_var_NS <= COMP_LOOP_C_487;
      WHEN COMP_LOOP_C_487 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101010000");
        state_var_NS <= COMP_LOOP_C_488;
      WHEN COMP_LOOP_C_488 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101010001");
        state_var_NS <= COMP_LOOP_C_489;
      WHEN COMP_LOOP_C_489 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101010010");
        state_var_NS <= COMP_LOOP_C_490;
      WHEN COMP_LOOP_C_490 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101010011");
        state_var_NS <= COMP_LOOP_C_491;
      WHEN COMP_LOOP_C_491 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101010100");
        state_var_NS <= COMP_LOOP_C_492;
      WHEN COMP_LOOP_C_492 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101010101");
        state_var_NS <= COMP_LOOP_C_493;
      WHEN COMP_LOOP_C_493 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101010110");
        state_var_NS <= COMP_LOOP_C_494;
      WHEN COMP_LOOP_C_494 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101010111");
        state_var_NS <= COMP_LOOP_C_495;
      WHEN COMP_LOOP_C_495 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101011000");
        state_var_NS <= COMP_LOOP_C_496;
      WHEN COMP_LOOP_C_496 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101011001");
        IF ( COMP_LOOP_C_496_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN VEC_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101011010");
        IF ( VEC_LOOP_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP_C_9;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN STAGE_LOOP_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101011011");
        IF ( STAGE_LOOP_C_9_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSE
          state_var_NS <= STAGE_LOOP_C_0;
        END IF;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101011100");
        state_var_NS <= main_C_0;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000");
        state_var_NS <= STAGE_LOOP_C_0;
    END CASE;
  END PROCESS inPlaceNTT_DIT_core_core_fsm_1;

  inPlaceNTT_DIT_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        state_var <= state_var_NS;
      END IF;
    END IF;
  END PROCESS inPlaceNTT_DIT_core_core_fsm_1_REG;

END v40;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC;
    vec_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_0_i_adra_d_pff : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    vec_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_1_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_2_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_3_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_4_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_5_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_6_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_7_i_wea_d_pff : OUT STD_LOGIC
  );
END inPlaceNTT_DIT_core;

ARCHITECTURE v40 OF inPlaceNTT_DIT_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL p_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL r_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_result_rem_cmp_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_result_rem_cmp_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_result_rem_cmp_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_b_9_0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL fsm_output : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL nor_tmp : STD_LOGIC;
  SIGNAL or_tmp : STD_LOGIC;
  SIGNAL or_tmp_92 : STD_LOGIC;
  SIGNAL nor_tmp_23 : STD_LOGIC;
  SIGNAL or_tmp_103 : STD_LOGIC;
  SIGNAL nor_tmp_27 : STD_LOGIC;
  SIGNAL mux_tmp_156 : STD_LOGIC;
  SIGNAL or_tmp_113 : STD_LOGIC;
  SIGNAL and_dcpl_4 : STD_LOGIC;
  SIGNAL or_tmp_154 : STD_LOGIC;
  SIGNAL and_dcpl_11 : STD_LOGIC;
  SIGNAL and_dcpl_14 : STD_LOGIC;
  SIGNAL and_dcpl_23 : STD_LOGIC;
  SIGNAL not_tmp_131 : STD_LOGIC;
  SIGNAL and_dcpl_46 : STD_LOGIC;
  SIGNAL and_dcpl_47 : STD_LOGIC;
  SIGNAL and_dcpl_48 : STD_LOGIC;
  SIGNAL and_dcpl_50 : STD_LOGIC;
  SIGNAL and_dcpl_51 : STD_LOGIC;
  SIGNAL and_dcpl_56 : STD_LOGIC;
  SIGNAL and_dcpl_57 : STD_LOGIC;
  SIGNAL and_dcpl_58 : STD_LOGIC;
  SIGNAL and_dcpl_59 : STD_LOGIC;
  SIGNAL and_dcpl_60 : STD_LOGIC;
  SIGNAL and_dcpl_63 : STD_LOGIC;
  SIGNAL and_dcpl_64 : STD_LOGIC;
  SIGNAL and_dcpl_65 : STD_LOGIC;
  SIGNAL and_dcpl_66 : STD_LOGIC;
  SIGNAL and_dcpl_67 : STD_LOGIC;
  SIGNAL and_dcpl_68 : STD_LOGIC;
  SIGNAL and_dcpl_69 : STD_LOGIC;
  SIGNAL and_dcpl_70 : STD_LOGIC;
  SIGNAL and_dcpl_73 : STD_LOGIC;
  SIGNAL and_dcpl_80 : STD_LOGIC;
  SIGNAL and_dcpl_82 : STD_LOGIC;
  SIGNAL and_dcpl_84 : STD_LOGIC;
  SIGNAL and_dcpl_89 : STD_LOGIC;
  SIGNAL and_dcpl_91 : STD_LOGIC;
  SIGNAL and_dcpl_93 : STD_LOGIC;
  SIGNAL and_dcpl_100 : STD_LOGIC;
  SIGNAL and_dcpl_102 : STD_LOGIC;
  SIGNAL and_dcpl_103 : STD_LOGIC;
  SIGNAL and_dcpl_108 : STD_LOGIC;
  SIGNAL and_dcpl_109 : STD_LOGIC;
  SIGNAL and_dcpl_110 : STD_LOGIC;
  SIGNAL and_dcpl_112 : STD_LOGIC;
  SIGNAL and_dcpl_121 : STD_LOGIC;
  SIGNAL and_dcpl_122 : STD_LOGIC;
  SIGNAL and_dcpl_123 : STD_LOGIC;
  SIGNAL and_dcpl_127 : STD_LOGIC;
  SIGNAL and_dcpl_128 : STD_LOGIC;
  SIGNAL and_dcpl_129 : STD_LOGIC;
  SIGNAL and_dcpl_130 : STD_LOGIC;
  SIGNAL and_dcpl_137 : STD_LOGIC;
  SIGNAL and_dcpl_138 : STD_LOGIC;
  SIGNAL or_tmp_268 : STD_LOGIC;
  SIGNAL or_tmp_273 : STD_LOGIC;
  SIGNAL not_tmp_165 : STD_LOGIC;
  SIGNAL or_tmp_335 : STD_LOGIC;
  SIGNAL or_tmp_340 : STD_LOGIC;
  SIGNAL or_tmp_395 : STD_LOGIC;
  SIGNAL nand_tmp_18 : STD_LOGIC;
  SIGNAL or_tmp_454 : STD_LOGIC;
  SIGNAL nand_tmp_21 : STD_LOGIC;
  SIGNAL or_tmp_525 : STD_LOGIC;
  SIGNAL or_tmp_535 : STD_LOGIC;
  SIGNAL or_tmp_590 : STD_LOGIC;
  SIGNAL or_tmp_600 : STD_LOGIC;
  SIGNAL or_tmp_655 : STD_LOGIC;
  SIGNAL nand_tmp_31 : STD_LOGIC;
  SIGNAL or_tmp_719 : STD_LOGIC;
  SIGNAL nand_tmp_35 : STD_LOGIC;
  SIGNAL and_dcpl_140 : STD_LOGIC;
  SIGNAL and_dcpl_147 : STD_LOGIC;
  SIGNAL mux_tmp_677 : STD_LOGIC;
  SIGNAL mux_tmp_688 : STD_LOGIC;
  SIGNAL mux_tmp_689 : STD_LOGIC;
  SIGNAL nor_tmp_146 : STD_LOGIC;
  SIGNAL mux_tmp_705 : STD_LOGIC;
  SIGNAL or_tmp_788 : STD_LOGIC;
  SIGNAL mux_tmp_718 : STD_LOGIC;
  SIGNAL mux_tmp_719 : STD_LOGIC;
  SIGNAL mux_tmp_722 : STD_LOGIC;
  SIGNAL or_tmp_792 : STD_LOGIC;
  SIGNAL nand_tmp_42 : STD_LOGIC;
  SIGNAL mux_tmp_731 : STD_LOGIC;
  SIGNAL not_tmp_274 : STD_LOGIC;
  SIGNAL not_tmp_280 : STD_LOGIC;
  SIGNAL or_tmp_810 : STD_LOGIC;
  SIGNAL mux_tmp_776 : STD_LOGIC;
  SIGNAL not_tmp_297 : STD_LOGIC;
  SIGNAL not_tmp_309 : STD_LOGIC;
  SIGNAL not_tmp_312 : STD_LOGIC;
  SIGNAL not_tmp_315 : STD_LOGIC;
  SIGNAL and_dcpl_152 : STD_LOGIC;
  SIGNAL and_dcpl_156 : STD_LOGIC;
  SIGNAL or_tmp_891 : STD_LOGIC;
  SIGNAL mux_tmp_845 : STD_LOGIC;
  SIGNAL not_tmp_347 : STD_LOGIC;
  SIGNAL and_dcpl_162 : STD_LOGIC;
  SIGNAL or_tmp_916 : STD_LOGIC;
  SIGNAL mux_tmp_886 : STD_LOGIC;
  SIGNAL or_tmp_918 : STD_LOGIC;
  SIGNAL and_tmp_28 : STD_LOGIC;
  SIGNAL and_dcpl_164 : STD_LOGIC;
  SIGNAL and_dcpl_167 : STD_LOGIC;
  SIGNAL and_dcpl_168 : STD_LOGIC;
  SIGNAL and_dcpl_171 : STD_LOGIC;
  SIGNAL and_dcpl_172 : STD_LOGIC;
  SIGNAL and_dcpl_176 : STD_LOGIC;
  SIGNAL and_dcpl_180 : STD_LOGIC;
  SIGNAL and_dcpl_184 : STD_LOGIC;
  SIGNAL and_dcpl_187 : STD_LOGIC;
  SIGNAL not_tmp_374 : STD_LOGIC;
  SIGNAL not_tmp_399 : STD_LOGIC;
  SIGNAL not_tmp_400 : STD_LOGIC;
  SIGNAL not_tmp_406 : STD_LOGIC;
  SIGNAL not_tmp_414 : STD_LOGIC;
  SIGNAL mux_tmp_997 : STD_LOGIC;
  SIGNAL mux_tmp_1006 : STD_LOGIC;
  SIGNAL not_tmp_436 : STD_LOGIC;
  SIGNAL not_tmp_462 : STD_LOGIC;
  SIGNAL and_dcpl_219 : STD_LOGIC;
  SIGNAL not_tmp_480 : STD_LOGIC;
  SIGNAL nor_tmp_240 : STD_LOGIC;
  SIGNAL mux_tmp_1159 : STD_LOGIC;
  SIGNAL nor_tmp_241 : STD_LOGIC;
  SIGNAL mux_tmp_1160 : STD_LOGIC;
  SIGNAL and_tmp_44 : STD_LOGIC;
  SIGNAL mux_tmp_1162 : STD_LOGIC;
  SIGNAL not_tmp_482 : STD_LOGIC;
  SIGNAL nor_tmp_244 : STD_LOGIC;
  SIGNAL mux_tmp_1164 : STD_LOGIC;
  SIGNAL mux_tmp_1170 : STD_LOGIC;
  SIGNAL or_tmp_1144 : STD_LOGIC;
  SIGNAL and_tmp_45 : STD_LOGIC;
  SIGNAL and_tmp_46 : STD_LOGIC;
  SIGNAL mux_tmp_1178 : STD_LOGIC;
  SIGNAL or_tmp_1159 : STD_LOGIC;
  SIGNAL or_tmp_1165 : STD_LOGIC;
  SIGNAL mux_tmp_1202 : STD_LOGIC;
  SIGNAL or_tmp_1174 : STD_LOGIC;
  SIGNAL or_tmp_1176 : STD_LOGIC;
  SIGNAL and_dcpl_226 : STD_LOGIC;
  SIGNAL not_tmp_513 : STD_LOGIC;
  SIGNAL not_tmp_523 : STD_LOGIC;
  SIGNAL or_tmp_1261 : STD_LOGIC;
  SIGNAL mux_tmp_1305 : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_11_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_145_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_1_cse_6_sva_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL VEC_LOOP_j_sva_11_0 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_k_9_3_sva_5_0 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL COMP_LOOP_k_9_3_sva_2 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_12_1_1_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_6_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_2_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_4_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_11_psp_sva : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_13_psp_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_14_psp_sva : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL tmp_10_lpi_4_dfm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_4_sva_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_2_sva_mx0w0 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL and_244_m1c : STD_LOGIC;
  SIGNAL mux_984_m1c : STD_LOGIC;
  SIGNAL and_224_m1c : STD_LOGIC;
  SIGNAL and_226_m1c : STD_LOGIC;
  SIGNAL and_229_m1c : STD_LOGIC;
  SIGNAL and_230_m1c : STD_LOGIC;
  SIGNAL and_233_m1c : STD_LOGIC;
  SIGNAL and_235_m1c : STD_LOGIC;
  SIGNAL and_237_m1c : STD_LOGIC;
  SIGNAL and_187_m1c : STD_LOGIC;
  SIGNAL and_416_cse : STD_LOGIC;
  SIGNAL nand_190_cse : STD_LOGIC;
  SIGNAL nand_168_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_triosy_0_7_obj_ld_cse : STD_LOGIC;
  SIGNAL and_389_cse : STD_LOGIC;
  SIGNAL or_838_cse : STD_LOGIC;
  SIGNAL or_1099_cse : STD_LOGIC;
  SIGNAL or_1385_cse : STD_LOGIC;
  SIGNAL or_1391_cse : STD_LOGIC;
  SIGNAL and_477_cse : STD_LOGIC;
  SIGNAL nor_425_cse : STD_LOGIC;
  SIGNAL or_247_cse : STD_LOGIC;
  SIGNAL and_483_cse : STD_LOGIC;
  SIGNAL or_245_cse : STD_LOGIC;
  SIGNAL and_314_cse : STD_LOGIC;
  SIGNAL nor_393_cse : STD_LOGIC;
  SIGNAL nand_100_cse : STD_LOGIC;
  SIGNAL or_1189_cse : STD_LOGIC;
  SIGNAL and_316_cse : STD_LOGIC;
  SIGNAL modulo_result_mux_1_cse : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL nand_97_cse : STD_LOGIC;
  SIGNAL or_81_cse : STD_LOGIC;
  SIGNAL or_83_cse : STD_LOGIC;
  SIGNAL or_171_cse : STD_LOGIC;
  SIGNAL or_216_cse : STD_LOGIC;
  SIGNAL or_1202_cse : STD_LOGIC;
  SIGNAL and_369_cse : STD_LOGIC;
  SIGNAL and_437_cse : STD_LOGIC;
  SIGNAL or_329_cse : STD_LOGIC;
  SIGNAL or_327_cse : STD_LOGIC;
  SIGNAL mux_392_cse : STD_LOGIC;
  SIGNAL or_320_cse : STD_LOGIC;
  SIGNAL nand_246_cse : STD_LOGIC;
  SIGNAL or_314_cse : STD_LOGIC;
  SIGNAL or_312_cse : STD_LOGIC;
  SIGNAL nand_194_cse : STD_LOGIC;
  SIGNAL nand_189_cse : STD_LOGIC;
  SIGNAL and_428_cse : STD_LOGIC;
  SIGNAL or_817_cse : STD_LOGIC;
  SIGNAL or_242_cse : STD_LOGIC;
  SIGNAL nor_601_cse : STD_LOGIC;
  SIGNAL mux_29_cse : STD_LOGIC;
  SIGNAL nand_230_cse : STD_LOGIC;
  SIGNAL and_502_cse : STD_LOGIC;
  SIGNAL or_816_cse : STD_LOGIC;
  SIGNAL or_210_cse : STD_LOGIC;
  SIGNAL or_1392_cse : STD_LOGIC;
  SIGNAL nand_89_cse : STD_LOGIC;
  SIGNAL nor_357_cse : STD_LOGIC;
  SIGNAL and_361_cse : STD_LOGIC;
  SIGNAL and_462_cse : STD_LOGIC;
  SIGNAL and_382_cse : STD_LOGIC;
  SIGNAL or_1394_cse : STD_LOGIC;
  SIGNAL or_1423_cse : STD_LOGIC;
  SIGNAL mux_331_cse : STD_LOGIC;
  SIGNAL mux_342_cse : STD_LOGIC;
  SIGNAL and_491_cse : STD_LOGIC;
  SIGNAL or_115_cse : STD_LOGIC;
  SIGNAL and_25_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_psp_sva_1 : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL mux_696_itm : STD_LOGIC;
  SIGNAL mux_1158_itm : STD_LOGIC;
  SIGNAL mux_1273_itm : STD_LOGIC;
  SIGNAL and_dcpl : STD_LOGIC;
  SIGNAL and_dcpl_236 : STD_LOGIC;
  SIGNAL and_dcpl_238 : STD_LOGIC;
  SIGNAL and_dcpl_240 : STD_LOGIC;
  SIGNAL and_dcpl_242 : STD_LOGIC;
  SIGNAL and_dcpl_243 : STD_LOGIC;
  SIGNAL and_dcpl_245 : STD_LOGIC;
  SIGNAL and_dcpl_247 : STD_LOGIC;
  SIGNAL and_dcpl_255 : STD_LOGIC;
  SIGNAL and_dcpl_260 : STD_LOGIC;
  SIGNAL and_dcpl_266 : STD_LOGIC;
  SIGNAL z_out : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL and_dcpl_268 : STD_LOGIC;
  SIGNAL and_dcpl_269 : STD_LOGIC;
  SIGNAL and_dcpl_276 : STD_LOGIC;
  SIGNAL and_dcpl_298 : STD_LOGIC;
  SIGNAL z_out_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL and_dcpl_324 : STD_LOGIC;
  SIGNAL and_dcpl_340 : STD_LOGIC;
  SIGNAL and_dcpl_345 : STD_LOGIC;
  SIGNAL z_out_2 : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL and_dcpl_347 : STD_LOGIC;
  SIGNAL and_dcpl_349 : STD_LOGIC;
  SIGNAL and_dcpl_354 : STD_LOGIC;
  SIGNAL or_tmp_1317 : STD_LOGIC;
  SIGNAL not_tmp_581 : STD_LOGIC;
  SIGNAL and_dcpl_357 : STD_LOGIC;
  SIGNAL and_dcpl_362 : STD_LOGIC;
  SIGNAL and_dcpl_364 : STD_LOGIC;
  SIGNAL and_dcpl_367 : STD_LOGIC;
  SIGNAL and_dcpl_368 : STD_LOGIC;
  SIGNAL and_dcpl_372 : STD_LOGIC;
  SIGNAL and_dcpl_379 : STD_LOGIC;
  SIGNAL and_dcpl_383 : STD_LOGIC;
  SIGNAL and_dcpl_385 : STD_LOGIC;
  SIGNAL and_dcpl_388 : STD_LOGIC;
  SIGNAL and_dcpl_394 : STD_LOGIC;
  SIGNAL and_dcpl_399 : STD_LOGIC;
  SIGNAL and_dcpl_404 : STD_LOGIC;
  SIGNAL and_dcpl_406 : STD_LOGIC;
  SIGNAL and_dcpl_409 : STD_LOGIC;
  SIGNAL and_dcpl_411 : STD_LOGIC;
  SIGNAL z_out_3 : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL or_tmp_1346 : STD_LOGIC;
  SIGNAL or_tmp_1348 : STD_LOGIC;
  SIGNAL or_tmp_1349 : STD_LOGIC;
  SIGNAL not_tmp_600 : STD_LOGIC;
  SIGNAL z_out_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL p_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL r_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_LOOP_i_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_psp_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL modExp_result_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modExp_exp_1_7_1_sva : STD_LOGIC;
  SIGNAL modExp_exp_1_6_1_sva : STD_LOGIC;
  SIGNAL modExp_exp_1_5_1_sva : STD_LOGIC;
  SIGNAL modExp_exp_1_4_1_sva : STD_LOGIC;
  SIGNAL modExp_exp_1_3_1_sva : STD_LOGIC;
  SIGNAL modExp_exp_1_2_1_sva : STD_LOGIC;
  SIGNAL modExp_exp_1_1_1_sva : STD_LOGIC;
  SIGNAL modExp_exp_1_0_1_sva_1 : STD_LOGIC;
  SIGNAL COMP_LOOP_1_mul_mut : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_1_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_12_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_8_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_4_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_30_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_32_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_33_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_34_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_86_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_89_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_124_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_125_itm : STD_LOGIC;
  SIGNAL STAGE_LOOP_i_3_0_sva_mx0c1 : STD_LOGIC;
  SIGNAL STAGE_LOOP_i_3_0_sva_2 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL modulo_qr_sva_1_mx0w1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_acc_5_mut_mx0w5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_psp_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL VEC_LOOP_j_sva_11_0_mx0c1 : STD_LOGIC;
  SIGNAL modExp_result_sva_mx0c0 : STD_LOGIC;
  SIGNAL operator_64_false_slc_modExp_exp_63_1_3 : STD_LOGIC_VECTOR (62 DOWNTO 0);
  SIGNAL modExp_while_and_3 : STD_LOGIC;
  SIGNAL modExp_while_and_5 : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_211 : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_213 : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_215 : STD_LOGIC;
  SIGNAL and_243_m1c : STD_LOGIC;
  SIGNAL modExp_result_and_rgt : STD_LOGIC;
  SIGNAL modExp_result_and_1_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_11_cse : STD_LOGIC;
  SIGNAL modExp_while_or_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_12_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_37_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_13_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_2_cse : STD_LOGIC;
  SIGNAL nor_473_cse : STD_LOGIC;
  SIGNAL nor_461_cse : STD_LOGIC;
  SIGNAL nor_447_cse : STD_LOGIC;
  SIGNAL and_494_cse : STD_LOGIC;
  SIGNAL operator_64_false_1_or_4_ssc : STD_LOGIC;
  SIGNAL operator_64_false_1_or_5_ssc : STD_LOGIC;
  SIGNAL and_511_cse : STD_LOGIC;
  SIGNAL or_tmp_1365 : STD_LOGIC;
  SIGNAL mux_tmp : STD_LOGIC;
  SIGNAL or_tmp_1367 : STD_LOGIC;
  SIGNAL nor_tmp_292 : STD_LOGIC;
  SIGNAL mux_tmp_1374 : STD_LOGIC;
  SIGNAL mux_tmp_1377 : STD_LOGIC;
  SIGNAL mux_tmp_1378 : STD_LOGIC;
  SIGNAL or_tmp_1370 : STD_LOGIC;
  SIGNAL nor_tmp_296 : STD_LOGIC;
  SIGNAL or_tmp_1374 : STD_LOGIC;
  SIGNAL mux_tmp_1399 : STD_LOGIC;
  SIGNAL or_tmp_1389 : STD_LOGIC;
  SIGNAL or_tmp_1394 : STD_LOGIC;
  SIGNAL nor_tmp_301 : STD_LOGIC;
  SIGNAL or_tmp_1401 : STD_LOGIC;
  SIGNAL operator_64_false_mux1h_2_rgt : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_64_false_acc_mut_64 : STD_LOGIC;
  SIGNAL operator_64_false_acc_mut_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL or_136_cse : STD_LOGIC;
  SIGNAL and_705_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_40_itm : STD_LOGIC;
  SIGNAL operator_64_false_1_or_1_itm : STD_LOGIC;
  SIGNAL STAGE_LOOP_acc_itm_2_1 : STD_LOGIC;
  SIGNAL or_1440_cse : STD_LOGIC;

  SIGNAL modulo_result_or_nl : STD_LOGIC;
  SIGNAL mux_782_nl : STD_LOGIC;
  SIGNAL and_388_nl : STD_LOGIC;
  SIGNAL mux_781_nl : STD_LOGIC;
  SIGNAL mux_780_nl : STD_LOGIC;
  SIGNAL or_864_nl : STD_LOGIC;
  SIGNAL or_862_nl : STD_LOGIC;
  SIGNAL nor_422_nl : STD_LOGIC;
  SIGNAL mux_779_nl : STD_LOGIC;
  SIGNAL mux_778_nl : STD_LOGIC;
  SIGNAL or_859_nl : STD_LOGIC;
  SIGNAL or_857_nl : STD_LOGIC;
  SIGNAL mux_777_nl : STD_LOGIC;
  SIGNAL or_855_nl : STD_LOGIC;
  SIGNAL mux_728_nl : STD_LOGIC;
  SIGNAL mux_727_nl : STD_LOGIC;
  SIGNAL mux_726_nl : STD_LOGIC;
  SIGNAL mux_725_nl : STD_LOGIC;
  SIGNAL mux_724_nl : STD_LOGIC;
  SIGNAL mux_723_nl : STD_LOGIC;
  SIGNAL mux_721_nl : STD_LOGIC;
  SIGNAL mux_720_nl : STD_LOGIC;
  SIGNAL mux_717_nl : STD_LOGIC;
  SIGNAL mux_716_nl : STD_LOGIC;
  SIGNAL mux_715_nl : STD_LOGIC;
  SIGNAL mux_714_nl : STD_LOGIC;
  SIGNAL mux_713_nl : STD_LOGIC;
  SIGNAL nand_41_nl : STD_LOGIC;
  SIGNAL mux_712_nl : STD_LOGIC;
  SIGNAL mux_711_nl : STD_LOGIC;
  SIGNAL mux_710_nl : STD_LOGIC;
  SIGNAL mux_709_nl : STD_LOGIC;
  SIGNAL mux_708_nl : STD_LOGIC;
  SIGNAL mux_707_nl : STD_LOGIC;
  SIGNAL mux_706_nl : STD_LOGIC;
  SIGNAL mux_704_nl : STD_LOGIC;
  SIGNAL mux_703_nl : STD_LOGIC;
  SIGNAL mux_702_nl : STD_LOGIC;
  SIGNAL mux_701_nl : STD_LOGIC;
  SIGNAL mux_700_nl : STD_LOGIC;
  SIGNAL mux_699_nl : STD_LOGIC;
  SIGNAL mux_698_nl : STD_LOGIC;
  SIGNAL mux_697_nl : STD_LOGIC;
  SIGNAL mux_695_nl : STD_LOGIC;
  SIGNAL mux_694_nl : STD_LOGIC;
  SIGNAL mux_693_nl : STD_LOGIC;
  SIGNAL mux_692_nl : STD_LOGIC;
  SIGNAL mux_691_nl : STD_LOGIC;
  SIGNAL or_819_nl : STD_LOGIC;
  SIGNAL mux_690_nl : STD_LOGIC;
  SIGNAL mux_687_nl : STD_LOGIC;
  SIGNAL mux_686_nl : STD_LOGIC;
  SIGNAL mux_685_nl : STD_LOGIC;
  SIGNAL mux_684_nl : STD_LOGIC;
  SIGNAL mux_683_nl : STD_LOGIC;
  SIGNAL nand_40_nl : STD_LOGIC;
  SIGNAL mux_682_nl : STD_LOGIC;
  SIGNAL nand_39_nl : STD_LOGIC;
  SIGNAL or_815_nl : STD_LOGIC;
  SIGNAL or_813_nl : STD_LOGIC;
  SIGNAL mux_681_nl : STD_LOGIC;
  SIGNAL mux_680_nl : STD_LOGIC;
  SIGNAL mux_679_nl : STD_LOGIC;
  SIGNAL mux_678_nl : STD_LOGIC;
  SIGNAL or_808_nl : STD_LOGIC;
  SIGNAL mux_775_nl : STD_LOGIC;
  SIGNAL mux_774_nl : STD_LOGIC;
  SIGNAL mux_773_nl : STD_LOGIC;
  SIGNAL mux_772_nl : STD_LOGIC;
  SIGNAL mux_771_nl : STD_LOGIC;
  SIGNAL mux_770_nl : STD_LOGIC;
  SIGNAL nand_130_nl : STD_LOGIC;
  SIGNAL mux_769_nl : STD_LOGIC;
  SIGNAL nand_44_nl : STD_LOGIC;
  SIGNAL mux_768_nl : STD_LOGIC;
  SIGNAL mux_767_nl : STD_LOGIC;
  SIGNAL nor_423_nl : STD_LOGIC;
  SIGNAL mux_766_nl : STD_LOGIC;
  SIGNAL mux_765_nl : STD_LOGIC;
  SIGNAL mux_764_nl : STD_LOGIC;
  SIGNAL or_850_nl : STD_LOGIC;
  SIGNAL mux_763_nl : STD_LOGIC;
  SIGNAL nor_424_nl : STD_LOGIC;
  SIGNAL mux_762_nl : STD_LOGIC;
  SIGNAL mux_761_nl : STD_LOGIC;
  SIGNAL and_167_nl : STD_LOGIC;
  SIGNAL mux_760_nl : STD_LOGIC;
  SIGNAL mux_759_nl : STD_LOGIC;
  SIGNAL mux_758_nl : STD_LOGIC;
  SIGNAL mux_757_nl : STD_LOGIC;
  SIGNAL mux_756_nl : STD_LOGIC;
  SIGNAL nand_249_nl : STD_LOGIC;
  SIGNAL or_848_nl : STD_LOGIC;
  SIGNAL mux_755_nl : STD_LOGIC;
  SIGNAL mux_754_nl : STD_LOGIC;
  SIGNAL mux_753_nl : STD_LOGIC;
  SIGNAL mux_752_nl : STD_LOGIC;
  SIGNAL mux_751_nl : STD_LOGIC;
  SIGNAL mux_750_nl : STD_LOGIC;
  SIGNAL or_847_nl : STD_LOGIC;
  SIGNAL mux_749_nl : STD_LOGIC;
  SIGNAL nand_43_nl : STD_LOGIC;
  SIGNAL mux_748_nl : STD_LOGIC;
  SIGNAL or_845_nl : STD_LOGIC;
  SIGNAL mux_747_nl : STD_LOGIC;
  SIGNAL mux_746_nl : STD_LOGIC;
  SIGNAL mux_745_nl : STD_LOGIC;
  SIGNAL mux_744_nl : STD_LOGIC;
  SIGNAL mux_743_nl : STD_LOGIC;
  SIGNAL or_843_nl : STD_LOGIC;
  SIGNAL mux_742_nl : STD_LOGIC;
  SIGNAL mux_741_nl : STD_LOGIC;
  SIGNAL or_842_nl : STD_LOGIC;
  SIGNAL mux_740_nl : STD_LOGIC;
  SIGNAL and_165_nl : STD_LOGIC;
  SIGNAL mux_739_nl : STD_LOGIC;
  SIGNAL mux_738_nl : STD_LOGIC;
  SIGNAL mux_737_nl : STD_LOGIC;
  SIGNAL nor_426_nl : STD_LOGIC;
  SIGNAL mux_736_nl : STD_LOGIC;
  SIGNAL mux_735_nl : STD_LOGIC;
  SIGNAL nor_427_nl : STD_LOGIC;
  SIGNAL mux_734_nl : STD_LOGIC;
  SIGNAL mux_733_nl : STD_LOGIC;
  SIGNAL mux_732_nl : STD_LOGIC;
  SIGNAL mux_730_nl : STD_LOGIC;
  SIGNAL mux_729_nl : STD_LOGIC;
  SIGNAL nor_428_nl : STD_LOGIC;
  SIGNAL nor_429_nl : STD_LOGIC;
  SIGNAL nor_430_nl : STD_LOGIC;
  SIGNAL mux_795_nl : STD_LOGIC;
  SIGNAL mux_794_nl : STD_LOGIC;
  SIGNAL mux_793_nl : STD_LOGIC;
  SIGNAL nor_411_nl : STD_LOGIC;
  SIGNAL mux_792_nl : STD_LOGIC;
  SIGNAL and_380_nl : STD_LOGIC;
  SIGNAL nor_412_nl : STD_LOGIC;
  SIGNAL mux_791_nl : STD_LOGIC;
  SIGNAL nor_414_nl : STD_LOGIC;
  SIGNAL mux_790_nl : STD_LOGIC;
  SIGNAL and_381_nl : STD_LOGIC;
  SIGNAL or_881_nl : STD_LOGIC;
  SIGNAL nor_415_nl : STD_LOGIC;
  SIGNAL mux_789_nl : STD_LOGIC;
  SIGNAL and_383_nl : STD_LOGIC;
  SIGNAL or_877_nl : STD_LOGIC;
  SIGNAL mux_788_nl : STD_LOGIC;
  SIGNAL nor_416_nl : STD_LOGIC;
  SIGNAL mux_787_nl : STD_LOGIC;
  SIGNAL nand_47_nl : STD_LOGIC;
  SIGNAL mux_786_nl : STD_LOGIC;
  SIGNAL nand_127_nl : STD_LOGIC;
  SIGNAL or_872_nl : STD_LOGIC;
  SIGNAL mux_785_nl : STD_LOGIC;
  SIGNAL mux_784_nl : STD_LOGIC;
  SIGNAL nor_417_nl : STD_LOGIC;
  SIGNAL nor_418_nl : STD_LOGIC;
  SIGNAL mux_783_nl : STD_LOGIC;
  SIGNAL nor_419_nl : STD_LOGIC;
  SIGNAL and_386_nl : STD_LOGIC;
  SIGNAL nor_659_nl : STD_LOGIC;
  SIGNAL and_704_nl : STD_LOGIC;
  SIGNAL mux_812_nl : STD_LOGIC;
  SIGNAL and_176_nl : STD_LOGIC;
  SIGNAL modExp_while_if_mux1h_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modExp_while_if_or_nl : STD_LOGIC;
  SIGNAL mux_1122_nl : STD_LOGIC;
  SIGNAL mux_1121_nl : STD_LOGIC;
  SIGNAL nor_340_nl : STD_LOGIC;
  SIGNAL mux_1120_nl : STD_LOGIC;
  SIGNAL or_1113_nl : STD_LOGIC;
  SIGNAL mux_1119_nl : STD_LOGIC;
  SIGNAL or_1111_nl : STD_LOGIC;
  SIGNAL or_1109_nl : STD_LOGIC;
  SIGNAL mux_1118_nl : STD_LOGIC;
  SIGNAL nor_341_nl : STD_LOGIC;
  SIGNAL and_324_nl : STD_LOGIC;
  SIGNAL mux_1117_nl : STD_LOGIC;
  SIGNAL nor_342_nl : STD_LOGIC;
  SIGNAL and_492_nl : STD_LOGIC;
  SIGNAL and_325_nl : STD_LOGIC;
  SIGNAL mux_1116_nl : STD_LOGIC;
  SIGNAL nor_344_nl : STD_LOGIC;
  SIGNAL nor_345_nl : STD_LOGIC;
  SIGNAL modExp_while_if_and_1_nl : STD_LOGIC;
  SIGNAL modExp_while_if_and_2_nl : STD_LOGIC;
  SIGNAL and_179_nl : STD_LOGIC;
  SIGNAL mux_856_nl : STD_LOGIC;
  SIGNAL mux_855_nl : STD_LOGIC;
  SIGNAL mux_854_nl : STD_LOGIC;
  SIGNAL mux_853_nl : STD_LOGIC;
  SIGNAL mux_852_nl : STD_LOGIC;
  SIGNAL mux_851_nl : STD_LOGIC;
  SIGNAL mux_850_nl : STD_LOGIC;
  SIGNAL mux_849_nl : STD_LOGIC;
  SIGNAL mux_848_nl : STD_LOGIC;
  SIGNAL mux_847_nl : STD_LOGIC;
  SIGNAL or_1388_nl : STD_LOGIC;
  SIGNAL mux_846_nl : STD_LOGIC;
  SIGNAL mux_844_nl : STD_LOGIC;
  SIGNAL or_928_nl : STD_LOGIC;
  SIGNAL mux_843_nl : STD_LOGIC;
  SIGNAL mux_842_nl : STD_LOGIC;
  SIGNAL mux_841_nl : STD_LOGIC;
  SIGNAL mux_840_nl : STD_LOGIC;
  SIGNAL and_372_nl : STD_LOGIC;
  SIGNAL mux_839_nl : STD_LOGIC;
  SIGNAL mux_838_nl : STD_LOGIC;
  SIGNAL and_373_nl : STD_LOGIC;
  SIGNAL nor_397_nl : STD_LOGIC;
  SIGNAL mux_836_nl : STD_LOGIC;
  SIGNAL mux_835_nl : STD_LOGIC;
  SIGNAL or_925_nl : STD_LOGIC;
  SIGNAL mux_834_nl : STD_LOGIC;
  SIGNAL mux_833_nl : STD_LOGIC;
  SIGNAL mux_832_nl : STD_LOGIC;
  SIGNAL mux_831_nl : STD_LOGIC;
  SIGNAL mux_830_nl : STD_LOGIC;
  SIGNAL mux_829_nl : STD_LOGIC;
  SIGNAL mux_828_nl : STD_LOGIC;
  SIGNAL mux_826_nl : STD_LOGIC;
  SIGNAL mux_825_nl : STD_LOGIC;
  SIGNAL mux_824_nl : STD_LOGIC;
  SIGNAL mux_823_nl : STD_LOGIC;
  SIGNAL mux_822_nl : STD_LOGIC;
  SIGNAL mux_821_nl : STD_LOGIC;
  SIGNAL mux_820_nl : STD_LOGIC;
  SIGNAL mux_819_nl : STD_LOGIC;
  SIGNAL mux_818_nl : STD_LOGIC;
  SIGNAL or_924_nl : STD_LOGIC;
  SIGNAL mux_817_nl : STD_LOGIC;
  SIGNAL mux_816_nl : STD_LOGIC;
  SIGNAL and_376_nl : STD_LOGIC;
  SIGNAL or_923_nl : STD_LOGIC;
  SIGNAL mux_815_nl : STD_LOGIC;
  SIGNAL mux_1423_nl : STD_LOGIC;
  SIGNAL mux_1422_nl : STD_LOGIC;
  SIGNAL mux_1421_nl : STD_LOGIC;
  SIGNAL mux_1420_nl : STD_LOGIC;
  SIGNAL mux_1419_nl : STD_LOGIC;
  SIGNAL or_1550_nl : STD_LOGIC;
  SIGNAL mux_1418_nl : STD_LOGIC;
  SIGNAL or_1499_nl : STD_LOGIC;
  SIGNAL mux_1417_nl : STD_LOGIC;
  SIGNAL mux_1416_nl : STD_LOGIC;
  SIGNAL mux_1415_nl : STD_LOGIC;
  SIGNAL and_707_nl : STD_LOGIC;
  SIGNAL mux_1414_nl : STD_LOGIC;
  SIGNAL mux_1413_nl : STD_LOGIC;
  SIGNAL and_706_nl : STD_LOGIC;
  SIGNAL or_1497_nl : STD_LOGIC;
  SIGNAL mux_1412_nl : STD_LOGIC;
  SIGNAL mux_1411_nl : STD_LOGIC;
  SIGNAL mux_1410_nl : STD_LOGIC;
  SIGNAL mux_1409_nl : STD_LOGIC;
  SIGNAL mux_1408_nl : STD_LOGIC;
  SIGNAL mux_1407_nl : STD_LOGIC;
  SIGNAL mux_1406_nl : STD_LOGIC;
  SIGNAL mux_1405_nl : STD_LOGIC;
  SIGNAL mux_1404_nl : STD_LOGIC;
  SIGNAL mux_1403_nl : STD_LOGIC;
  SIGNAL mux_1402_nl : STD_LOGIC;
  SIGNAL mux_1401_nl : STD_LOGIC;
  SIGNAL mux_1399_nl : STD_LOGIC;
  SIGNAL mux_1398_nl : STD_LOGIC;
  SIGNAL mux_1397_nl : STD_LOGIC;
  SIGNAL mux_1396_nl : STD_LOGIC;
  SIGNAL mux_1395_nl : STD_LOGIC;
  SIGNAL mux_1394_nl : STD_LOGIC;
  SIGNAL mux_1393_nl : STD_LOGIC;
  SIGNAL mux_1392_nl : STD_LOGIC;
  SIGNAL mux_1391_nl : STD_LOGIC;
  SIGNAL mux_1390_nl : STD_LOGIC;
  SIGNAL mux_1389_nl : STD_LOGIC;
  SIGNAL mux_1388_nl : STD_LOGIC;
  SIGNAL nand_275_nl : STD_LOGIC;
  SIGNAL mux_1387_nl : STD_LOGIC;
  SIGNAL mux_1386_nl : STD_LOGIC;
  SIGNAL mux_1385_nl : STD_LOGIC;
  SIGNAL nand_276_nl : STD_LOGIC;
  SIGNAL and_717_nl : STD_LOGIC;
  SIGNAL mux_1384_nl : STD_LOGIC;
  SIGNAL mux_1383_nl : STD_LOGIC;
  SIGNAL mux_1382_nl : STD_LOGIC;
  SIGNAL mux_1381_nl : STD_LOGIC;
  SIGNAL mux_1380_nl : STD_LOGIC;
  SIGNAL mux_1377_nl : STD_LOGIC;
  SIGNAL or_1489_nl : STD_LOGIC;
  SIGNAL mux_1376_nl : STD_LOGIC;
  SIGNAL mux_1374_nl : STD_LOGIC;
  SIGNAL and_718_nl : STD_LOGIC;
  SIGNAL or_1487_nl : STD_LOGIC;
  SIGNAL mux_1373_nl : STD_LOGIC;
  SIGNAL nand_266_nl : STD_LOGIC;
  SIGNAL or_1485_nl : STD_LOGIC;
  SIGNAL mux_1453_nl : STD_LOGIC;
  SIGNAL mux_1452_nl : STD_LOGIC;
  SIGNAL and_710_nl : STD_LOGIC;
  SIGNAL mux_1451_nl : STD_LOGIC;
  SIGNAL or_1540_nl : STD_LOGIC;
  SIGNAL mux_1450_nl : STD_LOGIC;
  SIGNAL or_1539_nl : STD_LOGIC;
  SIGNAL mux_1449_nl : STD_LOGIC;
  SIGNAL mux_1448_nl : STD_LOGIC;
  SIGNAL or_1537_nl : STD_LOGIC;
  SIGNAL nor_676_nl : STD_LOGIC;
  SIGNAL mux_1447_nl : STD_LOGIC;
  SIGNAL mux_1446_nl : STD_LOGIC;
  SIGNAL or_1535_nl : STD_LOGIC;
  SIGNAL or_1534_nl : STD_LOGIC;
  SIGNAL or_1533_nl : STD_LOGIC;
  SIGNAL mux_1445_nl : STD_LOGIC;
  SIGNAL mux_1444_nl : STD_LOGIC;
  SIGNAL mux_1443_nl : STD_LOGIC;
  SIGNAL mux_1442_nl : STD_LOGIC;
  SIGNAL mux_1441_nl : STD_LOGIC;
  SIGNAL nor_677_nl : STD_LOGIC;
  SIGNAL nor_678_nl : STD_LOGIC;
  SIGNAL and_711_nl : STD_LOGIC;
  SIGNAL nor_679_nl : STD_LOGIC;
  SIGNAL nor_680_nl : STD_LOGIC;
  SIGNAL mux_1440_nl : STD_LOGIC;
  SIGNAL mux_1439_nl : STD_LOGIC;
  SIGNAL nor_681_nl : STD_LOGIC;
  SIGNAL nor_682_nl : STD_LOGIC;
  SIGNAL nor_683_nl : STD_LOGIC;
  SIGNAL mux_1438_nl : STD_LOGIC;
  SIGNAL or_1524_nl : STD_LOGIC;
  SIGNAL mux_1437_nl : STD_LOGIC;
  SIGNAL mux_1436_nl : STD_LOGIC;
  SIGNAL mux_1435_nl : STD_LOGIC;
  SIGNAL nor_684_nl : STD_LOGIC;
  SIGNAL mux_1434_nl : STD_LOGIC;
  SIGNAL mux_1433_nl : STD_LOGIC;
  SIGNAL nor_685_nl : STD_LOGIC;
  SIGNAL and_712_nl : STD_LOGIC;
  SIGNAL mux_1432_nl : STD_LOGIC;
  SIGNAL mux_1431_nl : STD_LOGIC;
  SIGNAL mux_1430_nl : STD_LOGIC;
  SIGNAL or_1516_nl : STD_LOGIC;
  SIGNAL or_1513_nl : STD_LOGIC;
  SIGNAL mux_1429_nl : STD_LOGIC;
  SIGNAL and_713_nl : STD_LOGIC;
  SIGNAL mux_1428_nl : STD_LOGIC;
  SIGNAL or_1512_nl : STD_LOGIC;
  SIGNAL mux_1427_nl : STD_LOGIC;
  SIGNAL nand_278_nl : STD_LOGIC;
  SIGNAL nor_686_nl : STD_LOGIC;
  SIGNAL mux_1426_nl : STD_LOGIC;
  SIGNAL mux_1425_nl : STD_LOGIC;
  SIGNAL nand_274_nl : STD_LOGIC;
  SIGNAL or_1505_nl : STD_LOGIC;
  SIGNAL or_1504_nl : STD_LOGIC;
  SIGNAL mux_1424_nl : STD_LOGIC;
  SIGNAL or_1503_nl : STD_LOGIC;
  SIGNAL or_1501_nl : STD_LOGIC;
  SIGNAL nand_263_nl : STD_LOGIC;
  SIGNAL mux_865_nl : STD_LOGIC;
  SIGNAL nor_630_nl : STD_LOGIC;
  SIGNAL mux_864_nl : STD_LOGIC;
  SIGNAL or_940_nl : STD_LOGIC;
  SIGNAL nor_631_nl : STD_LOGIC;
  SIGNAL mux_1457_nl : STD_LOGIC;
  SIGNAL or_1549_nl : STD_LOGIC;
  SIGNAL mux_1456_nl : STD_LOGIC;
  SIGNAL or_1547_nl : STD_LOGIC;
  SIGNAL or_1545_nl : STD_LOGIC;
  SIGNAL nand_271_nl : STD_LOGIC;
  SIGNAL mux_1455_nl : STD_LOGIC;
  SIGNAL nor_674_nl : STD_LOGIC;
  SIGNAL nor_675_nl : STD_LOGIC;
  SIGNAL mux_885_nl : STD_LOGIC;
  SIGNAL mux_884_nl : STD_LOGIC;
  SIGNAL mux_883_nl : STD_LOGIC;
  SIGNAL mux_882_nl : STD_LOGIC;
  SIGNAL nor_389_nl : STD_LOGIC;
  SIGNAL nor_390_nl : STD_LOGIC;
  SIGNAL and_185_nl : STD_LOGIC;
  SIGNAL mux_881_nl : STD_LOGIC;
  SIGNAL and_360_nl : STD_LOGIC;
  SIGNAL mux_880_nl : STD_LOGIC;
  SIGNAL and_184_nl : STD_LOGIC;
  SIGNAL mux_879_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_15_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_16_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_17_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_18_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_19_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_20_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_21_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_22_nl : STD_LOGIC;
  SIGNAL mux_913_nl : STD_LOGIC;
  SIGNAL mux_912_nl : STD_LOGIC;
  SIGNAL mux_911_nl : STD_LOGIC;
  SIGNAL mux_910_nl : STD_LOGIC;
  SIGNAL mux_909_nl : STD_LOGIC;
  SIGNAL or_964_nl : STD_LOGIC;
  SIGNAL mux_908_nl : STD_LOGIC;
  SIGNAL nand_120_nl : STD_LOGIC;
  SIGNAL mux_907_nl : STD_LOGIC;
  SIGNAL mux_906_nl : STD_LOGIC;
  SIGNAL mux_905_nl : STD_LOGIC;
  SIGNAL mux_904_nl : STD_LOGIC;
  SIGNAL mux_903_nl : STD_LOGIC;
  SIGNAL mux_902_nl : STD_LOGIC;
  SIGNAL mux_901_nl : STD_LOGIC;
  SIGNAL nand_121_nl : STD_LOGIC;
  SIGNAL and_192_nl : STD_LOGIC;
  SIGNAL mux_900_nl : STD_LOGIC;
  SIGNAL nand_122_nl : STD_LOGIC;
  SIGNAL mux_899_nl : STD_LOGIC;
  SIGNAL mux_898_nl : STD_LOGIC;
  SIGNAL mux_897_nl : STD_LOGIC;
  SIGNAL nor_388_nl : STD_LOGIC;
  SIGNAL or_959_nl : STD_LOGIC;
  SIGNAL mux_896_nl : STD_LOGIC;
  SIGNAL mux_895_nl : STD_LOGIC;
  SIGNAL mux_894_nl : STD_LOGIC;
  SIGNAL mux_893_nl : STD_LOGIC;
  SIGNAL mux_892_nl : STD_LOGIC;
  SIGNAL mux_891_nl : STD_LOGIC;
  SIGNAL mux_890_nl : STD_LOGIC;
  SIGNAL mux_889_nl : STD_LOGIC;
  SIGNAL or_958_nl : STD_LOGIC;
  SIGNAL mux_888_nl : STD_LOGIC;
  SIGNAL mux_887_nl : STD_LOGIC;
  SIGNAL mux_34_nl : STD_LOGIC;
  SIGNAL mux_33_nl : STD_LOGIC;
  SIGNAL or_42_nl : STD_LOGIC;
  SIGNAL or_41_nl : STD_LOGIC;
  SIGNAL or_39_nl : STD_LOGIC;
  SIGNAL nor_604_nl : STD_LOGIC;
  SIGNAL nor_605_nl : STD_LOGIC;
  SIGNAL mux_915_nl : STD_LOGIC;
  SIGNAL nor_386_nl : STD_LOGIC;
  SIGNAL nor_387_nl : STD_LOGIC;
  SIGNAL and_238_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_26_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_27_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_7_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_8_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_9_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_11_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_12_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_13_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_14_nl : STD_LOGIC;
  SIGNAL mux_48_nl : STD_LOGIC;
  SIGNAL and_470_nl : STD_LOGIC;
  SIGNAL mux_47_nl : STD_LOGIC;
  SIGNAL mux_46_nl : STD_LOGIC;
  SIGNAL nor_591_nl : STD_LOGIC;
  SIGNAL nor_592_nl : STD_LOGIC;
  SIGNAL mux_45_nl : STD_LOGIC;
  SIGNAL nor_593_nl : STD_LOGIC;
  SIGNAL nor_594_nl : STD_LOGIC;
  SIGNAL nor_595_nl : STD_LOGIC;
  SIGNAL mux_44_nl : STD_LOGIC;
  SIGNAL or_62_nl : STD_LOGIC;
  SIGNAL mux_43_nl : STD_LOGIC;
  SIGNAL or_61_nl : STD_LOGIC;
  SIGNAL or_59_nl : STD_LOGIC;
  SIGNAL mux_42_nl : STD_LOGIC;
  SIGNAL nand_224_nl : STD_LOGIC;
  SIGNAL or_56_nl : STD_LOGIC;
  SIGNAL mux_971_nl : STD_LOGIC;
  SIGNAL mux_970_nl : STD_LOGIC;
  SIGNAL mux_349_nl : STD_LOGIC;
  SIGNAL mux_348_nl : STD_LOGIC;
  SIGNAL mux_347_nl : STD_LOGIC;
  SIGNAL or_248_nl : STD_LOGIC;
  SIGNAL nand_9_nl : STD_LOGIC;
  SIGNAL mux_346_nl : STD_LOGIC;
  SIGNAL mux_965_nl : STD_LOGIC;
  SIGNAL mux_964_nl : STD_LOGIC;
  SIGNAL mux_963_nl : STD_LOGIC;
  SIGNAL nor_371_nl : STD_LOGIC;
  SIGNAL or_246_nl : STD_LOGIC;
  SIGNAL mux_343_nl : STD_LOGIC;
  SIGNAL mux_341_nl : STD_LOGIC;
  SIGNAL mux_960_nl : STD_LOGIC;
  SIGNAL nand_56_nl : STD_LOGIC;
  SIGNAL mux_959_nl : STD_LOGIC;
  SIGNAL or_1009_nl : STD_LOGIC;
  SIGNAL mux_958_nl : STD_LOGIC;
  SIGNAL mux_957_nl : STD_LOGIC;
  SIGNAL mux_956_nl : STD_LOGIC;
  SIGNAL mux_955_nl : STD_LOGIC;
  SIGNAL and_246_nl : STD_LOGIC;
  SIGNAL mux_954_nl : STD_LOGIC;
  SIGNAL nor_190_nl : STD_LOGIC;
  SIGNAL mux_333_nl : STD_LOGIC;
  SIGNAL mux_332_nl : STD_LOGIC;
  SIGNAL mux_951_nl : STD_LOGIC;
  SIGNAL mux_950_nl : STD_LOGIC;
  SIGNAL nor_372_nl : STD_LOGIC;
  SIGNAL mux_328_nl : STD_LOGIC;
  SIGNAL mux_948_nl : STD_LOGIC;
  SIGNAL nor_560_nl : STD_LOGIC;
  SIGNAL mux_947_nl : STD_LOGIC;
  SIGNAL mux_334_nl : STD_LOGIC;
  SIGNAL or_1003_nl : STD_LOGIC;
  SIGNAL mux_945_nl : STD_LOGIC;
  SIGNAL mux_944_nl : STD_LOGIC;
  SIGNAL mux_943_nl : STD_LOGIC;
  SIGNAL mux_942_nl : STD_LOGIC;
  SIGNAL or_1002_nl : STD_LOGIC;
  SIGNAL mux_941_nl : STD_LOGIC;
  SIGNAL mux_940_nl : STD_LOGIC;
  SIGNAL or_999_nl : STD_LOGIC;
  SIGNAL mux_939_nl : STD_LOGIC;
  SIGNAL mux_938_nl : STD_LOGIC;
  SIGNAL mux_937_nl : STD_LOGIC;
  SIGNAL mux_936_nl : STD_LOGIC;
  SIGNAL or_1383_nl : STD_LOGIC;
  SIGNAL mux_935_nl : STD_LOGIC;
  SIGNAL mux_934_nl : STD_LOGIC;
  SIGNAL nand_117_nl : STD_LOGIC;
  SIGNAL mux_933_nl : STD_LOGIC;
  SIGNAL or_996_nl : STD_LOGIC;
  SIGNAL or_994_nl : STD_LOGIC;
  SIGNAL mux_932_nl : STD_LOGIC;
  SIGNAL or_231_nl : STD_LOGIC;
  SIGNAL mux_313_nl : STD_LOGIC;
  SIGNAL or_992_nl : STD_LOGIC;
  SIGNAL mux_930_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_31_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_12_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_and_76_nl : STD_LOGIC;
  SIGNAL mux_1032_nl : STD_LOGIC;
  SIGNAL mux_1031_nl : STD_LOGIC;
  SIGNAL mux_1030_nl : STD_LOGIC;
  SIGNAL mux_1029_nl : STD_LOGIC;
  SIGNAL mux_1028_nl : STD_LOGIC;
  SIGNAL mux_1027_nl : STD_LOGIC;
  SIGNAL mux_1026_nl : STD_LOGIC;
  SIGNAL mux_1025_nl : STD_LOGIC;
  SIGNAL nor_205_nl : STD_LOGIC;
  SIGNAL mux_1024_nl : STD_LOGIC;
  SIGNAL mux_1023_nl : STD_LOGIC;
  SIGNAL mux_1022_nl : STD_LOGIC;
  SIGNAL or_1072_nl : STD_LOGIC;
  SIGNAL mux_1021_nl : STD_LOGIC;
  SIGNAL mux_1020_nl : STD_LOGIC;
  SIGNAL mux_1019_nl : STD_LOGIC;
  SIGNAL and_252_nl : STD_LOGIC;
  SIGNAL mux_1018_nl : STD_LOGIC;
  SIGNAL mux_1017_nl : STD_LOGIC;
  SIGNAL mux_1016_nl : STD_LOGIC;
  SIGNAL mux_1015_nl : STD_LOGIC;
  SIGNAL and_340_nl : STD_LOGIC;
  SIGNAL nor_351_nl : STD_LOGIC;
  SIGNAL nor_352_nl : STD_LOGIC;
  SIGNAL mux_1014_nl : STD_LOGIC;
  SIGNAL mux_1013_nl : STD_LOGIC;
  SIGNAL and_251_nl : STD_LOGIC;
  SIGNAL mux_1012_nl : STD_LOGIC;
  SIGNAL mux_1011_nl : STD_LOGIC;
  SIGNAL mux_1010_nl : STD_LOGIC;
  SIGNAL mux_1009_nl : STD_LOGIC;
  SIGNAL mux_1008_nl : STD_LOGIC;
  SIGNAL mux_1007_nl : STD_LOGIC;
  SIGNAL mux_1005_nl : STD_LOGIC;
  SIGNAL mux_1004_nl : STD_LOGIC;
  SIGNAL mux_1003_nl : STD_LOGIC;
  SIGNAL mux_1002_nl : STD_LOGIC;
  SIGNAL or_1061_nl : STD_LOGIC;
  SIGNAL mux_1001_nl : STD_LOGIC;
  SIGNAL mux_1000_nl : STD_LOGIC;
  SIGNAL mux_999_nl : STD_LOGIC;
  SIGNAL or_1059_nl : STD_LOGIC;
  SIGNAL mux_998_nl : STD_LOGIC;
  SIGNAL mux_996_nl : STD_LOGIC;
  SIGNAL nor_353_nl : STD_LOGIC;
  SIGNAL nor_354_nl : STD_LOGIC;
  SIGNAL mux_995_nl : STD_LOGIC;
  SIGNAL mux_987_nl : STD_LOGIC;
  SIGNAL or_1432_nl : STD_LOGIC;
  SIGNAL or_1433_nl : STD_LOGIC;
  SIGNAL mux_986_nl : STD_LOGIC;
  SIGNAL mux_985_nl : STD_LOGIC;
  SIGNAL or_1040_nl : STD_LOGIC;
  SIGNAL or_1039_nl : STD_LOGIC;
  SIGNAL or_1037_nl : STD_LOGIC;
  SIGNAL mux_1035_nl : STD_LOGIC;
  SIGNAL nor_347_nl : STD_LOGIC;
  SIGNAL mux_1034_nl : STD_LOGIC;
  SIGNAL nand_108_nl : STD_LOGIC;
  SIGNAL or_1082_nl : STD_LOGIC;
  SIGNAL nor_348_nl : STD_LOGIC;
  SIGNAL mux_1033_nl : STD_LOGIC;
  SIGNAL or_1078_nl : STD_LOGIC;
  SIGNAL or_1077_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_8_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mux_1139_nl : STD_LOGIC;
  SIGNAL mux_1138_nl : STD_LOGIC;
  SIGNAL nor_334_nl : STD_LOGIC;
  SIGNAL mux_1137_nl : STD_LOGIC;
  SIGNAL or_1146_nl : STD_LOGIC;
  SIGNAL or_1145_nl : STD_LOGIC;
  SIGNAL mux_1136_nl : STD_LOGIC;
  SIGNAL nor_335_nl : STD_LOGIC;
  SIGNAL mux_1135_nl : STD_LOGIC;
  SIGNAL or_1142_nl : STD_LOGIC;
  SIGNAL or_1141_nl : STD_LOGIC;
  SIGNAL and_321_nl : STD_LOGIC;
  SIGNAL mux_1134_nl : STD_LOGIC;
  SIGNAL nor_336_nl : STD_LOGIC;
  SIGNAL mux_1133_nl : STD_LOGIC;
  SIGNAL or_1137_nl : STD_LOGIC;
  SIGNAL or_1136_nl : STD_LOGIC;
  SIGNAL and_322_nl : STD_LOGIC;
  SIGNAL mux_1132_nl : STD_LOGIC;
  SIGNAL nor_337_nl : STD_LOGIC;
  SIGNAL nor_338_nl : STD_LOGIC;
  SIGNAL mux_1156_nl : STD_LOGIC;
  SIGNAL mux_1155_nl : STD_LOGIC;
  SIGNAL nand_98_nl : STD_LOGIC;
  SIGNAL nand_99_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_145_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_nl : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL mux_1174_nl : STD_LOGIC;
  SIGNAL mux_1173_nl : STD_LOGIC;
  SIGNAL mux_1172_nl : STD_LOGIC;
  SIGNAL mux_1171_nl : STD_LOGIC;
  SIGNAL mux_1169_nl : STD_LOGIC;
  SIGNAL mux_1168_nl : STD_LOGIC;
  SIGNAL mux_1167_nl : STD_LOGIC;
  SIGNAL mux_1166_nl : STD_LOGIC;
  SIGNAL mux_1165_nl : STD_LOGIC;
  SIGNAL mux_1163_nl : STD_LOGIC;
  SIGNAL and_315_nl : STD_LOGIC;
  SIGNAL mux_1181_nl : STD_LOGIC;
  SIGNAL mux_1180_nl : STD_LOGIC;
  SIGNAL mux_1179_nl : STD_LOGIC;
  SIGNAL mux_1177_nl : STD_LOGIC;
  SIGNAL and_313_nl : STD_LOGIC;
  SIGNAL mux_1176_nl : STD_LOGIC;
  SIGNAL mux_1184_nl : STD_LOGIC;
  SIGNAL nand_234_nl : STD_LOGIC;
  SIGNAL mux_1183_nl : STD_LOGIC;
  SIGNAL or_1193_nl : STD_LOGIC;
  SIGNAL mux_1186_nl : STD_LOGIC;
  SIGNAL nor_328_nl : STD_LOGIC;
  SIGNAL mux_1185_nl : STD_LOGIC;
  SIGNAL and_272_nl : STD_LOGIC;
  SIGNAL and_271_nl : STD_LOGIC;
  SIGNAL or_1200_nl : STD_LOGIC;
  SIGNAL mux_1187_nl : STD_LOGIC;
  SIGNAL or_100_nl : STD_LOGIC;
  SIGNAL or_1197_nl : STD_LOGIC;
  SIGNAL or_1201_nl : STD_LOGIC;
  SIGNAL mux_1192_nl : STD_LOGIC;
  SIGNAL mux_1191_nl : STD_LOGIC;
  SIGNAL nor_327_nl : STD_LOGIC;
  SIGNAL mux_1190_nl : STD_LOGIC;
  SIGNAL and_274_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux_nl : STD_LOGIC;
  SIGNAL mux_1246_nl : STD_LOGIC;
  SIGNAL mux_1245_nl : STD_LOGIC;
  SIGNAL and_306_nl : STD_LOGIC;
  SIGNAL mux_1244_nl : STD_LOGIC;
  SIGNAL mux_1243_nl : STD_LOGIC;
  SIGNAL nor_316_nl : STD_LOGIC;
  SIGNAL nor_317_nl : STD_LOGIC;
  SIGNAL nor_318_nl : STD_LOGIC;
  SIGNAL nor_319_nl : STD_LOGIC;
  SIGNAL mux_1242_nl : STD_LOGIC;
  SIGNAL and_307_nl : STD_LOGIC;
  SIGNAL mux_1241_nl : STD_LOGIC;
  SIGNAL nor_320_nl : STD_LOGIC;
  SIGNAL and_493_nl : STD_LOGIC;
  SIGNAL nor_322_nl : STD_LOGIC;
  SIGNAL mux_1240_nl : STD_LOGIC;
  SIGNAL or_1229_nl : STD_LOGIC;
  SIGNAL nand_95_nl : STD_LOGIC;
  SIGNAL mux_1196_nl : STD_LOGIC;
  SIGNAL nor_324_nl : STD_LOGIC;
  SIGNAL mux_1195_nl : STD_LOGIC;
  SIGNAL or_1210_nl : STD_LOGIC;
  SIGNAL nor_325_nl : STD_LOGIC;
  SIGNAL mux_1194_nl : STD_LOGIC;
  SIGNAL or_1208_nl : STD_LOGIC;
  SIGNAL mux_1249_nl : STD_LOGIC;
  SIGNAL or_1430_nl : STD_LOGIC;
  SIGNAL or_1431_nl : STD_LOGIC;
  SIGNAL mux_1248_nl : STD_LOGIC;
  SIGNAL or_1245_nl : STD_LOGIC;
  SIGNAL mux_1247_nl : STD_LOGIC;
  SIGNAL or_1244_nl : STD_LOGIC;
  SIGNAL or_1243_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_52_nl : STD_LOGIC;
  SIGNAL mux_1285_nl : STD_LOGIC;
  SIGNAL mux_1284_nl : STD_LOGIC;
  SIGNAL nand_259_nl : STD_LOGIC;
  SIGNAL mux_1283_nl : STD_LOGIC;
  SIGNAL nor_304_nl : STD_LOGIC;
  SIGNAL nor_305_nl : STD_LOGIC;
  SIGNAL nand_260_nl : STD_LOGIC;
  SIGNAL mux_1282_nl : STD_LOGIC;
  SIGNAL nand_261_nl : STD_LOGIC;
  SIGNAL mux_1281_nl : STD_LOGIC;
  SIGNAL nor_306_nl : STD_LOGIC;
  SIGNAL nor_307_nl : STD_LOGIC;
  SIGNAL mux_1280_nl : STD_LOGIC;
  SIGNAL or_1283_nl : STD_LOGIC;
  SIGNAL nand_226_nl : STD_LOGIC;
  SIGNAL or_1483_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_66_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_68_nl : STD_LOGIC;
  SIGNAL mux_1320_nl : STD_LOGIC;
  SIGNAL mux_1319_nl : STD_LOGIC;
  SIGNAL mux_1318_nl : STD_LOGIC;
  SIGNAL mux_1317_nl : STD_LOGIC;
  SIGNAL nand_86_nl : STD_LOGIC;
  SIGNAL or_1323_nl : STD_LOGIC;
  SIGNAL mux_1316_nl : STD_LOGIC;
  SIGNAL mux_1315_nl : STD_LOGIC;
  SIGNAL mux_1314_nl : STD_LOGIC;
  SIGNAL nand_247_nl : STD_LOGIC;
  SIGNAL or_1366_nl : STD_LOGIC;
  SIGNAL or_1367_nl : STD_LOGIC;
  SIGNAL mux_1313_nl : STD_LOGIC;
  SIGNAL mux_1312_nl : STD_LOGIC;
  SIGNAL or_1316_nl : STD_LOGIC;
  SIGNAL mux_1311_nl : STD_LOGIC;
  SIGNAL mux_1310_nl : STD_LOGIC;
  SIGNAL mux_1309_nl : STD_LOGIC;
  SIGNAL mux_1308_nl : STD_LOGIC;
  SIGNAL mux_1307_nl : STD_LOGIC;
  SIGNAL mux_1306_nl : STD_LOGIC;
  SIGNAL or_1314_nl : STD_LOGIC;
  SIGNAL mux_1304_nl : STD_LOGIC;
  SIGNAL mux_1303_nl : STD_LOGIC;
  SIGNAL mux_1302_nl : STD_LOGIC;
  SIGNAL mux_1301_nl : STD_LOGIC;
  SIGNAL mux_1300_nl : STD_LOGIC;
  SIGNAL mux_1299_nl : STD_LOGIC;
  SIGNAL mux_1298_nl : STD_LOGIC;
  SIGNAL mux_1297_nl : STD_LOGIC;
  SIGNAL mux_1296_nl : STD_LOGIC;
  SIGNAL mux_1295_nl : STD_LOGIC;
  SIGNAL or_1311_nl : STD_LOGIC;
  SIGNAL mux_1294_nl : STD_LOGIC;
  SIGNAL mux_1293_nl : STD_LOGIC;
  SIGNAL or_1309_nl : STD_LOGIC;
  SIGNAL or_1307_nl : STD_LOGIC;
  SIGNAL mux_1323_nl : STD_LOGIC;
  SIGNAL or_1434_nl : STD_LOGIC;
  SIGNAL or_1435_nl : STD_LOGIC;
  SIGNAL mux_1322_nl : STD_LOGIC;
  SIGNAL or_1329_nl : STD_LOGIC;
  SIGNAL mux_1321_nl : STD_LOGIC;
  SIGNAL or_1328_nl : STD_LOGIC;
  SIGNAL or_1326_nl : STD_LOGIC;
  SIGNAL mux_1326_nl : STD_LOGIC;
  SIGNAL and_282_nl : STD_LOGIC;
  SIGNAL mux_1325_nl : STD_LOGIC;
  SIGNAL nor_292_nl : STD_LOGIC;
  SIGNAL mux_1324_nl : STD_LOGIC;
  SIGNAL nor_293_nl : STD_LOGIC;
  SIGNAL and_283_nl : STD_LOGIC;
  SIGNAL nor_294_nl : STD_LOGIC;
  SIGNAL nor_295_nl : STD_LOGIC;
  SIGNAL or_1402_nl : STD_LOGIC;
  SIGNAL nand_199_nl : STD_LOGIC;
  SIGNAL mux_361_nl : STD_LOGIC;
  SIGNAL and_432_nl : STD_LOGIC;
  SIGNAL mux_381_nl : STD_LOGIC;
  SIGNAL or_308_nl : STD_LOGIC;
  SIGNAL or_306_nl : STD_LOGIC;
  SIGNAL or_325_nl : STD_LOGIC;
  SIGNAL or_323_nl : STD_LOGIC;
  SIGNAL mux_418_nl : STD_LOGIC;
  SIGNAL or_375_nl : STD_LOGIC;
  SIGNAL or_373_nl : STD_LOGIC;
  SIGNAL mux_456_nl : STD_LOGIC;
  SIGNAL nor_512_nl : STD_LOGIC;
  SIGNAL nor_513_nl : STD_LOGIC;
  SIGNAL mux_494_nl : STD_LOGIC;
  SIGNAL nor_496_nl : STD_LOGIC;
  SIGNAL nor_497_nl : STD_LOGIC;
  SIGNAL mux_538_nl : STD_LOGIC;
  SIGNAL or_570_nl : STD_LOGIC;
  SIGNAL or_568_nl : STD_LOGIC;
  SIGNAL mux_575_nl : STD_LOGIC;
  SIGNAL or_635_nl : STD_LOGIC;
  SIGNAL or_633_nl : STD_LOGIC;
  SIGNAL mux_612_nl : STD_LOGIC;
  SIGNAL nor_458_nl : STD_LOGIC;
  SIGNAL nor_459_nl : STD_LOGIC;
  SIGNAL mux_649_nl : STD_LOGIC;
  SIGNAL nor_444_nl : STD_LOGIC;
  SIGNAL nor_445_nl : STD_LOGIC;
  SIGNAL or_854_nl : STD_LOGIC;
  SIGNAL or_853_nl : STD_LOGIC;
  SIGNAL nor_405_nl : STD_LOGIC;
  SIGNAL mux_801_nl : STD_LOGIC;
  SIGNAL mux_800_nl : STD_LOGIC;
  SIGNAL or_903_nl : STD_LOGIC;
  SIGNAL or_902_nl : STD_LOGIC;
  SIGNAL nand_49_nl : STD_LOGIC;
  SIGNAL mux_799_nl : STD_LOGIC;
  SIGNAL and_489_nl : STD_LOGIC;
  SIGNAL nor_407_nl : STD_LOGIC;
  SIGNAL mux_798_nl : STD_LOGIC;
  SIGNAL nor_408_nl : STD_LOGIC;
  SIGNAL mux_797_nl : STD_LOGIC;
  SIGNAL nor_409_nl : STD_LOGIC;
  SIGNAL mux_796_nl : STD_LOGIC;
  SIGNAL or_895_nl : STD_LOGIC;
  SIGNAL or_893_nl : STD_LOGIC;
  SIGNAL nor_410_nl : STD_LOGIC;
  SIGNAL mux_807_nl : STD_LOGIC;
  SIGNAL nor_400_nl : STD_LOGIC;
  SIGNAL mux_806_nl : STD_LOGIC;
  SIGNAL or_1362_nl : STD_LOGIC;
  SIGNAL or_913_nl : STD_LOGIC;
  SIGNAL mux_805_nl : STD_LOGIC;
  SIGNAL nor_401_nl : STD_LOGIC;
  SIGNAL and_377_nl : STD_LOGIC;
  SIGNAL mux_804_nl : STD_LOGIC;
  SIGNAL nor_402_nl : STD_LOGIC;
  SIGNAL and_378_nl : STD_LOGIC;
  SIGNAL mux_803_nl : STD_LOGIC;
  SIGNAL nor_403_nl : STD_LOGIC;
  SIGNAL nor_404_nl : STD_LOGIC;
  SIGNAL mux_811_nl : STD_LOGIC;
  SIGNAL mux_810_nl : STD_LOGIC;
  SIGNAL mux_809_nl : STD_LOGIC;
  SIGNAL or_916_nl : STD_LOGIC;
  SIGNAL mux_814_nl : STD_LOGIC;
  SIGNAL nor_398_nl : STD_LOGIC;
  SIGNAL nor_399_nl : STD_LOGIC;
  SIGNAL or_955_nl : STD_LOGIC;
  SIGNAL mux_919_nl : STD_LOGIC;
  SIGNAL mux_918_nl : STD_LOGIC;
  SIGNAL nor_382_nl : STD_LOGIC;
  SIGNAL and_474_nl : STD_LOGIC;
  SIGNAL mux_30_nl : STD_LOGIC;
  SIGNAL nor_603_nl : STD_LOGIC;
  SIGNAL and_475_nl : STD_LOGIC;
  SIGNAL mux_977_nl : STD_LOGIC;
  SIGNAL nor_366_nl : STD_LOGIC;
  SIGNAL mux_976_nl : STD_LOGIC;
  SIGNAL or_1026_nl : STD_LOGIC;
  SIGNAL or_1024_nl : STD_LOGIC;
  SIGNAL nor_367_nl : STD_LOGIC;
  SIGNAL mux_975_nl : STD_LOGIC;
  SIGNAL and_350_nl : STD_LOGIC;
  SIGNAL mux_974_nl : STD_LOGIC;
  SIGNAL nor_368_nl : STD_LOGIC;
  SIGNAL mux_973_nl : STD_LOGIC;
  SIGNAL and_351_nl : STD_LOGIC;
  SIGNAL nor_369_nl : STD_LOGIC;
  SIGNAL nor_370_nl : STD_LOGIC;
  SIGNAL mux_993_nl : STD_LOGIC;
  SIGNAL mux_992_nl : STD_LOGIC;
  SIGNAL and_344_nl : STD_LOGIC;
  SIGNAL mux_991_nl : STD_LOGIC;
  SIGNAL and_345_nl : STD_LOGIC;
  SIGNAL nor_355_nl : STD_LOGIC;
  SIGNAL nor_356_nl : STD_LOGIC;
  SIGNAL mux_990_nl : STD_LOGIC;
  SIGNAL and_346_nl : STD_LOGIC;
  SIGNAL mux_989_nl : STD_LOGIC;
  SIGNAL nor_358_nl : STD_LOGIC;
  SIGNAL mux_988_nl : STD_LOGIC;
  SIGNAL nand_111_nl : STD_LOGIC;
  SIGNAL or_1045_nl : STD_LOGIC;
  SIGNAL or_1183_nl : STD_LOGIC;
  SIGNAL mux_1157_nl : STD_LOGIC;
  SIGNAL and_320_nl : STD_LOGIC;
  SIGNAL and_263_nl : STD_LOGIC;
  SIGNAL mux_1161_nl : STD_LOGIC;
  SIGNAL nor_329_nl : STD_LOGIC;
  SIGNAL mux_1272_nl : STD_LOGIC;
  SIGNAL mux_1271_nl : STD_LOGIC;
  SIGNAL mux_1270_nl : STD_LOGIC;
  SIGNAL mux_1269_nl : STD_LOGIC;
  SIGNAL mux_1268_nl : STD_LOGIC;
  SIGNAL or_1268_nl : STD_LOGIC;
  SIGNAL mux_1267_nl : STD_LOGIC;
  SIGNAL or_1267_nl : STD_LOGIC;
  SIGNAL mux_1266_nl : STD_LOGIC;
  SIGNAL mux_1265_nl : STD_LOGIC;
  SIGNAL mux_1264_nl : STD_LOGIC;
  SIGNAL mux_1263_nl : STD_LOGIC;
  SIGNAL or_1263_nl : STD_LOGIC;
  SIGNAL mux_1262_nl : STD_LOGIC;
  SIGNAL mux_1261_nl : STD_LOGIC;
  SIGNAL mux_1260_nl : STD_LOGIC;
  SIGNAL mux_1259_nl : STD_LOGIC;
  SIGNAL mux_1258_nl : STD_LOGIC;
  SIGNAL mux_1257_nl : STD_LOGIC;
  SIGNAL nand_227_nl : STD_LOGIC;
  SIGNAL or_1258_nl : STD_LOGIC;
  SIGNAL mux_1256_nl : STD_LOGIC;
  SIGNAL or_1256_nl : STD_LOGIC;
  SIGNAL mux_1255_nl : STD_LOGIC;
  SIGNAL mux_1254_nl : STD_LOGIC;
  SIGNAL or_1254_nl : STD_LOGIC;
  SIGNAL mux_1253_nl : STD_LOGIC;
  SIGNAL mux_1252_nl : STD_LOGIC;
  SIGNAL mux_1250_nl : STD_LOGIC;
  SIGNAL or_1249_nl : STD_LOGIC;
  SIGNAL mux_1276_nl : STD_LOGIC;
  SIGNAL and_294_nl : STD_LOGIC;
  SIGNAL mux_1275_nl : STD_LOGIC;
  SIGNAL nor_310_nl : STD_LOGIC;
  SIGNAL and_295_nl : STD_LOGIC;
  SIGNAL mux_1291_nl : STD_LOGIC;
  SIGNAL mux_1290_nl : STD_LOGIC;
  SIGNAL nor_300_nl : STD_LOGIC;
  SIGNAL mux_1289_nl : STD_LOGIC;
  SIGNAL or_1304_nl : STD_LOGIC;
  SIGNAL or_1303_nl : STD_LOGIC;
  SIGNAL nor_628_nl : STD_LOGIC;
  SIGNAL and_289_nl : STD_LOGIC;
  SIGNAL mux_1288_nl : STD_LOGIC;
  SIGNAL nor_303_nl : STD_LOGIC;
  SIGNAL mux_1287_nl : STD_LOGIC;
  SIGNAL or_1295_nl : STD_LOGIC;
  SIGNAL mux_1286_nl : STD_LOGIC;
  SIGNAL or_1093_nl : STD_LOGIC;
  SIGNAL or_1292_nl : STD_LOGIC;
  SIGNAL mux_877_nl : STD_LOGIC;
  SIGNAL mux_876_nl : STD_LOGIC;
  SIGNAL mux_875_nl : STD_LOGIC;
  SIGNAL mux_874_nl : STD_LOGIC;
  SIGNAL and_363_nl : STD_LOGIC;
  SIGNAL and_364_nl : STD_LOGIC;
  SIGNAL STAGE_LOOP_acc_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_361_nl : STD_LOGIC;
  SIGNAL mux_983_nl : STD_LOGIC;
  SIGNAL mux_982_nl : STD_LOGIC;
  SIGNAL or_1381_nl : STD_LOGIC;
  SIGNAL or_1382_nl : STD_LOGIC;
  SIGNAL nand_113_nl : STD_LOGIC;
  SIGNAL mux_981_nl : STD_LOGIC;
  SIGNAL nor_362_nl : STD_LOGIC;
  SIGNAL and_348_nl : STD_LOGIC;
  SIGNAL and_349_nl : STD_LOGIC;
  SIGNAL mux_980_nl : STD_LOGIC;
  SIGNAL nor_363_nl : STD_LOGIC;
  SIGNAL mux_979_nl : STD_LOGIC;
  SIGNAL nor_364_nl : STD_LOGIC;
  SIGNAL nor_365_nl : STD_LOGIC;
  SIGNAL and_91_nl : STD_LOGIC;
  SIGNAL mux_370_nl : STD_LOGIC;
  SIGNAL mux_369_nl : STD_LOGIC;
  SIGNAL mux_368_nl : STD_LOGIC;
  SIGNAL and_419_nl : STD_LOGIC;
  SIGNAL mux_367_nl : STD_LOGIC;
  SIGNAL nor_553_nl : STD_LOGIC;
  SIGNAL nor_554_nl : STD_LOGIC;
  SIGNAL nor_555_nl : STD_LOGIC;
  SIGNAL and_420_nl : STD_LOGIC;
  SIGNAL mux_366_nl : STD_LOGIC;
  SIGNAL and_421_nl : STD_LOGIC;
  SIGNAL nor_556_nl : STD_LOGIC;
  SIGNAL and_422_nl : STD_LOGIC;
  SIGNAL mux_365_nl : STD_LOGIC;
  SIGNAL nor_557_nl : STD_LOGIC;
  SIGNAL nor_558_nl : STD_LOGIC;
  SIGNAL mux_364_nl : STD_LOGIC;
  SIGNAL or_269_nl : STD_LOGIC;
  SIGNAL or_268_nl : STD_LOGIC;
  SIGNAL and_96_nl : STD_LOGIC;
  SIGNAL mux_371_nl : STD_LOGIC;
  SIGNAL nor_551_nl : STD_LOGIC;
  SIGNAL nor_552_nl : STD_LOGIC;
  SIGNAL and_104_nl : STD_LOGIC;
  SIGNAL mux_372_nl : STD_LOGIC;
  SIGNAL nor_549_nl : STD_LOGIC;
  SIGNAL nor_550_nl : STD_LOGIC;
  SIGNAL and_115_nl : STD_LOGIC;
  SIGNAL mux_373_nl : STD_LOGIC;
  SIGNAL nor_547_nl : STD_LOGIC;
  SIGNAL nor_548_nl : STD_LOGIC;
  SIGNAL and_123_nl : STD_LOGIC;
  SIGNAL mux_374_nl : STD_LOGIC;
  SIGNAL nor_545_nl : STD_LOGIC;
  SIGNAL nor_546_nl : STD_LOGIC;
  SIGNAL and_136_nl : STD_LOGIC;
  SIGNAL mux_375_nl : STD_LOGIC;
  SIGNAL nor_544_nl : STD_LOGIC;
  SIGNAL and_143_nl : STD_LOGIC;
  SIGNAL mux_376_nl : STD_LOGIC;
  SIGNAL nor_542_nl : STD_LOGIC;
  SIGNAL nor_543_nl : STD_LOGIC;
  SIGNAL and_152_nl : STD_LOGIC;
  SIGNAL mux_377_nl : STD_LOGIC;
  SIGNAL and_500_nl : STD_LOGIC;
  SIGNAL nor_541_nl : STD_LOGIC;
  SIGNAL mux_399_nl : STD_LOGIC;
  SIGNAL mux_398_nl : STD_LOGIC;
  SIGNAL mux_397_nl : STD_LOGIC;
  SIGNAL mux_396_nl : STD_LOGIC;
  SIGNAL mux_395_nl : STD_LOGIC;
  SIGNAL or_331_nl : STD_LOGIC;
  SIGNAL mux_394_nl : STD_LOGIC;
  SIGNAL mux_393_nl : STD_LOGIC;
  SIGNAL or_326_nl : STD_LOGIC;
  SIGNAL mux_391_nl : STD_LOGIC;
  SIGNAL mux_390_nl : STD_LOGIC;
  SIGNAL mux_389_nl : STD_LOGIC;
  SIGNAL mux_388_nl : STD_LOGIC;
  SIGNAL or_321_nl : STD_LOGIC;
  SIGNAL mux_387_nl : STD_LOGIC;
  SIGNAL or_316_nl : STD_LOGIC;
  SIGNAL mux_386_nl : STD_LOGIC;
  SIGNAL mux_385_nl : STD_LOGIC;
  SIGNAL or_313_nl : STD_LOGIC;
  SIGNAL mux_384_nl : STD_LOGIC;
  SIGNAL mux_383_nl : STD_LOGIC;
  SIGNAL mux_382_nl : STD_LOGIC;
  SIGNAL or_311_nl : STD_LOGIC;
  SIGNAL or_305_nl : STD_LOGIC;
  SIGNAL mux_380_nl : STD_LOGIC;
  SIGNAL mux_379_nl : STD_LOGIC;
  SIGNAL mux_378_nl : STD_LOGIC;
  SIGNAL or_302_nl : STD_LOGIC;
  SIGNAL or_301_nl : STD_LOGIC;
  SIGNAL or_299_nl : STD_LOGIC;
  SIGNAL or_298_nl : STD_LOGIC;
  SIGNAL mux_413_nl : STD_LOGIC;
  SIGNAL nor_528_nl : STD_LOGIC;
  SIGNAL mux_412_nl : STD_LOGIC;
  SIGNAL nand_15_nl : STD_LOGIC;
  SIGNAL mux_411_nl : STD_LOGIC;
  SIGNAL nor_529_nl : STD_LOGIC;
  SIGNAL nor_530_nl : STD_LOGIC;
  SIGNAL or_359_nl : STD_LOGIC;
  SIGNAL mux_410_nl : STD_LOGIC;
  SIGNAL or_358_nl : STD_LOGIC;
  SIGNAL or_357_nl : STD_LOGIC;
  SIGNAL mux_409_nl : STD_LOGIC;
  SIGNAL and_417_nl : STD_LOGIC;
  SIGNAL mux_408_nl : STD_LOGIC;
  SIGNAL nor_531_nl : STD_LOGIC;
  SIGNAL nor_532_nl : STD_LOGIC;
  SIGNAL nor_533_nl : STD_LOGIC;
  SIGNAL mux_407_nl : STD_LOGIC;
  SIGNAL mux_406_nl : STD_LOGIC;
  SIGNAL mux_405_nl : STD_LOGIC;
  SIGNAL nor_534_nl : STD_LOGIC;
  SIGNAL nor_535_nl : STD_LOGIC;
  SIGNAL mux_404_nl : STD_LOGIC;
  SIGNAL or_347_nl : STD_LOGIC;
  SIGNAL or_345_nl : STD_LOGIC;
  SIGNAL nor_536_nl : STD_LOGIC;
  SIGNAL nor_537_nl : STD_LOGIC;
  SIGNAL mux_403_nl : STD_LOGIC;
  SIGNAL mux_402_nl : STD_LOGIC;
  SIGNAL or_340_nl : STD_LOGIC;
  SIGNAL mux_401_nl : STD_LOGIC;
  SIGNAL or_339_nl : STD_LOGIC;
  SIGNAL or_337_nl : STD_LOGIC;
  SIGNAL nand_13_nl : STD_LOGIC;
  SIGNAL mux_400_nl : STD_LOGIC;
  SIGNAL nor_538_nl : STD_LOGIC;
  SIGNAL nor_539_nl : STD_LOGIC;
  SIGNAL or_332_nl : STD_LOGIC;
  SIGNAL mux_436_nl : STD_LOGIC;
  SIGNAL mux_435_nl : STD_LOGIC;
  SIGNAL mux_434_nl : STD_LOGIC;
  SIGNAL mux_433_nl : STD_LOGIC;
  SIGNAL mux_432_nl : STD_LOGIC;
  SIGNAL or_398_nl : STD_LOGIC;
  SIGNAL mux_431_nl : STD_LOGIC;
  SIGNAL mux_430_nl : STD_LOGIC;
  SIGNAL or_393_nl : STD_LOGIC;
  SIGNAL mux_428_nl : STD_LOGIC;
  SIGNAL mux_427_nl : STD_LOGIC;
  SIGNAL mux_426_nl : STD_LOGIC;
  SIGNAL mux_425_nl : STD_LOGIC;
  SIGNAL or_388_nl : STD_LOGIC;
  SIGNAL mux_424_nl : STD_LOGIC;
  SIGNAL or_383_nl : STD_LOGIC;
  SIGNAL mux_423_nl : STD_LOGIC;
  SIGNAL mux_422_nl : STD_LOGIC;
  SIGNAL or_380_nl : STD_LOGIC;
  SIGNAL mux_421_nl : STD_LOGIC;
  SIGNAL mux_420_nl : STD_LOGIC;
  SIGNAL mux_419_nl : STD_LOGIC;
  SIGNAL or_378_nl : STD_LOGIC;
  SIGNAL or_372_nl : STD_LOGIC;
  SIGNAL mux_417_nl : STD_LOGIC;
  SIGNAL mux_416_nl : STD_LOGIC;
  SIGNAL mux_415_nl : STD_LOGIC;
  SIGNAL or_369_nl : STD_LOGIC;
  SIGNAL or_368_nl : STD_LOGIC;
  SIGNAL or_366_nl : STD_LOGIC;
  SIGNAL or_365_nl : STD_LOGIC;
  SIGNAL mux_451_nl : STD_LOGIC;
  SIGNAL mux_450_nl : STD_LOGIC;
  SIGNAL mux_449_nl : STD_LOGIC;
  SIGNAL nor_514_nl : STD_LOGIC;
  SIGNAL mux_448_nl : STD_LOGIC;
  SIGNAL or_423_nl : STD_LOGIC;
  SIGNAL or_421_nl : STD_LOGIC;
  SIGNAL nor_515_nl : STD_LOGIC;
  SIGNAL nor_516_nl : STD_LOGIC;
  SIGNAL mux_447_nl : STD_LOGIC;
  SIGNAL and_414_nl : STD_LOGIC;
  SIGNAL mux_446_nl : STD_LOGIC;
  SIGNAL nor_517_nl : STD_LOGIC;
  SIGNAL nor_518_nl : STD_LOGIC;
  SIGNAL nor_519_nl : STD_LOGIC;
  SIGNAL mux_445_nl : STD_LOGIC;
  SIGNAL or_411_nl : STD_LOGIC;
  SIGNAL or_410_nl : STD_LOGIC;
  SIGNAL mux_444_nl : STD_LOGIC;
  SIGNAL mux_443_nl : STD_LOGIC;
  SIGNAL nor_520_nl : STD_LOGIC;
  SIGNAL mux_442_nl : STD_LOGIC;
  SIGNAL nor_521_nl : STD_LOGIC;
  SIGNAL nor_522_nl : STD_LOGIC;
  SIGNAL mux_441_nl : STD_LOGIC;
  SIGNAL mux_440_nl : STD_LOGIC;
  SIGNAL mux_439_nl : STD_LOGIC;
  SIGNAL nor_523_nl : STD_LOGIC;
  SIGNAL nor_524_nl : STD_LOGIC;
  SIGNAL and_415_nl : STD_LOGIC;
  SIGNAL mux_438_nl : STD_LOGIC;
  SIGNAL mux_437_nl : STD_LOGIC;
  SIGNAL nor_525_nl : STD_LOGIC;
  SIGNAL nor_526_nl : STD_LOGIC;
  SIGNAL or_400_nl : STD_LOGIC;
  SIGNAL nor_527_nl : STD_LOGIC;
  SIGNAL mux_474_nl : STD_LOGIC;
  SIGNAL mux_473_nl : STD_LOGIC;
  SIGNAL mux_472_nl : STD_LOGIC;
  SIGNAL mux_471_nl : STD_LOGIC;
  SIGNAL mux_470_nl : STD_LOGIC;
  SIGNAL or_457_nl : STD_LOGIC;
  SIGNAL mux_469_nl : STD_LOGIC;
  SIGNAL mux_468_nl : STD_LOGIC;
  SIGNAL or_452_nl : STD_LOGIC;
  SIGNAL mux_466_nl : STD_LOGIC;
  SIGNAL mux_465_nl : STD_LOGIC;
  SIGNAL mux_464_nl : STD_LOGIC;
  SIGNAL mux_463_nl : STD_LOGIC;
  SIGNAL or_447_nl : STD_LOGIC;
  SIGNAL mux_462_nl : STD_LOGIC;
  SIGNAL or_442_nl : STD_LOGIC;
  SIGNAL mux_461_nl : STD_LOGIC;
  SIGNAL mux_460_nl : STD_LOGIC;
  SIGNAL or_439_nl : STD_LOGIC;
  SIGNAL mux_459_nl : STD_LOGIC;
  SIGNAL mux_458_nl : STD_LOGIC;
  SIGNAL mux_457_nl : STD_LOGIC;
  SIGNAL or_437_nl : STD_LOGIC;
  SIGNAL or_432_nl : STD_LOGIC;
  SIGNAL mux_455_nl : STD_LOGIC;
  SIGNAL mux_454_nl : STD_LOGIC;
  SIGNAL mux_453_nl : STD_LOGIC;
  SIGNAL or_429_nl : STD_LOGIC;
  SIGNAL or_428_nl : STD_LOGIC;
  SIGNAL or_426_nl : STD_LOGIC;
  SIGNAL or_425_nl : STD_LOGIC;
  SIGNAL mux_489_nl : STD_LOGIC;
  SIGNAL mux_488_nl : STD_LOGIC;
  SIGNAL mux_487_nl : STD_LOGIC;
  SIGNAL nor_498_nl : STD_LOGIC;
  SIGNAL mux_486_nl : STD_LOGIC;
  SIGNAL or_482_nl : STD_LOGIC;
  SIGNAL or_480_nl : STD_LOGIC;
  SIGNAL nor_499_nl : STD_LOGIC;
  SIGNAL nor_500_nl : STD_LOGIC;
  SIGNAL mux_485_nl : STD_LOGIC;
  SIGNAL and_411_nl : STD_LOGIC;
  SIGNAL mux_484_nl : STD_LOGIC;
  SIGNAL nor_501_nl : STD_LOGIC;
  SIGNAL nor_502_nl : STD_LOGIC;
  SIGNAL nor_503_nl : STD_LOGIC;
  SIGNAL mux_483_nl : STD_LOGIC;
  SIGNAL or_470_nl : STD_LOGIC;
  SIGNAL or_469_nl : STD_LOGIC;
  SIGNAL mux_482_nl : STD_LOGIC;
  SIGNAL mux_481_nl : STD_LOGIC;
  SIGNAL nor_504_nl : STD_LOGIC;
  SIGNAL mux_480_nl : STD_LOGIC;
  SIGNAL nor_505_nl : STD_LOGIC;
  SIGNAL nor_506_nl : STD_LOGIC;
  SIGNAL mux_479_nl : STD_LOGIC;
  SIGNAL mux_478_nl : STD_LOGIC;
  SIGNAL mux_477_nl : STD_LOGIC;
  SIGNAL nor_507_nl : STD_LOGIC;
  SIGNAL nor_508_nl : STD_LOGIC;
  SIGNAL and_412_nl : STD_LOGIC;
  SIGNAL mux_476_nl : STD_LOGIC;
  SIGNAL mux_475_nl : STD_LOGIC;
  SIGNAL nor_509_nl : STD_LOGIC;
  SIGNAL nor_510_nl : STD_LOGIC;
  SIGNAL or_459_nl : STD_LOGIC;
  SIGNAL nor_511_nl : STD_LOGIC;
  SIGNAL mux_512_nl : STD_LOGIC;
  SIGNAL mux_511_nl : STD_LOGIC;
  SIGNAL mux_510_nl : STD_LOGIC;
  SIGNAL mux_509_nl : STD_LOGIC;
  SIGNAL mux_508_nl : STD_LOGIC;
  SIGNAL or_516_nl : STD_LOGIC;
  SIGNAL mux_507_nl : STD_LOGIC;
  SIGNAL mux_506_nl : STD_LOGIC;
  SIGNAL or_511_nl : STD_LOGIC;
  SIGNAL mux_504_nl : STD_LOGIC;
  SIGNAL mux_503_nl : STD_LOGIC;
  SIGNAL mux_502_nl : STD_LOGIC;
  SIGNAL mux_501_nl : STD_LOGIC;
  SIGNAL or_506_nl : STD_LOGIC;
  SIGNAL mux_500_nl : STD_LOGIC;
  SIGNAL or_501_nl : STD_LOGIC;
  SIGNAL mux_499_nl : STD_LOGIC;
  SIGNAL mux_498_nl : STD_LOGIC;
  SIGNAL or_498_nl : STD_LOGIC;
  SIGNAL mux_497_nl : STD_LOGIC;
  SIGNAL mux_496_nl : STD_LOGIC;
  SIGNAL mux_495_nl : STD_LOGIC;
  SIGNAL or_496_nl : STD_LOGIC;
  SIGNAL or_491_nl : STD_LOGIC;
  SIGNAL mux_493_nl : STD_LOGIC;
  SIGNAL mux_492_nl : STD_LOGIC;
  SIGNAL mux_491_nl : STD_LOGIC;
  SIGNAL or_488_nl : STD_LOGIC;
  SIGNAL or_487_nl : STD_LOGIC;
  SIGNAL or_485_nl : STD_LOGIC;
  SIGNAL or_484_nl : STD_LOGIC;
  SIGNAL mux_526_nl : STD_LOGIC;
  SIGNAL nor_484_nl : STD_LOGIC;
  SIGNAL mux_525_nl : STD_LOGIC;
  SIGNAL nand_24_nl : STD_LOGIC;
  SIGNAL mux_524_nl : STD_LOGIC;
  SIGNAL nor_485_nl : STD_LOGIC;
  SIGNAL nor_486_nl : STD_LOGIC;
  SIGNAL or_544_nl : STD_LOGIC;
  SIGNAL mux_523_nl : STD_LOGIC;
  SIGNAL or_543_nl : STD_LOGIC;
  SIGNAL or_542_nl : STD_LOGIC;
  SIGNAL mux_522_nl : STD_LOGIC;
  SIGNAL and_410_nl : STD_LOGIC;
  SIGNAL mux_521_nl : STD_LOGIC;
  SIGNAL and_499_nl : STD_LOGIC;
  SIGNAL nor_488_nl : STD_LOGIC;
  SIGNAL nor_489_nl : STD_LOGIC;
  SIGNAL mux_520_nl : STD_LOGIC;
  SIGNAL mux_519_nl : STD_LOGIC;
  SIGNAL mux_518_nl : STD_LOGIC;
  SIGNAL nor_490_nl : STD_LOGIC;
  SIGNAL nor_491_nl : STD_LOGIC;
  SIGNAL mux_517_nl : STD_LOGIC;
  SIGNAL or_532_nl : STD_LOGIC;
  SIGNAL or_530_nl : STD_LOGIC;
  SIGNAL nor_492_nl : STD_LOGIC;
  SIGNAL nor_493_nl : STD_LOGIC;
  SIGNAL mux_516_nl : STD_LOGIC;
  SIGNAL mux_515_nl : STD_LOGIC;
  SIGNAL or_525_nl : STD_LOGIC;
  SIGNAL mux_514_nl : STD_LOGIC;
  SIGNAL nand_232_nl : STD_LOGIC;
  SIGNAL or_522_nl : STD_LOGIC;
  SIGNAL nand_22_nl : STD_LOGIC;
  SIGNAL mux_513_nl : STD_LOGIC;
  SIGNAL nor_494_nl : STD_LOGIC;
  SIGNAL nor_495_nl : STD_LOGIC;
  SIGNAL or_517_nl : STD_LOGIC;
  SIGNAL mux_549_nl : STD_LOGIC;
  SIGNAL mux_548_nl : STD_LOGIC;
  SIGNAL mux_547_nl : STD_LOGIC;
  SIGNAL mux_546_nl : STD_LOGIC;
  SIGNAL or_582_nl : STD_LOGIC;
  SIGNAL or_580_nl : STD_LOGIC;
  SIGNAL mux_545_nl : STD_LOGIC;
  SIGNAL mux_544_nl : STD_LOGIC;
  SIGNAL mux_543_nl : STD_LOGIC;
  SIGNAL or_579_nl : STD_LOGIC;
  SIGNAL or_578_nl : STD_LOGIC;
  SIGNAL or_576_nl : STD_LOGIC;
  SIGNAL mux_542_nl : STD_LOGIC;
  SIGNAL mux_541_nl : STD_LOGIC;
  SIGNAL mux_540_nl : STD_LOGIC;
  SIGNAL mux_539_nl : STD_LOGIC;
  SIGNAL or_575_nl : STD_LOGIC;
  SIGNAL mux_537_nl : STD_LOGIC;
  SIGNAL mux_536_nl : STD_LOGIC;
  SIGNAL or_566_nl : STD_LOGIC;
  SIGNAL mux_534_nl : STD_LOGIC;
  SIGNAL mux_533_nl : STD_LOGIC;
  SIGNAL mux_532_nl : STD_LOGIC;
  SIGNAL mux_531_nl : STD_LOGIC;
  SIGNAL or_559_nl : STD_LOGIC;
  SIGNAL mux_530_nl : STD_LOGIC;
  SIGNAL or_554_nl : STD_LOGIC;
  SIGNAL mux_529_nl : STD_LOGIC;
  SIGNAL mux_528_nl : STD_LOGIC;
  SIGNAL or_551_nl : STD_LOGIC;
  SIGNAL nor_114_nl : STD_LOGIC;
  SIGNAL mux_563_nl : STD_LOGIC;
  SIGNAL nor_472_nl : STD_LOGIC;
  SIGNAL mux_562_nl : STD_LOGIC;
  SIGNAL nand_27_nl : STD_LOGIC;
  SIGNAL mux_561_nl : STD_LOGIC;
  SIGNAL nor_474_nl : STD_LOGIC;
  SIGNAL or_609_nl : STD_LOGIC;
  SIGNAL mux_560_nl : STD_LOGIC;
  SIGNAL or_608_nl : STD_LOGIC;
  SIGNAL or_607_nl : STD_LOGIC;
  SIGNAL mux_559_nl : STD_LOGIC;
  SIGNAL and_409_nl : STD_LOGIC;
  SIGNAL mux_558_nl : STD_LOGIC;
  SIGNAL nor_475_nl : STD_LOGIC;
  SIGNAL nor_476_nl : STD_LOGIC;
  SIGNAL nor_477_nl : STD_LOGIC;
  SIGNAL mux_557_nl : STD_LOGIC;
  SIGNAL mux_556_nl : STD_LOGIC;
  SIGNAL mux_555_nl : STD_LOGIC;
  SIGNAL nor_478_nl : STD_LOGIC;
  SIGNAL nor_479_nl : STD_LOGIC;
  SIGNAL mux_554_nl : STD_LOGIC;
  SIGNAL or_598_nl : STD_LOGIC;
  SIGNAL or_596_nl : STD_LOGIC;
  SIGNAL nor_480_nl : STD_LOGIC;
  SIGNAL nor_481_nl : STD_LOGIC;
  SIGNAL mux_553_nl : STD_LOGIC;
  SIGNAL mux_552_nl : STD_LOGIC;
  SIGNAL or_591_nl : STD_LOGIC;
  SIGNAL mux_551_nl : STD_LOGIC;
  SIGNAL or_590_nl : STD_LOGIC;
  SIGNAL or_589_nl : STD_LOGIC;
  SIGNAL nand_25_nl : STD_LOGIC;
  SIGNAL mux_550_nl : STD_LOGIC;
  SIGNAL nor_482_nl : STD_LOGIC;
  SIGNAL or_583_nl : STD_LOGIC;
  SIGNAL mux_586_nl : STD_LOGIC;
  SIGNAL mux_585_nl : STD_LOGIC;
  SIGNAL mux_584_nl : STD_LOGIC;
  SIGNAL mux_583_nl : STD_LOGIC;
  SIGNAL or_647_nl : STD_LOGIC;
  SIGNAL or_645_nl : STD_LOGIC;
  SIGNAL mux_582_nl : STD_LOGIC;
  SIGNAL mux_581_nl : STD_LOGIC;
  SIGNAL mux_580_nl : STD_LOGIC;
  SIGNAL or_644_nl : STD_LOGIC;
  SIGNAL or_643_nl : STD_LOGIC;
  SIGNAL or_641_nl : STD_LOGIC;
  SIGNAL mux_579_nl : STD_LOGIC;
  SIGNAL mux_578_nl : STD_LOGIC;
  SIGNAL mux_577_nl : STD_LOGIC;
  SIGNAL mux_576_nl : STD_LOGIC;
  SIGNAL or_640_nl : STD_LOGIC;
  SIGNAL mux_574_nl : STD_LOGIC;
  SIGNAL mux_573_nl : STD_LOGIC;
  SIGNAL or_631_nl : STD_LOGIC;
  SIGNAL mux_571_nl : STD_LOGIC;
  SIGNAL mux_570_nl : STD_LOGIC;
  SIGNAL mux_569_nl : STD_LOGIC;
  SIGNAL mux_568_nl : STD_LOGIC;
  SIGNAL or_624_nl : STD_LOGIC;
  SIGNAL mux_567_nl : STD_LOGIC;
  SIGNAL or_619_nl : STD_LOGIC;
  SIGNAL mux_566_nl : STD_LOGIC;
  SIGNAL mux_565_nl : STD_LOGIC;
  SIGNAL or_616_nl : STD_LOGIC;
  SIGNAL nor_120_nl : STD_LOGIC;
  SIGNAL mux_600_nl : STD_LOGIC;
  SIGNAL nor_460_nl : STD_LOGIC;
  SIGNAL mux_599_nl : STD_LOGIC;
  SIGNAL nand_30_nl : STD_LOGIC;
  SIGNAL mux_598_nl : STD_LOGIC;
  SIGNAL nor_462_nl : STD_LOGIC;
  SIGNAL or_674_nl : STD_LOGIC;
  SIGNAL mux_597_nl : STD_LOGIC;
  SIGNAL or_673_nl : STD_LOGIC;
  SIGNAL or_672_nl : STD_LOGIC;
  SIGNAL mux_596_nl : STD_LOGIC;
  SIGNAL and_408_nl : STD_LOGIC;
  SIGNAL mux_595_nl : STD_LOGIC;
  SIGNAL and_498_nl : STD_LOGIC;
  SIGNAL nor_464_nl : STD_LOGIC;
  SIGNAL nor_465_nl : STD_LOGIC;
  SIGNAL mux_594_nl : STD_LOGIC;
  SIGNAL mux_593_nl : STD_LOGIC;
  SIGNAL mux_592_nl : STD_LOGIC;
  SIGNAL nor_466_nl : STD_LOGIC;
  SIGNAL nor_467_nl : STD_LOGIC;
  SIGNAL mux_591_nl : STD_LOGIC;
  SIGNAL or_663_nl : STD_LOGIC;
  SIGNAL or_661_nl : STD_LOGIC;
  SIGNAL nor_468_nl : STD_LOGIC;
  SIGNAL nor_469_nl : STD_LOGIC;
  SIGNAL mux_590_nl : STD_LOGIC;
  SIGNAL mux_589_nl : STD_LOGIC;
  SIGNAL or_656_nl : STD_LOGIC;
  SIGNAL mux_588_nl : STD_LOGIC;
  SIGNAL or_655_nl : STD_LOGIC;
  SIGNAL or_654_nl : STD_LOGIC;
  SIGNAL nand_28_nl : STD_LOGIC;
  SIGNAL mux_587_nl : STD_LOGIC;
  SIGNAL nor_470_nl : STD_LOGIC;
  SIGNAL or_648_nl : STD_LOGIC;
  SIGNAL mux_623_nl : STD_LOGIC;
  SIGNAL mux_622_nl : STD_LOGIC;
  SIGNAL mux_621_nl : STD_LOGIC;
  SIGNAL mux_620_nl : STD_LOGIC;
  SIGNAL or_711_nl : STD_LOGIC;
  SIGNAL or_709_nl : STD_LOGIC;
  SIGNAL mux_619_nl : STD_LOGIC;
  SIGNAL mux_618_nl : STD_LOGIC;
  SIGNAL mux_617_nl : STD_LOGIC;
  SIGNAL or_708_nl : STD_LOGIC;
  SIGNAL or_707_nl : STD_LOGIC;
  SIGNAL or_705_nl : STD_LOGIC;
  SIGNAL mux_616_nl : STD_LOGIC;
  SIGNAL mux_615_nl : STD_LOGIC;
  SIGNAL mux_614_nl : STD_LOGIC;
  SIGNAL mux_613_nl : STD_LOGIC;
  SIGNAL or_704_nl : STD_LOGIC;
  SIGNAL mux_611_nl : STD_LOGIC;
  SIGNAL mux_610_nl : STD_LOGIC;
  SIGNAL or_696_nl : STD_LOGIC;
  SIGNAL mux_608_nl : STD_LOGIC;
  SIGNAL mux_607_nl : STD_LOGIC;
  SIGNAL mux_606_nl : STD_LOGIC;
  SIGNAL mux_605_nl : STD_LOGIC;
  SIGNAL or_689_nl : STD_LOGIC;
  SIGNAL mux_604_nl : STD_LOGIC;
  SIGNAL or_684_nl : STD_LOGIC;
  SIGNAL mux_603_nl : STD_LOGIC;
  SIGNAL mux_602_nl : STD_LOGIC;
  SIGNAL or_681_nl : STD_LOGIC;
  SIGNAL nor_126_nl : STD_LOGIC;
  SIGNAL mux_637_nl : STD_LOGIC;
  SIGNAL nor_446_nl : STD_LOGIC;
  SIGNAL mux_636_nl : STD_LOGIC;
  SIGNAL nand_34_nl : STD_LOGIC;
  SIGNAL mux_635_nl : STD_LOGIC;
  SIGNAL nor_448_nl : STD_LOGIC;
  SIGNAL or_738_nl : STD_LOGIC;
  SIGNAL mux_634_nl : STD_LOGIC;
  SIGNAL or_737_nl : STD_LOGIC;
  SIGNAL or_736_nl : STD_LOGIC;
  SIGNAL mux_633_nl : STD_LOGIC;
  SIGNAL and_407_nl : STD_LOGIC;
  SIGNAL mux_632_nl : STD_LOGIC;
  SIGNAL and_497_nl : STD_LOGIC;
  SIGNAL nor_450_nl : STD_LOGIC;
  SIGNAL nor_451_nl : STD_LOGIC;
  SIGNAL mux_631_nl : STD_LOGIC;
  SIGNAL mux_630_nl : STD_LOGIC;
  SIGNAL mux_629_nl : STD_LOGIC;
  SIGNAL nor_452_nl : STD_LOGIC;
  SIGNAL nor_453_nl : STD_LOGIC;
  SIGNAL mux_628_nl : STD_LOGIC;
  SIGNAL or_727_nl : STD_LOGIC;
  SIGNAL or_725_nl : STD_LOGIC;
  SIGNAL nor_454_nl : STD_LOGIC;
  SIGNAL nor_455_nl : STD_LOGIC;
  SIGNAL mux_627_nl : STD_LOGIC;
  SIGNAL mux_626_nl : STD_LOGIC;
  SIGNAL or_720_nl : STD_LOGIC;
  SIGNAL mux_625_nl : STD_LOGIC;
  SIGNAL or_719_nl : STD_LOGIC;
  SIGNAL or_718_nl : STD_LOGIC;
  SIGNAL nand_32_nl : STD_LOGIC;
  SIGNAL mux_624_nl : STD_LOGIC;
  SIGNAL nor_456_nl : STD_LOGIC;
  SIGNAL or_712_nl : STD_LOGIC;
  SIGNAL mux_660_nl : STD_LOGIC;
  SIGNAL mux_659_nl : STD_LOGIC;
  SIGNAL mux_658_nl : STD_LOGIC;
  SIGNAL mux_657_nl : STD_LOGIC;
  SIGNAL nand_251_nl : STD_LOGIC;
  SIGNAL or_773_nl : STD_LOGIC;
  SIGNAL mux_656_nl : STD_LOGIC;
  SIGNAL mux_655_nl : STD_LOGIC;
  SIGNAL mux_654_nl : STD_LOGIC;
  SIGNAL or_772_nl : STD_LOGIC;
  SIGNAL nand_252_nl : STD_LOGIC;
  SIGNAL nand_144_nl : STD_LOGIC;
  SIGNAL mux_653_nl : STD_LOGIC;
  SIGNAL mux_652_nl : STD_LOGIC;
  SIGNAL mux_651_nl : STD_LOGIC;
  SIGNAL mux_650_nl : STD_LOGIC;
  SIGNAL nand_250_nl : STD_LOGIC;
  SIGNAL mux_648_nl : STD_LOGIC;
  SIGNAL mux_647_nl : STD_LOGIC;
  SIGNAL or_760_nl : STD_LOGIC;
  SIGNAL mux_645_nl : STD_LOGIC;
  SIGNAL mux_644_nl : STD_LOGIC;
  SIGNAL mux_643_nl : STD_LOGIC;
  SIGNAL mux_642_nl : STD_LOGIC;
  SIGNAL nand_147_nl : STD_LOGIC;
  SIGNAL mux_641_nl : STD_LOGIC;
  SIGNAL or_748_nl : STD_LOGIC;
  SIGNAL mux_640_nl : STD_LOGIC;
  SIGNAL mux_639_nl : STD_LOGIC;
  SIGNAL nand_149_nl : STD_LOGIC;
  SIGNAL and_406_nl : STD_LOGIC;
  SIGNAL mux_674_nl : STD_LOGIC;
  SIGNAL nor_433_nl : STD_LOGIC;
  SIGNAL mux_673_nl : STD_LOGIC;
  SIGNAL nand_38_nl : STD_LOGIC;
  SIGNAL mux_672_nl : STD_LOGIC;
  SIGNAL nor_435_nl : STD_LOGIC;
  SIGNAL or_802_nl : STD_LOGIC;
  SIGNAL mux_671_nl : STD_LOGIC;
  SIGNAL nand_134_nl : STD_LOGIC;
  SIGNAL or_800_nl : STD_LOGIC;
  SIGNAL mux_670_nl : STD_LOGIC;
  SIGNAL and_404_nl : STD_LOGIC;
  SIGNAL mux_669_nl : STD_LOGIC;
  SIGNAL and_495_nl : STD_LOGIC;
  SIGNAL nor_437_nl : STD_LOGIC;
  SIGNAL nor_438_nl : STD_LOGIC;
  SIGNAL mux_668_nl : STD_LOGIC;
  SIGNAL mux_667_nl : STD_LOGIC;
  SIGNAL mux_666_nl : STD_LOGIC;
  SIGNAL nor_439_nl : STD_LOGIC;
  SIGNAL nor_440_nl : STD_LOGIC;
  SIGNAL mux_665_nl : STD_LOGIC;
  SIGNAL nand_237_nl : STD_LOGIC;
  SIGNAL or_789_nl : STD_LOGIC;
  SIGNAL and_405_nl : STD_LOGIC;
  SIGNAL nor_441_nl : STD_LOGIC;
  SIGNAL mux_664_nl : STD_LOGIC;
  SIGNAL mux_663_nl : STD_LOGIC;
  SIGNAL or_784_nl : STD_LOGIC;
  SIGNAL mux_662_nl : STD_LOGIC;
  SIGNAL nand_139_nl : STD_LOGIC;
  SIGNAL nand_231_nl : STD_LOGIC;
  SIGNAL nand_36_nl : STD_LOGIC;
  SIGNAL mux_661_nl : STD_LOGIC;
  SIGNAL nor_442_nl : STD_LOGIC;
  SIGNAL or_776_nl : STD_LOGIC;
  SIGNAL mux_1347_nl : STD_LOGIC;
  SIGNAL nor_635_nl : STD_LOGIC;
  SIGNAL nor_636_nl : STD_LOGIC;
  SIGNAL mux_1346_nl : STD_LOGIC;
  SIGNAL nor_637_nl : STD_LOGIC;
  SIGNAL mux_1345_nl : STD_LOGIC;
  SIGNAL and_nl : STD_LOGIC;
  SIGNAL mux_1344_nl : STD_LOGIC;
  SIGNAL or_1438_nl : STD_LOGIC;
  SIGNAL mux_1372_nl : STD_LOGIC;
  SIGNAL or_1436_nl : STD_LOGIC;
  SIGNAL acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_7_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_mux_8_nl : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_or_44_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_mux_9_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_8_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_9_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_45_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL COMP_LOOP_mux1h_125_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL and_722_nl : STD_LOGIC;
  SIGNAL and_723_nl : STD_LOGIC;
  SIGNAL and_724_nl : STD_LOGIC;
  SIGNAL and_725_nl : STD_LOGIC;
  SIGNAL and_726_nl : STD_LOGIC;
  SIGNAL and_727_nl : STD_LOGIC;
  SIGNAL acc_2_nl : STD_LOGIC_VECTOR (65 DOWNTO 0);
  SIGNAL COMP_LOOP_mux1h_126_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_or_46_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_11_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_12_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL COMP_LOOP_and_85_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL COMP_LOOP_nor_107_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_13_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL COMP_LOOP_mux_41_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL operator_64_false_1_operator_64_false_1_or_53_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_54_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_55_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_51_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_56_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_52_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_57_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_53_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_58_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_54_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_59_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_55_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_60_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_56_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_61_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_57_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_62_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_58_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_63_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_59_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_64_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_60_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_65_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_61_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_66_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_62_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_67_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_63_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_68_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_64_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_69_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_65_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_70_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_66_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_71_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_67_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_72_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_68_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_73_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_69_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_74_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_70_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_75_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_71_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_76_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_72_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_77_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_73_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_78_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_74_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_79_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_75_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_80_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_76_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_81_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_77_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_82_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_78_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_83_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_79_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_84_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_80_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_85_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_81_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_86_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_82_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_87_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_83_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_88_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_84_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_89_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_85_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_90_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_86_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_91_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_87_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_92_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_88_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_93_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_89_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_94_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_90_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_95_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_91_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_96_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_92_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_97_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_93_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_98_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_94_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_99_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_95_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_100_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_96_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_101_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_97_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_102_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_98_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_103_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_99_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_104_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_100_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_operator_64_false_1_or_105_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_101_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_or_7_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL operator_64_false_1_operator_64_false_1_nor_105_nl : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL operator_64_false_1_mux1h_4_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL operator_64_false_1_or_8_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux1h_5_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL operator_64_false_1_and_53_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL operator_64_false_1_mux1h_6_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL operator_64_false_1_not_3_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux1h_7_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL operator_64_false_1_or_9_nl : STD_LOGIC;
  SIGNAL modExp_while_if_mux1h_2_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL and_728_nl : STD_LOGIC;
  SIGNAL mux_1459_nl : STD_LOGIC;
  SIGNAL mux_1460_nl : STD_LOGIC;
  SIGNAL mux_1461_nl : STD_LOGIC;
  SIGNAL nor_690_nl : STD_LOGIC;
  SIGNAL nor_691_nl : STD_LOGIC;
  SIGNAL mux_1462_nl : STD_LOGIC;
  SIGNAL or_1560_nl : STD_LOGIC;
  SIGNAL or_1561_nl : STD_LOGIC;
  SIGNAL mux_1463_nl : STD_LOGIC;
  SIGNAL nor_692_nl : STD_LOGIC;
  SIGNAL and_729_nl : STD_LOGIC;
  SIGNAL mux_1464_nl : STD_LOGIC;
  SIGNAL nor_693_nl : STD_LOGIC;
  SIGNAL mux_1465_nl : STD_LOGIC;
  SIGNAL or_1562_nl : STD_LOGIC;
  SIGNAL and_730_nl : STD_LOGIC;
  SIGNAL mux_1466_nl : STD_LOGIC;
  SIGNAL nor_694_nl : STD_LOGIC;
  SIGNAL nor_695_nl : STD_LOGIC;
  SIGNAL mux_1467_nl : STD_LOGIC;
  SIGNAL mux_1468_nl : STD_LOGIC;
  SIGNAL nand_279_nl : STD_LOGIC;
  SIGNAL mux_1469_nl : STD_LOGIC;
  SIGNAL nor_696_nl : STD_LOGIC;
  SIGNAL nor_697_nl : STD_LOGIC;
  SIGNAL mux_1470_nl : STD_LOGIC;
  SIGNAL mux_1471_nl : STD_LOGIC;
  SIGNAL mux_1472_nl : STD_LOGIC;
  SIGNAL or_1564_nl : STD_LOGIC;
  SIGNAL or_1565_nl : STD_LOGIC;
  SIGNAL or_1566_nl : STD_LOGIC;
  SIGNAL mux_1473_nl : STD_LOGIC;
  SIGNAL or_1567_nl : STD_LOGIC;
  SIGNAL or_1568_nl : STD_LOGIC;
  SIGNAL mux_1474_nl : STD_LOGIC;
  SIGNAL mux_1475_nl : STD_LOGIC;
  SIGNAL mux_1476_nl : STD_LOGIC;
  SIGNAL or_1569_nl : STD_LOGIC;
  SIGNAL mux_1477_nl : STD_LOGIC;
  SIGNAL or_1570_nl : STD_LOGIC;
  SIGNAL or_1571_nl : STD_LOGIC;
  SIGNAL mux_1478_nl : STD_LOGIC;
  SIGNAL mux_1479_nl : STD_LOGIC;
  SIGNAL nand_280_nl : STD_LOGIC;
  SIGNAL mux_1480_nl : STD_LOGIC;
  SIGNAL nand_281_nl : STD_LOGIC;
  SIGNAL mux_1481_nl : STD_LOGIC;
  SIGNAL or_1572_nl : STD_LOGIC;
  SIGNAL p_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL p_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL r_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL r_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL modulo_result_rem_cmp_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_result_rem_cmp_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_result_rem_cmp_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL operator_66_true_div_cmp_a_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_b : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL STAGE_LOOP_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_rg_z : STD_LOGIC_VECTOR (9 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      STAGE_LOOP_C_8_tr0 : IN STD_LOGIC;
      modExp_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_1_tr0 : IN STD_LOGIC;
      COMP_LOOP_1_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_62_tr0 : IN STD_LOGIC;
      COMP_LOOP_2_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_124_tr0 : IN STD_LOGIC;
      COMP_LOOP_3_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_186_tr0 : IN STD_LOGIC;
      COMP_LOOP_4_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_248_tr0 : IN STD_LOGIC;
      COMP_LOOP_5_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_310_tr0 : IN STD_LOGIC;
      COMP_LOOP_6_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_372_tr0 : IN STD_LOGIC;
      COMP_LOOP_7_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_434_tr0 : IN STD_LOGIC;
      COMP_LOOP_8_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_496_tr0 : IN STD_LOGIC;
      VEC_LOOP_C_0_tr0 : IN STD_LOGIC;
      STAGE_LOOP_C_9_tr0 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (9 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_62_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_124_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_186_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_248_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_310_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_372_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_434_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_s_1_3_2(input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_4_2(input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_7_2(input_6 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
      tmp := sel(6);
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_3_2(input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_6_2(input_5 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_3_2(input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_13_2(input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(12 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_3_2(input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_4_2(input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_5_2(input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_9_2(input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(8 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_65_3_2(input_2 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(64 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(64 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_7_3_2(input_2 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_8_6_2(input_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_9_11_2(input_10 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(10 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(8 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(8 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_10_2_2(input_0 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(9 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_12_2_2(input_0 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(11 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_3_2_2(input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_4_2_2(input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_63_2_2(input_0 : STD_LOGIC_VECTOR(62 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(62 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(62 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_64_2_2(input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_65_2_2(input_0 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(64 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_6_2_2(input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_7_2_2(input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_9_2_2(input_0 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(8 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  p_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 2,
      width => 64
      )
    PORT MAP(
      dat => p_rsci_dat,
      idat => p_rsci_idat_1
    );
  p_rsci_dat <= p_rsc_dat;
  p_rsci_idat <= p_rsci_idat_1;

  r_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 3,
      width => 64
      )
    PORT MAP(
      dat => r_rsci_dat,
      idat => r_rsci_idat_1
    );
  r_rsci_dat <= r_rsc_dat;
  r_rsci_idat <= r_rsci_idat_1;

  vec_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_7_obj_ld_cse,
      lz => vec_rsc_triosy_0_7_lz
    );
  vec_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_7_obj_ld_cse,
      lz => vec_rsc_triosy_0_6_lz
    );
  vec_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_7_obj_ld_cse,
      lz => vec_rsc_triosy_0_5_lz
    );
  vec_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_7_obj_ld_cse,
      lz => vec_rsc_triosy_0_4_lz
    );
  vec_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_7_obj_ld_cse,
      lz => vec_rsc_triosy_0_3_lz
    );
  vec_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_7_obj_ld_cse,
      lz => vec_rsc_triosy_0_2_lz
    );
  vec_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_7_obj_ld_cse,
      lz => vec_rsc_triosy_0_1_lz
    );
  vec_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_7_obj_ld_cse,
      lz => vec_rsc_triosy_0_0_lz
    );
  p_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_7_obj_ld_cse,
      lz => p_rsc_triosy_lz
    );
  r_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_7_obj_ld_cse,
      lz => r_rsc_triosy_lz
    );
  modulo_result_rem_cmp : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 1
      )
    PORT MAP(
      a => modulo_result_rem_cmp_a_1,
      b => modulo_result_rem_cmp_b_1,
      z => modulo_result_rem_cmp_z_1
    );
  modulo_result_rem_cmp_a_1 <= modulo_result_rem_cmp_a;
  modulo_result_rem_cmp_b_1 <= modulo_result_rem_cmp_b;
  modulo_result_rem_cmp_z <= modulo_result_rem_cmp_z_1;

  operator_66_true_div_cmp : work.mgc_comps.mgc_div
    GENERIC MAP(
      width_a => 65,
      width_b => 11,
      signd => 1
      )
    PORT MAP(
      a => operator_66_true_div_cmp_a_1,
      b => operator_66_true_div_cmp_b,
      z => operator_66_true_div_cmp_z_1
    );
  operator_66_true_div_cmp_a_1 <= operator_66_true_div_cmp_a;
  operator_66_true_div_cmp_b <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(operator_66_true_div_cmp_b_9_0));
  operator_66_true_div_cmp_z <= operator_66_true_div_cmp_z_1;

  STAGE_LOOP_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_l_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 0,
      width_s => 4,
      width_z => 10
      )
    PORT MAP(
      a => STAGE_LOOP_lshift_rg_a,
      s => STAGE_LOOP_lshift_rg_s,
      z => STAGE_LOOP_lshift_rg_z
    );
  STAGE_LOOP_lshift_rg_a(0) <= '1';
  STAGE_LOOP_lshift_rg_s <= STAGE_LOOP_i_3_0_sva;
  STAGE_LOOP_lshift_psp_sva_mx0w0 <= STAGE_LOOP_lshift_rg_z;

  inPlaceNTT_DIT_core_core_fsm_inst : inPlaceNTT_DIT_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      fsm_output => inPlaceNTT_DIT_core_core_fsm_inst_fsm_output,
      STAGE_LOOP_C_8_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0,
      modExp_while_C_38_tr0 => COMP_LOOP_COMP_LOOP_and_11_itm,
      COMP_LOOP_C_1_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0,
      COMP_LOOP_1_modExp_1_while_C_38_tr0 => COMP_LOOP_COMP_LOOP_and_11_itm,
      COMP_LOOP_C_62_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_62_tr0,
      COMP_LOOP_2_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_124_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_124_tr0,
      COMP_LOOP_3_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_186_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_186_tr0,
      COMP_LOOP_4_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_248_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_248_tr0,
      COMP_LOOP_5_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_310_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_310_tr0,
      COMP_LOOP_6_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_372_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_372_tr0,
      COMP_LOOP_7_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_434_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_434_tr0,
      COMP_LOOP_8_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_496_tr0 => COMP_LOOP_COMP_LOOP_and_145_itm,
      VEC_LOOP_C_0_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0,
      STAGE_LOOP_C_9_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0
    );
  fsm_output <= inPlaceNTT_DIT_core_core_fsm_inst_fsm_output;
  inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0 <= NOT (z_out_3(64));
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_62_tr0 <= NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_124_tr0 <= NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_186_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_248_tr0 <= NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_310_tr0 <= NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_372_tr0 <= NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_434_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 <= z_out_3(12);
  inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0 <= NOT STAGE_LOOP_acc_itm_2_1;

  nand_190_cse <= NOT((fsm_output(3)) AND (fsm_output(2)) AND (fsm_output(6)) AND
      (fsm_output(7)));
  and_416_cse <= (fsm_output(5)) AND (fsm_output(4)) AND (fsm_output(6)) AND (NOT
      (fsm_output(8)));
  nand_168_cse <= NOT((fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(7)));
  and_389_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  or_838_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"));
  or_1391_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"));
  nor_425_cse <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")));
  or_817_cse <= (NOT (fsm_output(5))) OR (fsm_output(3));
  or_816_cse <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("01"));
  or_1392_cse <= (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(9));
  and_382_cse <= or_838_cse AND (fsm_output(2));
  or_1394_cse <= and_389_cse OR (fsm_output(2));
  or_1099_cse <= (fsm_output(6)) OR (fsm_output(9));
  or_1113_nl <= (fsm_output(5)) OR (NOT (fsm_output(0))) OR (fsm_output(9)) OR not_tmp_462;
  or_1111_nl <= (fsm_output(0)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(7)))
      OR (fsm_output(3)) OR (NOT (fsm_output(4)));
  or_1109_nl <= (NOT (fsm_output(0))) OR (fsm_output(9)) OR (fsm_output(7)) OR (fsm_output(3))
      OR (NOT (fsm_output(4)));
  mux_1119_nl <= MUX_s_1_2_2(or_1111_nl, or_1109_nl, fsm_output(5));
  mux_1120_nl <= MUX_s_1_2_2(or_1113_nl, mux_1119_nl, fsm_output(1));
  nor_340_nl <= NOT((fsm_output(6)) OR mux_1120_nl);
  nor_341_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(0)))
      OR (NOT (fsm_output(9))) OR (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(4)));
  nor_342_nl <= NOT((fsm_output(9)) OR not_tmp_462);
  and_492_nl <= (fsm_output(9)) AND (fsm_output(7)) AND (NOT (fsm_output(3))) AND
      (fsm_output(4));
  mux_1117_nl <= MUX_s_1_2_2(nor_342_nl, and_492_nl, fsm_output(0));
  and_324_nl <= (fsm_output(1)) AND (fsm_output(5)) AND mux_1117_nl;
  mux_1118_nl <= MUX_s_1_2_2(nor_341_nl, and_324_nl, fsm_output(6));
  mux_1121_nl <= MUX_s_1_2_2(nor_340_nl, mux_1118_nl, fsm_output(2));
  nor_344_nl <= NOT((fsm_output(5)) OR (fsm_output(0)) OR (fsm_output(9)) OR (NOT
      (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(4)));
  nor_345_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(0))) OR (fsm_output(9))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(4)));
  mux_1116_nl <= MUX_s_1_2_2(nor_344_nl, nor_345_nl, fsm_output(1));
  and_325_nl <= (NOT((fsm_output(2)) OR (NOT (fsm_output(6))))) AND mux_1116_nl;
  mux_1122_nl <= MUX_s_1_2_2(mux_1121_nl, and_325_nl, fsm_output(8));
  modExp_while_if_or_nl <= and_dcpl_147 OR (mux_1122_nl AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  modExp_while_if_and_1_nl <= modExp_while_and_3 AND not_tmp_414;
  modExp_while_if_and_2_nl <= modExp_while_and_5 AND not_tmp_414;
  modExp_while_if_mux1h_nl <= MUX1HOT_v_64_5_2(z_out_4, STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000001"),
      modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w1, COMP_LOOP_1_acc_5_mut_mx0w5,
      STD_LOGIC_VECTOR'( modExp_while_if_or_nl & not_tmp_374 & modExp_while_if_and_1_nl
      & modExp_while_if_and_2_nl & not_tmp_312));
  and_179_nl <= and_dcpl_51 AND and_dcpl_58 AND and_dcpl_48;
  mux_851_nl <= MUX_s_1_2_2(or_tmp_113, nor_tmp_23, fsm_output(5));
  mux_852_nl <= MUX_s_1_2_2(mux_851_nl, or_247_cse, fsm_output(6));
  mux_849_nl <= MUX_s_1_2_2((NOT nor_tmp), or_tmp_788, fsm_output(5));
  mux_850_nl <= MUX_s_1_2_2(mux_tmp_677, mux_849_nl, fsm_output(6));
  mux_853_nl <= MUX_s_1_2_2(mux_852_nl, mux_850_nl, fsm_output(2));
  or_1388_nl <= (fsm_output(5)) OR mux_tmp_845;
  mux_846_nl <= MUX_s_1_2_2(mux_tmp_845, (NOT or_216_cse), fsm_output(5));
  mux_847_nl <= MUX_s_1_2_2(or_1388_nl, mux_846_nl, fsm_output(6));
  or_928_nl <= (fsm_output(5)) OR and_462_cse;
  mux_843_nl <= MUX_s_1_2_2((fsm_output(4)), mux_342_cse, fsm_output(5));
  mux_844_nl <= MUX_s_1_2_2(or_928_nl, mux_843_nl, fsm_output(6));
  mux_848_nl <= MUX_s_1_2_2(mux_847_nl, mux_844_nl, fsm_output(2));
  mux_854_nl <= MUX_s_1_2_2(mux_853_nl, mux_848_nl, fsm_output(7));
  and_372_nl <= (fsm_output(5)) AND (NOT mux_tmp_719);
  mux_839_nl <= MUX_s_1_2_2(or_tmp_788, (NOT or_tmp_891), fsm_output(5));
  mux_840_nl <= MUX_s_1_2_2(and_372_nl, mux_839_nl, fsm_output(6));
  and_373_nl <= (fsm_output(5)) AND (NOT mux_342_cse);
  nor_397_nl <= NOT((fsm_output(5)) OR and_dcpl_50);
  mux_838_nl <= MUX_s_1_2_2(and_373_nl, nor_397_nl, fsm_output(6));
  mux_841_nl <= MUX_s_1_2_2(mux_840_nl, mux_838_nl, fsm_output(2));
  or_925_nl <= ((NOT (fsm_output(5))) AND (fsm_output(0)) AND (fsm_output(1)) AND
      (fsm_output(3))) OR (fsm_output(4));
  mux_835_nl <= MUX_s_1_2_2(or_925_nl, mux_tmp_722, fsm_output(6));
  mux_833_nl <= MUX_s_1_2_2((NOT mux_tmp_688), (fsm_output(4)), fsm_output(5));
  mux_834_nl <= MUX_s_1_2_2(mux_833_nl, mux_tmp_718, fsm_output(6));
  mux_836_nl <= MUX_s_1_2_2(mux_835_nl, mux_834_nl, fsm_output(2));
  mux_842_nl <= MUX_s_1_2_2(mux_841_nl, mux_836_nl, fsm_output(7));
  mux_855_nl <= MUX_s_1_2_2((NOT mux_854_nl), mux_842_nl, fsm_output(8));
  mux_828_nl <= MUX_s_1_2_2(mux_331_cse, (NOT or_tmp_788), fsm_output(5));
  mux_826_nl <= MUX_s_1_2_2(nor_tmp, mux_tmp_688, fsm_output(5));
  mux_829_nl <= MUX_s_1_2_2(mux_828_nl, mux_826_nl, fsm_output(6));
  mux_824_nl <= MUX_s_1_2_2(and_705_cse, (NOT or_216_cse), fsm_output(5));
  mux_823_nl <= MUX_s_1_2_2(and_705_cse, mux_tmp_156, fsm_output(5));
  mux_825_nl <= MUX_s_1_2_2(mux_824_nl, mux_823_nl, fsm_output(6));
  mux_830_nl <= MUX_s_1_2_2(mux_829_nl, mux_825_nl, fsm_output(2));
  mux_820_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), and_dcpl_59, fsm_output(5));
  mux_821_nl <= MUX_s_1_2_2(mux_820_nl, (NOT nor_tmp_146), fsm_output(6));
  mux_818_nl <= MUX_s_1_2_2(mux_tmp_689, (NOT and_705_cse), fsm_output(5));
  mux_819_nl <= MUX_s_1_2_2(mux_tmp_705, mux_818_nl, fsm_output(6));
  mux_822_nl <= MUX_s_1_2_2(mux_821_nl, mux_819_nl, fsm_output(2));
  mux_831_nl <= MUX_s_1_2_2(mux_830_nl, mux_822_nl, fsm_output(7));
  and_376_nl <= (fsm_output(5)) AND (NOT nor_tmp_23);
  mux_816_nl <= MUX_s_1_2_2(and_376_nl, or_1202_cse, fsm_output(6));
  mux_815_nl <= MUX_s_1_2_2(and_428_cse, (NOT (fsm_output(4))), fsm_output(5));
  or_923_nl <= (fsm_output(6)) OR mux_815_nl;
  mux_817_nl <= MUX_s_1_2_2(mux_816_nl, or_923_nl, fsm_output(2));
  or_924_nl <= (fsm_output(7)) OR mux_817_nl;
  mux_832_nl <= MUX_s_1_2_2(mux_831_nl, or_924_nl, fsm_output(8));
  mux_856_nl <= MUX_s_1_2_2(mux_855_nl, mux_832_nl, fsm_output(9));
  operator_64_false_mux1h_2_rgt <= MUX1HOT_v_65_3_2(z_out_2, (STD_LOGIC_VECTOR'(
      "00") & operator_64_false_slc_modExp_exp_63_1_3), ('0' & modExp_while_if_mux1h_nl),
      STD_LOGIC_VECTOR'( and_179_nl & and_dcpl_156 & (NOT mux_856_nl)));
  and_705_cse <= (fsm_output(4)) AND or_136_cse;
  or_1385_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  nor_393_cse <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("00")));
  and_369_cse <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)=STD_LOGIC_VECTOR'("11"));
  and_187_m1c <= and_dcpl_137 AND and_dcpl_89 AND nor_393_cse;
  and_491_cse <= (fsm_output(6)) AND or_tmp;
  modExp_result_and_rgt <= (NOT modExp_while_and_5) AND and_187_m1c;
  modExp_result_and_1_rgt <= modExp_while_and_5 AND and_187_m1c;
  and_477_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"));
  and_483_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"));
  or_1423_cse <= and_477_cse OR (fsm_output(9));
  or_245_cse <= (fsm_output(1)) OR (fsm_output(3));
  or_247_cse <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10"));
  modulo_result_mux_1_cse <= MUX_v_64_2_2(modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w1,
      modulo_result_rem_cmp_z(63));
  and_428_cse <= (fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(3)) AND (fsm_output(4));
  or_242_cse <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(3)) OR (NOT (fsm_output(4)));
  or_42_nl <= (fsm_output(6)) OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  or_41_nl <= (NOT (fsm_output(6))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (fsm_output(4)) OR (NOT (fsm_output(8)));
  mux_33_nl <= MUX_s_1_2_2(or_42_nl, or_41_nl, fsm_output(1));
  or_39_nl <= (NOT (fsm_output(1))) OR (fsm_output(6)) OR (NOT (fsm_output(2))) OR
      (NOT (fsm_output(7))) OR (fsm_output(9)) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_34_nl <= MUX_s_1_2_2(mux_33_nl, or_39_nl, fsm_output(0));
  nor_601_cse <= NOT((fsm_output(3)) OR mux_34_nl);
  nor_604_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(2)))
      OR (NOT (fsm_output(7))) OR (fsm_output(9)) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  nor_605_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(6)) OR (fsm_output(2)) OR
      (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_29_cse <= MUX_s_1_2_2(nor_604_nl, nor_605_nl, fsm_output(0));
  mux_331_cse <= MUX_s_1_2_2(mux_tmp_156, nor_tmp, and_389_cse);
  mux_342_cse <= MUX_s_1_2_2(mux_tmp_156, nor_tmp, fsm_output(1));
  and_25_cse <= (fsm_output(5)) AND nor_tmp_23;
  nor_386_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(0)) OR (fsm_output(3)));
  nor_387_nl <= NOT((fsm_output(5)) OR (NOT((fsm_output(0)) AND (fsm_output(3)))));
  mux_915_nl <= MUX_s_1_2_2(nor_386_nl, nor_387_nl, fsm_output(6));
  and_243_m1c <= mux_915_nl AND (fsm_output(4)) AND (NOT (fsm_output(1))) AND (NOT
      (fsm_output(2))) AND (NOT (fsm_output(7))) AND nor_393_cse;
  and_462_cse <= (and_389_cse OR (fsm_output(3))) AND (fsm_output(4));
  or_115_cse <= (or_838_cse AND (fsm_output(3))) OR (fsm_output(4));
  and_502_cse <= (fsm_output(6)) AND (fsm_output(3)) AND (fsm_output(7)) AND (fsm_output(2))
      AND (fsm_output(8)) AND (NOT (fsm_output(9))) AND (NOT (fsm_output(4)));
  COMP_LOOP_COMP_LOOP_and_11_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)=STD_LOGIC_VECTOR'("101"));
  modExp_while_or_cse <= and_dcpl_84 OR and_dcpl_93 OR and_dcpl_103 OR and_dcpl_112
      OR and_dcpl_123 OR and_dcpl_130 OR and_dcpl_138;
  COMP_LOOP_COMP_LOOP_and_37_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)=STD_LOGIC_VECTOR'("011"));
  nand_100_cse <= NOT((fsm_output(8)) AND (fsm_output(4)));
  or_1189_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"));
  and_316_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"));
  and_314_cse <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"));
  and_437_cse <= (fsm_output(0)) AND (fsm_output(4));
  or_171_cse <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00"));
  or_210_cse <= (fsm_output(4)) OR (NOT (fsm_output(8)));
  or_216_cse <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"));
  or_1202_cse <= CONV_SL_1_1(fsm_output(5 DOWNTO 3)/=STD_LOGIC_VECTOR'("000"));
  nand_97_cse <= NOT((fsm_output(6)) AND (fsm_output(8)));
  nand_230_cse <= NOT((fsm_output(9)) AND (fsm_output(4)));
  nand_89_cse <= NOT((fsm_output(9)) AND (fsm_output(8)) AND (fsm_output(4)));
  COMP_LOOP_or_2_cse <= and_dcpl_69 OR and_dcpl_84 OR and_dcpl_93 OR and_dcpl_103
      OR and_dcpl_112 OR and_dcpl_123 OR and_dcpl_130 OR and_dcpl_138;
  COMP_LOOP_COMP_LOOP_and_12_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)=STD_LOGIC_VECTOR'("110"));
  COMP_LOOP_COMP_LOOP_and_13_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111"));
  STAGE_LOOP_i_3_0_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_LOOP_i_3_0_sva)
      + UNSIGNED'( "0001"), 4));
  COMP_LOOP_acc_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0(11
      DOWNTO 3)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_3_sva_5_0),
      6), 9), 9));
  modulo_qr_sva_1_mx0w1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_result_rem_cmp_z)
      + UNSIGNED(p_sva), 64));
  COMP_LOOP_1_acc_5_mut_mx0w5 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_10_lpi_4_dfm)
      + SIGNED(modulo_result_mux_1_cse), 64));
  operator_64_false_slc_modExp_exp_63_1_3 <= MUX_v_63_2_2((operator_66_true_div_cmp_z(63
      DOWNTO 1)), (tmp_10_lpi_4_dfm(63 DOWNTO 1)), and_dcpl_162);
  COMP_LOOP_acc_1_cse_2_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_3_sva_5_0 & STD_LOGIC_VECTOR'(
      "001")), 9), 12), 12));
  COMP_LOOP_acc_1_cse_6_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_3_sva_5_0 & STD_LOGIC_VECTOR'(
      "101")), 9), 12), 12));
  COMP_LOOP_acc_1_cse_4_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_3_sva_5_0 & STD_LOGIC_VECTOR'(
      "011")), 9), 12), 12));
  COMP_LOOP_k_9_3_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_3_sva_5_0),
      6), 7) + UNSIGNED'( "0000001"), 7));
  modExp_while_and_3 <= (NOT (modulo_result_rem_cmp_z(63))) AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  modExp_while_and_5 <= (modulo_result_rem_cmp_z(63)) AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  COMP_LOOP_COMP_LOOP_and_211 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO
      0)=STD_LOGIC_VECTOR'("001"));
  COMP_LOOP_COMP_LOOP_and_213 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO
      0)=STD_LOGIC_VECTOR'("010"));
  COMP_LOOP_COMP_LOOP_and_215 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO
      0)=STD_LOGIC_VECTOR'("100"));
  nor_tmp <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11"));
  or_tmp <= (fsm_output(5)) OR nor_tmp;
  or_81_cse <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("01"));
  or_83_cse <= (fsm_output(4)) OR (fsm_output(9));
  or_tmp_92 <= NOT((fsm_output(0)) AND (fsm_output(1)) AND (NOT (fsm_output(3)))
      AND (fsm_output(4)));
  or_136_cse <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(3));
  nor_tmp_23 <= or_245_cse AND (fsm_output(4));
  or_tmp_103 <= and_389_cse OR CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"));
  nor_tmp_27 <= or_838_cse AND CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11"));
  mux_tmp_156 <= MUX_s_1_2_2((NOT (fsm_output(4))), (fsm_output(4)), fsm_output(3));
  or_tmp_113 <= ((fsm_output(1)) AND (fsm_output(3))) OR (fsm_output(4));
  and_dcpl_4 <= (fsm_output(0)) AND (fsm_output(5));
  or_tmp_154 <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  and_dcpl_11 <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_14 <= NOT((fsm_output(0)) OR (fsm_output(5)));
  and_dcpl_23 <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)=STD_LOGIC_VECTOR'("10"));
  or_1402_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000000"));
  and_432_nl <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("11"));
  mux_361_nl <= MUX_s_1_2_2(and_432_nl, and_491_cse, fsm_output(2));
  nand_199_nl <= NOT((fsm_output(8)) AND ((fsm_output(7)) OR mux_361_nl));
  not_tmp_131 <= MUX_s_1_2_2(or_1402_nl, nand_199_nl, fsm_output(9));
  and_dcpl_46 <= NOT((fsm_output(6)) OR (fsm_output(2)));
  and_dcpl_47 <= and_dcpl_46 AND (NOT (fsm_output(7)));
  and_dcpl_48 <= and_dcpl_47 AND nor_393_cse;
  and_dcpl_50 <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_51 <= and_dcpl_50 AND (NOT (fsm_output(1)));
  and_dcpl_56 <= (fsm_output(6)) AND (NOT (fsm_output(2))) AND (NOT (fsm_output(7)));
  and_dcpl_57 <= and_dcpl_56 AND and_369_cse;
  and_dcpl_58 <= (fsm_output(0)) AND (NOT (fsm_output(5)));
  and_dcpl_59 <= nor_tmp AND (fsm_output(1));
  and_dcpl_60 <= and_dcpl_59 AND and_dcpl_58;
  and_dcpl_63 <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_64 <= and_dcpl_63 AND (NOT (fsm_output(1)));
  and_dcpl_65 <= and_dcpl_64 AND and_dcpl_4;
  and_dcpl_66 <= and_dcpl_65 AND and_dcpl_48;
  and_dcpl_67 <= and_dcpl_56 AND nor_393_cse;
  and_dcpl_68 <= and_dcpl_59 AND and_dcpl_14;
  and_dcpl_69 <= and_dcpl_68 AND and_dcpl_67;
  and_dcpl_70 <= and_dcpl_46 AND (fsm_output(7));
  and_dcpl_73 <= and_dcpl_50 AND (fsm_output(1)) AND and_dcpl_14;
  and_dcpl_80 <= (NOT (fsm_output(6))) AND (fsm_output(2));
  and_dcpl_82 <= and_dcpl_80 AND (fsm_output(7)) AND nor_393_cse;
  and_dcpl_84 <= and_dcpl_59 AND and_dcpl_4 AND and_dcpl_82;
  and_dcpl_89 <= and_dcpl_80 AND (NOT (fsm_output(7)));
  and_dcpl_91 <= (NOT (fsm_output(0))) AND (fsm_output(5));
  and_dcpl_93 <= and_dcpl_51 AND and_dcpl_91 AND and_dcpl_89 AND and_dcpl_11;
  and_dcpl_100 <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_102 <= and_dcpl_100 AND (NOT (fsm_output(1))) AND and_dcpl_58;
  and_dcpl_103 <= and_dcpl_102 AND and_dcpl_70 AND and_dcpl_11;
  and_dcpl_108 <= (fsm_output(6)) AND (fsm_output(2)) AND (fsm_output(7));
  and_dcpl_109 <= and_dcpl_108 AND and_dcpl_11;
  and_dcpl_110 <= and_dcpl_100 AND (fsm_output(1));
  and_dcpl_112 <= and_dcpl_110 AND and_dcpl_91 AND and_dcpl_109;
  and_dcpl_121 <= and_dcpl_63 AND (fsm_output(1));
  and_dcpl_122 <= and_dcpl_121 AND and_dcpl_58;
  and_dcpl_123 <= and_dcpl_122 AND and_dcpl_56 AND and_dcpl_23;
  and_dcpl_127 <= and_dcpl_70 AND and_dcpl_23;
  and_dcpl_128 <= nor_tmp AND (NOT (fsm_output(1)));
  and_dcpl_129 <= and_dcpl_128 AND and_dcpl_91;
  and_dcpl_130 <= and_dcpl_129 AND and_dcpl_127;
  and_dcpl_137 <= and_dcpl_128 AND and_dcpl_58;
  and_dcpl_138 <= and_dcpl_137 AND and_dcpl_89 AND and_369_cse;
  nand_194_cse <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11")));
  or_tmp_268 <= (NOT (fsm_output(4))) OR (fsm_output(9)) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR nand_194_cse;
  or_308_nl <= (fsm_output(4)) OR (VEC_LOOP_j_sva_11_0(0)) OR (VEC_LOOP_j_sva_11_0(2))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00100"));
  or_306_nl <= (NOT (fsm_output(4))) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (COMP_LOOP_acc_13_psp_sva(0)) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("000"));
  mux_381_nl <= MUX_s_1_2_2(or_308_nl, or_306_nl, fsm_output(2));
  or_tmp_273 <= (VEC_LOOP_j_sva_11_0(1)) OR mux_381_nl;
  or_329_cse <= CONV_SL_1_1(fsm_output(9 DOWNTO 4)/=STD_LOGIC_VECTOR'("011100"));
  or_327_cse <= CONV_SL_1_1(fsm_output(9 DOWNTO 4)/=STD_LOGIC_VECTOR'("110101"));
  or_325_nl <= CONV_SL_1_1(fsm_output(9 DOWNTO 4)/=STD_LOGIC_VECTOR'("001111"));
  or_323_nl <= CONV_SL_1_1(fsm_output(9 DOWNTO 4)/=STD_LOGIC_VECTOR'("101000"));
  mux_392_cse <= MUX_s_1_2_2(or_325_nl, or_323_nl, fsm_output(2));
  or_320_cse <= CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00100"));
  nand_246_cse <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 4)=STD_LOGIC_VECTOR'("101111")));
  or_314_cse <= (fsm_output(2)) OR (fsm_output(4)) OR (NOT (fsm_output(9))) OR (NOT
      (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(8)) OR (fsm_output(7));
  or_312_cse <= CONV_SL_1_1(fsm_output(9 DOWNTO 4)/=STD_LOGIC_VECTOR'("010101"));
  not_tmp_165 <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11")));
  nand_189_cse <= NOT((COMP_LOOP_acc_1_cse_4_sva(0)) AND CONV_SL_1_1(fsm_output(8
      DOWNTO 7)=STD_LOGIC_VECTOR'("11")));
  or_tmp_335 <= (NOT (fsm_output(4))) OR (fsm_output(9)) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))
      OR nand_189_cse;
  or_375_nl <= (fsm_output(4)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (VEC_LOOP_j_sva_11_0(2))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00100"));
  or_373_nl <= (NOT (fsm_output(4))) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (COMP_LOOP_acc_13_psp_sva(0)) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("000"));
  mux_418_nl <= MUX_s_1_2_2(or_375_nl, or_373_nl, fsm_output(2));
  or_tmp_340 <= (VEC_LOOP_j_sva_11_0(1)) OR mux_418_nl;
  or_tmp_395 <= (NOT (fsm_output(4))) OR (fsm_output(9)) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR nand_194_cse;
  nor_512_nl <= NOT((fsm_output(4)) OR (VEC_LOOP_j_sva_11_0(0)) OR (VEC_LOOP_j_sva_11_0(2))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00100")));
  nor_513_nl <= NOT((NOT (fsm_output(4))) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (COMP_LOOP_acc_13_psp_sva(0)) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_456_nl <= MUX_s_1_2_2(nor_512_nl, nor_513_nl, fsm_output(2));
  nand_tmp_18 <= NOT((VEC_LOOP_j_sva_11_0(1)) AND mux_456_nl);
  or_tmp_454 <= (NOT (fsm_output(4))) OR (fsm_output(9)) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR (COMP_LOOP_acc_1_cse_4_sva(2)) OR (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11"))));
  nor_496_nl <= NOT((fsm_output(4)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (VEC_LOOP_j_sva_11_0(2))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00100")));
  nor_497_nl <= NOT((NOT (fsm_output(4))) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT
      (fsm_output(9))) OR (fsm_output(5)) OR (COMP_LOOP_acc_13_psp_sva(0)) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_494_nl <= MUX_s_1_2_2(nor_496_nl, nor_497_nl, fsm_output(2));
  nand_tmp_21 <= NOT((VEC_LOOP_j_sva_11_0(1)) AND mux_494_nl);
  or_tmp_525 <= (NOT (fsm_output(4))) OR (fsm_output(9)) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR nand_194_cse;
  or_570_nl <= (fsm_output(4)) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (VEC_LOOP_j_sva_11_0(2)))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00100"));
  or_568_nl <= (NOT (fsm_output(4))) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (NOT (COMP_LOOP_acc_13_psp_sva(0))) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("000"));
  mux_538_nl <= MUX_s_1_2_2(or_570_nl, or_568_nl, fsm_output(2));
  or_tmp_535 <= (VEC_LOOP_j_sva_11_0(1)) OR mux_538_nl;
  or_tmp_590 <= (NOT (fsm_output(4))) OR (fsm_output(9)) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("10"))
      OR nand_189_cse;
  or_635_nl <= (fsm_output(4)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (VEC_LOOP_j_sva_11_0(2)))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00100"));
  or_633_nl <= (NOT (fsm_output(4))) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (NOT (COMP_LOOP_acc_13_psp_sva(0))) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("000"));
  mux_575_nl <= MUX_s_1_2_2(or_635_nl, or_633_nl, fsm_output(2));
  or_tmp_600 <= (VEC_LOOP_j_sva_11_0(1)) OR mux_575_nl;
  or_tmp_655 <= (NOT (fsm_output(4))) OR (fsm_output(9)) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR nand_194_cse;
  nor_458_nl <= NOT((fsm_output(4)) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (VEC_LOOP_j_sva_11_0(2)))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00100")));
  nor_459_nl <= NOT((NOT (fsm_output(4))) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (NOT (COMP_LOOP_acc_13_psp_sva(0))) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_612_nl <= MUX_s_1_2_2(nor_458_nl, nor_459_nl, fsm_output(2));
  nand_tmp_31 <= NOT((VEC_LOOP_j_sva_11_0(1)) AND mux_612_nl);
  or_tmp_719 <= (NOT (fsm_output(4))) OR (fsm_output(9)) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11"))));
  nor_444_nl <= NOT((fsm_output(4)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (VEC_LOOP_j_sva_11_0(2)))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00100")));
  nor_445_nl <= NOT((NOT (fsm_output(4))) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT
      (fsm_output(9))) OR (fsm_output(5)) OR (NOT (COMP_LOOP_acc_13_psp_sva(0)))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_649_nl <= MUX_s_1_2_2(nor_444_nl, nor_445_nl, fsm_output(2));
  nand_tmp_35 <= NOT((VEC_LOOP_j_sva_11_0(1)) AND mux_649_nl);
  and_dcpl_140 <= NOT((fsm_output(2)) OR (fsm_output(7)));
  and_dcpl_147 <= and_dcpl_110 AND and_dcpl_14 AND and_dcpl_48;
  mux_tmp_677 <= MUX_s_1_2_2((NOT mux_tmp_156), (fsm_output(4)), fsm_output(5));
  mux_tmp_688 <= MUX_s_1_2_2(and_dcpl_50, mux_tmp_156, fsm_output(1));
  mux_tmp_689 <= MUX_s_1_2_2((NOT or_tmp_113), mux_tmp_688, fsm_output(0));
  mux_696_itm <= MUX_s_1_2_2(and_dcpl_50, mux_tmp_156, and_389_cse);
  nor_tmp_146 <= or_817_cse AND (fsm_output(4));
  mux_tmp_705 <= MUX_s_1_2_2((NOT (fsm_output(4))), nor_tmp, fsm_output(5));
  or_tmp_788 <= ((fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(3))) OR (fsm_output(4));
  mux_tmp_718 <= MUX_s_1_2_2(and_dcpl_51, (fsm_output(4)), fsm_output(5));
  mux_tmp_719 <= MUX_s_1_2_2(and_dcpl_50, mux_tmp_156, or_838_cse);
  mux_tmp_722 <= MUX_s_1_2_2(and_dcpl_50, (fsm_output(4)), fsm_output(5));
  or_tmp_792 <= (fsm_output(6)) OR (NOT or_1385_cse);
  nand_tmp_42 <= NOT((fsm_output(6)) AND (NOT and_382_cse));
  mux_tmp_731 <= MUX_s_1_2_2((NOT (fsm_output(6))), (fsm_output(6)), fsm_output(5));
  not_tmp_274 <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111")));
  not_tmp_280 <= NOT((fsm_output(6)) OR (NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")))));
  or_tmp_810 <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("10"));
  or_854_nl <= (NOT (fsm_output(0))) OR (fsm_output(5)) OR (fsm_output(2)) OR (NOT
      (fsm_output(7))) OR (fsm_output(4));
  or_853_nl <= (NOT (fsm_output(0))) OR (fsm_output(5)) OR (NOT (fsm_output(2)))
      OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_tmp_776 <= MUX_s_1_2_2(or_854_nl, or_853_nl, fsm_output(9));
  not_tmp_297 <= NOT((fsm_output(7)) AND (fsm_output(4)));
  not_tmp_309 <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11")));
  or_903_nl <= (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(1)))
      OR (NOT (fsm_output(9))) OR (fsm_output(3)) OR (fsm_output(4));
  or_902_nl <= (NOT (fsm_output(5))) OR (fsm_output(0)) OR (fsm_output(1)) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(3))) OR (fsm_output(4));
  mux_800_nl <= MUX_s_1_2_2(or_903_nl, or_902_nl, fsm_output(6));
  and_489_nl <= (fsm_output(1)) AND (fsm_output(9)) AND (NOT (fsm_output(3))) AND
      (fsm_output(4));
  nor_407_nl <= NOT((fsm_output(1)) OR (fsm_output(9)) OR not_tmp_309);
  mux_799_nl <= MUX_s_1_2_2(and_489_nl, nor_407_nl, fsm_output(0));
  nand_49_nl <= NOT(nor_425_cse AND mux_799_nl);
  mux_801_nl <= MUX_s_1_2_2(mux_800_nl, nand_49_nl, fsm_output(8));
  nor_405_nl <= NOT((fsm_output(7)) OR mux_801_nl);
  nor_408_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(1))) OR (fsm_output(9)) OR (NOT
      (fsm_output(3))) OR (fsm_output(4)));
  or_895_nl <= (fsm_output(1)) OR (fsm_output(9)) OR (fsm_output(3)) OR (NOT (fsm_output(4)));
  or_893_nl <= (fsm_output(1)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(3)))
      OR (fsm_output(4));
  mux_796_nl <= MUX_s_1_2_2(or_895_nl, or_893_nl, fsm_output(0));
  nor_409_nl <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("10"))
      OR mux_796_nl);
  nor_410_nl <= NOT((fsm_output(6)) OR (fsm_output(5)) OR (fsm_output(0)) OR (NOT
      (fsm_output(1))) OR (fsm_output(9)) OR not_tmp_309);
  mux_797_nl <= MUX_s_1_2_2(nor_409_nl, nor_410_nl, fsm_output(8));
  mux_798_nl <= MUX_s_1_2_2(nor_408_nl, mux_797_nl, fsm_output(7));
  not_tmp_312 <= MUX_s_1_2_2(nor_405_nl, mux_798_nl, fsm_output(2));
  or_1362_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(4))) OR (fsm_output(8));
  or_913_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(4)))
      OR (fsm_output(3)) OR (fsm_output(8));
  mux_806_nl <= MUX_s_1_2_2(or_1362_nl, or_913_nl, fsm_output(0));
  nor_400_nl <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00"))
      OR mux_806_nl);
  nor_401_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(0)) OR (fsm_output(7)) OR
      (NOT (fsm_output(9))) OR (fsm_output(4)) OR (NOT (fsm_output(3))) OR (fsm_output(8)));
  and_377_nl <= (fsm_output(5)) AND (fsm_output(0)) AND (fsm_output(7)) AND (NOT
      (fsm_output(9))) AND (fsm_output(4)) AND (fsm_output(3)) AND (NOT (fsm_output(8)));
  mux_805_nl <= MUX_s_1_2_2(nor_401_nl, and_377_nl, fsm_output(6));
  mux_807_nl <= MUX_s_1_2_2(nor_400_nl, mux_805_nl, fsm_output(2));
  nor_402_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(5))) OR (fsm_output(0))
      OR (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(4)) OR (fsm_output(3))
      OR (NOT (fsm_output(8))));
  nor_403_nl <= NOT((NOT (fsm_output(0))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (fsm_output(4)) OR (fsm_output(3)) OR (NOT (fsm_output(8))));
  nor_404_nl <= NOT((fsm_output(0)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(4))) OR (fsm_output(3)) OR (fsm_output(8)));
  mux_803_nl <= MUX_s_1_2_2(nor_403_nl, nor_404_nl, fsm_output(5));
  and_378_nl <= (fsm_output(6)) AND mux_803_nl;
  mux_804_nl <= MUX_s_1_2_2(nor_402_nl, and_378_nl, fsm_output(2));
  not_tmp_315 <= MUX_s_1_2_2(mux_807_nl, mux_804_nl, fsm_output(1));
  mux_809_nl <= MUX_s_1_2_2((NOT (fsm_output(3))), (fsm_output(3)), fsm_output(1));
  or_916_nl <= (NOT (fsm_output(1))) OR (fsm_output(3));
  mux_810_nl <= MUX_s_1_2_2(mux_809_nl, or_916_nl, fsm_output(0));
  mux_811_nl <= MUX_s_1_2_2(mux_810_nl, (fsm_output(3)), fsm_output(2));
  and_dcpl_152 <= NOT(mux_811_nl OR CONV_SL_1_1(fsm_output(7 DOWNTO 4)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT nor_393_cse));
  nor_398_nl <= NOT((NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(4)));
  nor_399_nl <= NOT((fsm_output(0)) OR (fsm_output(3)) OR (NOT (fsm_output(4))));
  mux_814_nl <= MUX_s_1_2_2(nor_398_nl, nor_399_nl, fsm_output(5));
  and_dcpl_156 <= mux_814_nl AND (NOT (fsm_output(1))) AND and_dcpl_48;
  or_tmp_891 <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(4));
  mux_tmp_845 <= MUX_s_1_2_2(mux_tmp_156, nor_tmp, or_838_cse);
  not_tmp_347 <= NOT((fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(8)) OR (fsm_output(9)));
  and_361_cse <= (fsm_output(6)) AND (fsm_output(8)) AND (fsm_output(9));
  and_dcpl_162 <= and_dcpl_64 AND and_dcpl_91 AND and_dcpl_48;
  or_tmp_916 <= (fsm_output(6)) OR and_314_cse;
  or_955_nl <= (fsm_output(6)) OR and_25_cse;
  mux_tmp_886 <= MUX_s_1_2_2(or_955_nl, or_tmp_916, fsm_output(2));
  or_tmp_918 <= (fsm_output(7)) OR mux_tmp_886;
  and_tmp_28 <= (fsm_output(5)) AND or_216_cse;
  and_dcpl_164 <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 7)/=STD_LOGIC_VECTOR'("000")));
  and_dcpl_167 <= NOT(CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(2)) OR (NOT and_dcpl_164));
  and_dcpl_168 <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_171 <= and_dcpl_63 AND CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_172 <= and_dcpl_171 AND and_dcpl_168 AND (NOT (VEC_LOOP_j_sva_11_0(2)));
  and_dcpl_176 <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND (NOT (fsm_output(2))) AND and_dcpl_164;
  and_dcpl_180 <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND (NOT (fsm_output(2))) AND and_dcpl_164;
  and_dcpl_184 <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (NOT (fsm_output(2))) AND and_dcpl_164;
  and_dcpl_187 <= and_dcpl_171 AND and_dcpl_168 AND (VEC_LOOP_j_sva_11_0(2));
  nor_382_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(6)) OR (fsm_output(2)) OR
      (fsm_output(7)) OR (fsm_output(9)) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  nor_603_nl <= NOT((fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(4)) OR (NOT
      (fsm_output(8))));
  and_475_nl <= (fsm_output(7)) AND (fsm_output(9)) AND (fsm_output(4)) AND (NOT
      (fsm_output(8)));
  mux_30_nl <= MUX_s_1_2_2(nor_603_nl, and_475_nl, fsm_output(2));
  and_474_nl <= (NOT((fsm_output(1)) OR (NOT (fsm_output(6))))) AND mux_30_nl;
  mux_918_nl <= MUX_s_1_2_2(nor_382_nl, and_474_nl, fsm_output(0));
  mux_919_nl <= MUX_s_1_2_2(mux_918_nl, mux_29_cse, fsm_output(3));
  not_tmp_374 <= MUX_s_1_2_2(nor_601_cse, mux_919_nl, fsm_output(5));
  or_1026_nl <= (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(5)) OR nand_100_cse;
  or_1024_nl <= (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(5)))
      OR (fsm_output(8)) OR (fsm_output(4));
  mux_976_nl <= MUX_s_1_2_2(or_1026_nl, or_1024_nl, fsm_output(7));
  nor_366_nl <= NOT((fsm_output(3)) OR (fsm_output(1)) OR mux_976_nl);
  nor_367_nl <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(5)) OR nand_100_cse);
  mux_977_nl <= MUX_s_1_2_2(nor_366_nl, nor_367_nl, fsm_output(6));
  nor_368_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(2)) OR
      (fsm_output(5)) OR (NOT (fsm_output(8))) OR (fsm_output(4)));
  and_351_nl <= (fsm_output(9)) AND (fsm_output(2)) AND (fsm_output(5)) AND (NOT
      (fsm_output(8))) AND (fsm_output(4));
  nor_369_nl <= NOT((fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(5))) OR
      (fsm_output(8)) OR (fsm_output(4)));
  mux_973_nl <= MUX_s_1_2_2(and_351_nl, nor_369_nl, fsm_output(7));
  mux_974_nl <= MUX_s_1_2_2(nor_368_nl, mux_973_nl, fsm_output(1));
  and_350_nl <= (fsm_output(3)) AND mux_974_nl;
  nor_370_nl <= NOT((fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(7)) OR (fsm_output(9))
      OR (NOT((fsm_output(2)) AND (fsm_output(5)) AND (fsm_output(8)) AND (fsm_output(4)))));
  mux_975_nl <= MUX_s_1_2_2(and_350_nl, nor_370_nl, fsm_output(6));
  not_tmp_399 <= MUX_s_1_2_2(mux_977_nl, mux_975_nl, fsm_output(0));
  not_tmp_400 <= NOT((fsm_output(0)) AND (fsm_output(5)));
  not_tmp_406 <= NOT((fsm_output(7)) AND (fsm_output(2)) AND (fsm_output(6)));
  nor_357_cse <= NOT((NOT (fsm_output(1))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(8)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(2))) OR (fsm_output(9))
      OR (NOT (fsm_output(4))));
  and_345_nl <= (fsm_output(2)) AND (fsm_output(9)) AND (fsm_output(4));
  nor_355_nl <= NOT((fsm_output(2)) OR (fsm_output(9)) OR (fsm_output(4)));
  mux_991_nl <= MUX_s_1_2_2(and_345_nl, nor_355_nl, fsm_output(7));
  and_344_nl <= (NOT((NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(8)))))
      AND mux_991_nl;
  mux_990_nl <= MUX_s_1_2_2(nand_230_cse, or_83_cse, fsm_output(2));
  nor_356_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(8)) OR
      (fsm_output(7)) OR mux_990_nl);
  mux_992_nl <= MUX_s_1_2_2(and_344_nl, nor_356_nl, fsm_output(1));
  mux_993_nl <= MUX_s_1_2_2(mux_992_nl, nor_357_cse, fsm_output(5));
  nand_111_nl <= NOT((fsm_output(7)) AND (fsm_output(2)) AND (fsm_output(9)) AND
      (fsm_output(4)));
  or_1045_nl <= (fsm_output(7)) OR (fsm_output(2)) OR (fsm_output(9)) OR (fsm_output(4));
  mux_988_nl <= MUX_s_1_2_2(nand_111_nl, or_1045_nl, fsm_output(8));
  nor_358_nl <= NOT((fsm_output(3)) OR (fsm_output(6)) OR mux_988_nl);
  mux_989_nl <= MUX_s_1_2_2(and_502_cse, nor_358_nl, fsm_output(1));
  and_346_nl <= (fsm_output(5)) AND mux_989_nl;
  not_tmp_414 <= MUX_s_1_2_2(mux_993_nl, and_346_nl, fsm_output(0));
  mux_tmp_997 <= MUX_s_1_2_2((NOT (fsm_output(4))), (fsm_output(4)), fsm_output(5));
  mux_tmp_1006 <= MUX_s_1_2_2((fsm_output(5)), or_171_cse, or_1391_cse);
  not_tmp_436 <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("11")));
  not_tmp_462 <= NOT((fsm_output(7)) AND (fsm_output(3)) AND (fsm_output(4)));
  and_dcpl_219 <= and_dcpl_121 AND and_dcpl_4 AND and_dcpl_48;
  not_tmp_480 <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_886);
  and_320_nl <= CONV_SL_1_1(fsm_output(6 DOWNTO 3)=STD_LOGIC_VECTOR'("1111"));
  and_263_nl <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("11")) AND and_705_cse;
  mux_1157_nl <= MUX_s_1_2_2(and_320_nl, and_263_nl, fsm_output(2));
  or_1183_nl <= (fsm_output(8)) OR ((fsm_output(7)) AND mux_1157_nl);
  mux_1158_itm <= MUX_s_1_2_2(not_tmp_480, or_1183_nl, fsm_output(9));
  nor_tmp_240 <= (fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(9));
  mux_tmp_1159 <= MUX_s_1_2_2(nor_tmp_240, (fsm_output(9)), fsm_output(8));
  nor_tmp_241 <= ((fsm_output(5)) OR (fsm_output(7))) AND (fsm_output(9));
  mux_tmp_1160 <= MUX_s_1_2_2(nor_tmp_240, nor_tmp_241, fsm_output(8));
  and_tmp_44 <= (fsm_output(8)) AND nor_tmp_241;
  mux_1161_nl <= MUX_s_1_2_2(and_tmp_44, mux_tmp_1160, fsm_output(2));
  mux_tmp_1162 <= MUX_s_1_2_2(mux_1161_nl, mux_tmp_1159, fsm_output(3));
  not_tmp_482 <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (fsm_output(9)));
  nor_tmp_244 <= ((NOT (fsm_output(5))) OR (fsm_output(7))) AND (fsm_output(9));
  mux_tmp_1164 <= MUX_s_1_2_2(not_tmp_482, nor_tmp_244, fsm_output(8));
  nor_329_nl <= NOT((fsm_output(7)) OR (fsm_output(9)));
  mux_tmp_1170 <= MUX_s_1_2_2(nor_329_nl, nor_tmp_244, fsm_output(8));
  or_tmp_1144 <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000"));
  and_tmp_45 <= (fsm_output(9)) AND or_tmp_1144;
  and_tmp_46 <= (fsm_output(9)) AND or_tmp_154;
  mux_tmp_1178 <= MUX_s_1_2_2((NOT or_tmp_1144), or_tmp_154, fsm_output(9));
  or_tmp_1159 <= (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(4))) OR (fsm_output(6))
      OR (fsm_output(8));
  or_tmp_1165 <= (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_tmp_1202 <= MUX_s_1_2_2(or_210_cse, or_tmp_1165, fsm_output(9));
  or_tmp_1174 <= (fsm_output(9)) OR nand_100_cse;
  or_tmp_1176 <= (fsm_output(9)) OR (fsm_output(4)) OR (NOT (fsm_output(8)));
  and_dcpl_226 <= and_dcpl_121 AND and_dcpl_91 AND and_dcpl_48;
  or_1268_nl <= (NOT (fsm_output(9))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1268_nl <= MUX_s_1_2_2(mux_tmp_1202, or_1268_nl, and_389_cse);
  mux_1269_nl <= MUX_s_1_2_2(mux_1268_nl, or_tmp_1165, fsm_output(2));
  mux_1270_nl <= MUX_s_1_2_2((NOT (fsm_output(8))), mux_1269_nl, fsm_output(5));
  or_1267_nl <= (or_1391_cse AND (fsm_output(9)) AND (fsm_output(4))) OR (fsm_output(8));
  mux_1266_nl <= MUX_s_1_2_2(or_tmp_1174, or_81_cse, or_1391_cse);
  mux_1267_nl <= MUX_s_1_2_2(or_1267_nl, mux_1266_nl, fsm_output(5));
  mux_1271_nl <= MUX_s_1_2_2(mux_1270_nl, mux_1267_nl, fsm_output(6));
  mux_1263_nl <= MUX_s_1_2_2(or_tmp_1176, mux_tmp_1202, or_1385_cse);
  or_1263_nl <= ((fsm_output(2)) AND (fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(9))
      AND (fsm_output(4))) OR (fsm_output(8));
  mux_1264_nl <= MUX_s_1_2_2(mux_1263_nl, or_1263_nl, fsm_output(5));
  mux_1261_nl <= MUX_s_1_2_2(or_tmp_1174, or_81_cse, and_477_cse);
  mux_1260_nl <= MUX_s_1_2_2(or_tmp_1176, mux_tmp_1202, and_483_cse);
  mux_1262_nl <= MUX_s_1_2_2(mux_1261_nl, mux_1260_nl, fsm_output(5));
  mux_1265_nl <= MUX_s_1_2_2(mux_1264_nl, mux_1262_nl, fsm_output(6));
  mux_1272_nl <= MUX_s_1_2_2(mux_1271_nl, mux_1265_nl, fsm_output(7));
  nand_227_nl <= NOT((NOT((fsm_output(2)) AND (fsm_output(9)) AND (fsm_output(4))))
      AND (fsm_output(8)));
  or_1258_nl <= (NOT(((fsm_output(2)) AND (fsm_output(9))) OR (fsm_output(4)))) OR
      (fsm_output(8));
  mux_1257_nl <= MUX_s_1_2_2(nand_227_nl, or_1258_nl, fsm_output(5));
  or_1256_nl <= (or_1392_cse AND (fsm_output(4))) OR (fsm_output(8));
  mux_1256_nl <= MUX_s_1_2_2(or_1256_nl, or_81_cse, fsm_output(5));
  mux_1258_nl <= MUX_s_1_2_2(mux_1257_nl, mux_1256_nl, fsm_output(6));
  or_1254_nl <= ((and_483_cse OR (fsm_output(9))) AND (fsm_output(4))) OR (fsm_output(8));
  mux_1254_nl <= MUX_s_1_2_2(or_tmp_1165, or_1254_nl, fsm_output(5));
  or_1249_nl <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(9));
  mux_1250_nl <= MUX_s_1_2_2(or_210_cse, or_tmp_1165, or_1249_nl);
  mux_1252_nl <= MUX_s_1_2_2(mux_tmp_1202, mux_1250_nl, fsm_output(2));
  mux_1253_nl <= MUX_s_1_2_2(or_81_cse, mux_1252_nl, fsm_output(5));
  mux_1255_nl <= MUX_s_1_2_2(mux_1254_nl, mux_1253_nl, fsm_output(6));
  mux_1259_nl <= MUX_s_1_2_2(mux_1258_nl, mux_1255_nl, fsm_output(7));
  mux_1273_itm <= MUX_s_1_2_2(mux_1272_nl, mux_1259_nl, fsm_output(3));
  nor_310_nl <= NOT((fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (NOT
      (fsm_output(8))));
  and_295_nl <= (fsm_output(2)) AND (fsm_output(7)) AND (fsm_output(4)) AND (NOT
      (fsm_output(8)));
  mux_1275_nl <= MUX_s_1_2_2(nor_310_nl, and_295_nl, fsm_output(9));
  and_294_nl <= (NOT((NOT (fsm_output(0))) OR (fsm_output(1)) OR (NOT (fsm_output(6)))))
      AND mux_1275_nl;
  mux_1276_nl <= MUX_s_1_2_2(and_294_nl, mux_29_cse, fsm_output(3));
  not_tmp_513 <= MUX_s_1_2_2(nor_601_cse, mux_1276_nl, fsm_output(5));
  or_1304_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(8))) OR (fsm_output(9))
      OR (fsm_output(4));
  or_1303_nl <= (fsm_output(7)) OR nand_89_cse;
  mux_1289_nl <= MUX_s_1_2_2(or_1304_nl, or_1303_nl, fsm_output(2));
  nor_300_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(6)) OR mux_1289_nl);
  nor_628_nl <= NOT((NOT (fsm_output(6))) OR (fsm_output(3)) OR (fsm_output(7)) OR
      (fsm_output(2)) OR (fsm_output(8)) OR nand_230_cse);
  mux_1290_nl <= MUX_s_1_2_2(nor_300_nl, nor_628_nl, fsm_output(1));
  mux_1291_nl <= MUX_s_1_2_2(mux_1290_nl, nor_357_cse, fsm_output(5));
  or_1093_nl <= (fsm_output(9)) OR (NOT (fsm_output(4)));
  mux_1286_nl <= MUX_s_1_2_2(or_1093_nl, or_83_cse, fsm_output(8));
  or_1295_nl <= (fsm_output(7)) OR mux_1286_nl;
  or_1292_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01")) OR nand_230_cse;
  mux_1287_nl <= MUX_s_1_2_2(or_1295_nl, or_1292_nl, fsm_output(2));
  nor_303_nl <= NOT((fsm_output(3)) OR (fsm_output(6)) OR mux_1287_nl);
  mux_1288_nl <= MUX_s_1_2_2(and_502_cse, nor_303_nl, fsm_output(1));
  and_289_nl <= (fsm_output(5)) AND mux_1288_nl;
  not_tmp_523 <= MUX_s_1_2_2(mux_1291_nl, and_289_nl, fsm_output(0));
  or_tmp_1261 <= (fsm_output(9)) OR (NOT (fsm_output(6)));
  mux_tmp_1305 <= MUX_s_1_2_2((NOT (fsm_output(6))), (fsm_output(6)), fsm_output(9));
  STAGE_LOOP_i_3_0_sva_mx0c1 <= and_dcpl_60 AND and_dcpl_57;
  VEC_LOOP_j_sva_11_0_mx0c1 <= and_dcpl_68 AND and_dcpl_57;
  and_363_nl <= (fsm_output(0)) AND (fsm_output(4)) AND (fsm_output(6)) AND (fsm_output(8))
      AND (fsm_output(9));
  mux_874_nl <= MUX_s_1_2_2(not_tmp_347, and_363_nl, fsm_output(1));
  and_364_nl <= (fsm_output(4)) AND (fsm_output(6)) AND (fsm_output(8)) AND (fsm_output(9));
  mux_875_nl <= MUX_s_1_2_2(mux_874_nl, and_364_nl, fsm_output(2));
  mux_876_nl <= MUX_s_1_2_2(not_tmp_347, mux_875_nl, fsm_output(3));
  mux_877_nl <= MUX_s_1_2_2(mux_876_nl, and_361_cse, fsm_output(5));
  modExp_result_sva_mx0c0 <= MUX_s_1_2_2(mux_877_nl, and_369_cse, fsm_output(7));
  STAGE_LOOP_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(STAGE_LOOP_i_3_0_sva_2(3
      DOWNTO 1)) + SIGNED'( "011"), 3));
  STAGE_LOOP_acc_itm_2_1 <= STAGE_LOOP_acc_nl(2);
  and_224_m1c <= and_dcpl_122 AND and_dcpl_82;
  and_226_m1c <= and_dcpl_129 AND and_dcpl_108 AND nor_393_cse;
  and_229_m1c <= and_dcpl_51 AND and_dcpl_4 AND and_dcpl_56 AND and_dcpl_11;
  and_230_m1c <= and_dcpl_73 AND and_dcpl_109;
  and_233_m1c <= and_dcpl_110 AND and_dcpl_4 AND and_dcpl_47 AND and_dcpl_23;
  and_235_m1c <= and_dcpl_64 AND and_dcpl_14 AND and_dcpl_127;
  and_237_m1c <= and_dcpl_65 AND and_dcpl_108 AND and_dcpl_23;
  and_244_m1c <= and_dcpl_60 AND and_dcpl_67;
  or_1381_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(8))) OR (fsm_output(1))
      OR (fsm_output(6)) OR not_tmp_400;
  or_1382_nl <= (fsm_output(2)) OR (fsm_output(8)) OR (fsm_output(1)) OR (NOT (fsm_output(6)))
      OR (fsm_output(0)) OR (fsm_output(5));
  mux_982_nl <= MUX_s_1_2_2(or_1381_nl, or_1382_nl, fsm_output(7));
  nor_362_nl <= NOT((NOT (fsm_output(8))) OR (NOT (fsm_output(1))) OR (fsm_output(6))
      OR (fsm_output(0)) OR (fsm_output(5)));
  and_348_nl <= (fsm_output(8)) AND (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(0))
      AND (fsm_output(5));
  mux_981_nl <= MUX_s_1_2_2(nor_362_nl, and_348_nl, fsm_output(2));
  nand_113_nl <= NOT((fsm_output(7)) AND mux_981_nl);
  mux_983_nl <= MUX_s_1_2_2(mux_982_nl, nand_113_nl, fsm_output(3));
  nor_361_nl <= NOT((fsm_output(9)) OR mux_983_nl);
  nor_363_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(2))) OR (fsm_output(8)) OR
      (fsm_output(1)) OR (NOT (fsm_output(6))) OR (fsm_output(0)) OR (fsm_output(5)));
  nor_364_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(8))) OR (NOT (fsm_output(1)))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (fsm_output(5)));
  nor_365_nl <= NOT((fsm_output(2)) OR (fsm_output(8)) OR (fsm_output(1)) OR (fsm_output(6))
      OR not_tmp_400);
  mux_979_nl <= MUX_s_1_2_2(nor_364_nl, nor_365_nl, fsm_output(7));
  mux_980_nl <= MUX_s_1_2_2(nor_363_nl, mux_979_nl, fsm_output(3));
  and_349_nl <= (fsm_output(9)) AND mux_980_nl;
  mux_984_m1c <= MUX_s_1_2_2(nor_361_nl, and_349_nl, fsm_output(4));
  and_91_nl <= and_dcpl_73 AND and_dcpl_70 AND nor_393_cse;
  nor_553_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(0)))
      OR (NOT (fsm_output(5))) OR (fsm_output(2)));
  nor_554_nl <= NOT((NOT (fsm_output(1))) OR (NOT (fsm_output(9))) OR (fsm_output(0))
      OR (fsm_output(5)) OR (NOT (fsm_output(2))));
  mux_367_nl <= MUX_s_1_2_2(nor_553_nl, nor_554_nl, fsm_output(7));
  and_419_nl <= (fsm_output(3)) AND mux_367_nl;
  nor_555_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(7))) OR (fsm_output(1)) OR
      (fsm_output(9)) OR (NOT (fsm_output(0))) OR (fsm_output(5)) OR (NOT (fsm_output(2))));
  mux_368_nl <= MUX_s_1_2_2(and_419_nl, nor_555_nl, fsm_output(4));
  and_421_nl <= (fsm_output(7)) AND (fsm_output(1)) AND (fsm_output(9)) AND (fsm_output(0))
      AND (fsm_output(5)) AND (NOT (fsm_output(2)));
  nor_556_nl <= NOT((NOT (fsm_output(7))) OR (NOT (fsm_output(1))) OR (fsm_output(9))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(2)));
  mux_366_nl <= MUX_s_1_2_2(and_421_nl, nor_556_nl, fsm_output(3));
  and_420_nl <= (fsm_output(4)) AND mux_366_nl;
  mux_369_nl <= MUX_s_1_2_2(mux_368_nl, and_420_nl, fsm_output(6));
  nor_557_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(7))) OR (fsm_output(1)) OR
      (fsm_output(9)) OR (fsm_output(0)) OR (fsm_output(5)) OR (NOT (fsm_output(2))));
  or_269_nl <= (NOT (fsm_output(9))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(2));
  or_268_nl <= (fsm_output(9)) OR (NOT (fsm_output(0))) OR (fsm_output(5)) OR (NOT
      (fsm_output(2)));
  mux_364_nl <= MUX_s_1_2_2(or_269_nl, or_268_nl, fsm_output(1));
  nor_558_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(7)) OR mux_364_nl);
  mux_365_nl <= MUX_s_1_2_2(nor_557_nl, nor_558_nl, fsm_output(4));
  and_422_nl <= (fsm_output(6)) AND mux_365_nl;
  mux_370_nl <= MUX_s_1_2_2(mux_369_nl, and_422_nl, fsm_output(8));
  nor_551_nl <= NOT((fsm_output(5)) OR (fsm_output(0)) OR (NOT (fsm_output(4))));
  nor_552_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(0))) OR (fsm_output(4)));
  mux_371_nl <= MUX_s_1_2_2(nor_551_nl, nor_552_nl, fsm_output(6));
  and_96_nl <= mux_371_nl AND (NOT (fsm_output(3))) AND (fsm_output(1)) AND (fsm_output(2))
      AND (fsm_output(7)) AND nor_393_cse;
  nor_549_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(2)) OR (NOT((fsm_output(5))
      AND (fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(4)))));
  nor_550_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(2))) OR (fsm_output(5)) OR
      (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(4)));
  mux_372_nl <= MUX_s_1_2_2(nor_549_nl, nor_550_nl, fsm_output(8));
  and_104_nl <= mux_372_nl AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(9)));
  nor_547_nl <= NOT((NOT (fsm_output(6))) OR (fsm_output(0)) OR (fsm_output(4)));
  nor_548_nl <= NOT((fsm_output(6)) OR (NOT and_437_cse));
  mux_373_nl <= MUX_s_1_2_2(nor_547_nl, nor_548_nl, fsm_output(7));
  and_115_nl <= mux_373_nl AND (NOT (fsm_output(3))) AND (NOT (fsm_output(1))) AND
      (fsm_output(5)) AND (NOT (fsm_output(2))) AND and_dcpl_11;
  nor_545_nl <= NOT((NOT (fsm_output(8))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(0))) OR (fsm_output(1)) OR (fsm_output(4)));
  nor_546_nl <= NOT((fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(0))
      OR (NOT((fsm_output(1)) AND (fsm_output(4)))));
  mux_374_nl <= MUX_s_1_2_2(nor_545_nl, nor_546_nl, fsm_output(9));
  and_123_nl <= mux_374_nl AND (NOT (fsm_output(3))) AND (NOT (fsm_output(5))) AND
      (fsm_output(2));
  nor_544_nl <= NOT((fsm_output(0)) OR (fsm_output(4)));
  mux_375_nl <= MUX_s_1_2_2(nor_544_nl, and_437_cse, fsm_output(6));
  and_136_nl <= mux_375_nl AND (fsm_output(3)) AND (fsm_output(1)) AND (fsm_output(5))
      AND (NOT (fsm_output(2))) AND (NOT (fsm_output(7))) AND and_dcpl_23;
  nor_542_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(5))) OR (fsm_output(0))
      OR (fsm_output(1)) OR (fsm_output(3)));
  nor_543_nl <= NOT((fsm_output(6)) OR (fsm_output(5)) OR (NOT((fsm_output(0)) AND
      (fsm_output(1)) AND (fsm_output(3)))));
  mux_376_nl <= MUX_s_1_2_2(nor_542_nl, nor_543_nl, fsm_output(2));
  and_143_nl <= mux_376_nl AND (NOT (fsm_output(4))) AND (fsm_output(7)) AND and_dcpl_23;
  and_500_nl <= (fsm_output(7)) AND (fsm_output(5)) AND (NOT (fsm_output(0))) AND
      (fsm_output(4));
  nor_541_nl <= NOT((fsm_output(7)) OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR
      (fsm_output(4)));
  mux_377_nl <= MUX_s_1_2_2(and_500_nl, nor_541_nl, fsm_output(8));
  and_152_nl <= mux_377_nl AND (NOT (fsm_output(3))) AND (NOT (fsm_output(1))) AND
      (fsm_output(6)) AND (fsm_output(2)) AND (fsm_output(9));
  vec_rsc_0_0_i_adra_d_pff <= MUX1HOT_v_9_11_2(COMP_LOOP_acc_psp_sva_1, (z_out_3(12
      DOWNTO 4)), COMP_LOOP_acc_psp_sva, (COMP_LOOP_acc_10_cse_12_1_1_sva(11 DOWNTO
      3)), (COMP_LOOP_acc_1_cse_2_sva(11 DOWNTO 3)), (COMP_LOOP_acc_11_psp_sva(10
      DOWNTO 2)), (COMP_LOOP_acc_1_cse_4_sva(11 DOWNTO 3)), (COMP_LOOP_acc_13_psp_sva(9
      DOWNTO 1)), (COMP_LOOP_acc_1_cse_6_sva(11 DOWNTO 3)), (COMP_LOOP_acc_14_psp_sva(10
      DOWNTO 2)), (COMP_LOOP_acc_1_cse_sva(11 DOWNTO 3)), STD_LOGIC_VECTOR'( and_dcpl_66
      & COMP_LOOP_or_2_cse & and_91_nl & mux_370_nl & and_96_nl & and_104_nl & and_115_nl
      & and_123_nl & and_136_nl & and_143_nl & and_152_nl));
  vec_rsc_0_0_i_da_d_pff <= modulo_result_mux_1_cse;
  or_331_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("10111"));
  mux_395_nl <= MUX_s_1_2_2(or_331_nl, or_329_cse, fsm_output(2));
  mux_396_nl <= MUX_s_1_2_2(mux_395_nl, or_tmp_273, fsm_output(1));
  or_326_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("01010"));
  mux_393_nl <= MUX_s_1_2_2(or_327_cse, or_326_nl, fsm_output(2));
  mux_394_nl <= MUX_s_1_2_2(mux_393_nl, mux_392_cse, fsm_output(1));
  mux_397_nl <= MUX_s_1_2_2(mux_396_nl, mux_394_nl, fsm_output(3));
  or_321_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("11010"));
  mux_388_nl <= MUX_s_1_2_2(or_321_nl, or_320_cse, fsm_output(4));
  mux_389_nl <= MUX_s_1_2_2(or_tmp_268, mux_388_nl, fsm_output(2));
  or_316_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("000")) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00111"));
  mux_387_nl <= MUX_s_1_2_2(nand_246_cse, or_316_nl, fsm_output(2));
  mux_390_nl <= MUX_s_1_2_2(mux_389_nl, mux_387_nl, fsm_output(1));
  or_313_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(6))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("000")) OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_385_nl <= MUX_s_1_2_2(or_313_nl, or_312_cse, fsm_output(2));
  mux_386_nl <= MUX_s_1_2_2(or_314_cse, mux_385_nl, fsm_output(1));
  mux_391_nl <= MUX_s_1_2_2(mux_390_nl, mux_386_nl, fsm_output(3));
  mux_398_nl <= MUX_s_1_2_2(mux_397_nl, mux_391_nl, fsm_output(0));
  or_311_nl <= (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(9
      DOWNTO 5)/=STD_LOGIC_VECTOR'("10111"));
  mux_382_nl <= MUX_s_1_2_2(or_311_nl, or_tmp_273, fsm_output(1));
  or_305_nl <= (fsm_output(1)) OR (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(9
      DOWNTO 5)/=STD_LOGIC_VECTOR'("01010"));
  mux_383_nl <= MUX_s_1_2_2(mux_382_nl, or_305_nl, fsm_output(3));
  or_302_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("11010"));
  mux_378_nl <= MUX_s_1_2_2(or_tmp_268, or_302_nl, fsm_output(2));
  or_301_nl <= (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00111"));
  mux_379_nl <= MUX_s_1_2_2(mux_378_nl, or_301_nl, fsm_output(1));
  or_299_nl <= (NOT (fsm_output(1))) OR (fsm_output(2)) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_380_nl <= MUX_s_1_2_2(mux_379_nl, or_299_nl, fsm_output(3));
  mux_384_nl <= MUX_s_1_2_2(mux_383_nl, mux_380_nl, fsm_output(0));
  or_298_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_399_nl <= MUX_s_1_2_2(mux_398_nl, mux_384_nl, or_298_nl);
  vec_rsc_0_0_i_wea_d_pff <= NOT mux_399_nl;
  nor_529_nl <= NOT((COMP_LOOP_acc_13_psp_sva(0)) OR (VEC_LOOP_j_sva_11_0(1)) OR
      (NOT (fsm_output(2))) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      OR not_tmp_165);
  nor_530_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")) OR
      (fsm_output(2)) OR (fsm_output(6)) OR (NOT (fsm_output(7))));
  mux_411_nl <= MUX_s_1_2_2(nor_529_nl, nor_530_nl, fsm_output(3));
  nand_15_nl <= NOT((fsm_output(0)) AND mux_411_nl);
  or_358_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  or_357_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")) OR CONV_SL_1_1(fsm_output(7
      DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_410_nl <= MUX_s_1_2_2(or_358_nl, or_357_nl, fsm_output(2));
  or_359_nl <= (fsm_output(0)) OR (fsm_output(3)) OR mux_410_nl;
  mux_412_nl <= MUX_s_1_2_2(nand_15_nl, or_359_nl, fsm_output(5));
  nor_528_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("01"))
      OR mux_412_nl);
  nor_531_nl <= NOT((NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT (fsm_output(2))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10")));
  nor_532_nl <= NOT((fsm_output(0)) OR (NOT (fsm_output(3))) OR (fsm_output(2)) OR
      (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_408_nl <= MUX_s_1_2_2(nor_531_nl, nor_532_nl, fsm_output(5));
  and_417_nl <= (fsm_output(9)) AND mux_408_nl;
  nor_533_nl <= NOT((fsm_output(9)) OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR nand_190_cse);
  mux_409_nl <= MUX_s_1_2_2(and_417_nl, nor_533_nl, fsm_output(8));
  mux_413_nl <= MUX_s_1_2_2(nor_528_nl, mux_409_nl, fsm_output(1));
  nor_534_nl <= NOT((VEC_LOOP_j_sva_11_0(2)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(0)))
      OR (fsm_output(3)) OR (VEC_LOOP_j_sva_11_0(1)) OR (fsm_output(2)) OR (VEC_LOOP_j_sva_11_0(0))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  or_347_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(2))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR not_tmp_165;
  or_345_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")) OR (fsm_output(2))
      OR (fsm_output(6)) OR (NOT (fsm_output(7)));
  mux_404_nl <= MUX_s_1_2_2(or_347_nl, or_345_nl, fsm_output(3));
  nor_535_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(0)) OR mux_404_nl);
  mux_405_nl <= MUX_s_1_2_2(nor_534_nl, nor_535_nl, fsm_output(9));
  nor_536_nl <= NOT((NOT (fsm_output(9))) OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_406_nl <= MUX_s_1_2_2(mux_405_nl, nor_536_nl, fsm_output(8));
  or_339_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(2))) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(fsm_output(7
      DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_337_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")) OR (fsm_output(2))
      OR (NOT (fsm_output(6))) OR (fsm_output(7));
  mux_401_nl <= MUX_s_1_2_2(or_339_nl, or_337_nl, fsm_output(3));
  or_340_nl <= (fsm_output(0)) OR mux_401_nl;
  nor_538_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) OR
      not_tmp_165);
  nor_539_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")) OR
      CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  mux_400_nl <= MUX_s_1_2_2(nor_538_nl, nor_539_nl, fsm_output(2));
  nand_13_nl <= NOT((fsm_output(0)) AND (fsm_output(3)) AND mux_400_nl);
  mux_402_nl <= MUX_s_1_2_2(or_340_nl, nand_13_nl, fsm_output(5));
  or_332_nl <= (fsm_output(5)) OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR CONV_SL_1_1(z_out_3(3
      DOWNTO 1)/=STD_LOGIC_VECTOR'("000")) OR (fsm_output(2)) OR (NOT (fsm_output(6)))
      OR (fsm_output(7));
  mux_403_nl <= MUX_s_1_2_2(mux_402_nl, or_332_nl, fsm_output(9));
  nor_537_nl <= NOT((fsm_output(8)) OR mux_403_nl);
  mux_407_nl <= MUX_s_1_2_2(mux_406_nl, nor_537_nl, fsm_output(1));
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_413_nl, mux_407_nl,
      fsm_output(4));
  or_398_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("10111"));
  mux_432_nl <= MUX_s_1_2_2(or_398_nl, or_329_cse, fsm_output(2));
  mux_433_nl <= MUX_s_1_2_2(mux_432_nl, or_tmp_340, fsm_output(1));
  or_393_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("01010"));
  mux_430_nl <= MUX_s_1_2_2(or_327_cse, or_393_nl, fsm_output(2));
  mux_431_nl <= MUX_s_1_2_2(mux_430_nl, mux_392_cse, fsm_output(1));
  mux_434_nl <= MUX_s_1_2_2(mux_433_nl, mux_431_nl, fsm_output(3));
  or_388_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("11010"));
  mux_425_nl <= MUX_s_1_2_2(or_388_nl, or_320_cse, fsm_output(4));
  mux_426_nl <= MUX_s_1_2_2(or_tmp_335, mux_425_nl, fsm_output(2));
  or_383_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("001")) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00111"));
  mux_424_nl <= MUX_s_1_2_2(nand_246_cse, or_383_nl, fsm_output(2));
  mux_427_nl <= MUX_s_1_2_2(mux_426_nl, mux_424_nl, fsm_output(1));
  or_380_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(6))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("001")) OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_422_nl <= MUX_s_1_2_2(or_380_nl, or_312_cse, fsm_output(2));
  mux_423_nl <= MUX_s_1_2_2(or_314_cse, mux_422_nl, fsm_output(1));
  mux_428_nl <= MUX_s_1_2_2(mux_427_nl, mux_423_nl, fsm_output(3));
  mux_435_nl <= MUX_s_1_2_2(mux_434_nl, mux_428_nl, fsm_output(0));
  or_378_nl <= (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(9
      DOWNTO 5)/=STD_LOGIC_VECTOR'("10111"));
  mux_419_nl <= MUX_s_1_2_2(or_378_nl, or_tmp_340, fsm_output(1));
  or_372_nl <= (fsm_output(1)) OR (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(9
      DOWNTO 5)/=STD_LOGIC_VECTOR'("01010"));
  mux_420_nl <= MUX_s_1_2_2(mux_419_nl, or_372_nl, fsm_output(3));
  or_369_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("11010"));
  mux_415_nl <= MUX_s_1_2_2(or_tmp_335, or_369_nl, fsm_output(2));
  or_368_nl <= (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00111"));
  mux_416_nl <= MUX_s_1_2_2(mux_415_nl, or_368_nl, fsm_output(1));
  or_366_nl <= (NOT (fsm_output(1))) OR (fsm_output(2)) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_417_nl <= MUX_s_1_2_2(mux_416_nl, or_366_nl, fsm_output(3));
  mux_421_nl <= MUX_s_1_2_2(mux_420_nl, mux_417_nl, fsm_output(0));
  or_365_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_436_nl <= MUX_s_1_2_2(mux_435_nl, mux_421_nl, or_365_nl);
  vec_rsc_0_1_i_wea_d_pff <= NOT mux_436_nl;
  or_423_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR CONV_SL_1_1(fsm_output(5 DOWNTO
      4)/=STD_LOGIC_VECTOR'("10")) OR nand_97_cse;
  or_421_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("001")) OR (NOT
      (fsm_output(5))) OR (fsm_output(4)) OR (fsm_output(6)) OR (NOT (fsm_output(8)));
  mux_448_nl <= MUX_s_1_2_2(or_423_nl, or_421_nl, fsm_output(2));
  nor_514_nl <= NOT((fsm_output(3)) OR mux_448_nl);
  nor_515_nl <= NOT((VEC_LOOP_j_sva_11_0(2)) OR (fsm_output(3)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(2)) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(4))) OR (fsm_output(6)) OR (fsm_output(8)));
  mux_449_nl <= MUX_s_1_2_2(nor_514_nl, nor_515_nl, fsm_output(0));
  nor_516_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("001")) OR
      (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(2))) OR
      (fsm_output(5)) OR (NOT (fsm_output(4))) OR (fsm_output(6)) OR (NOT (fsm_output(8))));
  mux_450_nl <= MUX_s_1_2_2(mux_449_nl, nor_516_nl, fsm_output(9));
  nor_517_nl <= NOT((COMP_LOOP_acc_13_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(2))) OR (fsm_output(5)) OR (fsm_output(4)) OR nand_97_cse);
  nor_518_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("001")) OR
      (fsm_output(2)) OR (fsm_output(5)) OR (fsm_output(4)) OR (fsm_output(6)) OR
      (NOT (fsm_output(8))));
  mux_446_nl <= MUX_s_1_2_2(nor_517_nl, nor_518_nl, fsm_output(3));
  and_414_nl <= (fsm_output(0)) AND mux_446_nl;
  or_411_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(2))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT
      (fsm_output(5))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(8));
  or_410_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("001")) OR (fsm_output(2))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(4))) OR (fsm_output(6)) OR (fsm_output(8));
  mux_445_nl <= MUX_s_1_2_2(or_411_nl, or_410_nl, fsm_output(3));
  nor_519_nl <= NOT((fsm_output(0)) OR mux_445_nl);
  mux_447_nl <= MUX_s_1_2_2(and_414_nl, nor_519_nl, fsm_output(9));
  mux_451_nl <= MUX_s_1_2_2(mux_450_nl, mux_447_nl, fsm_output(7));
  nor_520_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("001")) OR
      (fsm_output(0)) OR (NOT (fsm_output(3))) OR (fsm_output(2)) OR (fsm_output(5))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_521_nl <= NOT((NOT (fsm_output(3))) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(2)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (fsm_output(4)) OR (fsm_output(6))
      OR (fsm_output(8)));
  nor_522_nl <= NOT((fsm_output(3)) OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(2)) OR (fsm_output(5)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6)))
      OR (fsm_output(8)));
  mux_442_nl <= MUX_s_1_2_2(nor_521_nl, nor_522_nl, fsm_output(0));
  mux_443_nl <= MUX_s_1_2_2(nor_520_nl, mux_442_nl, fsm_output(9));
  nor_523_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(2))) OR (fsm_output(5))
      OR (NOT (fsm_output(4))) OR (fsm_output(6)) OR (fsm_output(8)));
  nor_524_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("001")) OR
      (NOT (fsm_output(2))) OR (NOT (fsm_output(5))) OR (fsm_output(4)) OR nand_97_cse);
  mux_439_nl <= MUX_s_1_2_2(nor_523_nl, nor_524_nl, fsm_output(3));
  nor_525_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("001")) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(4))) OR (fsm_output(6)) OR (fsm_output(8)));
  mux_437_nl <= MUX_s_1_2_2(and_416_cse, nor_525_nl, fsm_output(2));
  nor_526_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(4))) OR (fsm_output(6)) OR (fsm_output(8)));
  or_400_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm);
  mux_438_nl <= MUX_s_1_2_2(mux_437_nl, nor_526_nl, or_400_nl);
  and_415_nl <= (fsm_output(3)) AND mux_438_nl;
  mux_440_nl <= MUX_s_1_2_2(mux_439_nl, and_415_nl, fsm_output(0));
  nor_527_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(2))) OR (fsm_output(5))
      OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(8)));
  mux_441_nl <= MUX_s_1_2_2(mux_440_nl, nor_527_nl, fsm_output(9));
  mux_444_nl <= MUX_s_1_2_2(mux_443_nl, mux_441_nl, fsm_output(7));
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_451_nl, mux_444_nl,
      fsm_output(1));
  or_457_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("10111"));
  mux_470_nl <= MUX_s_1_2_2(or_457_nl, or_329_cse, fsm_output(2));
  mux_471_nl <= MUX_s_1_2_2(mux_470_nl, nand_tmp_18, fsm_output(1));
  or_452_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("01010"));
  mux_468_nl <= MUX_s_1_2_2(or_327_cse, or_452_nl, fsm_output(2));
  mux_469_nl <= MUX_s_1_2_2(mux_468_nl, mux_392_cse, fsm_output(1));
  mux_472_nl <= MUX_s_1_2_2(mux_471_nl, mux_469_nl, fsm_output(3));
  or_447_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("11010"));
  mux_463_nl <= MUX_s_1_2_2(or_447_nl, or_320_cse, fsm_output(4));
  mux_464_nl <= MUX_s_1_2_2(or_tmp_395, mux_463_nl, fsm_output(2));
  or_442_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("010")) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00111"));
  mux_462_nl <= MUX_s_1_2_2(nand_246_cse, or_442_nl, fsm_output(2));
  mux_465_nl <= MUX_s_1_2_2(mux_464_nl, mux_462_nl, fsm_output(1));
  or_439_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(6))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("010")) OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_460_nl <= MUX_s_1_2_2(or_439_nl, or_312_cse, fsm_output(2));
  mux_461_nl <= MUX_s_1_2_2(or_314_cse, mux_460_nl, fsm_output(1));
  mux_466_nl <= MUX_s_1_2_2(mux_465_nl, mux_461_nl, fsm_output(3));
  mux_473_nl <= MUX_s_1_2_2(mux_472_nl, mux_466_nl, fsm_output(0));
  or_437_nl <= (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(9
      DOWNTO 5)/=STD_LOGIC_VECTOR'("10111"));
  mux_457_nl <= MUX_s_1_2_2(or_437_nl, nand_tmp_18, fsm_output(1));
  or_432_nl <= (fsm_output(1)) OR (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(9
      DOWNTO 5)/=STD_LOGIC_VECTOR'("01010"));
  mux_458_nl <= MUX_s_1_2_2(mux_457_nl, or_432_nl, fsm_output(3));
  or_429_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("11010"));
  mux_453_nl <= MUX_s_1_2_2(or_tmp_395, or_429_nl, fsm_output(2));
  or_428_nl <= (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00111"));
  mux_454_nl <= MUX_s_1_2_2(mux_453_nl, or_428_nl, fsm_output(1));
  or_426_nl <= (NOT (fsm_output(1))) OR (fsm_output(2)) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_455_nl <= MUX_s_1_2_2(mux_454_nl, or_426_nl, fsm_output(3));
  mux_459_nl <= MUX_s_1_2_2(mux_458_nl, mux_455_nl, fsm_output(0));
  or_425_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_474_nl <= MUX_s_1_2_2(mux_473_nl, mux_459_nl, or_425_nl);
  vec_rsc_0_2_i_wea_d_pff <= NOT mux_474_nl;
  or_482_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR CONV_SL_1_1(fsm_output(5 DOWNTO
      4)/=STD_LOGIC_VECTOR'("10")) OR nand_97_cse;
  or_480_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010")) OR (NOT
      (fsm_output(5))) OR (fsm_output(4)) OR (fsm_output(6)) OR (NOT (fsm_output(8)));
  mux_486_nl <= MUX_s_1_2_2(or_482_nl, or_480_nl, fsm_output(2));
  nor_498_nl <= NOT((fsm_output(3)) OR mux_486_nl);
  nor_499_nl <= NOT((VEC_LOOP_j_sva_11_0(2)) OR (fsm_output(3)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(2)) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(4))) OR (fsm_output(6)) OR (fsm_output(8)));
  mux_487_nl <= MUX_s_1_2_2(nor_498_nl, nor_499_nl, fsm_output(0));
  nor_500_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010")) OR
      (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(2))) OR
      (fsm_output(5)) OR (NOT (fsm_output(4))) OR (fsm_output(6)) OR (NOT (fsm_output(8))));
  mux_488_nl <= MUX_s_1_2_2(mux_487_nl, nor_500_nl, fsm_output(9));
  nor_501_nl <= NOT((COMP_LOOP_acc_13_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(2))) OR (fsm_output(5)) OR (fsm_output(4)) OR nand_97_cse);
  nor_502_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010")) OR
      (fsm_output(2)) OR (fsm_output(5)) OR (fsm_output(4)) OR (fsm_output(6)) OR
      (NOT (fsm_output(8))));
  mux_484_nl <= MUX_s_1_2_2(nor_501_nl, nor_502_nl, fsm_output(3));
  and_411_nl <= (fsm_output(0)) AND mux_484_nl;
  or_470_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(2))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (NOT
      (fsm_output(5))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(8));
  or_469_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010")) OR (fsm_output(2))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(4))) OR (fsm_output(6)) OR (fsm_output(8));
  mux_483_nl <= MUX_s_1_2_2(or_470_nl, or_469_nl, fsm_output(3));
  nor_503_nl <= NOT((fsm_output(0)) OR mux_483_nl);
  mux_485_nl <= MUX_s_1_2_2(and_411_nl, nor_503_nl, fsm_output(9));
  mux_489_nl <= MUX_s_1_2_2(mux_488_nl, mux_485_nl, fsm_output(7));
  nor_504_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010")) OR
      (fsm_output(0)) OR (NOT (fsm_output(3))) OR (fsm_output(2)) OR (fsm_output(5))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_505_nl <= NOT((NOT (fsm_output(3))) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(2)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (fsm_output(4)) OR (fsm_output(6))
      OR (fsm_output(8)));
  nor_506_nl <= NOT((fsm_output(3)) OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(2)) OR (fsm_output(5)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6)))
      OR (fsm_output(8)));
  mux_480_nl <= MUX_s_1_2_2(nor_505_nl, nor_506_nl, fsm_output(0));
  mux_481_nl <= MUX_s_1_2_2(nor_504_nl, mux_480_nl, fsm_output(9));
  nor_507_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(2))) OR (fsm_output(5))
      OR (NOT (fsm_output(4))) OR (fsm_output(6)) OR (fsm_output(8)));
  nor_508_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010")) OR
      (NOT (fsm_output(2))) OR (NOT (fsm_output(5))) OR (fsm_output(4)) OR nand_97_cse);
  mux_477_nl <= MUX_s_1_2_2(nor_507_nl, nor_508_nl, fsm_output(3));
  nor_509_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010")) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(4))) OR (fsm_output(6)) OR (fsm_output(8)));
  mux_475_nl <= MUX_s_1_2_2(and_416_cse, nor_509_nl, fsm_output(2));
  nor_510_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(4))) OR (fsm_output(6)) OR (fsm_output(8)));
  or_459_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm);
  mux_476_nl <= MUX_s_1_2_2(mux_475_nl, nor_510_nl, or_459_nl);
  and_412_nl <= (fsm_output(3)) AND mux_476_nl;
  mux_478_nl <= MUX_s_1_2_2(mux_477_nl, and_412_nl, fsm_output(0));
  nor_511_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(2))) OR (fsm_output(5))
      OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(8)));
  mux_479_nl <= MUX_s_1_2_2(mux_478_nl, nor_511_nl, fsm_output(9));
  mux_482_nl <= MUX_s_1_2_2(mux_481_nl, mux_479_nl, fsm_output(7));
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_489_nl, mux_482_nl,
      fsm_output(1));
  or_516_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("10111"));
  mux_508_nl <= MUX_s_1_2_2(or_516_nl, or_329_cse, fsm_output(2));
  mux_509_nl <= MUX_s_1_2_2(mux_508_nl, nand_tmp_21, fsm_output(1));
  or_511_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("01010"));
  mux_506_nl <= MUX_s_1_2_2(or_327_cse, or_511_nl, fsm_output(2));
  mux_507_nl <= MUX_s_1_2_2(mux_506_nl, mux_392_cse, fsm_output(1));
  mux_510_nl <= MUX_s_1_2_2(mux_509_nl, mux_507_nl, fsm_output(3));
  or_506_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("11010"));
  mux_501_nl <= MUX_s_1_2_2(or_506_nl, or_320_cse, fsm_output(4));
  mux_502_nl <= MUX_s_1_2_2(or_tmp_454, mux_501_nl, fsm_output(2));
  or_501_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("011")) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00111"));
  mux_500_nl <= MUX_s_1_2_2(nand_246_cse, or_501_nl, fsm_output(2));
  mux_503_nl <= MUX_s_1_2_2(mux_502_nl, mux_500_nl, fsm_output(1));
  or_498_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(6))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("011")) OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_498_nl <= MUX_s_1_2_2(or_498_nl, or_312_cse, fsm_output(2));
  mux_499_nl <= MUX_s_1_2_2(or_314_cse, mux_498_nl, fsm_output(1));
  mux_504_nl <= MUX_s_1_2_2(mux_503_nl, mux_499_nl, fsm_output(3));
  mux_511_nl <= MUX_s_1_2_2(mux_510_nl, mux_504_nl, fsm_output(0));
  or_496_nl <= (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(9
      DOWNTO 5)/=STD_LOGIC_VECTOR'("10111"));
  mux_495_nl <= MUX_s_1_2_2(or_496_nl, nand_tmp_21, fsm_output(1));
  or_491_nl <= (fsm_output(1)) OR (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(9
      DOWNTO 5)/=STD_LOGIC_VECTOR'("01010"));
  mux_496_nl <= MUX_s_1_2_2(mux_495_nl, or_491_nl, fsm_output(3));
  or_488_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("11010"));
  mux_491_nl <= MUX_s_1_2_2(or_tmp_454, or_488_nl, fsm_output(2));
  or_487_nl <= (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00111"));
  mux_492_nl <= MUX_s_1_2_2(mux_491_nl, or_487_nl, fsm_output(1));
  or_485_nl <= (NOT (fsm_output(1))) OR (fsm_output(2)) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_493_nl <= MUX_s_1_2_2(mux_492_nl, or_485_nl, fsm_output(3));
  mux_497_nl <= MUX_s_1_2_2(mux_496_nl, mux_493_nl, fsm_output(0));
  or_484_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"));
  mux_512_nl <= MUX_s_1_2_2(mux_511_nl, mux_497_nl, or_484_nl);
  vec_rsc_0_3_i_wea_d_pff <= NOT mux_512_nl;
  nor_485_nl <= NOT((NOT((NOT (COMP_LOOP_acc_13_psp_sva(0))) AND (VEC_LOOP_j_sva_11_0(1))
      AND (fsm_output(2)) AND (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm))
      OR not_tmp_165);
  nor_486_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("011")) OR
      (fsm_output(2)) OR (fsm_output(6)) OR (NOT (fsm_output(7))));
  mux_524_nl <= MUX_s_1_2_2(nor_485_nl, nor_486_nl, fsm_output(3));
  nand_24_nl <= NOT((fsm_output(0)) AND mux_524_nl);
  or_543_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  or_542_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("011")) OR CONV_SL_1_1(fsm_output(7
      DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_523_nl <= MUX_s_1_2_2(or_543_nl, or_542_nl, fsm_output(2));
  or_544_nl <= (fsm_output(0)) OR (fsm_output(3)) OR mux_523_nl;
  mux_525_nl <= MUX_s_1_2_2(nand_24_nl, or_544_nl, fsm_output(5));
  nor_484_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("01"))
      OR mux_525_nl);
  and_499_nl <= (fsm_output(0)) AND (fsm_output(3)) AND CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("01")) AND (fsm_output(2)) AND (VEC_LOOP_j_sva_11_0(0))
      AND COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("10"));
  nor_488_nl <= NOT((fsm_output(0)) OR (NOT (fsm_output(3))) OR (fsm_output(2)) OR
      (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_521_nl <= MUX_s_1_2_2(and_499_nl, nor_488_nl, fsm_output(5));
  and_410_nl <= (fsm_output(9)) AND mux_521_nl;
  nor_489_nl <= NOT((fsm_output(9)) OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR nand_190_cse);
  mux_522_nl <= MUX_s_1_2_2(and_410_nl, nor_489_nl, fsm_output(8));
  mux_526_nl <= MUX_s_1_2_2(nor_484_nl, mux_522_nl, fsm_output(1));
  nor_490_nl <= NOT((VEC_LOOP_j_sva_11_0(2)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(0)))
      OR (fsm_output(3)) OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR (fsm_output(2)) OR
      (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  or_532_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))
      AND (fsm_output(2)) AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)) OR not_tmp_165;
  or_530_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("011")) OR (fsm_output(2))
      OR (fsm_output(6)) OR (NOT (fsm_output(7)));
  mux_517_nl <= MUX_s_1_2_2(or_532_nl, or_530_nl, fsm_output(3));
  nor_491_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(0)) OR mux_517_nl);
  mux_518_nl <= MUX_s_1_2_2(nor_490_nl, nor_491_nl, fsm_output(9));
  nor_492_nl <= NOT((NOT (fsm_output(9))) OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_519_nl <= MUX_s_1_2_2(mux_518_nl, nor_492_nl, fsm_output(8));
  nand_232_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))
      AND (fsm_output(2)) AND COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm AND CONV_SL_1_1(fsm_output(7
      DOWNTO 6)=STD_LOGIC_VECTOR'("10")));
  or_522_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("011")) OR (fsm_output(2))
      OR (NOT (fsm_output(6))) OR (fsm_output(7));
  mux_514_nl <= MUX_s_1_2_2(nand_232_nl, or_522_nl, fsm_output(3));
  or_525_nl <= (fsm_output(0)) OR mux_514_nl;
  nor_494_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)) OR not_tmp_165);
  nor_495_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("011")) OR
      CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  mux_513_nl <= MUX_s_1_2_2(nor_494_nl, nor_495_nl, fsm_output(2));
  nand_22_nl <= NOT((fsm_output(0)) AND (fsm_output(3)) AND mux_513_nl);
  mux_515_nl <= MUX_s_1_2_2(or_525_nl, nand_22_nl, fsm_output(5));
  or_517_nl <= (fsm_output(5)) OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR CONV_SL_1_1(z_out_3(3
      DOWNTO 1)/=STD_LOGIC_VECTOR'("011")) OR (fsm_output(2)) OR (NOT (fsm_output(6)))
      OR (fsm_output(7));
  mux_516_nl <= MUX_s_1_2_2(mux_515_nl, or_517_nl, fsm_output(9));
  nor_493_nl <= NOT((fsm_output(8)) OR mux_516_nl);
  mux_520_nl <= MUX_s_1_2_2(mux_519_nl, nor_493_nl, fsm_output(1));
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_526_nl, mux_520_nl,
      fsm_output(4));
  or_582_nl <= (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(9
      DOWNTO 5)/=STD_LOGIC_VECTOR'("10111"));
  mux_546_nl <= MUX_s_1_2_2(or_582_nl, or_tmp_535, fsm_output(1));
  or_580_nl <= (fsm_output(1)) OR (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(9
      DOWNTO 5)/=STD_LOGIC_VECTOR'("01010"));
  mux_547_nl <= MUX_s_1_2_2(mux_546_nl, or_580_nl, fsm_output(3));
  or_579_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("11010"));
  mux_543_nl <= MUX_s_1_2_2(or_tmp_525, or_579_nl, fsm_output(2));
  or_578_nl <= (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00111"));
  mux_544_nl <= MUX_s_1_2_2(mux_543_nl, or_578_nl, fsm_output(1));
  or_576_nl <= (NOT (fsm_output(1))) OR (fsm_output(2)) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_545_nl <= MUX_s_1_2_2(mux_544_nl, or_576_nl, fsm_output(3));
  mux_548_nl <= MUX_s_1_2_2(mux_547_nl, mux_545_nl, fsm_output(0));
  or_575_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("10111"));
  mux_539_nl <= MUX_s_1_2_2(or_575_nl, or_329_cse, fsm_output(2));
  mux_540_nl <= MUX_s_1_2_2(mux_539_nl, or_tmp_535, fsm_output(1));
  or_566_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("01010"));
  mux_536_nl <= MUX_s_1_2_2(or_327_cse, or_566_nl, fsm_output(2));
  mux_537_nl <= MUX_s_1_2_2(mux_536_nl, mux_392_cse, fsm_output(1));
  mux_541_nl <= MUX_s_1_2_2(mux_540_nl, mux_537_nl, fsm_output(3));
  or_559_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("11010"));
  mux_531_nl <= MUX_s_1_2_2(or_559_nl, or_320_cse, fsm_output(4));
  mux_532_nl <= MUX_s_1_2_2(or_tmp_525, mux_531_nl, fsm_output(2));
  or_554_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("100")) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00111"));
  mux_530_nl <= MUX_s_1_2_2(nand_246_cse, or_554_nl, fsm_output(2));
  mux_533_nl <= MUX_s_1_2_2(mux_532_nl, mux_530_nl, fsm_output(1));
  or_551_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(6))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("100")) OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_528_nl <= MUX_s_1_2_2(or_551_nl, or_312_cse, fsm_output(2));
  mux_529_nl <= MUX_s_1_2_2(or_314_cse, mux_528_nl, fsm_output(1));
  mux_534_nl <= MUX_s_1_2_2(mux_533_nl, mux_529_nl, fsm_output(3));
  mux_542_nl <= MUX_s_1_2_2(mux_541_nl, mux_534_nl, fsm_output(0));
  nor_114_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100")));
  mux_549_nl <= MUX_s_1_2_2(mux_548_nl, mux_542_nl, nor_114_nl);
  vec_rsc_0_4_i_wea_d_pff <= NOT mux_549_nl;
  nor_473_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("100")) OR
      (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(7))));
  nor_474_nl <= NOT((NOT (COMP_LOOP_acc_13_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR not_tmp_165);
  mux_561_nl <= MUX_s_1_2_2(nor_473_cse, nor_474_nl, fsm_output(2));
  nand_27_nl <= NOT((fsm_output(0)) AND mux_561_nl);
  or_608_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR (fsm_output(7));
  or_607_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("100")) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(7));
  mux_560_nl <= MUX_s_1_2_2(or_608_nl, or_607_nl, fsm_output(2));
  or_609_nl <= (fsm_output(0)) OR mux_560_nl;
  mux_562_nl <= MUX_s_1_2_2(nand_27_nl, or_609_nl, fsm_output(5));
  nor_472_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("01"))
      OR mux_562_nl);
  nor_475_nl <= NOT((NOT (fsm_output(0))) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(7))));
  nor_476_nl <= NOT((fsm_output(0)) OR (fsm_output(2)) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(3))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("100")) OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_558_nl <= MUX_s_1_2_2(nor_475_nl, nor_476_nl, fsm_output(5));
  and_409_nl <= (fsm_output(9)) AND mux_558_nl;
  nor_477_nl <= NOT((fsm_output(9)) OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR nand_190_cse);
  mux_559_nl <= MUX_s_1_2_2(and_409_nl, nor_477_nl, fsm_output(8));
  mux_563_nl <= MUX_s_1_2_2(nor_472_nl, mux_559_nl, fsm_output(1));
  nor_478_nl <= NOT((NOT (VEC_LOOP_j_sva_11_0(2))) OR (NOT (fsm_output(5))) OR (NOT
      (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(7)));
  or_598_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("100")) OR (NOT
      (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(7)));
  or_596_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(3)) OR not_tmp_165;
  mux_554_nl <= MUX_s_1_2_2(or_598_nl, or_596_nl, fsm_output(2));
  nor_479_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(0)) OR mux_554_nl);
  mux_555_nl <= MUX_s_1_2_2(nor_478_nl, nor_479_nl, fsm_output(9));
  nor_480_nl <= NOT((NOT (fsm_output(9))) OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(2))) OR (NOT
      (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_556_nl <= MUX_s_1_2_2(mux_555_nl, nor_480_nl, fsm_output(8));
  or_590_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("100")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(7));
  or_589_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(7)));
  mux_551_nl <= MUX_s_1_2_2(or_590_nl, or_589_nl, fsm_output(2));
  or_591_nl <= (fsm_output(0)) OR mux_551_nl;
  nor_482_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) OR
      nand_168_cse);
  mux_550_nl <= MUX_s_1_2_2(nor_482_nl, nor_473_cse, fsm_output(2));
  nand_25_nl <= NOT((fsm_output(0)) AND mux_550_nl);
  mux_552_nl <= MUX_s_1_2_2(or_591_nl, nand_25_nl, fsm_output(5));
  or_583_nl <= (fsm_output(5)) OR (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(3))
      OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("100")) OR CONV_SL_1_1(fsm_output(7
      DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_553_nl <= MUX_s_1_2_2(mux_552_nl, or_583_nl, fsm_output(9));
  nor_481_nl <= NOT((fsm_output(8)) OR mux_553_nl);
  mux_557_nl <= MUX_s_1_2_2(mux_556_nl, nor_481_nl, fsm_output(1));
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_563_nl, mux_557_nl,
      fsm_output(4));
  or_647_nl <= (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(9
      DOWNTO 5)/=STD_LOGIC_VECTOR'("10111"));
  mux_583_nl <= MUX_s_1_2_2(or_647_nl, or_tmp_600, fsm_output(1));
  or_645_nl <= (fsm_output(1)) OR (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(9
      DOWNTO 5)/=STD_LOGIC_VECTOR'("01010"));
  mux_584_nl <= MUX_s_1_2_2(mux_583_nl, or_645_nl, fsm_output(3));
  or_644_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("11010"));
  mux_580_nl <= MUX_s_1_2_2(or_tmp_590, or_644_nl, fsm_output(2));
  or_643_nl <= (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00111"));
  mux_581_nl <= MUX_s_1_2_2(mux_580_nl, or_643_nl, fsm_output(1));
  or_641_nl <= (NOT (fsm_output(1))) OR (fsm_output(2)) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_582_nl <= MUX_s_1_2_2(mux_581_nl, or_641_nl, fsm_output(3));
  mux_585_nl <= MUX_s_1_2_2(mux_584_nl, mux_582_nl, fsm_output(0));
  or_640_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("10111"));
  mux_576_nl <= MUX_s_1_2_2(or_640_nl, or_329_cse, fsm_output(2));
  mux_577_nl <= MUX_s_1_2_2(mux_576_nl, or_tmp_600, fsm_output(1));
  or_631_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("01010"));
  mux_573_nl <= MUX_s_1_2_2(or_327_cse, or_631_nl, fsm_output(2));
  mux_574_nl <= MUX_s_1_2_2(mux_573_nl, mux_392_cse, fsm_output(1));
  mux_578_nl <= MUX_s_1_2_2(mux_577_nl, mux_574_nl, fsm_output(3));
  or_624_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("11010"));
  mux_568_nl <= MUX_s_1_2_2(or_624_nl, or_320_cse, fsm_output(4));
  mux_569_nl <= MUX_s_1_2_2(or_tmp_590, mux_568_nl, fsm_output(2));
  or_619_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("101")) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00111"));
  mux_567_nl <= MUX_s_1_2_2(nand_246_cse, or_619_nl, fsm_output(2));
  mux_570_nl <= MUX_s_1_2_2(mux_569_nl, mux_567_nl, fsm_output(1));
  or_616_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(6))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("101")) OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_565_nl <= MUX_s_1_2_2(or_616_nl, or_312_cse, fsm_output(2));
  mux_566_nl <= MUX_s_1_2_2(or_314_cse, mux_565_nl, fsm_output(1));
  mux_571_nl <= MUX_s_1_2_2(mux_570_nl, mux_566_nl, fsm_output(3));
  mux_579_nl <= MUX_s_1_2_2(mux_578_nl, mux_571_nl, fsm_output(0));
  nor_120_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101")));
  mux_586_nl <= MUX_s_1_2_2(mux_585_nl, mux_579_nl, nor_120_nl);
  vec_rsc_0_5_i_wea_d_pff <= NOT mux_586_nl;
  nor_461_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("101")) OR
      (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(7))));
  nor_462_nl <= NOT((NOT (COMP_LOOP_acc_13_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR not_tmp_165);
  mux_598_nl <= MUX_s_1_2_2(nor_461_cse, nor_462_nl, fsm_output(2));
  nand_30_nl <= NOT((fsm_output(0)) AND mux_598_nl);
  or_673_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR (fsm_output(7));
  or_672_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("101")) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(7));
  mux_597_nl <= MUX_s_1_2_2(or_673_nl, or_672_nl, fsm_output(2));
  or_674_nl <= (fsm_output(0)) OR mux_597_nl;
  mux_599_nl <= MUX_s_1_2_2(nand_30_nl, or_674_nl, fsm_output(5));
  nor_460_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("01"))
      OR mux_599_nl);
  and_498_nl <= (fsm_output(0)) AND (fsm_output(2)) AND CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("10")) AND (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(7));
  nor_464_nl <= NOT((fsm_output(0)) OR (fsm_output(2)) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(3))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("101")) OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_595_nl <= MUX_s_1_2_2(and_498_nl, nor_464_nl, fsm_output(5));
  and_408_nl <= (fsm_output(9)) AND mux_595_nl;
  nor_465_nl <= NOT((fsm_output(9)) OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR nand_190_cse);
  mux_596_nl <= MUX_s_1_2_2(and_408_nl, nor_465_nl, fsm_output(8));
  mux_600_nl <= MUX_s_1_2_2(nor_460_nl, mux_596_nl, fsm_output(1));
  nor_466_nl <= NOT((NOT (VEC_LOOP_j_sva_11_0(2))) OR (NOT (fsm_output(5))) OR (NOT
      (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(7)));
  or_663_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("101")) OR (NOT
      (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(7)));
  or_661_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(3)) OR not_tmp_165;
  mux_591_nl <= MUX_s_1_2_2(or_663_nl, or_661_nl, fsm_output(2));
  nor_467_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(0)) OR mux_591_nl);
  mux_592_nl <= MUX_s_1_2_2(nor_466_nl, nor_467_nl, fsm_output(9));
  nor_468_nl <= NOT((NOT (fsm_output(9))) OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(2))) OR (NOT
      (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_593_nl <= MUX_s_1_2_2(mux_592_nl, nor_468_nl, fsm_output(8));
  or_655_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("101")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(7));
  or_654_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(7)));
  mux_588_nl <= MUX_s_1_2_2(or_655_nl, or_654_nl, fsm_output(2));
  or_656_nl <= (fsm_output(0)) OR mux_588_nl;
  nor_470_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)) OR nand_168_cse);
  mux_587_nl <= MUX_s_1_2_2(nor_470_nl, nor_461_cse, fsm_output(2));
  nand_28_nl <= NOT((fsm_output(0)) AND mux_587_nl);
  mux_589_nl <= MUX_s_1_2_2(or_656_nl, nand_28_nl, fsm_output(5));
  or_648_nl <= (fsm_output(5)) OR (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(3))
      OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("101")) OR CONV_SL_1_1(fsm_output(7
      DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_590_nl <= MUX_s_1_2_2(mux_589_nl, or_648_nl, fsm_output(9));
  nor_469_nl <= NOT((fsm_output(8)) OR mux_590_nl);
  mux_594_nl <= MUX_s_1_2_2(mux_593_nl, nor_469_nl, fsm_output(1));
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_600_nl, mux_594_nl,
      fsm_output(4));
  or_711_nl <= (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(9
      DOWNTO 5)/=STD_LOGIC_VECTOR'("10111"));
  mux_620_nl <= MUX_s_1_2_2(or_711_nl, nand_tmp_31, fsm_output(1));
  or_709_nl <= (fsm_output(1)) OR (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(9
      DOWNTO 5)/=STD_LOGIC_VECTOR'("01010"));
  mux_621_nl <= MUX_s_1_2_2(mux_620_nl, or_709_nl, fsm_output(3));
  or_708_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("11010"));
  mux_617_nl <= MUX_s_1_2_2(or_tmp_655, or_708_nl, fsm_output(2));
  or_707_nl <= (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00111"));
  mux_618_nl <= MUX_s_1_2_2(mux_617_nl, or_707_nl, fsm_output(1));
  or_705_nl <= (NOT (fsm_output(1))) OR (fsm_output(2)) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_619_nl <= MUX_s_1_2_2(mux_618_nl, or_705_nl, fsm_output(3));
  mux_622_nl <= MUX_s_1_2_2(mux_621_nl, mux_619_nl, fsm_output(0));
  or_704_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("10111"));
  mux_613_nl <= MUX_s_1_2_2(or_704_nl, or_329_cse, fsm_output(2));
  mux_614_nl <= MUX_s_1_2_2(mux_613_nl, nand_tmp_31, fsm_output(1));
  or_696_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("01010"));
  mux_610_nl <= MUX_s_1_2_2(or_327_cse, or_696_nl, fsm_output(2));
  mux_611_nl <= MUX_s_1_2_2(mux_610_nl, mux_392_cse, fsm_output(1));
  mux_615_nl <= MUX_s_1_2_2(mux_614_nl, mux_611_nl, fsm_output(3));
  or_689_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("11010"));
  mux_605_nl <= MUX_s_1_2_2(or_689_nl, or_320_cse, fsm_output(4));
  mux_606_nl <= MUX_s_1_2_2(or_tmp_655, mux_605_nl, fsm_output(2));
  or_684_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("110")) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00111"));
  mux_604_nl <= MUX_s_1_2_2(nand_246_cse, or_684_nl, fsm_output(2));
  mux_607_nl <= MUX_s_1_2_2(mux_606_nl, mux_604_nl, fsm_output(1));
  or_681_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(6))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("110")) OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_602_nl <= MUX_s_1_2_2(or_681_nl, or_312_cse, fsm_output(2));
  mux_603_nl <= MUX_s_1_2_2(or_314_cse, mux_602_nl, fsm_output(1));
  mux_608_nl <= MUX_s_1_2_2(mux_607_nl, mux_603_nl, fsm_output(3));
  mux_616_nl <= MUX_s_1_2_2(mux_615_nl, mux_608_nl, fsm_output(0));
  nor_126_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110")));
  mux_623_nl <= MUX_s_1_2_2(mux_622_nl, mux_616_nl, nor_126_nl);
  vec_rsc_0_6_i_wea_d_pff <= NOT mux_623_nl;
  nor_447_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("110")) OR
      (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(7))));
  nor_448_nl <= NOT((NOT (COMP_LOOP_acc_13_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR not_tmp_165);
  mux_635_nl <= MUX_s_1_2_2(nor_447_cse, nor_448_nl, fsm_output(2));
  nand_34_nl <= NOT((fsm_output(0)) AND mux_635_nl);
  or_737_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR (fsm_output(7));
  or_736_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("110")) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(7));
  mux_634_nl <= MUX_s_1_2_2(or_737_nl, or_736_nl, fsm_output(2));
  or_738_nl <= (fsm_output(0)) OR mux_634_nl;
  mux_636_nl <= MUX_s_1_2_2(nand_34_nl, or_738_nl, fsm_output(5));
  nor_446_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("01"))
      OR mux_636_nl);
  and_497_nl <= (fsm_output(0)) AND (fsm_output(2)) AND CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (NOT (VEC_LOOP_j_sva_11_0(0))) AND COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(7));
  nor_450_nl <= NOT((fsm_output(0)) OR (fsm_output(2)) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(3))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("110")) OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_632_nl <= MUX_s_1_2_2(and_497_nl, nor_450_nl, fsm_output(5));
  and_407_nl <= (fsm_output(9)) AND mux_632_nl;
  nor_451_nl <= NOT((fsm_output(9)) OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR nand_190_cse);
  mux_633_nl <= MUX_s_1_2_2(and_407_nl, nor_451_nl, fsm_output(8));
  mux_637_nl <= MUX_s_1_2_2(nor_446_nl, mux_633_nl, fsm_output(1));
  nor_452_nl <= NOT((NOT (VEC_LOOP_j_sva_11_0(2))) OR (NOT (fsm_output(5))) OR (NOT
      (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(7)));
  or_727_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("110")) OR (NOT
      (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(7)));
  or_725_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(3)) OR not_tmp_165;
  mux_628_nl <= MUX_s_1_2_2(or_727_nl, or_725_nl, fsm_output(2));
  nor_453_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(0)) OR mux_628_nl);
  mux_629_nl <= MUX_s_1_2_2(nor_452_nl, nor_453_nl, fsm_output(9));
  nor_454_nl <= NOT((NOT (fsm_output(9))) OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(2))) OR (NOT
      (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_630_nl <= MUX_s_1_2_2(mux_629_nl, nor_454_nl, fsm_output(8));
  or_719_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("110")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(7));
  or_718_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(7)));
  mux_625_nl <= MUX_s_1_2_2(or_719_nl, or_718_nl, fsm_output(2));
  or_720_nl <= (fsm_output(0)) OR mux_625_nl;
  nor_456_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (NOT (VEC_LOOP_j_sva_11_0(0))) AND COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm))
      OR nand_168_cse);
  mux_624_nl <= MUX_s_1_2_2(nor_456_nl, nor_447_cse, fsm_output(2));
  nand_32_nl <= NOT((fsm_output(0)) AND mux_624_nl);
  mux_626_nl <= MUX_s_1_2_2(or_720_nl, nand_32_nl, fsm_output(5));
  or_712_nl <= (fsm_output(5)) OR (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(3))
      OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("110")) OR CONV_SL_1_1(fsm_output(7
      DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_627_nl <= MUX_s_1_2_2(mux_626_nl, or_712_nl, fsm_output(9));
  nor_455_nl <= NOT((fsm_output(8)) OR mux_627_nl);
  mux_631_nl <= MUX_s_1_2_2(mux_630_nl, nor_455_nl, fsm_output(1));
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_637_nl, mux_631_nl,
      fsm_output(4));
  nand_251_nl <= NOT((NOT (fsm_output(2))) AND (NOT (fsm_output(4))) AND CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (VEC_LOOP_j_sva_11_0(0)) AND CONV_SL_1_1(fsm_output(9
      DOWNTO 5)=STD_LOGIC_VECTOR'("10111")));
  mux_657_nl <= MUX_s_1_2_2(nand_251_nl, nand_tmp_35, fsm_output(1));
  or_773_nl <= (fsm_output(1)) OR (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(9
      DOWNTO 5)/=STD_LOGIC_VECTOR'("01010"));
  mux_658_nl <= MUX_s_1_2_2(mux_657_nl, or_773_nl, fsm_output(3));
  or_772_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("11010"));
  mux_654_nl <= MUX_s_1_2_2(or_tmp_719, or_772_nl, fsm_output(2));
  nand_252_nl <= NOT((fsm_output(2)) AND (NOT (fsm_output(4))) AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND CONV_SL_1_1(fsm_output(9 DOWNTO 5)=STD_LOGIC_VECTOR'("00111")));
  mux_655_nl <= MUX_s_1_2_2(mux_654_nl, nand_252_nl, fsm_output(1));
  nand_144_nl <= NOT((fsm_output(1)) AND (NOT (fsm_output(2))) AND (fsm_output(4))
      AND (fsm_output(9)) AND (fsm_output(5)) AND (fsm_output(6)) AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("00")));
  mux_656_nl <= MUX_s_1_2_2(mux_655_nl, nand_144_nl, fsm_output(3));
  mux_659_nl <= MUX_s_1_2_2(mux_658_nl, mux_656_nl, fsm_output(0));
  nand_250_nl <= NOT((NOT (fsm_output(4))) AND CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (VEC_LOOP_j_sva_11_0(0)) AND CONV_SL_1_1(fsm_output(9
      DOWNTO 5)=STD_LOGIC_VECTOR'("10111")));
  mux_650_nl <= MUX_s_1_2_2(nand_250_nl, or_329_cse, fsm_output(2));
  mux_651_nl <= MUX_s_1_2_2(mux_650_nl, nand_tmp_35, fsm_output(1));
  or_760_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("01010"));
  mux_647_nl <= MUX_s_1_2_2(or_327_cse, or_760_nl, fsm_output(2));
  mux_648_nl <= MUX_s_1_2_2(mux_647_nl, mux_392_cse, fsm_output(1));
  mux_652_nl <= MUX_s_1_2_2(mux_651_nl, mux_648_nl, fsm_output(3));
  nand_147_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND CONV_SL_1_1(fsm_output(9 DOWNTO 5)=STD_LOGIC_VECTOR'("11010")));
  mux_642_nl <= MUX_s_1_2_2(nand_147_nl, or_320_cse, fsm_output(4));
  mux_643_nl <= MUX_s_1_2_2(or_tmp_719, mux_642_nl, fsm_output(2));
  or_748_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("111")) OR CONV_SL_1_1(fsm_output(9 DOWNTO 5)/=STD_LOGIC_VECTOR'("00111"));
  mux_641_nl <= MUX_s_1_2_2(nand_246_cse, or_748_nl, fsm_output(2));
  mux_644_nl <= MUX_s_1_2_2(mux_643_nl, mux_641_nl, fsm_output(1));
  nand_149_nl <= NOT((fsm_output(4)) AND (fsm_output(9)) AND (fsm_output(5)) AND
      (fsm_output(6)) AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("00")));
  mux_639_nl <= MUX_s_1_2_2(nand_149_nl, or_312_cse, fsm_output(2));
  mux_640_nl <= MUX_s_1_2_2(or_314_cse, mux_639_nl, fsm_output(1));
  mux_645_nl <= MUX_s_1_2_2(mux_644_nl, mux_640_nl, fsm_output(3));
  mux_653_nl <= MUX_s_1_2_2(mux_652_nl, mux_645_nl, fsm_output(0));
  and_406_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"));
  mux_660_nl <= MUX_s_1_2_2(mux_659_nl, mux_653_nl, and_406_nl);
  vec_rsc_0_7_i_wea_d_pff <= NOT mux_660_nl;
  and_494_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111")) AND (fsm_output(3))
      AND (NOT (fsm_output(6))) AND (fsm_output(7));
  nor_435_nl <= NOT((NOT((COMP_LOOP_acc_13_psp_sva(0)) AND CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm
      AND (NOT (fsm_output(3))))) OR not_tmp_165);
  mux_672_nl <= MUX_s_1_2_2(and_494_cse, nor_435_nl, fsm_output(2));
  nand_38_nl <= NOT((fsm_output(0)) AND mux_672_nl);
  nand_134_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND (NOT (fsm_output(3))) AND (fsm_output(6))
      AND (NOT (fsm_output(7))));
  or_800_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("111")) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(7));
  mux_671_nl <= MUX_s_1_2_2(nand_134_nl, or_800_nl, fsm_output(2));
  or_802_nl <= (fsm_output(0)) OR mux_671_nl;
  mux_673_nl <= MUX_s_1_2_2(nand_38_nl, or_802_nl, fsm_output(5));
  nor_433_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("01"))
      OR mux_673_nl);
  and_495_nl <= (fsm_output(0)) AND (fsm_output(2)) AND CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(7));
  nor_437_nl <= NOT((fsm_output(0)) OR (fsm_output(2)) OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(3))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("111")) OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_669_nl <= MUX_s_1_2_2(and_495_nl, nor_437_nl, fsm_output(5));
  and_404_nl <= (fsm_output(9)) AND mux_669_nl;
  nor_438_nl <= NOT((fsm_output(9)) OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("111"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR nand_190_cse);
  mux_670_nl <= MUX_s_1_2_2(and_404_nl, nor_438_nl, fsm_output(8));
  mux_674_nl <= MUX_s_1_2_2(nor_433_nl, mux_670_nl, fsm_output(1));
  nor_439_nl <= NOT((NOT (VEC_LOOP_j_sva_11_0(2))) OR (NOT (fsm_output(5))) OR (NOT
      (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(7)));
  nand_237_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111")) AND
      (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(7)));
  or_789_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND (NOT (fsm_output(3))))) OR not_tmp_165;
  mux_665_nl <= MUX_s_1_2_2(nand_237_nl, or_789_nl, fsm_output(2));
  nor_440_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(0)) OR mux_665_nl);
  mux_666_nl <= MUX_s_1_2_2(nor_439_nl, nor_440_nl, fsm_output(9));
  and_405_nl <= (fsm_output(9)) AND CONV_SL_1_1(z_out_3(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111"))
      AND (NOT (fsm_output(5))) AND (fsm_output(0)) AND (fsm_output(2)) AND (fsm_output(3))
      AND (NOT (fsm_output(6))) AND (NOT (fsm_output(7)));
  mux_667_nl <= MUX_s_1_2_2(mux_666_nl, and_405_nl, fsm_output(8));
  nand_139_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111")) AND
      (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(7))));
  nand_231_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm AND (NOT (fsm_output(3))) AND (NOT
      (fsm_output(6))) AND (fsm_output(7)));
  mux_662_nl <= MUX_s_1_2_2(nand_139_nl, nand_231_nl, fsm_output(2));
  or_784_nl <= (fsm_output(0)) OR mux_662_nl;
  nor_442_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)) OR nand_168_cse);
  mux_661_nl <= MUX_s_1_2_2(nor_442_nl, and_494_cse, fsm_output(2));
  nand_36_nl <= NOT((fsm_output(0)) AND mux_661_nl);
  mux_663_nl <= MUX_s_1_2_2(or_784_nl, nand_36_nl, fsm_output(5));
  or_776_nl <= (fsm_output(5)) OR (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(3))
      OR CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("111")) OR CONV_SL_1_1(fsm_output(7
      DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_664_nl <= MUX_s_1_2_2(mux_663_nl, or_776_nl, fsm_output(9));
  nor_441_nl <= NOT((fsm_output(8)) OR mux_664_nl);
  mux_668_nl <= MUX_s_1_2_2(mux_667_nl, nor_441_nl, fsm_output(1));
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_674_nl, mux_668_nl,
      fsm_output(4));
  and_dcpl <= (NOT (fsm_output(6))) AND (fsm_output(0));
  and_511_cse <= (fsm_output(4)) AND (NOT (fsm_output(1))) AND (NOT (fsm_output(3)))
      AND nor_393_cse AND (NOT (fsm_output(7))) AND (fsm_output(5)) AND (NOT (fsm_output(2)))
      AND and_dcpl;
  and_dcpl_236 <= (fsm_output(6)) AND (NOT (fsm_output(0)));
  and_dcpl_238 <= NOT((fsm_output(7)) OR (fsm_output(5)) OR (fsm_output(2)));
  and_dcpl_240 <= (fsm_output(4)) AND (fsm_output(1));
  and_dcpl_242 <= and_dcpl_240 AND (fsm_output(3)) AND nor_393_cse;
  and_dcpl_243 <= and_dcpl_242 AND and_dcpl_238 AND and_dcpl_236;
  and_dcpl_245 <= (fsm_output(7)) AND (fsm_output(5)) AND (fsm_output(2));
  and_dcpl_247 <= and_dcpl_242 AND and_dcpl_245 AND and_dcpl;
  and_dcpl_255 <= (NOT (fsm_output(4))) AND (NOT (fsm_output(1))) AND (fsm_output(3))
      AND and_dcpl_11 AND (fsm_output(7)) AND (NOT (fsm_output(5))) AND (NOT (fsm_output(2)))
      AND and_dcpl;
  and_dcpl_260 <= (NOT (fsm_output(4))) AND (fsm_output(1)) AND (fsm_output(3)) AND
      and_dcpl_11 AND and_dcpl_245 AND and_dcpl_236;
  and_dcpl_266 <= and_dcpl_240 AND (NOT (fsm_output(3))) AND (fsm_output(9)) AND
      (NOT (fsm_output(8))) AND and_dcpl_238 AND (fsm_output(6)) AND (fsm_output(0));
  and_dcpl_268 <= (fsm_output(7)) AND (fsm_output(5));
  and_dcpl_269 <= and_dcpl_268 AND (fsm_output(2));
  and_dcpl_276 <= NOT((fsm_output(6)) OR (fsm_output(0)));
  and_dcpl_298 <= NOT((fsm_output(7)) OR (fsm_output(5)));
  and_dcpl_324 <= nor_tmp AND (NOT (fsm_output(1))) AND (fsm_output(9)) AND (NOT
      (fsm_output(8))) AND (fsm_output(7)) AND (fsm_output(5)) AND (NOT (fsm_output(2)))
      AND (NOT (fsm_output(6))) AND (NOT (fsm_output(0)));
  and_dcpl_340 <= (NOT (fsm_output(4))) AND (NOT (fsm_output(3))) AND (NOT (fsm_output(1)))
      AND nor_393_cse AND and_dcpl_238 AND and_dcpl;
  and_dcpl_345 <= nor_tmp AND (fsm_output(1)) AND nor_393_cse AND and_dcpl_238 AND
      (fsm_output(6)) AND (NOT (fsm_output(0)));
  and_dcpl_347 <= (NOT (fsm_output(7))) AND (fsm_output(5));
  and_dcpl_349 <= and_dcpl_347 AND (NOT (fsm_output(2))) AND and_dcpl;
  and_dcpl_354 <= and_dcpl_63 AND (NOT (fsm_output(1))) AND nor_393_cse AND and_dcpl_349;
  or_tmp_1317 <= (fsm_output(1)) OR (fsm_output(9)) OR (NOT (fsm_output(4))) OR (NOT
      (fsm_output(3))) OR (fsm_output(8));
  or_1440_cse <= (fsm_output(1)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(4)))
      OR (fsm_output(3)) OR (fsm_output(8));
  nor_635_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(5))) OR (fsm_output(0))
      OR (NOT (fsm_output(1))) OR (fsm_output(9)) OR (fsm_output(4)) OR (fsm_output(3))
      OR (NOT (fsm_output(8))));
  nor_636_nl <= NOT((fsm_output(6)) OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR
      (fsm_output(1)) OR (NOT (fsm_output(9))) OR (fsm_output(4)) OR (NOT (fsm_output(3)))
      OR (fsm_output(8)));
  mux_1347_nl <= MUX_s_1_2_2(nor_635_nl, nor_636_nl, fsm_output(2));
  mux_1345_nl <= MUX_s_1_2_2(or_tmp_1317, or_1440_cse, fsm_output(0));
  nor_637_nl <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1345_nl);
  or_1438_nl <= (NOT (fsm_output(0))) OR (NOT (fsm_output(1))) OR (fsm_output(9))
      OR (fsm_output(4)) OR (fsm_output(3)) OR (NOT (fsm_output(8)));
  or_1436_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(4)))
      OR (fsm_output(3)) OR (fsm_output(8));
  mux_1372_nl <= MUX_s_1_2_2(or_1436_nl, or_tmp_1317, fsm_output(0));
  mux_1344_nl <= MUX_s_1_2_2(or_1438_nl, mux_1372_nl, fsm_output(5));
  and_nl <= (fsm_output(6)) AND (NOT mux_1344_nl);
  mux_1346_nl <= MUX_s_1_2_2(nor_637_nl, and_nl, fsm_output(2));
  not_tmp_581 <= MUX_s_1_2_2(mux_1347_nl, mux_1346_nl, fsm_output(7));
  and_dcpl_357 <= and_dcpl_298 AND (NOT (fsm_output(2)));
  and_dcpl_362 <= and_dcpl_110 AND nor_393_cse AND and_dcpl_357 AND and_dcpl_276;
  and_dcpl_364 <= and_dcpl_357 AND and_dcpl_236;
  and_dcpl_367 <= and_dcpl_59 AND nor_393_cse;
  and_dcpl_368 <= and_dcpl_367 AND and_dcpl_364;
  and_dcpl_372 <= and_dcpl_367 AND and_dcpl_269 AND and_dcpl;
  and_dcpl_379 <= (NOT (fsm_output(3))) AND (NOT (fsm_output(4))) AND (NOT (fsm_output(1)))
      AND and_dcpl_11 AND and_dcpl_347 AND (fsm_output(2)) AND and_dcpl_276;
  and_dcpl_383 <= and_dcpl_100 AND (NOT (fsm_output(1)));
  and_dcpl_385 <= and_dcpl_383 AND and_dcpl_11 AND (fsm_output(7)) AND (NOT (fsm_output(5)))
      AND (NOT (fsm_output(2))) AND and_dcpl;
  and_dcpl_388 <= and_dcpl_110 AND and_dcpl_11 AND and_dcpl_269 AND and_dcpl_236;
  and_dcpl_394 <= and_dcpl_121 AND and_dcpl_23 AND and_dcpl_357 AND (fsm_output(6))
      AND (fsm_output(0));
  and_dcpl_399 <= and_dcpl_128 AND and_dcpl_23 AND and_dcpl_268 AND (NOT (fsm_output(2)))
      AND and_dcpl_276;
  and_dcpl_404 <= and_dcpl_128 AND and_369_cse AND and_dcpl_298 AND (fsm_output(2))
      AND and_dcpl;
  and_dcpl_406 <= and_dcpl_59 AND and_369_cse AND and_dcpl_364;
  and_dcpl_409 <= and_dcpl_383 AND nor_393_cse AND and_dcpl_357 AND and_dcpl;
  and_dcpl_411 <= and_dcpl_121 AND nor_393_cse AND and_dcpl_349;
  or_tmp_1346 <= (fsm_output(8)) OR (NOT((fsm_output(2)) AND (fsm_output(9)) AND
      (fsm_output(4)) AND (fsm_output(0))));
  or_tmp_1348 <= (NOT (fsm_output(8))) OR (fsm_output(2)) OR (fsm_output(9)) OR (fsm_output(4))
      OR (NOT (fsm_output(0)));
  or_tmp_1349 <= (NOT (fsm_output(7))) OR (fsm_output(8)) OR (fsm_output(2)) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(4))) OR (fsm_output(0));
  not_tmp_600 <= NOT((fsm_output(4)) AND (fsm_output(0)));
  operator_64_false_1_or_4_ssc <= and_dcpl_354 OR not_tmp_581 OR and_dcpl_362 OR
      and_dcpl_409 OR and_dcpl_411;
  operator_64_false_1_or_5_ssc <= and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385 OR
      and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404;
  or_tmp_1365 <= (fsm_output(6)) OR (NOT (fsm_output(3)));
  mux_tmp <= MUX_s_1_2_2(or_tmp_1365, (fsm_output(6)), fsm_output(1));
  or_tmp_1367 <= (fsm_output(6)) OR (fsm_output(3));
  nor_tmp_292 <= (fsm_output(6)) AND (fsm_output(3));
  mux_tmp_1374 <= MUX_s_1_2_2(nor_tmp_292, (fsm_output(6)), fsm_output(4));
  mux_tmp_1377 <= MUX_s_1_2_2((NOT (fsm_output(3))), (fsm_output(3)), fsm_output(6));
  mux_tmp_1378 <= MUX_s_1_2_2(mux_tmp_1377, or_tmp_1365, or_838_cse);
  or_tmp_1370 <= (NOT (fsm_output(6))) OR (fsm_output(3));
  nor_tmp_296 <= (fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(3));
  or_tmp_1374 <= and_389_cse OR (fsm_output(6)) OR (fsm_output(3));
  mux_tmp_1399 <= MUX_s_1_2_2((fsm_output(6)), or_tmp_1367, fsm_output(1));
  or_tmp_1389 <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 5)=STD_LOGIC_VECTOR'("0111")));
  or_tmp_1394 <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 7)/=STD_LOGIC_VECTOR'("01"));
  nor_tmp_301 <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11"));
  or_tmp_1401 <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100"));
  COMP_LOOP_or_40_itm <= and_dcpl_243 OR and_dcpl_247 OR and_dcpl_255 OR and_dcpl_260
      OR and_dcpl_266;
  operator_64_false_1_or_1_itm <= and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR
      and_dcpl_385 OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404
      OR and_dcpl_406;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( not_tmp_131 = '0' ) THEN
        p_sva <= p_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( ((and_dcpl_51 AND and_dcpl_14 AND and_dcpl_48) OR STAGE_LOOP_i_3_0_sva_mx0c1)
          = '1' ) THEN
        STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'( "0001"), STAGE_LOOP_i_3_0_sva_2,
            STAGE_LOOP_i_3_0_sva_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( not_tmp_131 = '0' ) THEN
        r_sva <= r_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_vec_rsc_triosy_0_7_obj_ld_cse <= '0';
        COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= '0';
        modExp_exp_1_0_1_sva_1 <= '0';
        modExp_exp_1_7_1_sva <= '0';
        modExp_exp_1_2_1_sva <= '0';
        modExp_exp_1_1_1_sva <= '0';
        COMP_LOOP_COMP_LOOP_nor_1_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_12_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_124_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_125_itm <= '0';
      ELSE
        reg_vec_rsc_triosy_0_7_obj_ld_cse <= and_dcpl_59 AND and_dcpl_58 AND (fsm_output(6))
            AND and_dcpl_140 AND CONV_SL_1_1(fsm_output(9 DOWNTO 8)=STD_LOGIC_VECTOR'("11"))
            AND (NOT STAGE_LOOP_acc_itm_2_1);
        COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= (COMP_LOOP_mux1h_31_nl AND (mux_987_nl
            OR (fsm_output(0)))) OR (mux_1035_nl AND (fsm_output(0)));
        modExp_exp_1_0_1_sva_1 <= (COMP_LOOP_mux_nl AND (NOT(mux_1196_nl AND (fsm_output(1)))))
            OR (NOT(mux_1249_nl OR (fsm_output(1))));
        modExp_exp_1_7_1_sva <= COMP_LOOP_mux1h_52_nl AND mux_1285_nl;
        modExp_exp_1_2_1_sva <= COMP_LOOP_mux1h_66_nl AND (NOT and_dcpl_226);
        modExp_exp_1_1_1_sva <= (COMP_LOOP_mux1h_68_nl AND (mux_1323_nl OR (fsm_output(9))))
            OR mux_1326_nl;
        COMP_LOOP_COMP_LOOP_nor_1_itm <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_12_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_12_cse,
            COMP_LOOP_COMP_LOOP_and_11_cse, modExp_while_or_cse);
        COMP_LOOP_COMP_LOOP_and_124_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_13_cse,
            COMP_LOOP_COMP_LOOP_and_12_cse, modExp_while_or_cse);
        COMP_LOOP_COMP_LOOP_and_125_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_37_cse,
            COMP_LOOP_COMP_LOOP_and_13_cse, modExp_while_or_cse);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      modulo_result_rem_cmp_a <= MUX1HOT_v_64_5_2(z_out_4, operator_64_false_acc_mut_63_0,
          COMP_LOOP_1_acc_8_itm, COMP_LOOP_1_mul_mut, COMP_LOOP_1_acc_5_mut_mx0w5,
          STD_LOGIC_VECTOR'( modulo_result_or_nl & (NOT mux_728_nl) & mux_775_nl
          & mux_795_nl & not_tmp_312));
      modulo_result_rem_cmp_b <= p_sva;
      operator_66_true_div_cmp_a <= MUX_v_65_2_2(z_out_2, (operator_64_false_acc_mut_64
          & operator_64_false_acc_mut_63_0), and_dcpl_152);
      operator_66_true_div_cmp_b_9_0 <= MUX_v_10_2_2(STAGE_LOOP_lshift_psp_sva_mx0w0,
          STAGE_LOOP_lshift_psp_sva, and_dcpl_152);
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(nor_659_nl, and_704_nl, fsm_output(9))) = '1' ) THEN
        STAGE_LOOP_lshift_psp_sva <= STAGE_LOOP_lshift_psp_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mux_1423_nl = '0' ) THEN
        operator_64_false_acc_mut_64 <= operator_64_false_mux1h_2_rgt(64);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_1453_nl, mux_1437_nl, fsm_output(2))) = '1' ) THEN
        operator_64_false_acc_mut_63_0 <= operator_64_false_mux1h_2_rgt(63 DOWNTO
            0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        VEC_LOOP_j_sva_11_0 <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (and_dcpl_156 OR VEC_LOOP_j_sva_11_0_mx0c1) = '1' ) THEN
        VEC_LOOP_j_sva_11_0 <= MUX_v_12_2_2(STD_LOGIC_VECTOR'("000000000000"), (z_out_3(11
            DOWNTO 0)), VEC_LOOP_j_sva_11_0_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_k_9_3_sva_5_0 <= STD_LOGIC_VECTOR'( "000000");
      ELSIF ( (NOT(mux_1457_nl OR (fsm_output(7)))) = '1' ) THEN
        COMP_LOOP_k_9_3_sva_5_0 <= MUX_v_6_2_2(STD_LOGIC_VECTOR'("000000"), (COMP_LOOP_k_9_3_sva_2(5
            DOWNTO 0)), nand_263_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( ((modExp_while_and_3 OR modExp_while_and_5 OR modExp_result_sva_mx0c0
          OR (NOT mux_885_nl)) AND (modExp_result_sva_mx0c0 OR modExp_result_and_rgt
          OR modExp_result_and_1_rgt)) = '1' ) THEN
        modExp_result_sva <= MUX1HOT_v_64_3_2(STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000001"),
            modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w1, STD_LOGIC_VECTOR'( modExp_result_sva_mx0c0
            & modExp_result_and_rgt & modExp_result_and_1_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        tmp_10_lpi_4_dfm <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
      ELSIF ( (MUX_s_1_2_2((NOT mux_913_nl), mux_896_nl, fsm_output(9))) = '1' )
          THEN
        tmp_10_lpi_4_dfm <= MUX1HOT_v_64_9_2(('0' & operator_64_false_slc_modExp_exp_63_1_3),
            vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d,
            vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_6_i_qa_d, vec_rsc_0_7_i_qa_d,
            STD_LOGIC_VECTOR'( and_dcpl_156 & COMP_LOOP_or_15_nl & COMP_LOOP_or_16_nl
            & COMP_LOOP_or_17_nl & COMP_LOOP_or_18_nl & COMP_LOOP_or_19_nl & COMP_LOOP_or_20_nl
            & COMP_LOOP_or_21_nl & COMP_LOOP_or_22_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_971_nl, mux_945_nl, fsm_output(9))) = '1' ) THEN
        COMP_LOOP_1_mul_mut <= MUX1HOT_v_64_13_2(r_sva, modulo_result_rem_cmp_z,
            modulo_qr_sva_1_mx0w1, modExp_result_sva, vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d,
            vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d, vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d,
            vec_rsc_0_6_i_qa_d, vec_rsc_0_7_i_qa_d, z_out_4, STD_LOGIC_VECTOR'( and_238_nl
            & COMP_LOOP_or_26_nl & COMP_LOOP_or_27_nl & not_tmp_374 & COMP_LOOP_or_7_nl
            & COMP_LOOP_or_8_nl & COMP_LOOP_or_9_nl & COMP_LOOP_or_10_nl & COMP_LOOP_or_11_nl
            & COMP_LOOP_or_12_nl & COMP_LOOP_or_13_nl & COMP_LOOP_or_14_nl & mux_48_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_11_itm <= '0';
      ELSIF ( (and_dcpl_147 OR and_dcpl_219 OR and_dcpl_69 OR and_dcpl_84 OR and_dcpl_93
          OR and_dcpl_103 OR and_dcpl_112 OR and_dcpl_123 OR and_dcpl_130 OR and_dcpl_138)
          = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_11_itm <= MUX1HOT_s_1_4_2((NOT (z_out_3(63))), (NOT
            (z_out_3(8))), COMP_LOOP_COMP_LOOP_and_11_cse, COMP_LOOP_COMP_LOOP_and_37_cse,
            STD_LOGIC_VECTOR'( and_dcpl_147 & and_dcpl_219 & and_dcpl_69 & modExp_while_or_cse));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_1139_nl OR not_tmp_312) = '1' ) THEN
        COMP_LOOP_1_acc_8_itm <= MUX_v_64_2_2(z_out_4, STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(COMP_LOOP_1_acc_8_nl),
            64)), not_tmp_312);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (NOT(CONV_SL_1_1(fsm_output/=STD_LOGIC_VECTOR'("0000110001")))) = '1'
          ) THEN
        COMP_LOOP_acc_psp_sva <= COMP_LOOP_acc_psp_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_2_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (NOT(mux_1156_nl AND nor_393_cse)) = '1' ) THEN
        COMP_LOOP_acc_1_cse_2_sva <= COMP_LOOP_acc_1_cse_2_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_4_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_86_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_30_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_89_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_32_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_33_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_34_itm <= '0';
      ELSIF ( mux_1158_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_4_itm <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_86_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva_1(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("011"));
        COMP_LOOP_COMP_LOOP_and_30_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_mx0w0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("011"));
        COMP_LOOP_COMP_LOOP_and_89_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva_1(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("110"));
        COMP_LOOP_COMP_LOOP_and_32_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_mx0w0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("101"));
        COMP_LOOP_COMP_LOOP_and_33_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_mx0w0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("110"));
        COMP_LOOP_COMP_LOOP_and_34_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_mx0w0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_145_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_1174_nl, mux_1173_nl, fsm_output(4))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_145_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_145_nl,
            (NOT (COMP_LOOP_1_acc_nl(9))), and_dcpl_138);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_6_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (MUX_s_1_2_2(mux_tmp_1178, mux_1181_nl, and_314_cse)) = '1' ) THEN
        COMP_LOOP_acc_1_cse_6_sva <= COMP_LOOP_acc_1_cse_6_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_4_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (NOT(mux_1184_nl AND (NOT (fsm_output(9))))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_4_sva <= COMP_LOOP_acc_1_cse_4_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_11_psp_sva <= STD_LOGIC_VECTOR'( "00000000000");
      ELSIF ( (NOT(mux_1186_nl AND (NOT (fsm_output(9))))) = '1' ) THEN
        COMP_LOOP_acc_11_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0(11
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_3_sva_5_0
            & STD_LOGIC_VECTOR'( "01")), 8), 11), 11));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_13_psp_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(not_tmp_480, or_1200_nl, fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_13_psp_sva <= z_out;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_14_psp_sva <= STD_LOGIC_VECTOR'( "00000000000");
      ELSIF ( (MUX_s_1_2_2(not_tmp_480, or_1201_nl, fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_14_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0(11
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_3_sva_5_0
            & STD_LOGIC_VECTOR'( "11")), 8), 11), 11));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (MUX_s_1_2_2(mux_1192_nl, and_369_cse, fsm_output(7))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_sva <= z_out_2(11 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        modExp_exp_1_6_1_sva <= '0';
        modExp_exp_1_5_1_sva <= '0';
        modExp_exp_1_4_1_sva <= '0';
        modExp_exp_1_3_1_sva <= '0';
      ELSIF ( mux_1273_itm = '1' ) THEN
        modExp_exp_1_6_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_3_sva_5_0(3)), modExp_exp_1_7_1_sva,
            (COMP_LOOP_k_9_3_sva_5_0(4)), STD_LOGIC_VECTOR'( and_dcpl_226 & not_tmp_523
            & not_tmp_513));
        modExp_exp_1_5_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_3_sva_5_0(2)), modExp_exp_1_6_1_sva,
            (COMP_LOOP_k_9_3_sva_5_0(3)), STD_LOGIC_VECTOR'( and_dcpl_226 & not_tmp_523
            & not_tmp_513));
        modExp_exp_1_4_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_3_sva_5_0(1)), modExp_exp_1_5_1_sva,
            (COMP_LOOP_k_9_3_sva_5_0(2)), STD_LOGIC_VECTOR'( and_dcpl_226 & not_tmp_523
            & not_tmp_513));
        modExp_exp_1_3_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_3_sva_5_0(0)), modExp_exp_1_4_1_sva,
            (COMP_LOOP_k_9_3_sva_5_0(1)), STD_LOGIC_VECTOR'( and_dcpl_226 & not_tmp_523
            & not_tmp_513));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_12_1_1_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( COMP_LOOP_or_2_cse = '1' ) THEN
        COMP_LOOP_acc_10_cse_12_1_1_sva <= z_out_3(12 DOWNTO 1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (and_dcpl_69 OR not_tmp_315 OR and_dcpl_84 OR and_dcpl_103 OR and_dcpl_112
          OR and_dcpl_123) = '1' ) THEN
        COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm <= MUX_s_1_2_2((z_out(9)), (z_out_3(8)),
            not_tmp_315);
      END IF;
    END IF;
  END PROCESS;
  or_864_nl <= (fsm_output(9)) OR (fsm_output(0)) OR (fsm_output(5)) OR (NOT (fsm_output(2)))
      OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_780_nl <= MUX_s_1_2_2(mux_tmp_776, or_864_nl, fsm_output(3));
  or_862_nl <= (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(0)) OR (NOT (fsm_output(5)))
      OR (fsm_output(2)) OR not_tmp_297;
  mux_781_nl <= MUX_s_1_2_2(mux_780_nl, or_862_nl, fsm_output(8));
  and_388_nl <= (fsm_output(6)) AND (NOT mux_781_nl);
  or_859_nl <= (fsm_output(9)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5)))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_857_nl <= (NOT (fsm_output(9))) OR (fsm_output(0)) OR (NOT (fsm_output(5)))
      OR (fsm_output(2)) OR not_tmp_297;
  mux_778_nl <= MUX_s_1_2_2(or_859_nl, or_857_nl, fsm_output(3));
  or_855_nl <= (fsm_output(9)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT
      (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(4));
  mux_777_nl <= MUX_s_1_2_2(or_855_nl, mux_tmp_776, fsm_output(3));
  mux_779_nl <= MUX_s_1_2_2(mux_778_nl, mux_777_nl, fsm_output(8));
  nor_422_nl <= NOT((fsm_output(6)) OR mux_779_nl);
  mux_782_nl <= MUX_s_1_2_2(and_388_nl, nor_422_nl, fsm_output(1));
  modulo_result_or_nl <= and_dcpl_147 OR not_tmp_315 OR mux_782_nl;
  mux_723_nl <= MUX_s_1_2_2(or_tmp_788, nor_tmp, fsm_output(5));
  mux_724_nl <= MUX_s_1_2_2(mux_723_nl, mux_tmp_722, fsm_output(6));
  mux_720_nl <= MUX_s_1_2_2((NOT mux_tmp_719), (fsm_output(4)), fsm_output(5));
  mux_721_nl <= MUX_s_1_2_2(mux_720_nl, mux_tmp_718, fsm_output(6));
  mux_725_nl <= MUX_s_1_2_2(mux_724_nl, mux_721_nl, fsm_output(2));
  mux_715_nl <= MUX_s_1_2_2(and_dcpl_51, or_tmp_788, fsm_output(5));
  mux_714_nl <= MUX_s_1_2_2((NOT nor_tmp), or_216_cse, fsm_output(5));
  mux_716_nl <= MUX_s_1_2_2((NOT mux_715_nl), mux_714_nl, fsm_output(6));
  nand_41_nl <= NOT((fsm_output(5)) AND (NOT mux_tmp_688));
  mux_712_nl <= MUX_s_1_2_2((NOT and_705_cse), or_tmp_103, fsm_output(5));
  mux_713_nl <= MUX_s_1_2_2(nand_41_nl, mux_712_nl, fsm_output(6));
  mux_717_nl <= MUX_s_1_2_2(mux_716_nl, mux_713_nl, fsm_output(2));
  mux_726_nl <= MUX_s_1_2_2((NOT mux_725_nl), mux_717_nl, fsm_output(7));
  mux_706_nl <= MUX_s_1_2_2(and_dcpl_50, nor_tmp, fsm_output(1));
  mux_707_nl <= MUX_s_1_2_2(mux_tmp_688, mux_706_nl, fsm_output(0));
  mux_708_nl <= MUX_s_1_2_2((fsm_output(4)), mux_707_nl, fsm_output(5));
  mux_709_nl <= MUX_s_1_2_2(mux_708_nl, mux_tmp_705, fsm_output(6));
  mux_703_nl <= MUX_s_1_2_2(and_dcpl_50, and_705_cse, fsm_output(5));
  mux_704_nl <= MUX_s_1_2_2(nor_tmp_146, mux_703_nl, fsm_output(6));
  mux_710_nl <= MUX_s_1_2_2(mux_709_nl, mux_704_nl, fsm_output(2));
  mux_700_nl <= MUX_s_1_2_2(or_216_cse, and_705_cse, fsm_output(5));
  mux_699_nl <= MUX_s_1_2_2((NOT and_dcpl_59), (fsm_output(4)), fsm_output(5));
  mux_701_nl <= MUX_s_1_2_2(mux_700_nl, mux_699_nl, fsm_output(6));
  mux_697_nl <= MUX_s_1_2_2((NOT mux_696_itm), (fsm_output(4)), fsm_output(5));
  mux_695_nl <= MUX_s_1_2_2((NOT nor_tmp), or_115_cse, fsm_output(5));
  mux_698_nl <= MUX_s_1_2_2(mux_697_nl, mux_695_nl, fsm_output(6));
  mux_702_nl <= MUX_s_1_2_2(mux_701_nl, mux_698_nl, fsm_output(2));
  mux_711_nl <= MUX_s_1_2_2((NOT mux_710_nl), mux_702_nl, fsm_output(7));
  mux_727_nl <= MUX_s_1_2_2(mux_726_nl, mux_711_nl, fsm_output(8));
  or_819_nl <= (fsm_output(5)) OR mux_tmp_156;
  mux_690_nl <= MUX_s_1_2_2(nor_tmp_23, mux_tmp_689, fsm_output(5));
  mux_691_nl <= MUX_s_1_2_2(or_819_nl, mux_690_nl, fsm_output(6));
  mux_686_nl <= MUX_s_1_2_2(nor_tmp_23, (NOT and_428_cse), fsm_output(5));
  mux_685_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), (fsm_output(4)), or_817_cse);
  mux_687_nl <= MUX_s_1_2_2(mux_686_nl, mux_685_nl, fsm_output(6));
  mux_692_nl <= MUX_s_1_2_2(mux_691_nl, mux_687_nl, fsm_output(2));
  nand_40_nl <= NOT((fsm_output(5)) AND (NOT mux_tmp_156));
  mux_683_nl <= MUX_s_1_2_2(nand_40_nl, or_816_cse, fsm_output(6));
  nand_39_nl <= NOT((fsm_output(5)) AND (NOT and_462_cse));
  or_815_nl <= (fsm_output(5)) OR (NOT or_tmp_113);
  mux_682_nl <= MUX_s_1_2_2(nand_39_nl, or_815_nl, fsm_output(6));
  mux_684_nl <= MUX_s_1_2_2(mux_683_nl, mux_682_nl, fsm_output(2));
  mux_693_nl <= MUX_s_1_2_2(mux_692_nl, mux_684_nl, fsm_output(7));
  mux_679_nl <= MUX_s_1_2_2(or_115_cse, and_462_cse, fsm_output(5));
  mux_680_nl <= MUX_s_1_2_2((NOT mux_679_nl), or_1202_cse, fsm_output(6));
  or_808_nl <= (fsm_output(5)) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(4));
  mux_678_nl <= MUX_s_1_2_2((NOT mux_tmp_677), or_808_nl, fsm_output(6));
  mux_681_nl <= MUX_s_1_2_2(mux_680_nl, mux_678_nl, fsm_output(2));
  or_813_nl <= (fsm_output(7)) OR mux_681_nl;
  mux_694_nl <= MUX_s_1_2_2(mux_693_nl, or_813_nl, fsm_output(8));
  mux_728_nl <= MUX_s_1_2_2(mux_727_nl, mux_694_nl, fsm_output(9));
  nand_130_nl <= NOT((fsm_output(6)) AND (fsm_output(1)) AND (fsm_output(2)));
  mux_770_nl <= MUX_s_1_2_2(nand_130_nl, (fsm_output(6)), fsm_output(5));
  nand_44_nl <= NOT((fsm_output(6)) AND not_tmp_274);
  mux_769_nl <= MUX_s_1_2_2(not_tmp_280, nand_44_nl, fsm_output(5));
  mux_771_nl <= MUX_s_1_2_2((NOT mux_770_nl), mux_769_nl, fsm_output(7));
  nor_423_nl <= NOT((fsm_output(6)) OR and_382_cse);
  mux_767_nl <= MUX_s_1_2_2(nor_423_nl, (fsm_output(6)), fsm_output(5));
  mux_768_nl <= MUX_s_1_2_2((NOT or_tmp_810), mux_767_nl, fsm_output(7));
  mux_772_nl <= MUX_s_1_2_2(mux_771_nl, mux_768_nl, fsm_output(4));
  or_850_nl <= (fsm_output(6)) OR (NOT or_1394_cse);
  mux_764_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), or_850_nl, fsm_output(5));
  mux_765_nl <= MUX_s_1_2_2((NOT mux_tmp_731), mux_764_nl, fsm_output(7));
  mux_762_nl <= MUX_s_1_2_2((NOT and_382_cse), or_1385_cse, fsm_output(6));
  nor_424_nl <= NOT((fsm_output(5)) OR mux_762_nl);
  mux_760_nl <= MUX_s_1_2_2((NOT (fsm_output(2))), (fsm_output(2)), fsm_output(1));
  and_167_nl <= (fsm_output(6)) AND mux_760_nl;
  mux_761_nl <= MUX_s_1_2_2((NOT or_tmp_792), and_167_nl, fsm_output(5));
  mux_763_nl <= MUX_s_1_2_2(nor_424_nl, mux_761_nl, fsm_output(7));
  mux_766_nl <= MUX_s_1_2_2(mux_765_nl, mux_763_nl, fsm_output(4));
  mux_773_nl <= MUX_s_1_2_2(mux_772_nl, mux_766_nl, fsm_output(3));
  nand_249_nl <= NOT((fsm_output(6)) AND or_1394_cse);
  mux_756_nl <= MUX_s_1_2_2((fsm_output(6)), nand_249_nl, fsm_output(5));
  or_848_nl <= (fsm_output(5)) OR (NOT (fsm_output(6))) OR (fsm_output(2));
  mux_757_nl <= MUX_s_1_2_2(mux_756_nl, or_848_nl, fsm_output(7));
  mux_754_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), nand_tmp_42, fsm_output(5));
  mux_753_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), or_tmp_792, fsm_output(5));
  mux_755_nl <= MUX_s_1_2_2(mux_754_nl, mux_753_nl, fsm_output(7));
  mux_758_nl <= MUX_s_1_2_2(mux_757_nl, mux_755_nl, fsm_output(4));
  or_847_nl <= (NOT (fsm_output(6))) OR (fsm_output(2));
  mux_750_nl <= MUX_s_1_2_2(or_847_nl, (fsm_output(6)), fsm_output(5));
  mux_751_nl <= MUX_s_1_2_2((NOT mux_750_nl), or_tmp_810, fsm_output(7));
  nand_43_nl <= NOT((NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("10"))))
      AND not_tmp_274);
  or_845_nl <= (NOT (fsm_output(6))) OR (fsm_output(1)) OR (fsm_output(2));
  mux_748_nl <= MUX_s_1_2_2(or_845_nl, (fsm_output(6)), fsm_output(5));
  mux_749_nl <= MUX_s_1_2_2(nand_43_nl, mux_748_nl, fsm_output(7));
  mux_752_nl <= MUX_s_1_2_2(mux_751_nl, mux_749_nl, fsm_output(4));
  mux_759_nl <= MUX_s_1_2_2(mux_758_nl, mux_752_nl, fsm_output(3));
  mux_774_nl <= MUX_s_1_2_2(mux_773_nl, (NOT mux_759_nl), fsm_output(8));
  or_843_nl <= (fsm_output(6)) OR (NOT (fsm_output(2)));
  mux_743_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), or_843_nl, fsm_output(5));
  mux_744_nl <= MUX_s_1_2_2(nor_425_cse, mux_743_nl, fsm_output(7));
  or_842_nl <= (fsm_output(6)) OR (NOT and_483_cse);
  mux_741_nl <= MUX_s_1_2_2(or_842_nl, (fsm_output(6)), fsm_output(5));
  mux_739_nl <= MUX_s_1_2_2((NOT (fsm_output(2))), (fsm_output(2)), and_389_cse);
  and_165_nl <= (fsm_output(6)) AND mux_739_nl;
  mux_740_nl <= MUX_s_1_2_2(not_tmp_280, and_165_nl, fsm_output(5));
  mux_742_nl <= MUX_s_1_2_2((NOT mux_741_nl), mux_740_nl, fsm_output(7));
  mux_745_nl <= MUX_s_1_2_2(mux_744_nl, mux_742_nl, fsm_output(4));
  mux_736_nl <= MUX_s_1_2_2((fsm_output(2)), (NOT (fsm_output(2))), or_838_cse);
  nor_426_nl <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01"))
      OR mux_736_nl);
  nor_427_nl <= NOT((fsm_output(6)) OR and_483_cse);
  mux_735_nl <= MUX_s_1_2_2(nor_427_nl, (fsm_output(6)), fsm_output(5));
  mux_737_nl <= MUX_s_1_2_2(nor_426_nl, mux_735_nl, fsm_output(7));
  mux_732_nl <= MUX_s_1_2_2(not_tmp_274, or_1394_cse, fsm_output(6));
  mux_733_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), mux_732_nl, fsm_output(5));
  mux_734_nl <= MUX_s_1_2_2(mux_733_nl, mux_tmp_731, fsm_output(7));
  mux_738_nl <= MUX_s_1_2_2(mux_737_nl, mux_734_nl, fsm_output(4));
  mux_746_nl <= MUX_s_1_2_2(mux_745_nl, mux_738_nl, fsm_output(3));
  nor_428_nl <= NOT((fsm_output(7)) OR (fsm_output(5)) OR (NOT nand_tmp_42));
  nor_429_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 5)/=STD_LOGIC_VECTOR'("010")));
  mux_729_nl <= MUX_s_1_2_2(nor_428_nl, nor_429_nl, fsm_output(4));
  nor_430_nl <= NOT((fsm_output(4)) OR (fsm_output(7)) OR (fsm_output(5)) OR (NOT
      or_tmp_792));
  mux_730_nl <= MUX_s_1_2_2(mux_729_nl, nor_430_nl, fsm_output(3));
  mux_747_nl <= MUX_s_1_2_2(mux_746_nl, mux_730_nl, fsm_output(8));
  mux_775_nl <= MUX_s_1_2_2(mux_774_nl, mux_747_nl, fsm_output(9));
  nor_411_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR (fsm_output(3)) OR and_389_cse
      OR (fsm_output(2)) OR (NOT (fsm_output(9))));
  and_380_nl <= (fsm_output(6)) AND (NOT((fsm_output(3)) AND or_1423_cse));
  nor_412_nl <= NOT((fsm_output(6)) OR (NOT((fsm_output(3)) OR or_1423_cse)));
  mux_792_nl <= MUX_s_1_2_2(and_380_nl, nor_412_nl, fsm_output(8));
  mux_793_nl <= MUX_s_1_2_2(nor_411_nl, mux_792_nl, fsm_output(5));
  and_381_nl <= (fsm_output(1)) AND (fsm_output(2)) AND (fsm_output(9));
  or_881_nl <= and_382_cse OR (fsm_output(9));
  mux_790_nl <= MUX_s_1_2_2(and_381_nl, or_881_nl, fsm_output(3));
  nor_414_nl <= NOT((fsm_output(8)) OR (NOT((fsm_output(6)) AND mux_790_nl)));
  and_383_nl <= or_1391_cse AND (fsm_output(9));
  or_877_nl <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(9));
  mux_789_nl <= MUX_s_1_2_2(and_383_nl, or_877_nl, fsm_output(3));
  nor_415_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(6)) OR mux_789_nl);
  mux_791_nl <= MUX_s_1_2_2(nor_414_nl, nor_415_nl, fsm_output(5));
  mux_794_nl <= MUX_s_1_2_2(mux_793_nl, mux_791_nl, fsm_output(4));
  nand_127_nl <= NOT(or_838_cse AND (fsm_output(2)) AND (fsm_output(9)));
  mux_786_nl <= MUX_s_1_2_2(or_1392_cse, nand_127_nl, fsm_output(3));
  nand_47_nl <= NOT((fsm_output(6)) AND mux_786_nl);
  or_872_nl <= (fsm_output(6)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(2)))
      OR (fsm_output(9));
  mux_787_nl <= MUX_s_1_2_2(nand_47_nl, or_872_nl, fsm_output(8));
  nor_416_nl <= NOT((fsm_output(5)) OR mux_787_nl);
  nor_417_nl <= NOT((NOT (fsm_output(6))) OR (fsm_output(3)) OR (fsm_output(2)) OR
      (fsm_output(9)));
  nor_418_nl <= NOT((fsm_output(6)) OR (CONV_SL_1_1(fsm_output(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111")))
      OR (fsm_output(9)));
  mux_784_nl <= MUX_s_1_2_2(nor_417_nl, nor_418_nl, fsm_output(8));
  nor_419_nl <= NOT((fsm_output(6)) OR (NOT((fsm_output(3)) AND or_1394_cse AND (fsm_output(9)))));
  and_386_nl <= (fsm_output(6)) AND (NOT((NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))))
      OR (fsm_output(9))));
  mux_783_nl <= MUX_s_1_2_2(nor_419_nl, and_386_nl, fsm_output(8));
  mux_785_nl <= MUX_s_1_2_2(mux_784_nl, mux_783_nl, fsm_output(5));
  mux_788_nl <= MUX_s_1_2_2(nor_416_nl, mux_785_nl, fsm_output(4));
  mux_795_nl <= MUX_s_1_2_2(mux_794_nl, mux_788_nl, fsm_output(7));
  COMP_LOOP_acc_12_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(9
      DOWNTO 3)))) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_3_sva_5_0
      & '0'), 7), 8) + UNSIGNED'( "00000001"), 8));
  COMP_LOOP_and_76_nl <= (NOT and_dcpl_162) AND and_dcpl_156;
  mux_1026_nl <= MUX_s_1_2_2((NOT or_816_cse), (fsm_output(4)), and_389_cse);
  mux_1027_nl <= MUX_s_1_2_2(mux_1026_nl, (fsm_output(4)), fsm_output(2));
  nor_205_nl <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110")));
  mux_1025_nl <= MUX_s_1_2_2((fsm_output(5)), or_816_cse, nor_205_nl);
  mux_1028_nl <= MUX_s_1_2_2(mux_1027_nl, (NOT mux_1025_nl), fsm_output(6));
  mux_1029_nl <= MUX_s_1_2_2(mux_1028_nl, nor_425_cse, fsm_output(7));
  or_1072_nl <= (NOT((NOT (fsm_output(1))) OR (fsm_output(5)))) OR (fsm_output(4));
  mux_1021_nl <= MUX_s_1_2_2(or_247_cse, mux_tmp_997, or_838_cse);
  mux_1022_nl <= MUX_s_1_2_2(or_1072_nl, mux_1021_nl, fsm_output(2));
  mux_1023_nl <= MUX_s_1_2_2(mux_1022_nl, (NOT mux_tmp_1006), fsm_output(6));
  mux_1019_nl <= MUX_s_1_2_2(or_171_cse, (NOT mux_tmp_997), and_483_cse);
  and_252_nl <= (fsm_output(2)) AND or_838_cse AND CONV_SL_1_1(fsm_output(5 DOWNTO
      4)=STD_LOGIC_VECTOR'("11"));
  mux_1020_nl <= MUX_s_1_2_2(mux_1019_nl, and_252_nl, fsm_output(6));
  mux_1024_nl <= MUX_s_1_2_2(mux_1023_nl, mux_1020_nl, fsm_output(7));
  mux_1030_nl <= MUX_s_1_2_2(mux_1029_nl, mux_1024_nl, fsm_output(3));
  and_340_nl <= (fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(5)) AND (NOT
      (fsm_output(4)));
  nor_351_nl <= NOT((fsm_output(0)) OR (fsm_output(1)) OR (NOT (fsm_output(5))) OR
      (fsm_output(4)));
  mux_1015_nl <= MUX_s_1_2_2(and_340_nl, nor_351_nl, fsm_output(2));
  nor_352_nl <= NOT((fsm_output(2)) OR (fsm_output(1)) OR (NOT (fsm_output(5))) OR
      (fsm_output(4)));
  mux_1016_nl <= MUX_s_1_2_2(mux_1015_nl, nor_352_nl, fsm_output(6));
  mux_1013_nl <= MUX_s_1_2_2(mux_tmp_997, and_314_cse, and_477_cse);
  mux_1014_nl <= MUX_s_1_2_2(or_171_cse, mux_1013_nl, fsm_output(6));
  mux_1017_nl <= MUX_s_1_2_2(mux_1016_nl, mux_1014_nl, fsm_output(7));
  mux_1011_nl <= MUX_s_1_2_2(and_314_cse, (fsm_output(5)), or_838_cse);
  mux_1012_nl <= MUX_s_1_2_2(and_314_cse, mux_1011_nl, fsm_output(2));
  and_251_nl <= (fsm_output(7)) AND (NOT((fsm_output(6)) AND (NOT mux_1012_nl)));
  mux_1018_nl <= MUX_s_1_2_2(mux_1017_nl, and_251_nl, fsm_output(3));
  mux_1031_nl <= MUX_s_1_2_2(mux_1030_nl, (NOT mux_1018_nl), fsm_output(8));
  mux_1007_nl <= MUX_s_1_2_2(and_314_cse, (NOT mux_tmp_1006), fsm_output(6));
  mux_1003_nl <= MUX_s_1_2_2((fsm_output(5)), or_171_cse, or_838_cse);
  mux_1002_nl <= MUX_s_1_2_2(or_171_cse, (NOT mux_tmp_997), and_389_cse);
  mux_1004_nl <= MUX_s_1_2_2(mux_1003_nl, mux_1002_nl, fsm_output(2));
  or_1061_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("10")) OR (NOT
      and_314_cse);
  mux_1005_nl <= MUX_s_1_2_2(mux_1004_nl, or_1061_nl, fsm_output(6));
  mux_1008_nl <= MUX_s_1_2_2(mux_1007_nl, mux_1005_nl, fsm_output(7));
  mux_999_nl <= MUX_s_1_2_2(and_314_cse, (fsm_output(5)), fsm_output(2));
  mux_1000_nl <= MUX_s_1_2_2(mux_999_nl, (NOT or_171_cse), fsm_output(6));
  mux_998_nl <= MUX_s_1_2_2((NOT mux_tmp_997), or_171_cse, or_1385_cse);
  or_1059_nl <= (fsm_output(6)) OR mux_998_nl;
  mux_1001_nl <= MUX_s_1_2_2(mux_1000_nl, or_1059_nl, fsm_output(7));
  mux_1009_nl <= MUX_s_1_2_2(mux_1008_nl, mux_1001_nl, fsm_output(3));
  nor_353_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 5)/=STD_LOGIC_VECTOR'("000")));
  mux_995_nl <= MUX_s_1_2_2((fsm_output(5)), or_171_cse, fsm_output(2));
  nor_354_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"))
      OR mux_995_nl);
  mux_996_nl <= MUX_s_1_2_2(nor_353_nl, nor_354_nl, fsm_output(3));
  mux_1010_nl <= MUX_s_1_2_2(mux_1009_nl, mux_996_nl, fsm_output(8));
  mux_1032_nl <= MUX_s_1_2_2(mux_1031_nl, mux_1010_nl, fsm_output(9));
  COMP_LOOP_mux1h_31_nl <= MUX1HOT_s_1_7_2((operator_66_true_div_cmp_z(0)), (tmp_10_lpi_4_dfm(0)),
      (z_out_3(6)), modExp_exp_1_0_1_sva_1, COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm,
      (COMP_LOOP_acc_12_nl(7)), (z_out_2(6)), STD_LOGIC_VECTOR'( COMP_LOOP_and_76_nl
      & and_dcpl_162 & and_dcpl_66 & not_tmp_414 & mux_1032_nl & and_dcpl_93 & and_dcpl_130));
  or_1432_nl <= (NOT (fsm_output(8))) OR (NOT (fsm_output(1))) OR (fsm_output(5))
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_406;
  or_1040_nl <= (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(7)))
      OR (fsm_output(2)) OR (fsm_output(6));
  or_1039_nl <= (NOT (fsm_output(3))) OR (fsm_output(9)) OR not_tmp_406;
  mux_985_nl <= MUX_s_1_2_2(or_1040_nl, or_1039_nl, fsm_output(5));
  or_1037_nl <= (NOT (fsm_output(5))) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(7))
      OR (fsm_output(2)) OR (fsm_output(6));
  mux_986_nl <= MUX_s_1_2_2(mux_985_nl, or_1037_nl, fsm_output(1));
  or_1433_nl <= (fsm_output(8)) OR mux_986_nl;
  mux_987_nl <= MUX_s_1_2_2(or_1432_nl, or_1433_nl, fsm_output(4));
  nand_108_nl <= NOT((fsm_output(9)) AND (fsm_output(3)) AND (fsm_output(1)) AND
      (NOT (fsm_output(6))) AND (fsm_output(5)));
  or_1082_nl <= (fsm_output(9)) OR (fsm_output(3)) OR (fsm_output(1)) OR not_tmp_436;
  mux_1034_nl <= MUX_s_1_2_2(nand_108_nl, or_1082_nl, fsm_output(8));
  nor_347_nl <= NOT((fsm_output(4)) OR (fsm_output(7)) OR mux_1034_nl);
  or_1078_nl <= (fsm_output(3)) OR (NOT (fsm_output(1))) OR (fsm_output(6)) OR (fsm_output(5));
  or_1077_nl <= (fsm_output(3)) OR (fsm_output(1)) OR not_tmp_436;
  mux_1033_nl <= MUX_s_1_2_2(or_1078_nl, or_1077_nl, fsm_output(9));
  nor_348_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(7))) OR (fsm_output(8))
      OR mux_1033_nl);
  mux_1035_nl <= MUX_s_1_2_2(nor_347_nl, nor_348_nl, fsm_output(2));
  nor_316_nl <= NOT((fsm_output(5)) OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR
      (NOT (fsm_output(8))) OR (fsm_output(4)));
  nor_317_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR
      nand_100_cse);
  mux_1243_nl <= MUX_s_1_2_2(nor_316_nl, nor_317_nl, fsm_output(9));
  nor_318_nl <= NOT((fsm_output(9)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(2)))
      OR (NOT (fsm_output(7))) OR (fsm_output(8)) OR (NOT (fsm_output(4))));
  mux_1244_nl <= MUX_s_1_2_2(mux_1243_nl, nor_318_nl, fsm_output(1));
  and_306_nl <= (fsm_output(3)) AND mux_1244_nl;
  nor_319_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(8))
      OR (NOT (fsm_output(4))));
  mux_1245_nl <= MUX_s_1_2_2(and_306_nl, nor_319_nl, fsm_output(6));
  nor_320_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(2)) OR (fsm_output(7)) OR
      (NOT (fsm_output(8))) OR (fsm_output(4)));
  and_493_nl <= (fsm_output(5)) AND (fsm_output(2)) AND (fsm_output(7)) AND (NOT
      (fsm_output(8))) AND (fsm_output(4));
  mux_1241_nl <= MUX_s_1_2_2(nor_320_nl, and_493_nl, fsm_output(9));
  and_307_nl <= (NOT((fsm_output(3)) OR (NOT (fsm_output(1))))) AND mux_1241_nl;
  or_1229_nl <= (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(8)) OR (NOT (fsm_output(4)));
  nand_95_nl <= NOT((fsm_output(2)) AND (fsm_output(7)) AND (fsm_output(8)) AND (NOT
      (fsm_output(4))));
  mux_1240_nl <= MUX_s_1_2_2(or_1229_nl, nand_95_nl, fsm_output(5));
  nor_322_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(1)) OR (fsm_output(9)) OR
      mux_1240_nl);
  mux_1242_nl <= MUX_s_1_2_2(and_307_nl, nor_322_nl, fsm_output(6));
  mux_1246_nl <= MUX_s_1_2_2(mux_1245_nl, mux_1242_nl, fsm_output(0));
  COMP_LOOP_mux_nl <= MUX_s_1_2_2(modExp_exp_1_0_1_sva_1, modExp_exp_1_1_1_sva, mux_1246_nl);
  or_1210_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(4))
      OR (fsm_output(6)) OR (fsm_output(8));
  mux_1195_nl <= MUX_s_1_2_2(or_tmp_1159, or_1210_nl, fsm_output(0));
  nor_324_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR mux_1195_nl);
  or_1208_nl <= (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(4)) OR nand_97_cse;
  mux_1194_nl <= MUX_s_1_2_2(or_1208_nl, or_tmp_1159, fsm_output(0));
  nor_325_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR mux_1194_nl);
  mux_1196_nl <= MUX_s_1_2_2(nor_324_nl, nor_325_nl, fsm_output(2));
  or_1430_nl <= (fsm_output(7)) OR (NOT (fsm_output(8))) OR (fsm_output(9)) OR (NOT
      (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(3)) OR not_tmp_436;
  or_1245_nl <= (fsm_output(0)) OR (NOT((fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(5))
      AND (fsm_output(6))));
  or_1244_nl <= (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(5)) OR (fsm_output(6));
  or_1243_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_436;
  mux_1247_nl <= MUX_s_1_2_2(or_1244_nl, or_1243_nl, fsm_output(0));
  mux_1248_nl <= MUX_s_1_2_2(or_1245_nl, mux_1247_nl, fsm_output(9));
  or_1431_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01")) OR mux_1248_nl;
  mux_1249_nl <= MUX_s_1_2_2(or_1430_nl, or_1431_nl, fsm_output(4));
  COMP_LOOP_mux1h_52_nl <= MUX1HOT_s_1_4_2((COMP_LOOP_k_9_3_sva_5_0(4)), modExp_exp_1_1_1_sva,
      modExp_exp_1_7_1_sva, (COMP_LOOP_k_9_3_sva_5_0(5)), STD_LOGIC_VECTOR'( and_dcpl_226
      & and_dcpl_219 & (NOT mux_1273_itm) & not_tmp_513));
  nor_304_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(9)) OR (NOT (fsm_output(8)))
      OR (fsm_output(4)));
  nor_305_nl <= NOT((fsm_output(7)) OR nand_89_cse);
  mux_1283_nl <= MUX_s_1_2_2(nor_304_nl, nor_305_nl, fsm_output(2));
  nand_259_nl <= NOT((NOT((fsm_output(5)) OR (fsm_output(0)) OR (NOT (fsm_output(3)))))
      AND mux_1283_nl);
  nand_260_nl <= NOT((fsm_output(5)) AND (fsm_output(0)) AND (fsm_output(3)) AND
      (fsm_output(2)) AND (fsm_output(7)) AND (NOT (fsm_output(9))) AND (fsm_output(8))
      AND (NOT (fsm_output(4))));
  mux_1284_nl <= MUX_s_1_2_2(nand_259_nl, nand_260_nl, fsm_output(6));
  nor_306_nl <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(4))));
  or_1283_nl <= (fsm_output(7)) OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(4));
  nand_226_nl <= NOT((fsm_output(7)) AND (fsm_output(9)) AND (NOT (fsm_output(8)))
      AND (fsm_output(4)));
  mux_1280_nl <= MUX_s_1_2_2(or_1283_nl, nand_226_nl, fsm_output(2));
  nor_307_nl <= NOT((fsm_output(3)) OR mux_1280_nl);
  mux_1281_nl <= MUX_s_1_2_2(nor_306_nl, nor_307_nl, fsm_output(0));
  nand_261_nl <= NOT((fsm_output(5)) AND mux_1281_nl);
  or_1483_nl <= (fsm_output(5)) OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(2))
      OR (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(4)));
  mux_1282_nl <= MUX_s_1_2_2(nand_261_nl, or_1483_nl, fsm_output(6));
  mux_1285_nl <= MUX_s_1_2_2(mux_1284_nl, mux_1282_nl, fsm_output(1));
  COMP_LOOP_mux1h_66_nl <= MUX1HOT_s_1_3_2(modExp_exp_1_3_1_sva, modExp_exp_1_2_1_sva,
      (COMP_LOOP_k_9_3_sva_5_0(0)), STD_LOGIC_VECTOR'( not_tmp_523 & (NOT mux_1273_itm)
      & not_tmp_513));
  nand_86_nl <= NOT((fsm_output(3)) AND (fsm_output(2)) AND (fsm_output(9)) AND (NOT
      (fsm_output(6))));
  mux_1317_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), nand_86_nl, fsm_output(5));
  or_1323_nl <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01"));
  mux_1318_nl <= MUX_s_1_2_2(mux_1317_nl, or_1323_nl, fsm_output(7));
  nand_247_nl <= NOT((NOT(or_1391_cse AND (fsm_output(9)))) AND (fsm_output(6)));
  or_1366_nl <= (fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(0)) OR (fsm_output(9))
      OR (NOT (fsm_output(6)));
  mux_1314_nl <= MUX_s_1_2_2(nand_247_nl, or_1366_nl, fsm_output(3));
  or_1367_nl <= (NOT((fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(9)))) OR (fsm_output(6));
  mux_1315_nl <= MUX_s_1_2_2(mux_1314_nl, or_1367_nl, fsm_output(5));
  or_1316_nl <= (NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))))
      OR (NOT (fsm_output(9))) OR (fsm_output(6));
  mux_1312_nl <= MUX_s_1_2_2(or_1316_nl, (fsm_output(6)), fsm_output(3));
  mux_1309_nl <= MUX_s_1_2_2(or_tmp_1261, mux_tmp_1305, fsm_output(0));
  mux_1310_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), mux_1309_nl, and_483_cse);
  or_1314_nl <= (NOT (fsm_output(9))) OR (fsm_output(6));
  mux_1306_nl <= MUX_s_1_2_2(mux_tmp_1305, or_1314_nl, fsm_output(0));
  mux_1307_nl <= MUX_s_1_2_2(mux_1306_nl, (fsm_output(6)), fsm_output(1));
  mux_1308_nl <= MUX_s_1_2_2(mux_tmp_1305, mux_1307_nl, fsm_output(2));
  mux_1311_nl <= MUX_s_1_2_2(mux_1310_nl, mux_1308_nl, fsm_output(3));
  mux_1313_nl <= MUX_s_1_2_2(mux_1312_nl, (NOT mux_1311_nl), fsm_output(5));
  mux_1316_nl <= MUX_s_1_2_2(mux_1315_nl, mux_1313_nl, fsm_output(7));
  mux_1319_nl <= MUX_s_1_2_2(mux_1318_nl, mux_1316_nl, fsm_output(4));
  mux_1299_nl <= MUX_s_1_2_2((fsm_output(9)), or_tmp_1261, fsm_output(0));
  mux_1300_nl <= MUX_s_1_2_2(or_1099_cse, mux_1299_nl, fsm_output(1));
  mux_1301_nl <= MUX_s_1_2_2(mux_1300_nl, or_tmp_1261, or_1189_cse);
  mux_1302_nl <= MUX_s_1_2_2((fsm_output(6)), mux_1301_nl, fsm_output(5));
  mux_1296_nl <= MUX_s_1_2_2(or_1099_cse, (fsm_output(9)), and_477_cse);
  mux_1297_nl <= MUX_s_1_2_2(mux_1296_nl, or_tmp_1261, fsm_output(3));
  or_1311_nl <= (fsm_output(1)) OR (fsm_output(0)) OR (fsm_output(9)) OR (NOT (fsm_output(6)));
  mux_1295_nl <= MUX_s_1_2_2(or_tmp_1261, or_1311_nl, and_316_cse);
  mux_1298_nl <= MUX_s_1_2_2(mux_1297_nl, mux_1295_nl, fsm_output(5));
  mux_1303_nl <= MUX_s_1_2_2(mux_1302_nl, mux_1298_nl, fsm_output(7));
  or_1309_nl <= ((fsm_output(3)) AND (fsm_output(2)) AND (fsm_output(9))) OR (fsm_output(6));
  mux_1293_nl <= MUX_s_1_2_2(or_1309_nl, or_tmp_1261, fsm_output(5));
  or_1307_nl <= (fsm_output(5)) OR (fsm_output(9)) OR (NOT (fsm_output(6)));
  mux_1294_nl <= MUX_s_1_2_2(mux_1293_nl, or_1307_nl, fsm_output(7));
  mux_1304_nl <= MUX_s_1_2_2(mux_1303_nl, mux_1294_nl, fsm_output(4));
  mux_1320_nl <= MUX_s_1_2_2(mux_1319_nl, mux_1304_nl, fsm_output(8));
  COMP_LOOP_mux1h_68_nl <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_3_sva_5_0(5)), modExp_exp_1_2_1_sva,
      modExp_exp_1_1_1_sva, STD_LOGIC_VECTOR'( and_dcpl_226 & not_tmp_523 & (NOT
      mux_1320_nl)));
  or_1434_nl <= (NOT (fsm_output(8))) OR (fsm_output(3)) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(1))
      OR (NOT (fsm_output(6)));
  or_1329_nl <= (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(2)))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(1))) OR (fsm_output(6));
  or_1328_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(1))
      OR (NOT (fsm_output(6)));
  or_1326_nl <= (fsm_output(0)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR (fsm_output(1)) OR (NOT (fsm_output(6)));
  mux_1321_nl <= MUX_s_1_2_2(or_1328_nl, or_1326_nl, fsm_output(5));
  mux_1322_nl <= MUX_s_1_2_2(or_1329_nl, mux_1321_nl, fsm_output(3));
  or_1435_nl <= (fsm_output(8)) OR mux_1322_nl;
  mux_1323_nl <= MUX_s_1_2_2(or_1434_nl, or_1435_nl, fsm_output(4));
  nor_293_nl <= NOT((fsm_output(5)) OR (fsm_output(2)) OR (fsm_output(6)));
  and_283_nl <= (fsm_output(5)) AND (fsm_output(2)) AND (fsm_output(6));
  mux_1324_nl <= MUX_s_1_2_2(nor_293_nl, and_283_nl, fsm_output(0));
  nor_292_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT((fsm_output(7)) AND mux_1324_nl)));
  nor_294_nl <= NOT((fsm_output(4)) OR (NOT (fsm_output(3))) OR (fsm_output(7)) OR
      (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(2)) OR (fsm_output(6)));
  mux_1325_nl <= MUX_s_1_2_2(nor_292_nl, nor_294_nl, fsm_output(1));
  and_282_nl <= (fsm_output(9)) AND mux_1325_nl;
  nor_295_nl <= NOT((fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(4)) OR
      (fsm_output(3)) OR (NOT (fsm_output(7))) OR (fsm_output(0)) OR (fsm_output(5))
      OR (NOT((fsm_output(2)) AND (fsm_output(6)))));
  mux_1326_nl <= MUX_s_1_2_2(and_282_nl, nor_295_nl, fsm_output(8));
  nor_659_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 1)/=STD_LOGIC_VECTOR'("00000000")));
  and_176_nl <= (fsm_output(6)) AND ((fsm_output(5)) OR and_428_cse);
  mux_812_nl <= MUX_s_1_2_2(and_176_nl, and_491_cse, fsm_output(2));
  and_704_nl <= (fsm_output(8)) AND ((fsm_output(7)) OR mux_812_nl);
  or_1499_nl <= (NOT (fsm_output(1))) OR (fsm_output(6)) OR (fsm_output(3));
  mux_1418_nl <= MUX_s_1_2_2(mux_tmp_1399, or_1499_nl, fsm_output(0));
  or_1550_nl <= (fsm_output(4)) OR mux_1418_nl;
  mux_1417_nl <= MUX_s_1_2_2(or_tmp_1367, (NOT (fsm_output(3))), fsm_output(4));
  mux_1419_nl <= MUX_s_1_2_2(or_1550_nl, mux_1417_nl, fsm_output(2));
  mux_1415_nl <= MUX_s_1_2_2((NOT or_136_cse), (fsm_output(3)), fsm_output(4));
  and_707_nl <= (fsm_output(4)) AND or_tmp_1374;
  mux_1416_nl <= MUX_s_1_2_2(mux_1415_nl, and_707_nl, fsm_output(2));
  mux_1420_nl <= MUX_s_1_2_2(mux_1419_nl, mux_1416_nl, fsm_output(7));
  and_706_nl <= (fsm_output(4)) AND ((NOT (fsm_output(0))) OR (fsm_output(1)) OR
      (fsm_output(6)) OR (fsm_output(3)));
  or_1497_nl <= (fsm_output(4)) OR nor_tmp_296;
  mux_1413_nl <= MUX_s_1_2_2(and_706_nl, or_1497_nl, fsm_output(2));
  mux_1410_nl <= MUX_s_1_2_2(nor_tmp_292, (fsm_output(6)), fsm_output(1));
  mux_1411_nl <= MUX_s_1_2_2((NOT mux_1410_nl), or_tmp_1370, fsm_output(4));
  mux_1412_nl <= MUX_s_1_2_2((NOT mux_tmp_1374), mux_1411_nl, fsm_output(2));
  mux_1414_nl <= MUX_s_1_2_2(mux_1413_nl, mux_1412_nl, fsm_output(7));
  mux_1421_nl <= MUX_s_1_2_2(mux_1420_nl, mux_1414_nl, fsm_output(5));
  mux_1406_nl <= MUX_s_1_2_2(nor_tmp_296, (fsm_output(6)), fsm_output(4));
  mux_1407_nl <= MUX_s_1_2_2(mux_1406_nl, mux_tmp_1374, fsm_output(2));
  mux_1403_nl <= MUX_s_1_2_2(or_tmp_1370, mux_tmp_1377, and_389_cse);
  mux_1404_nl <= MUX_s_1_2_2(mux_1403_nl, (fsm_output(6)), fsm_output(4));
  mux_1401_nl <= MUX_s_1_2_2(mux_tmp_1377, or_tmp_1365, fsm_output(1));
  mux_1402_nl <= MUX_s_1_2_2(mux_1401_nl, mux_tmp_1399, fsm_output(4));
  mux_1405_nl <= MUX_s_1_2_2(mux_1404_nl, mux_1402_nl, fsm_output(2));
  mux_1408_nl <= MUX_s_1_2_2(mux_1407_nl, (NOT mux_1405_nl), fsm_output(7));
  mux_1396_nl <= MUX_s_1_2_2((fsm_output(6)), or_tmp_1367, or_838_cse);
  mux_1397_nl <= MUX_s_1_2_2(mux_tmp_1378, mux_1396_nl, fsm_output(4));
  mux_1395_nl <= MUX_s_1_2_2(mux_tmp, or_tmp_1367, fsm_output(4));
  mux_1398_nl <= MUX_s_1_2_2(mux_1397_nl, mux_1395_nl, fsm_output(2));
  mux_1399_nl <= MUX_s_1_2_2((NOT mux_1398_nl), (fsm_output(4)), fsm_output(7));
  mux_1409_nl <= MUX_s_1_2_2(mux_1408_nl, mux_1399_nl, fsm_output(5));
  mux_1422_nl <= MUX_s_1_2_2((NOT mux_1421_nl), mux_1409_nl, fsm_output(8));
  mux_1390_nl <= MUX_s_1_2_2((NOT or_tmp_1374), (fsm_output(3)), fsm_output(4));
  mux_1391_nl <= MUX_s_1_2_2(mux_1390_nl, and_705_cse, fsm_output(2));
  nand_275_nl <= NOT(or_838_cse AND (fsm_output(6)) AND (fsm_output(3)));
  mux_1388_nl <= MUX_s_1_2_2(nand_275_nl, nor_tmp_296, fsm_output(4));
  mux_1389_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), mux_1388_nl, fsm_output(2));
  mux_1392_nl <= MUX_s_1_2_2(mux_1391_nl, mux_1389_nl, fsm_output(7));
  nand_276_nl <= NOT((and_389_cse OR (fsm_output(6))) AND (fsm_output(3)));
  and_717_nl <= (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(3));
  mux_1385_nl <= MUX_s_1_2_2(nand_276_nl, and_717_nl, fsm_output(4));
  mux_1384_nl <= MUX_s_1_2_2((NOT (fsm_output(3))), nor_tmp_292, fsm_output(4));
  mux_1386_nl <= MUX_s_1_2_2(mux_1385_nl, mux_1384_nl, fsm_output(2));
  mux_1381_nl <= MUX_s_1_2_2(or_tmp_1370, mux_tmp_1377, fsm_output(1));
  mux_1382_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), mux_1381_nl, fsm_output(4));
  mux_1380_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), mux_tmp_1378, fsm_output(4));
  mux_1383_nl <= MUX_s_1_2_2(mux_1382_nl, mux_1380_nl, fsm_output(2));
  mux_1387_nl <= MUX_s_1_2_2(mux_1386_nl, (NOT mux_1383_nl), fsm_output(7));
  mux_1393_nl <= MUX_s_1_2_2(mux_1392_nl, mux_1387_nl, fsm_output(5));
  and_718_nl <= (fsm_output(4)) AND (fsm_output(0)) AND (fsm_output(1));
  mux_1374_nl <= MUX_s_1_2_2((fsm_output(6)), or_tmp_1367, and_718_nl);
  mux_1376_nl <= MUX_s_1_2_2(mux_tmp_1374, mux_1374_nl, fsm_output(2));
  or_1489_nl <= (fsm_output(7)) OR mux_1376_nl;
  nand_266_nl <= NOT((fsm_output(4)) AND (NOT mux_tmp));
  or_1485_nl <= (NOT (fsm_output(4))) OR (fsm_output(6));
  mux_1373_nl <= MUX_s_1_2_2(nand_266_nl, or_1485_nl, fsm_output(2));
  or_1487_nl <= (fsm_output(7)) OR mux_1373_nl;
  mux_1377_nl <= MUX_s_1_2_2(or_1489_nl, or_1487_nl, fsm_output(5));
  mux_1394_nl <= MUX_s_1_2_2(mux_1393_nl, mux_1377_nl, fsm_output(8));
  mux_1423_nl <= MUX_s_1_2_2(mux_1422_nl, mux_1394_nl, fsm_output(9));
  or_1540_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 5)/=STD_LOGIC_VECTOR'("0001"));
  or_1539_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 5)/=STD_LOGIC_VECTOR'("0100"));
  or_1537_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_1448_nl <= MUX_s_1_2_2(or_tmp_1394, or_1537_nl, fsm_output(6));
  mux_1449_nl <= MUX_s_1_2_2(mux_1448_nl, or_tmp_1401, fsm_output(5));
  mux_1450_nl <= MUX_s_1_2_2(or_1539_nl, mux_1449_nl, fsm_output(1));
  mux_1451_nl <= MUX_s_1_2_2(or_1540_nl, mux_1450_nl, fsm_output(9));
  and_710_nl <= (fsm_output(4)) AND (NOT mux_1451_nl);
  or_1535_nl <= (fsm_output(5)) OR (NOT(COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND
      CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11"))));
  or_1534_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 5)/=STD_LOGIC_VECTOR'("0000"));
  mux_1446_nl <= MUX_s_1_2_2(or_1535_nl, or_1534_nl, fsm_output(1));
  or_1533_nl <= (fsm_output(1)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR (fsm_output(8)) OR (fsm_output(7));
  mux_1447_nl <= MUX_s_1_2_2(mux_1446_nl, or_1533_nl, fsm_output(9));
  nor_676_nl <= NOT((fsm_output(4)) OR mux_1447_nl);
  mux_1452_nl <= MUX_s_1_2_2(and_710_nl, nor_676_nl, fsm_output(3));
  nor_677_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  nor_678_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("101")));
  mux_1441_nl <= MUX_s_1_2_2(nor_677_nl, nor_678_nl, fsm_output(5));
  and_711_nl <= (fsm_output(5)) AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND CONV_SL_1_1(fsm_output(8
      DOWNTO 7)=STD_LOGIC_VECTOR'("10"));
  mux_1442_nl <= MUX_s_1_2_2(mux_1441_nl, and_711_nl, fsm_output(1));
  nor_679_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(6)) OR
      (fsm_output(8)) OR (fsm_output(7)));
  mux_1443_nl <= MUX_s_1_2_2(mux_1442_nl, nor_679_nl, fsm_output(9));
  nor_680_nl <= NOT((fsm_output(9)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 7)/=STD_LOGIC_VECTOR'("00")));
  mux_1444_nl <= MUX_s_1_2_2(mux_1443_nl, nor_680_nl, fsm_output(4));
  nor_681_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(8))
      OR (fsm_output(7)));
  nor_682_nl <= NOT((NOT (fsm_output(1))) OR (NOT (fsm_output(5))) OR (fsm_output(6))
      OR (fsm_output(8)) OR (fsm_output(7)));
  mux_1439_nl <= MUX_s_1_2_2(nor_681_nl, nor_682_nl, fsm_output(9));
  or_1524_nl <= (fsm_output(6)) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR
      CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"));
  mux_1438_nl <= MUX_s_1_2_2(or_1524_nl, or_tmp_1401, fsm_output(5));
  nor_683_nl <= NOT((fsm_output(9)) OR (fsm_output(1)) OR mux_1438_nl);
  mux_1440_nl <= MUX_s_1_2_2(mux_1439_nl, nor_683_nl, fsm_output(4));
  mux_1445_nl <= MUX_s_1_2_2(mux_1444_nl, mux_1440_nl, fsm_output(3));
  mux_1453_nl <= MUX_s_1_2_2(mux_1452_nl, mux_1445_nl, fsm_output(0));
  mux_1433_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), (fsm_output(7)), fsm_output(8));
  mux_1434_nl <= MUX_s_1_2_2(nor_tmp_301, mux_1433_nl, COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  nor_684_nl <= NOT((fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(5)) OR
      (NOT((fsm_output(6)) AND mux_1434_nl)));
  nor_685_nl <= NOT((fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(5)) OR (NOT
      (fsm_output(6))) OR (fsm_output(8)) OR (NOT (fsm_output(7))));
  mux_1435_nl <= MUX_s_1_2_2(nor_684_nl, nor_685_nl, fsm_output(4));
  or_1516_nl <= (fsm_output(6)) OR (NOT nor_tmp_301);
  mux_1430_nl <= MUX_s_1_2_2(or_1516_nl, or_tmp_1394, fsm_output(5));
  mux_1431_nl <= MUX_s_1_2_2(or_tmp_1389, mux_1430_nl, fsm_output(1));
  or_1513_nl <= (fsm_output(1)) OR (fsm_output(5)) OR (fsm_output(6)) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"));
  mux_1432_nl <= MUX_s_1_2_2(mux_1431_nl, or_1513_nl, fsm_output(9));
  and_712_nl <= (fsm_output(4)) AND (NOT mux_1432_nl);
  mux_1436_nl <= MUX_s_1_2_2(mux_1435_nl, and_712_nl, fsm_output(3));
  or_1512_nl <= (NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(8))
      OR (NOT (fsm_output(7)));
  nand_278_nl <= NOT((fsm_output(5)) AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND
      CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("01")));
  mux_1427_nl <= MUX_s_1_2_2(or_tmp_1389, nand_278_nl, fsm_output(1));
  mux_1428_nl <= MUX_s_1_2_2(or_1512_nl, mux_1427_nl, fsm_output(9));
  and_713_nl <= (fsm_output(4)) AND (NOT mux_1428_nl);
  nand_274_nl <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND CONV_SL_1_1(fsm_output(8 DOWNTO
      7)=STD_LOGIC_VECTOR'("11")));
  or_1505_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 5)/=STD_LOGIC_VECTOR'("0011"));
  mux_1425_nl <= MUX_s_1_2_2(nand_274_nl, or_1505_nl, fsm_output(1));
  or_1503_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011"));
  or_1501_nl <= (fsm_output(6)) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR
      CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_1424_nl <= MUX_s_1_2_2(or_1503_nl, or_1501_nl, fsm_output(5));
  or_1504_nl <= (fsm_output(1)) OR mux_1424_nl;
  mux_1426_nl <= MUX_s_1_2_2(mux_1425_nl, or_1504_nl, fsm_output(9));
  nor_686_nl <= NOT((fsm_output(4)) OR mux_1426_nl);
  mux_1429_nl <= MUX_s_1_2_2(and_713_nl, nor_686_nl, fsm_output(3));
  mux_1437_nl <= MUX_s_1_2_2(mux_1436_nl, mux_1429_nl, fsm_output(0));
  or_940_nl <= (NOT (fsm_output(0))) OR (fsm_output(1)) OR (NOT (fsm_output(3)))
      OR (fsm_output(4));
  mux_864_nl <= MUX_s_1_2_2(or_940_nl, or_242_cse, fsm_output(5));
  nor_630_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_864_nl);
  nor_631_nl <= NOT((NOT (fsm_output(8))) OR (NOT (fsm_output(6))) OR (fsm_output(5))
      OR (fsm_output(0)) OR (NOT and_dcpl_59));
  mux_865_nl <= MUX_s_1_2_2(nor_630_nl, nor_631_nl, fsm_output(9));
  nand_263_nl <= NOT(mux_865_nl AND and_dcpl_140);
  or_1547_nl <= (fsm_output(2)) OR (NOT (fsm_output(0))) OR (fsm_output(6)) OR (fsm_output(1))
      OR (fsm_output(5)) OR (NOT (fsm_output(3)));
  or_1545_nl <= (fsm_output(2)) OR (fsm_output(0)) OR (fsm_output(6)) OR (fsm_output(1))
      OR (NOT (fsm_output(5))) OR (fsm_output(3));
  mux_1456_nl <= MUX_s_1_2_2(or_1547_nl, or_1545_nl, fsm_output(4));
  or_1549_nl <= (fsm_output(8)) OR mux_1456_nl;
  nor_674_nl <= NOT((fsm_output(0)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(1)))
      OR (fsm_output(5)) OR (NOT (fsm_output(3))));
  nor_675_nl <= NOT((NOT (fsm_output(0))) OR (fsm_output(6)) OR (fsm_output(1)) OR
      (fsm_output(5)) OR (NOT (fsm_output(3))));
  mux_1455_nl <= MUX_s_1_2_2(nor_674_nl, nor_675_nl, fsm_output(2));
  nand_271_nl <= NOT((fsm_output(8)) AND (fsm_output(4)) AND mux_1455_nl);
  mux_1457_nl <= MUX_s_1_2_2(or_1549_nl, nand_271_nl, fsm_output(9));
  nor_389_nl <= NOT((fsm_output(6)) OR (fsm_output(8)) OR (fsm_output(9)));
  nor_390_nl <= NOT((fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(8))
      OR (fsm_output(9)));
  mux_882_nl <= MUX_s_1_2_2(nor_389_nl, nor_390_nl, fsm_output(3));
  and_360_nl <= (fsm_output(2)) AND (fsm_output(6)) AND (fsm_output(8)) AND (fsm_output(9));
  mux_879_nl <= MUX_s_1_2_2(nor_393_cse, and_369_cse, fsm_output(6));
  and_184_nl <= (fsm_output(2)) AND mux_879_nl;
  mux_880_nl <= MUX_s_1_2_2(and_184_nl, and_361_cse, fsm_output(1));
  mux_881_nl <= MUX_s_1_2_2(and_360_nl, mux_880_nl, fsm_output(0));
  and_185_nl <= (fsm_output(3)) AND mux_881_nl;
  mux_883_nl <= MUX_s_1_2_2(mux_882_nl, and_185_nl, fsm_output(4));
  mux_884_nl <= MUX_s_1_2_2(mux_883_nl, and_361_cse, fsm_output(5));
  mux_885_nl <= MUX_s_1_2_2(mux_884_nl, and_369_cse, fsm_output(7));
  COMP_LOOP_or_15_nl <= (and_dcpl_172 AND and_dcpl_167) OR (COMP_LOOP_COMP_LOOP_nor_4_itm
      AND and_224_m1c) OR (COMP_LOOP_COMP_LOOP_and_34_itm AND and_226_m1c) OR (COMP_LOOP_COMP_LOOP_and_33_itm
      AND and_229_m1c) OR (COMP_LOOP_COMP_LOOP_and_32_itm AND and_230_m1c) OR (COMP_LOOP_COMP_LOOP_and_89_itm
      AND and_233_m1c) OR (COMP_LOOP_COMP_LOOP_and_30_itm AND and_235_m1c) OR (COMP_LOOP_COMP_LOOP_and_145_itm
      AND and_237_m1c);
  COMP_LOOP_or_16_nl <= (and_dcpl_172 AND and_dcpl_176) OR (COMP_LOOP_COMP_LOOP_and_86_itm
      AND and_224_m1c) OR (COMP_LOOP_COMP_LOOP_nor_4_itm AND and_226_m1c) OR (COMP_LOOP_COMP_LOOP_and_34_itm
      AND and_229_m1c) OR (COMP_LOOP_COMP_LOOP_and_33_itm AND and_230_m1c) OR (COMP_LOOP_COMP_LOOP_and_32_itm
      AND and_233_m1c) OR (COMP_LOOP_COMP_LOOP_and_89_itm AND and_235_m1c) OR (COMP_LOOP_COMP_LOOP_and_30_itm
      AND and_237_m1c);
  COMP_LOOP_or_17_nl <= (and_dcpl_172 AND and_dcpl_180) OR (COMP_LOOP_COMP_LOOP_and_145_itm
      AND and_224_m1c) OR (COMP_LOOP_COMP_LOOP_and_86_itm AND and_226_m1c) OR (COMP_LOOP_COMP_LOOP_nor_4_itm
      AND and_229_m1c) OR (COMP_LOOP_COMP_LOOP_and_34_itm AND and_230_m1c) OR (COMP_LOOP_COMP_LOOP_and_33_itm
      AND and_233_m1c) OR (COMP_LOOP_COMP_LOOP_and_32_itm AND and_235_m1c) OR (COMP_LOOP_COMP_LOOP_and_89_itm
      AND and_237_m1c);
  COMP_LOOP_or_18_nl <= (and_dcpl_172 AND and_dcpl_184) OR (COMP_LOOP_COMP_LOOP_and_30_itm
      AND and_224_m1c) OR (COMP_LOOP_COMP_LOOP_and_145_itm AND and_226_m1c) OR (COMP_LOOP_COMP_LOOP_and_86_itm
      AND and_229_m1c) OR (COMP_LOOP_COMP_LOOP_nor_4_itm AND and_230_m1c) OR (COMP_LOOP_COMP_LOOP_and_34_itm
      AND and_233_m1c) OR (COMP_LOOP_COMP_LOOP_and_33_itm AND and_235_m1c) OR (COMP_LOOP_COMP_LOOP_and_32_itm
      AND and_237_m1c);
  COMP_LOOP_or_19_nl <= (and_dcpl_187 AND and_dcpl_167) OR (COMP_LOOP_COMP_LOOP_and_89_itm
      AND and_224_m1c) OR (COMP_LOOP_COMP_LOOP_and_30_itm AND and_226_m1c) OR (COMP_LOOP_COMP_LOOP_and_145_itm
      AND and_229_m1c) OR (COMP_LOOP_COMP_LOOP_and_86_itm AND and_230_m1c) OR (COMP_LOOP_COMP_LOOP_nor_4_itm
      AND and_233_m1c) OR (COMP_LOOP_COMP_LOOP_and_34_itm AND and_235_m1c) OR (COMP_LOOP_COMP_LOOP_and_33_itm
      AND and_237_m1c);
  COMP_LOOP_or_20_nl <= (and_dcpl_187 AND and_dcpl_176) OR (COMP_LOOP_COMP_LOOP_and_32_itm
      AND and_224_m1c) OR (COMP_LOOP_COMP_LOOP_and_89_itm AND and_226_m1c) OR (COMP_LOOP_COMP_LOOP_and_30_itm
      AND and_229_m1c) OR (COMP_LOOP_COMP_LOOP_and_145_itm AND and_230_m1c) OR (COMP_LOOP_COMP_LOOP_and_86_itm
      AND and_233_m1c) OR (COMP_LOOP_COMP_LOOP_nor_4_itm AND and_235_m1c) OR (COMP_LOOP_COMP_LOOP_and_34_itm
      AND and_237_m1c);
  COMP_LOOP_or_21_nl <= (and_dcpl_187 AND and_dcpl_180) OR (COMP_LOOP_COMP_LOOP_and_33_itm
      AND and_224_m1c) OR (COMP_LOOP_COMP_LOOP_and_32_itm AND and_226_m1c) OR (COMP_LOOP_COMP_LOOP_and_89_itm
      AND and_229_m1c) OR (COMP_LOOP_COMP_LOOP_and_30_itm AND and_230_m1c) OR (COMP_LOOP_COMP_LOOP_and_145_itm
      AND and_233_m1c) OR (COMP_LOOP_COMP_LOOP_and_86_itm AND and_235_m1c) OR (COMP_LOOP_COMP_LOOP_nor_4_itm
      AND and_237_m1c);
  COMP_LOOP_or_22_nl <= (and_dcpl_187 AND and_dcpl_184) OR (COMP_LOOP_COMP_LOOP_and_34_itm
      AND and_224_m1c) OR (COMP_LOOP_COMP_LOOP_and_33_itm AND and_226_m1c) OR (COMP_LOOP_COMP_LOOP_and_32_itm
      AND and_229_m1c) OR (COMP_LOOP_COMP_LOOP_and_89_itm AND and_230_m1c) OR (COMP_LOOP_COMP_LOOP_and_30_itm
      AND and_233_m1c) OR (COMP_LOOP_COMP_LOOP_and_145_itm AND and_235_m1c) OR (COMP_LOOP_COMP_LOOP_and_86_itm
      AND and_237_m1c);
  or_964_nl <= and_389_cse OR CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10"));
  mux_909_nl <= MUX_s_1_2_2(or_tmp_113, or_964_nl, fsm_output(5));
  mux_910_nl <= MUX_s_1_2_2(mux_909_nl, (NOT and_314_cse), fsm_output(6));
  nand_120_nl <= NOT((fsm_output(5)) AND or_tmp_788);
  mux_908_nl <= MUX_s_1_2_2(or_1202_cse, nand_120_nl, fsm_output(6));
  mux_911_nl <= MUX_s_1_2_2(mux_910_nl, mux_908_nl, fsm_output(2));
  mux_906_nl <= MUX_s_1_2_2(or_tmp, (NOT or_tmp), fsm_output(6));
  mux_904_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), nor_tmp_27, fsm_output(5));
  mux_905_nl <= MUX_s_1_2_2(or_tmp, mux_904_nl, fsm_output(6));
  mux_907_nl <= MUX_s_1_2_2(mux_906_nl, mux_905_nl, fsm_output(2));
  mux_912_nl <= MUX_s_1_2_2(mux_911_nl, mux_907_nl, fsm_output(7));
  nand_121_nl <= NOT((fsm_output(5)) AND nor_tmp_27);
  and_192_nl <= (fsm_output(5)) AND ((fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(4)));
  mux_901_nl <= MUX_s_1_2_2(nand_121_nl, and_192_nl, fsm_output(6));
  nand_122_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 3)=STD_LOGIC_VECTOR'("111")));
  mux_900_nl <= MUX_s_1_2_2(nand_122_nl, (fsm_output(5)), fsm_output(6));
  mux_902_nl <= MUX_s_1_2_2(mux_901_nl, mux_900_nl, fsm_output(2));
  mux_898_nl <= MUX_s_1_2_2((NOT (fsm_output(5))), or_1202_cse, fsm_output(6));
  nor_388_nl <= NOT((fsm_output(5)) OR and_dcpl_59);
  or_959_nl <= (fsm_output(5)) OR or_tmp_103;
  mux_897_nl <= MUX_s_1_2_2(nor_388_nl, or_959_nl, fsm_output(6));
  mux_899_nl <= MUX_s_1_2_2(mux_898_nl, mux_897_nl, fsm_output(2));
  mux_903_nl <= MUX_s_1_2_2(mux_902_nl, mux_899_nl, fsm_output(7));
  mux_913_nl <= MUX_s_1_2_2(mux_912_nl, mux_903_nl, fsm_output(8));
  mux_892_nl <= MUX_s_1_2_2(or_tmp_103, (NOT (fsm_output(4))), fsm_output(5));
  mux_893_nl <= MUX_s_1_2_2(mux_892_nl, and_tmp_28, fsm_output(6));
  mux_891_nl <= MUX_s_1_2_2((NOT and_tmp_28), and_tmp_28, fsm_output(6));
  mux_894_nl <= MUX_s_1_2_2(mux_893_nl, mux_891_nl, fsm_output(2));
  or_958_nl <= (fsm_output(5)) OR and_705_cse;
  mux_889_nl <= MUX_s_1_2_2(or_958_nl, mux_tmp_705, fsm_output(6));
  mux_887_nl <= MUX_s_1_2_2((NOT or_115_cse), nor_tmp_23, fsm_output(5));
  mux_888_nl <= MUX_s_1_2_2(or_171_cse, mux_887_nl, fsm_output(6));
  mux_890_nl <= MUX_s_1_2_2(mux_889_nl, mux_888_nl, fsm_output(2));
  mux_895_nl <= MUX_s_1_2_2(mux_894_nl, (NOT mux_890_nl), fsm_output(7));
  mux_896_nl <= MUX_s_1_2_2(mux_895_nl, or_tmp_918, fsm_output(8));
  and_238_nl <= and_dcpl_102 AND and_dcpl_48;
  COMP_LOOP_or_26_nl <= ((NOT (modulo_result_rem_cmp_z(63))) AND and_243_m1c) OR
      (not_tmp_399 AND (NOT (modulo_result_rem_cmp_z(63))));
  COMP_LOOP_or_27_nl <= ((modulo_result_rem_cmp_z(63)) AND and_243_m1c) OR (not_tmp_399
      AND (modulo_result_rem_cmp_z(63)));
  COMP_LOOP_or_7_nl <= (COMP_LOOP_COMP_LOOP_nor_1_itm AND and_244_m1c) OR (COMP_LOOP_COMP_LOOP_nor_1_itm
      AND mux_984_m1c);
  COMP_LOOP_or_8_nl <= (COMP_LOOP_COMP_LOOP_and_211 AND and_244_m1c) OR (COMP_LOOP_COMP_LOOP_and_211
      AND mux_984_m1c);
  COMP_LOOP_or_9_nl <= (COMP_LOOP_COMP_LOOP_and_213 AND and_244_m1c) OR (COMP_LOOP_COMP_LOOP_and_213
      AND mux_984_m1c);
  COMP_LOOP_or_10_nl <= (COMP_LOOP_COMP_LOOP_and_125_itm AND and_244_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND mux_984_m1c);
  COMP_LOOP_or_11_nl <= (COMP_LOOP_COMP_LOOP_and_215 AND and_244_m1c) OR (COMP_LOOP_COMP_LOOP_and_215
      AND mux_984_m1c);
  COMP_LOOP_or_12_nl <= (COMP_LOOP_COMP_LOOP_and_11_itm AND and_244_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND mux_984_m1c);
  COMP_LOOP_or_13_nl <= (COMP_LOOP_COMP_LOOP_and_12_itm AND and_244_m1c) OR (COMP_LOOP_COMP_LOOP_and_124_itm
      AND mux_984_m1c);
  COMP_LOOP_or_14_nl <= (COMP_LOOP_COMP_LOOP_and_124_itm AND and_244_m1c) OR (COMP_LOOP_COMP_LOOP_and_125_itm
      AND mux_984_m1c);
  nor_591_nl <= NOT((NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(9)) OR
      (fsm_output(4)) OR (fsm_output(1)) OR (NOT (fsm_output(6))));
  nor_592_nl <= NOT((fsm_output(0)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(1))) OR (fsm_output(6)));
  mux_46_nl <= MUX_s_1_2_2(nor_591_nl, nor_592_nl, fsm_output(5));
  nor_593_nl <= NOT((NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(4)) OR (NOT (fsm_output(1))) OR (fsm_output(6)));
  nor_594_nl <= NOT((fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT
      (fsm_output(4))) OR (fsm_output(1)) OR (NOT (fsm_output(6))));
  mux_45_nl <= MUX_s_1_2_2(nor_593_nl, nor_594_nl, fsm_output(5));
  mux_47_nl <= MUX_s_1_2_2(mux_46_nl, mux_45_nl, fsm_output(8));
  and_470_nl <= (fsm_output(7)) AND mux_47_nl;
  or_61_nl <= (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(4))) OR
      (fsm_output(1)) OR (NOT (fsm_output(6)));
  or_59_nl <= (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(4))) OR
      (fsm_output(1)) OR (NOT (fsm_output(6)));
  mux_43_nl <= MUX_s_1_2_2(or_61_nl, or_59_nl, fsm_output(0));
  or_62_nl <= (fsm_output(5)) OR mux_43_nl;
  nand_224_nl <= NOT((fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(9)) AND
      (fsm_output(4)) AND (fsm_output(1)) AND (NOT (fsm_output(6))));
  or_56_nl <= (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(4))
      OR (NOT (fsm_output(1))) OR (fsm_output(6));
  mux_42_nl <= MUX_s_1_2_2(nand_224_nl, or_56_nl, fsm_output(5));
  mux_44_nl <= MUX_s_1_2_2(or_62_nl, mux_42_nl, fsm_output(8));
  nor_595_nl <= NOT((fsm_output(7)) OR mux_44_nl);
  mux_48_nl <= MUX_s_1_2_2(and_470_nl, nor_595_nl, fsm_output(2));
  or_248_nl <= (fsm_output(0)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(3)))
      OR (fsm_output(4));
  mux_347_nl <= MUX_s_1_2_2(or_248_nl, or_tmp_92, fsm_output(5));
  mux_348_nl <= MUX_s_1_2_2(mux_347_nl, or_247_cse, fsm_output(6));
  mux_346_nl <= MUX_s_1_2_2(nor_tmp_27, (NOT or_tmp_113), fsm_output(5));
  nand_9_nl <= NOT((fsm_output(6)) AND mux_346_nl);
  mux_349_nl <= MUX_s_1_2_2(mux_348_nl, nand_9_nl, fsm_output(2));
  nor_371_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT nor_tmp));
  mux_963_nl <= MUX_s_1_2_2(nor_371_nl, (fsm_output(4)), fsm_output(5));
  mux_341_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), (fsm_output(4)), or_245_cse);
  mux_343_nl <= MUX_s_1_2_2(mux_342_cse, mux_341_nl, fsm_output(0));
  or_246_nl <= (fsm_output(5)) OR mux_343_nl;
  mux_964_nl <= MUX_s_1_2_2((NOT mux_963_nl), or_246_nl, fsm_output(6));
  nand_56_nl <= NOT((fsm_output(5)) AND (NOT mux_696_itm));
  or_1009_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (NOT
      nor_tmp);
  mux_959_nl <= MUX_s_1_2_2((fsm_output(4)), or_1009_nl, fsm_output(5));
  mux_960_nl <= MUX_s_1_2_2(nand_56_nl, mux_959_nl, fsm_output(6));
  mux_965_nl <= MUX_s_1_2_2(mux_964_nl, mux_960_nl, fsm_output(2));
  mux_970_nl <= MUX_s_1_2_2(mux_349_nl, mux_965_nl, fsm_output(7));
  mux_955_nl <= MUX_s_1_2_2(and_705_cse, (NOT nor_tmp), fsm_output(5));
  nor_190_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")));
  mux_954_nl <= MUX_s_1_2_2(nor_tmp, mux_tmp_156, nor_190_nl);
  and_246_nl <= (fsm_output(5)) AND mux_954_nl;
  mux_956_nl <= MUX_s_1_2_2(mux_955_nl, and_246_nl, fsm_output(6));
  mux_332_nl <= MUX_s_1_2_2((fsm_output(4)), (NOT mux_331_cse), fsm_output(5));
  mux_333_nl <= MUX_s_1_2_2(mux_332_nl, and_25_cse, fsm_output(6));
  mux_957_nl <= MUX_s_1_2_2(mux_956_nl, mux_333_nl, fsm_output(2));
  nor_372_nl <= NOT((fsm_output(5)) OR (NOT((NOT(CONV_SL_1_1(fsm_output(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("00")))) OR CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("01")))));
  mux_328_nl <= MUX_s_1_2_2(and_428_cse, or_242_cse, fsm_output(5));
  mux_950_nl <= MUX_s_1_2_2(nor_372_nl, mux_328_nl, fsm_output(6));
  nor_560_nl <= NOT((fsm_output(5)) OR nor_tmp_27);
  mux_334_nl <= MUX_s_1_2_2(nor_tmp, mux_tmp_156, and_389_cse);
  or_1003_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(3))) OR (fsm_output(4));
  mux_947_nl <= MUX_s_1_2_2(mux_334_nl, or_1003_nl, fsm_output(5));
  mux_948_nl <= MUX_s_1_2_2(nor_560_nl, mux_947_nl, fsm_output(6));
  mux_951_nl <= MUX_s_1_2_2(mux_950_nl, mux_948_nl, fsm_output(2));
  mux_958_nl <= MUX_s_1_2_2(mux_957_nl, mux_951_nl, fsm_output(7));
  mux_971_nl <= MUX_s_1_2_2(mux_970_nl, (NOT mux_958_nl), fsm_output(8));
  or_1002_nl <= (fsm_output(5)) OR (fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(4));
  mux_941_nl <= MUX_s_1_2_2((NOT or_tmp_92), or_216_cse, fsm_output(5));
  mux_942_nl <= MUX_s_1_2_2(or_1002_nl, mux_941_nl, fsm_output(6));
  or_999_nl <= (NOT (fsm_output(5))) OR (fsm_output(0)) OR (fsm_output(1)) OR (NOT
      (fsm_output(3))) OR (fsm_output(4));
  mux_939_nl <= MUX_s_1_2_2(and_dcpl_64, or_tmp_103, fsm_output(5));
  mux_940_nl <= MUX_s_1_2_2(or_999_nl, mux_939_nl, fsm_output(6));
  mux_943_nl <= MUX_s_1_2_2(mux_942_nl, mux_940_nl, fsm_output(2));
  or_1383_nl <= (NOT (fsm_output(0))) OR (fsm_output(1)) OR (fsm_output(3)) OR (NOT
      (fsm_output(4)));
  mux_935_nl <= MUX_s_1_2_2(mux_tmp_156, (NOT or_216_cse), and_389_cse);
  mux_936_nl <= MUX_s_1_2_2(or_1383_nl, mux_935_nl, fsm_output(5));
  mux_937_nl <= MUX_s_1_2_2(mux_936_nl, or_171_cse, fsm_output(6));
  nand_117_nl <= NOT((fsm_output(5)) AND or_tmp_891);
  or_996_nl <= (fsm_output(0)) OR (NOT (fsm_output(1))) OR (fsm_output(3)) OR (NOT
      (fsm_output(4)));
  mux_933_nl <= MUX_s_1_2_2(or_216_cse, or_996_nl, fsm_output(5));
  mux_934_nl <= MUX_s_1_2_2(nand_117_nl, mux_933_nl, fsm_output(6));
  mux_938_nl <= MUX_s_1_2_2(mux_937_nl, mux_934_nl, fsm_output(2));
  mux_944_nl <= MUX_s_1_2_2(mux_943_nl, mux_938_nl, fsm_output(7));
  mux_313_nl <= MUX_s_1_2_2((NOT or_tmp_113), and_705_cse, fsm_output(5));
  or_231_nl <= (fsm_output(6)) OR mux_313_nl;
  mux_930_nl <= MUX_s_1_2_2(mux_tmp_719, (fsm_output(4)), fsm_output(5));
  or_992_nl <= (fsm_output(6)) OR mux_930_nl;
  mux_932_nl <= MUX_s_1_2_2(or_231_nl, or_992_nl, fsm_output(2));
  or_994_nl <= (fsm_output(7)) OR mux_932_nl;
  mux_945_nl <= MUX_s_1_2_2(mux_944_nl, or_994_nl, fsm_output(8));
  COMP_LOOP_1_acc_8_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_10_lpi_4_dfm) -
      SIGNED(modulo_result_mux_1_cse), 64));
  or_1146_nl <= (fsm_output(9)) OR (NOT (fsm_output(4))) OR (fsm_output(6)) OR (NOT
      (fsm_output(3))) OR (fsm_output(8));
  or_1145_nl <= (NOT (fsm_output(9))) OR (NOT (fsm_output(4))) OR (fsm_output(6))
      OR (fsm_output(3)) OR (fsm_output(8));
  mux_1137_nl <= MUX_s_1_2_2(or_1146_nl, or_1145_nl, fsm_output(0));
  nor_334_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(5)) OR mux_1137_nl);
  or_1142_nl <= (NOT (fsm_output(4))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(8));
  or_1141_nl <= (fsm_output(4)) OR (fsm_output(6)) OR (NOT (fsm_output(3))) OR (fsm_output(8));
  mux_1135_nl <= MUX_s_1_2_2(or_1142_nl, or_1141_nl, fsm_output(9));
  nor_335_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(0)) OR mux_1135_nl);
  and_321_nl <= (fsm_output(5)) AND (fsm_output(0)) AND (NOT (fsm_output(9))) AND
      (fsm_output(4)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(8)));
  mux_1136_nl <= MUX_s_1_2_2(nor_335_nl, and_321_nl, fsm_output(7));
  mux_1138_nl <= MUX_s_1_2_2(nor_334_nl, mux_1136_nl, fsm_output(2));
  or_1137_nl <= (NOT (fsm_output(0))) OR (fsm_output(9)) OR (fsm_output(4)) OR (fsm_output(6))
      OR (NOT (fsm_output(3))) OR (fsm_output(8));
  or_1136_nl <= (fsm_output(0)) OR (fsm_output(9)) OR (fsm_output(4)) OR (NOT (fsm_output(6)))
      OR (fsm_output(3)) OR (NOT (fsm_output(8)));
  mux_1133_nl <= MUX_s_1_2_2(or_1137_nl, or_1136_nl, fsm_output(5));
  nor_336_nl <= NOT((fsm_output(7)) OR mux_1133_nl);
  nor_337_nl <= NOT((NOT (fsm_output(0))) OR (fsm_output(9)) OR (fsm_output(4)) OR
      (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT (fsm_output(8))));
  nor_338_nl <= NOT((fsm_output(0)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (fsm_output(8)));
  mux_1132_nl <= MUX_s_1_2_2(nor_337_nl, nor_338_nl, fsm_output(5));
  and_322_nl <= (fsm_output(7)) AND mux_1132_nl;
  mux_1134_nl <= MUX_s_1_2_2(nor_336_nl, and_322_nl, fsm_output(2));
  mux_1139_nl <= MUX_s_1_2_2(mux_1138_nl, mux_1134_nl, fsm_output(1));
  nand_98_nl <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("11")) AND
      or_216_cse);
  nand_99_nl <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("11")) AND
      or_tmp_103);
  mux_1155_nl <= MUX_s_1_2_2(nand_98_nl, nand_99_nl, fsm_output(2));
  mux_1156_nl <= MUX_s_1_2_2(mux_tmp_886, mux_1155_nl, fsm_output(7));
  COMP_LOOP_COMP_LOOP_and_145_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva_1(2 DOWNTO
      0)=STD_LOGIC_VECTOR'("110"));
  COMP_LOOP_1_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(COMP_LOOP_k_9_3_sva_2
      & STD_LOGIC_VECTOR'( "000")) + SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(9
      DOWNTO 1)))) + SIGNED'( "0000000001"), 10));
  mux_1174_nl <= MUX_s_1_2_2(mux_tmp_1170, and_tmp_44, fsm_output(6));
  mux_1171_nl <= MUX_s_1_2_2(mux_tmp_1170, mux_tmp_1164, or_1189_cse);
  mux_1167_nl <= MUX_s_1_2_2(mux_tmp_1160, mux_tmp_1159, fsm_output(2));
  mux_1168_nl <= MUX_s_1_2_2(and_tmp_44, mux_1167_nl, fsm_output(3));
  mux_1169_nl <= MUX_s_1_2_2(mux_1168_nl, mux_tmp_1162, fsm_output(0));
  mux_1172_nl <= MUX_s_1_2_2(mux_1171_nl, mux_1169_nl, fsm_output(6));
  and_315_nl <= (fsm_output(7)) AND (fsm_output(9));
  mux_1163_nl <= MUX_s_1_2_2(not_tmp_482, and_315_nl, fsm_output(8));
  mux_1165_nl <= MUX_s_1_2_2(mux_tmp_1164, mux_1163_nl, and_316_cse);
  mux_1166_nl <= MUX_s_1_2_2(mux_1165_nl, mux_tmp_1162, fsm_output(6));
  mux_1173_nl <= MUX_s_1_2_2(mux_1172_nl, mux_1166_nl, fsm_output(1));
  mux_1179_nl <= MUX_s_1_2_2(mux_tmp_1178, and_tmp_46, fsm_output(3));
  and_313_nl <= (fsm_output(0)) AND (fsm_output(3));
  mux_1177_nl <= MUX_s_1_2_2(and_tmp_46, and_tmp_45, and_313_nl);
  mux_1180_nl <= MUX_s_1_2_2(mux_1179_nl, mux_1177_nl, fsm_output(1));
  mux_1176_nl <= MUX_s_1_2_2(and_tmp_46, and_tmp_45, fsm_output(3));
  mux_1181_nl <= MUX_s_1_2_2(mux_1180_nl, mux_1176_nl, fsm_output(2));
  or_1193_nl <= (fsm_output(6)) OR ((fsm_output(5)) AND and_705_cse);
  mux_1183_nl <= MUX_s_1_2_2(or_1193_nl, or_tmp_916, fsm_output(2));
  nand_234_nl <= NOT((fsm_output(7)) AND mux_1183_nl);
  mux_1184_nl <= MUX_s_1_2_2(or_tmp_918, nand_234_nl, fsm_output(8));
  and_272_nl <= (fsm_output(6)) AND or_171_cse;
  and_271_nl <= (fsm_output(6)) AND or_1202_cse;
  mux_1185_nl <= MUX_s_1_2_2(and_272_nl, and_271_nl, fsm_output(2));
  nor_328_nl <= NOT((fsm_output(7)) OR mux_1185_nl);
  mux_1186_nl <= MUX_s_1_2_2(or_tmp_918, nor_328_nl, fsm_output(8));
  or_100_nl <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00")) OR nor_tmp;
  or_1197_nl <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00")) OR nor_tmp_23;
  mux_1187_nl <= MUX_s_1_2_2(or_100_nl, or_1197_nl, fsm_output(2));
  or_1200_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00")) OR mux_1187_nl;
  or_1201_nl <= (fsm_output(8)) OR (CONV_SL_1_1(fsm_output(7 DOWNTO 5)=STD_LOGIC_VECTOR'("111")));
  nor_327_nl <= NOT((fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(8))
      OR (fsm_output(9)));
  mux_1191_nl <= MUX_s_1_2_2(nor_393_cse, nor_327_nl, and_314_cse);
  and_274_nl <= (fsm_output(2)) AND or_838_cse AND CONV_SL_1_1(fsm_output(9 DOWNTO
      8)=STD_LOGIC_VECTOR'("11"));
  mux_1190_nl <= MUX_s_1_2_2(and_274_nl, and_369_cse, or_1202_cse);
  mux_1192_nl <= MUX_s_1_2_2(mux_1191_nl, mux_1190_nl, fsm_output(6));
  COMP_LOOP_COMP_LOOP_or_7_nl <= (VEC_LOOP_j_sva_11_0(11)) OR and_dcpl_243 OR and_dcpl_247
      OR and_dcpl_255 OR and_dcpl_260 OR and_dcpl_266;
  COMP_LOOP_COMP_LOOP_mux_8_nl <= MUX_v_9_2_2((VEC_LOOP_j_sva_11_0(10 DOWNTO 2)),
      (NOT (STAGE_LOOP_lshift_psp_sva(9 DOWNTO 1))), COMP_LOOP_or_40_itm);
  COMP_LOOP_or_44_nl <= (NOT and_511_cse) OR and_dcpl_243 OR and_dcpl_247 OR and_dcpl_255
      OR and_dcpl_260 OR and_dcpl_266;
  COMP_LOOP_COMP_LOOP_mux_9_nl <= MUX_v_6_2_2((STD_LOGIC_VECTOR'( "00") & (COMP_LOOP_k_9_3_sva_5_0(5
      DOWNTO 2))), COMP_LOOP_k_9_3_sva_5_0, COMP_LOOP_or_40_itm);
  COMP_LOOP_COMP_LOOP_or_8_nl <= ((COMP_LOOP_k_9_3_sva_5_0(1)) AND (NOT(and_dcpl_243
      OR and_dcpl_247))) OR and_dcpl_255 OR and_dcpl_260 OR and_dcpl_266;
  COMP_LOOP_COMP_LOOP_or_9_nl <= ((COMP_LOOP_k_9_3_sva_5_0(0)) AND (NOT(and_dcpl_243
      OR and_dcpl_255 OR and_dcpl_260))) OR and_dcpl_247 OR and_dcpl_266;
  COMP_LOOP_COMP_LOOP_or_10_nl <= (NOT(and_dcpl_247 OR and_dcpl_255 OR and_dcpl_266))
      OR and_511_cse OR and_dcpl_243 OR and_dcpl_260;
  acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_or_7_nl &
      COMP_LOOP_COMP_LOOP_mux_8_nl & COMP_LOOP_or_44_nl) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_mux_9_nl
      & COMP_LOOP_COMP_LOOP_or_8_nl & COMP_LOOP_COMP_LOOP_or_9_nl & COMP_LOOP_COMP_LOOP_or_10_nl
      & '1'), 10), 11), 11));
  z_out <= acc_nl(10 DOWNTO 1);
  and_722_nl <= nor_tmp AND (fsm_output(1)) AND (NOT (fsm_output(9))) AND (NOT (fsm_output(8)))
      AND and_dcpl_269 AND and_dcpl;
  and_723_nl <= (NOT (fsm_output(3))) AND (NOT (fsm_output(4))) AND (NOT (fsm_output(1)))
      AND and_dcpl_11 AND (NOT (fsm_output(7))) AND (fsm_output(5)) AND (fsm_output(2))
      AND and_dcpl_276;
  and_724_nl <= and_dcpl_100 AND (NOT (fsm_output(1))) AND and_dcpl_11 AND (fsm_output(7))
      AND (NOT (fsm_output(5))) AND (NOT (fsm_output(2))) AND and_dcpl;
  and_725_nl <= and_dcpl_100 AND (fsm_output(1)) AND and_dcpl_11 AND and_dcpl_269
      AND (fsm_output(6)) AND (NOT (fsm_output(0)));
  and_726_nl <= (NOT (fsm_output(3))) AND (fsm_output(4)) AND (fsm_output(1)) AND
      and_dcpl_23 AND and_dcpl_298 AND (NOT (fsm_output(2))) AND (fsm_output(6))
      AND (fsm_output(0));
  COMP_LOOP_mux1h_125_nl <= MUX1HOT_v_3_6_2(STD_LOGIC_VECTOR'( "001"), STD_LOGIC_VECTOR'(
      "010"), STD_LOGIC_VECTOR'( "011"), STD_LOGIC_VECTOR'( "100"), STD_LOGIC_VECTOR'(
      "101"), STD_LOGIC_VECTOR'( "110"), STD_LOGIC_VECTOR'( and_722_nl & and_723_nl
      & and_724_nl & and_725_nl & and_726_nl & and_dcpl_399));
  and_727_nl <= and_dcpl_128 AND CONV_SL_1_1(fsm_output(9 DOWNTO 8)=STD_LOGIC_VECTOR'("11"))
      AND and_dcpl_298 AND (fsm_output(2)) AND and_dcpl;
  COMP_LOOP_or_45_nl <= MUX_v_3_2_2(COMP_LOOP_mux1h_125_nl, STD_LOGIC_VECTOR'("111"),
      and_727_nl);
  z_out_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_LOOP_lshift_psp_sva) +
      CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_3_sva_5_0 & COMP_LOOP_or_45_nl),
      9), 10), 10));
  COMP_LOOP_mux1h_126_nl <= MUX1HOT_v_64_4_2((STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000001")
      & (NOT (STAGE_LOOP_lshift_psp_sva(9 DOWNTO 4)))), (STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000")
      & VEC_LOOP_j_sva_11_0), p_sva, (STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000000000000000000000")
      & (STAGE_LOOP_lshift_psp_sva(9 DOWNTO 3))), STD_LOGIC_VECTOR'( and_dcpl_324
      & and_511_cse & and_dcpl_340 & and_dcpl_345));
  COMP_LOOP_or_46_nl <= (NOT(and_511_cse OR and_dcpl_340 OR and_dcpl_345)) OR and_dcpl_324;
  COMP_LOOP_COMP_LOOP_or_11_nl <= (NOT(and_dcpl_324 OR and_511_cse OR and_dcpl_345))
      OR and_dcpl_340;
  COMP_LOOP_nor_107_nl <= NOT(and_dcpl_324 OR and_dcpl_345);
  COMP_LOOP_and_85_nl <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), (COMP_LOOP_k_9_3_sva_5_0(5
      DOWNTO 3)), COMP_LOOP_nor_107_nl);
  COMP_LOOP_COMP_LOOP_or_12_nl <= MUX_v_3_2_2(COMP_LOOP_and_85_nl, STD_LOGIC_VECTOR'("111"),
      and_dcpl_340);
  COMP_LOOP_mux_41_nl <= MUX_v_6_2_2(COMP_LOOP_k_9_3_sva_5_0, ((COMP_LOOP_k_9_3_sva_5_0(2
      DOWNTO 0)) & STD_LOGIC_VECTOR'( "111")), and_511_cse);
  COMP_LOOP_COMP_LOOP_or_13_nl <= MUX_v_6_2_2(COMP_LOOP_mux_41_nl, STD_LOGIC_VECTOR'("111111"),
      and_dcpl_340);
  acc_2_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux1h_126_nl
      & COMP_LOOP_or_46_nl), 65), 66) + CONV_UNSIGNED(CONV_SIGNED(SIGNED(COMP_LOOP_COMP_LOOP_or_11_nl
      & COMP_LOOP_COMP_LOOP_or_12_nl & COMP_LOOP_COMP_LOOP_or_13_nl & '1'), 11),
      66), 66));
  z_out_2 <= acc_2_nl(65 DOWNTO 1);
  operator_64_false_1_operator_64_false_1_or_53_nl <= (NOT(and_dcpl_354 OR and_dcpl_368
      OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385 OR and_dcpl_388 OR and_dcpl_394
      OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406)) OR not_tmp_581 OR and_dcpl_362
      OR and_dcpl_411 OR and_dcpl_409;
  operator_64_false_1_operator_64_false_1_or_54_nl <= (NOT((operator_66_true_div_cmp_z(63))
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_362 OR and_dcpl_411;
  operator_64_false_1_mux_51_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(62)),
      (operator_66_true_div_cmp_z(62)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_55_nl <= (NOT(operator_64_false_1_mux_51_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_52_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(61)),
      (operator_66_true_div_cmp_z(61)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_56_nl <= (NOT(operator_64_false_1_mux_52_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_53_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(60)),
      (operator_66_true_div_cmp_z(60)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_57_nl <= (NOT(operator_64_false_1_mux_53_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_54_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(59)),
      (operator_66_true_div_cmp_z(59)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_58_nl <= (NOT(operator_64_false_1_mux_54_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_55_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(58)),
      (operator_66_true_div_cmp_z(58)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_59_nl <= (NOT(operator_64_false_1_mux_55_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_56_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(57)),
      (operator_66_true_div_cmp_z(57)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_60_nl <= (NOT(operator_64_false_1_mux_56_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_57_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(56)),
      (operator_66_true_div_cmp_z(56)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_61_nl <= (NOT(operator_64_false_1_mux_57_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_58_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(55)),
      (operator_66_true_div_cmp_z(55)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_62_nl <= (NOT(operator_64_false_1_mux_58_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_59_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(54)),
      (operator_66_true_div_cmp_z(54)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_63_nl <= (NOT(operator_64_false_1_mux_59_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_60_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(53)),
      (operator_66_true_div_cmp_z(53)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_64_nl <= (NOT(operator_64_false_1_mux_60_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_61_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(52)),
      (operator_66_true_div_cmp_z(52)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_65_nl <= (NOT(operator_64_false_1_mux_61_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_62_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(51)),
      (operator_66_true_div_cmp_z(51)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_66_nl <= (NOT(operator_64_false_1_mux_62_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_63_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(50)),
      (operator_66_true_div_cmp_z(50)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_67_nl <= (NOT(operator_64_false_1_mux_63_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_64_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(49)),
      (operator_66_true_div_cmp_z(49)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_68_nl <= (NOT(operator_64_false_1_mux_64_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_65_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(48)),
      (operator_66_true_div_cmp_z(48)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_69_nl <= (NOT(operator_64_false_1_mux_65_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_66_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(47)),
      (operator_66_true_div_cmp_z(47)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_70_nl <= (NOT(operator_64_false_1_mux_66_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_67_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(46)),
      (operator_66_true_div_cmp_z(46)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_71_nl <= (NOT(operator_64_false_1_mux_67_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_68_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(45)),
      (operator_66_true_div_cmp_z(45)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_72_nl <= (NOT(operator_64_false_1_mux_68_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_69_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(44)),
      (operator_66_true_div_cmp_z(44)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_73_nl <= (NOT(operator_64_false_1_mux_69_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_70_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(43)),
      (operator_66_true_div_cmp_z(43)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_74_nl <= (NOT(operator_64_false_1_mux_70_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_71_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(42)),
      (operator_66_true_div_cmp_z(42)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_75_nl <= (NOT(operator_64_false_1_mux_71_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_72_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(41)),
      (operator_66_true_div_cmp_z(41)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_76_nl <= (NOT(operator_64_false_1_mux_72_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_73_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(40)),
      (operator_66_true_div_cmp_z(40)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_77_nl <= (NOT(operator_64_false_1_mux_73_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_74_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(39)),
      (operator_66_true_div_cmp_z(39)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_78_nl <= (NOT(operator_64_false_1_mux_74_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_75_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(38)),
      (operator_66_true_div_cmp_z(38)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_79_nl <= (NOT(operator_64_false_1_mux_75_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_76_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(37)),
      (operator_66_true_div_cmp_z(37)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_80_nl <= (NOT(operator_64_false_1_mux_76_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_77_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(36)),
      (operator_66_true_div_cmp_z(36)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_81_nl <= (NOT(operator_64_false_1_mux_77_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_78_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(35)),
      (operator_66_true_div_cmp_z(35)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_82_nl <= (NOT(operator_64_false_1_mux_78_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_79_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(34)),
      (operator_66_true_div_cmp_z(34)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_83_nl <= (NOT(operator_64_false_1_mux_79_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_80_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(33)),
      (operator_66_true_div_cmp_z(33)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_84_nl <= (NOT(operator_64_false_1_mux_80_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_81_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(32)),
      (operator_66_true_div_cmp_z(32)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_85_nl <= (NOT(operator_64_false_1_mux_81_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_82_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(31)),
      (operator_66_true_div_cmp_z(31)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_86_nl <= (NOT(operator_64_false_1_mux_82_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_83_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(30)),
      (operator_66_true_div_cmp_z(30)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_87_nl <= (NOT(operator_64_false_1_mux_83_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_84_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(29)),
      (operator_66_true_div_cmp_z(29)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_88_nl <= (NOT(operator_64_false_1_mux_84_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_85_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(28)),
      (operator_66_true_div_cmp_z(28)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_89_nl <= (NOT(operator_64_false_1_mux_85_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_86_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(27)),
      (operator_66_true_div_cmp_z(27)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_90_nl <= (NOT(operator_64_false_1_mux_86_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_87_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(26)),
      (operator_66_true_div_cmp_z(26)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_91_nl <= (NOT(operator_64_false_1_mux_87_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_88_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(25)),
      (operator_66_true_div_cmp_z(25)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_92_nl <= (NOT(operator_64_false_1_mux_88_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_89_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(24)),
      (operator_66_true_div_cmp_z(24)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_93_nl <= (NOT(operator_64_false_1_mux_89_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_90_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(23)),
      (operator_66_true_div_cmp_z(23)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_94_nl <= (NOT(operator_64_false_1_mux_90_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_91_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(22)),
      (operator_66_true_div_cmp_z(22)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_95_nl <= (NOT(operator_64_false_1_mux_91_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_92_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(21)),
      (operator_66_true_div_cmp_z(21)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_96_nl <= (NOT(operator_64_false_1_mux_92_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_93_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(20)),
      (operator_66_true_div_cmp_z(20)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_97_nl <= (NOT(operator_64_false_1_mux_93_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_94_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(19)),
      (operator_66_true_div_cmp_z(19)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_98_nl <= (NOT(operator_64_false_1_mux_94_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_95_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(18)),
      (operator_66_true_div_cmp_z(18)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_99_nl <= (NOT(operator_64_false_1_mux_95_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_96_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(17)),
      (operator_66_true_div_cmp_z(17)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_100_nl <= (NOT(operator_64_false_1_mux_96_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_97_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(16)),
      (operator_66_true_div_cmp_z(16)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_101_nl <= (NOT(operator_64_false_1_mux_97_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_98_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(15)),
      (operator_66_true_div_cmp_z(15)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_102_nl <= (NOT(operator_64_false_1_mux_98_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_99_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(14)),
      (operator_66_true_div_cmp_z(14)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_103_nl <= (NOT(operator_64_false_1_mux_99_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_100_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(13)),
      (operator_66_true_div_cmp_z(13)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_104_nl <= (NOT(operator_64_false_1_mux_100_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux_101_nl <= MUX_s_1_2_2((operator_64_false_acc_mut_63_0(12)),
      (operator_66_true_div_cmp_z(12)), and_dcpl_409);
  operator_64_false_1_operator_64_false_1_or_105_nl <= (NOT(operator_64_false_1_mux_101_nl
      OR and_dcpl_354 OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_379 OR and_dcpl_385
      OR and_dcpl_388 OR and_dcpl_394 OR and_dcpl_399 OR and_dcpl_404 OR and_dcpl_406))
      OR not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_mux1h_4_nl <= MUX1HOT_v_4_3_2((operator_64_false_acc_mut_63_0(11
      DOWNTO 8)), (NOT (VEC_LOOP_j_sva_11_0(11 DOWNTO 8))), (operator_66_true_div_cmp_z(11
      DOWNTO 8)), STD_LOGIC_VECTOR'( and_dcpl_362 & operator_64_false_1_or_1_itm
      & and_dcpl_409));
  operator_64_false_1_operator_64_false_1_nor_105_nl <= NOT(MUX_v_4_2_2(operator_64_false_1_mux1h_4_nl,
      STD_LOGIC_VECTOR'("1111"), and_dcpl_354));
  operator_64_false_1_or_8_nl <= not_tmp_581 OR and_dcpl_411;
  operator_64_false_1_or_7_nl <= MUX_v_4_2_2(operator_64_false_1_operator_64_false_1_nor_105_nl,
      STD_LOGIC_VECTOR'("1111"), operator_64_false_1_or_8_nl);
  operator_64_false_1_mux1h_5_nl <= MUX1HOT_v_8_6_2((STD_LOGIC_VECTOR'( "01") & (NOT
      COMP_LOOP_k_9_3_sva_5_0)), STD_LOGIC_VECTOR'( (NOT modExp_exp_1_7_1_sva) &
      (NOT modExp_exp_1_6_1_sva) & (NOT modExp_exp_1_5_1_sva) & (NOT modExp_exp_1_4_1_sva)
      & (NOT modExp_exp_1_3_1_sva) & (NOT modExp_exp_1_2_1_sva) & (NOT modExp_exp_1_1_1_sva)
      & (NOT modExp_exp_1_0_1_sva_1)), (NOT (operator_64_false_acc_mut_63_0(7 DOWNTO
      0))), (VEC_LOOP_j_sva_11_0(7 DOWNTO 0)), (NOT (operator_66_true_div_cmp_z(7
      DOWNTO 0))), STD_LOGIC_VECTOR'( (NOT modExp_exp_1_1_1_sva) & (NOT modExp_exp_1_7_1_sva)
      & (NOT modExp_exp_1_6_1_sva) & (NOT modExp_exp_1_5_1_sva) & (NOT modExp_exp_1_4_1_sva)
      & (NOT modExp_exp_1_3_1_sva) & (NOT modExp_exp_1_2_1_sva) & (NOT modExp_exp_1_0_1_sva_1)),
      STD_LOGIC_VECTOR'( and_dcpl_354 & not_tmp_581 & and_dcpl_362 & operator_64_false_1_or_1_itm
      & and_dcpl_409 & and_dcpl_411));
  operator_64_false_1_mux1h_6_nl <= MUX1HOT_v_7_3_2((z_out_2(6 DOWNTO 0)), (z_out_1(9
      DOWNTO 3)), (STAGE_LOOP_lshift_psp_sva(9 DOWNTO 3)), STD_LOGIC_VECTOR'( and_dcpl_368
      & operator_64_false_1_or_5_ssc & and_dcpl_406));
  operator_64_false_1_not_3_nl <= NOT operator_64_false_1_or_4_ssc;
  operator_64_false_1_and_53_nl <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"), operator_64_false_1_mux1h_6_nl,
      operator_64_false_1_not_3_nl);
  operator_64_false_1_or_9_nl <= and_dcpl_368 OR and_dcpl_406;
  operator_64_false_1_mux1h_7_nl <= MUX1HOT_v_3_3_2(STD_LOGIC_VECTOR'( "001"), (STAGE_LOOP_lshift_psp_sva(2
      DOWNTO 0)), (z_out_1(2 DOWNTO 0)), STD_LOGIC_VECTOR'( operator_64_false_1_or_4_ssc
      & operator_64_false_1_or_9_nl & operator_64_false_1_or_5_ssc));
  z_out_3 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(operator_64_false_1_operator_64_false_1_or_53_nl
      & operator_64_false_1_operator_64_false_1_or_54_nl & operator_64_false_1_operator_64_false_1_or_55_nl
      & operator_64_false_1_operator_64_false_1_or_56_nl & operator_64_false_1_operator_64_false_1_or_57_nl
      & operator_64_false_1_operator_64_false_1_or_58_nl & operator_64_false_1_operator_64_false_1_or_59_nl
      & operator_64_false_1_operator_64_false_1_or_60_nl & operator_64_false_1_operator_64_false_1_or_61_nl
      & operator_64_false_1_operator_64_false_1_or_62_nl & operator_64_false_1_operator_64_false_1_or_63_nl
      & operator_64_false_1_operator_64_false_1_or_64_nl & operator_64_false_1_operator_64_false_1_or_65_nl
      & operator_64_false_1_operator_64_false_1_or_66_nl & operator_64_false_1_operator_64_false_1_or_67_nl
      & operator_64_false_1_operator_64_false_1_or_68_nl & operator_64_false_1_operator_64_false_1_or_69_nl
      & operator_64_false_1_operator_64_false_1_or_70_nl & operator_64_false_1_operator_64_false_1_or_71_nl
      & operator_64_false_1_operator_64_false_1_or_72_nl & operator_64_false_1_operator_64_false_1_or_73_nl
      & operator_64_false_1_operator_64_false_1_or_74_nl & operator_64_false_1_operator_64_false_1_or_75_nl
      & operator_64_false_1_operator_64_false_1_or_76_nl & operator_64_false_1_operator_64_false_1_or_77_nl
      & operator_64_false_1_operator_64_false_1_or_78_nl & operator_64_false_1_operator_64_false_1_or_79_nl
      & operator_64_false_1_operator_64_false_1_or_80_nl & operator_64_false_1_operator_64_false_1_or_81_nl
      & operator_64_false_1_operator_64_false_1_or_82_nl & operator_64_false_1_operator_64_false_1_or_83_nl
      & operator_64_false_1_operator_64_false_1_or_84_nl & operator_64_false_1_operator_64_false_1_or_85_nl
      & operator_64_false_1_operator_64_false_1_or_86_nl & operator_64_false_1_operator_64_false_1_or_87_nl
      & operator_64_false_1_operator_64_false_1_or_88_nl & operator_64_false_1_operator_64_false_1_or_89_nl
      & operator_64_false_1_operator_64_false_1_or_90_nl & operator_64_false_1_operator_64_false_1_or_91_nl
      & operator_64_false_1_operator_64_false_1_or_92_nl & operator_64_false_1_operator_64_false_1_or_93_nl
      & operator_64_false_1_operator_64_false_1_or_94_nl & operator_64_false_1_operator_64_false_1_or_95_nl
      & operator_64_false_1_operator_64_false_1_or_96_nl & operator_64_false_1_operator_64_false_1_or_97_nl
      & operator_64_false_1_operator_64_false_1_or_98_nl & operator_64_false_1_operator_64_false_1_or_99_nl
      & operator_64_false_1_operator_64_false_1_or_100_nl & operator_64_false_1_operator_64_false_1_or_101_nl
      & operator_64_false_1_operator_64_false_1_or_102_nl & operator_64_false_1_operator_64_false_1_or_103_nl
      & operator_64_false_1_operator_64_false_1_or_104_nl & operator_64_false_1_operator_64_false_1_or_105_nl
      & operator_64_false_1_or_7_nl & operator_64_false_1_mux1h_5_nl) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(operator_64_false_1_and_53_nl
      & operator_64_false_1_mux1h_7_nl), 10), 65), 65));
  and_728_nl <= (NOT (fsm_output(4))) AND (fsm_output(3)) AND (fsm_output(1)) AND
      nor_393_cse AND and_dcpl_238 AND and_dcpl_276;
  nor_690_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(8)) OR
      (fsm_output(9)) OR (fsm_output(1)) OR not_tmp_309);
  or_1560_nl <= (fsm_output(1)) OR (fsm_output(3)) OR (NOT (fsm_output(4)));
  or_1561_nl <= (fsm_output(1)) OR (NOT (fsm_output(3))) OR (fsm_output(4));
  mux_1462_nl <= MUX_s_1_2_2(or_1560_nl, or_1561_nl, fsm_output(9));
  nor_691_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(8)) OR
      mux_1462_nl);
  mux_1461_nl <= MUX_s_1_2_2(nor_690_nl, nor_691_nl, fsm_output(2));
  nor_692_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(8)))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(4)));
  and_729_nl <= (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(8))) AND
      (fsm_output(9)) AND (fsm_output(1)) AND (NOT (fsm_output(3))) AND (fsm_output(4));
  mux_1463_nl <= MUX_s_1_2_2(nor_692_nl, and_729_nl, fsm_output(2));
  mux_1460_nl <= MUX_s_1_2_2(mux_1461_nl, mux_1463_nl, fsm_output(6));
  or_1562_nl <= (fsm_output(8)) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (NOT
      (fsm_output(3))) OR (fsm_output(4));
  mux_1465_nl <= MUX_s_1_2_2(or_1562_nl, or_1440_cse, fsm_output(7));
  nor_693_nl <= NOT((fsm_output(2)) OR (fsm_output(5)) OR mux_1465_nl);
  nor_694_nl <= NOT((NOT (fsm_output(7))) OR (NOT (fsm_output(8))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(4)));
  nor_695_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(8)) OR (fsm_output(9)) OR
      (fsm_output(1)) OR not_tmp_309);
  mux_1466_nl <= MUX_s_1_2_2(nor_694_nl, nor_695_nl, fsm_output(5));
  and_730_nl <= (fsm_output(2)) AND mux_1466_nl;
  mux_1464_nl <= MUX_s_1_2_2(nor_693_nl, and_730_nl, fsm_output(6));
  mux_1459_nl <= MUX_s_1_2_2(mux_1460_nl, mux_1464_nl, fsm_output(0));
  nor_696_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(8)) OR (fsm_output(2)) OR
      (fsm_output(9)) OR not_tmp_600);
  nor_697_nl <= NOT((fsm_output(7)) OR (fsm_output(8)) OR (NOT (fsm_output(2))) OR
      (NOT (fsm_output(9))) OR (fsm_output(4)) OR (NOT (fsm_output(0))));
  mux_1469_nl <= MUX_s_1_2_2(nor_696_nl, nor_697_nl, fsm_output(5));
  nand_279_nl <= NOT((fsm_output(3)) AND mux_1469_nl);
  or_1564_nl <= (fsm_output(8)) OR (fsm_output(2)) OR (fsm_output(9)) OR (fsm_output(4))
      OR (NOT (fsm_output(0)));
  mux_1472_nl <= MUX_s_1_2_2(or_tmp_1346, or_1564_nl, fsm_output(7));
  or_1565_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(8))) OR (fsm_output(2))
      OR (fsm_output(9)) OR (NOT (fsm_output(4))) OR (fsm_output(0));
  mux_1471_nl <= MUX_s_1_2_2(mux_1472_nl, or_1565_nl, fsm_output(5));
  or_1567_nl <= (fsm_output(8)) OR (NOT (fsm_output(2))) OR (fsm_output(9)) OR (NOT
      (fsm_output(4))) OR (fsm_output(0));
  or_1568_nl <= (NOT (fsm_output(8))) OR (fsm_output(2)) OR (fsm_output(9)) OR (fsm_output(4))
      OR (fsm_output(0));
  mux_1473_nl <= MUX_s_1_2_2(or_1567_nl, or_1568_nl, fsm_output(7));
  or_1566_nl <= (fsm_output(5)) OR mux_1473_nl;
  mux_1470_nl <= MUX_s_1_2_2(mux_1471_nl, or_1566_nl, fsm_output(3));
  mux_1468_nl <= MUX_s_1_2_2(nand_279_nl, mux_1470_nl, fsm_output(6));
  or_1570_nl <= (fsm_output(2)) OR (fsm_output(9)) OR not_tmp_600;
  or_1571_nl <= (NOT (fsm_output(2))) OR (fsm_output(9)) OR (fsm_output(4)) OR (fsm_output(0));
  mux_1477_nl <= MUX_s_1_2_2(or_1570_nl, or_1571_nl, fsm_output(8));
  or_1569_nl <= (fsm_output(7)) OR mux_1477_nl;
  mux_1476_nl <= MUX_s_1_2_2(or_tmp_1349, or_1569_nl, fsm_output(5));
  nand_280_nl <= NOT((fsm_output(8)) AND (fsm_output(2)) AND (fsm_output(9)) AND
      (fsm_output(4)) AND (fsm_output(0)));
  mux_1479_nl <= MUX_s_1_2_2(nand_280_nl, or_tmp_1348, fsm_output(7));
  mux_1478_nl <= MUX_s_1_2_2(mux_1479_nl, or_tmp_1349, fsm_output(5));
  mux_1475_nl <= MUX_s_1_2_2(mux_1476_nl, mux_1478_nl, fsm_output(3));
  mux_1481_nl <= MUX_s_1_2_2(or_tmp_1348, or_tmp_1346, fsm_output(7));
  nand_281_nl <= NOT((fsm_output(5)) AND (NOT mux_1481_nl));
  or_1572_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(8))
      OR (NOT (fsm_output(2))) OR (fsm_output(9)) OR (NOT (fsm_output(4))) OR (fsm_output(0));
  mux_1480_nl <= MUX_s_1_2_2(nand_281_nl, or_1572_nl, fsm_output(3));
  mux_1474_nl <= MUX_s_1_2_2(mux_1475_nl, mux_1480_nl, fsm_output(6));
  mux_1467_nl <= MUX_s_1_2_2(mux_1468_nl, mux_1474_nl, fsm_output(1));
  modExp_while_if_mux1h_2_nl <= MUX1HOT_v_64_3_2(modExp_result_sva, COMP_LOOP_1_mul_mut,
      operator_64_false_acc_mut_63_0, STD_LOGIC_VECTOR'( and_728_nl & mux_1459_nl
      & (NOT mux_1467_nl)));
  z_out_4 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(modExp_while_if_mux1h_2_nl)
      * SIGNED(COMP_LOOP_1_mul_mut)), 64));
END v40;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_0_adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    vec_rsc_0_0_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_wea : OUT STD_LOGIC;
    vec_rsc_0_0_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_0_1_adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    vec_rsc_0_1_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_wea : OUT STD_LOGIC;
    vec_rsc_0_1_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_0_2_adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    vec_rsc_0_2_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_wea : OUT STD_LOGIC;
    vec_rsc_0_2_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_0_3_adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    vec_rsc_0_3_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_wea : OUT STD_LOGIC;
    vec_rsc_0_3_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_0_4_adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    vec_rsc_0_4_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_wea : OUT STD_LOGIC;
    vec_rsc_0_4_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_0_5_adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    vec_rsc_0_5_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_wea : OUT STD_LOGIC;
    vec_rsc_0_5_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_0_6_adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    vec_rsc_0_6_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_wea : OUT STD_LOGIC;
    vec_rsc_0_6_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_0_7_adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    vec_rsc_0_7_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_wea : OUT STD_LOGIC;
    vec_rsc_0_7_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC
  );
END inPlaceNTT_DIT;

ARCHITECTURE v40 OF inPlaceNTT_DIT IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_adra_d_iff : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da_d_iff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_wea_d_iff : STD_LOGIC;

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_9_64_512_512_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_0_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_adra : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_9_64_512_512_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_1_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_adra : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_9_64_512_512_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_2_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_adra : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_9_64_512_512_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_3_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_adra : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_9_64_512_512_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_4_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_adra : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_9_64_512_512_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_5_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_adra : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_9_64_512_512_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_6_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_adra : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_9_64_512_512_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_7_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_adra : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      p_rsc_triosy_lz : OUT STD_LOGIC;
      r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      r_rsc_triosy_lz : OUT STD_LOGIC;
      vec_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_0_i_adra_d_pff : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
      vec_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_1_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_2_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_3_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_4_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_5_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_6_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_7_i_wea_d_pff : OUT STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIT_core_inst_p_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIT_core_inst_r_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_adra_d_pff : STD_LOGIC_VECTOR (8
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_da_d_pff : STD_LOGIC_VECTOR (63 DOWNTO
      0);

BEGIN
  vec_rsc_0_0_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_9_64_512_512_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_0_i_qa,
      wea => vec_rsc_0_0_wea,
      da => vec_rsc_0_0_i_da,
      adra => vec_rsc_0_0_i_adra,
      adra_d => vec_rsc_0_0_i_adra_d,
      da_d => vec_rsc_0_0_i_da_d,
      qa_d => vec_rsc_0_0_i_qa_d_1,
      wea_d => vec_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_0_i_wea_d_iff
    );
  vec_rsc_0_0_i_qa <= vec_rsc_0_0_qa;
  vec_rsc_0_0_da <= vec_rsc_0_0_i_da;
  vec_rsc_0_0_adra <= vec_rsc_0_0_i_adra;
  vec_rsc_0_0_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_0_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_0_i_qa_d <= vec_rsc_0_0_i_qa_d_1;

  vec_rsc_0_1_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_9_64_512_512_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_1_i_qa,
      wea => vec_rsc_0_1_wea,
      da => vec_rsc_0_1_i_da,
      adra => vec_rsc_0_1_i_adra,
      adra_d => vec_rsc_0_1_i_adra_d,
      da_d => vec_rsc_0_1_i_da_d,
      qa_d => vec_rsc_0_1_i_qa_d_1,
      wea_d => vec_rsc_0_1_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_1_i_wea_d_iff
    );
  vec_rsc_0_1_i_qa <= vec_rsc_0_1_qa;
  vec_rsc_0_1_da <= vec_rsc_0_1_i_da;
  vec_rsc_0_1_adra <= vec_rsc_0_1_i_adra;
  vec_rsc_0_1_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_1_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_1_i_qa_d <= vec_rsc_0_1_i_qa_d_1;

  vec_rsc_0_2_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_9_64_512_512_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_2_i_qa,
      wea => vec_rsc_0_2_wea,
      da => vec_rsc_0_2_i_da,
      adra => vec_rsc_0_2_i_adra,
      adra_d => vec_rsc_0_2_i_adra_d,
      da_d => vec_rsc_0_2_i_da_d,
      qa_d => vec_rsc_0_2_i_qa_d_1,
      wea_d => vec_rsc_0_2_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_2_i_wea_d_iff
    );
  vec_rsc_0_2_i_qa <= vec_rsc_0_2_qa;
  vec_rsc_0_2_da <= vec_rsc_0_2_i_da;
  vec_rsc_0_2_adra <= vec_rsc_0_2_i_adra;
  vec_rsc_0_2_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_2_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_2_i_qa_d <= vec_rsc_0_2_i_qa_d_1;

  vec_rsc_0_3_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_9_64_512_512_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_3_i_qa,
      wea => vec_rsc_0_3_wea,
      da => vec_rsc_0_3_i_da,
      adra => vec_rsc_0_3_i_adra,
      adra_d => vec_rsc_0_3_i_adra_d,
      da_d => vec_rsc_0_3_i_da_d,
      qa_d => vec_rsc_0_3_i_qa_d_1,
      wea_d => vec_rsc_0_3_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_3_i_wea_d_iff
    );
  vec_rsc_0_3_i_qa <= vec_rsc_0_3_qa;
  vec_rsc_0_3_da <= vec_rsc_0_3_i_da;
  vec_rsc_0_3_adra <= vec_rsc_0_3_i_adra;
  vec_rsc_0_3_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_3_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_3_i_qa_d <= vec_rsc_0_3_i_qa_d_1;

  vec_rsc_0_4_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_9_64_512_512_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_4_i_qa,
      wea => vec_rsc_0_4_wea,
      da => vec_rsc_0_4_i_da,
      adra => vec_rsc_0_4_i_adra,
      adra_d => vec_rsc_0_4_i_adra_d,
      da_d => vec_rsc_0_4_i_da_d,
      qa_d => vec_rsc_0_4_i_qa_d_1,
      wea_d => vec_rsc_0_4_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_4_i_wea_d_iff
    );
  vec_rsc_0_4_i_qa <= vec_rsc_0_4_qa;
  vec_rsc_0_4_da <= vec_rsc_0_4_i_da;
  vec_rsc_0_4_adra <= vec_rsc_0_4_i_adra;
  vec_rsc_0_4_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_4_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_4_i_qa_d <= vec_rsc_0_4_i_qa_d_1;

  vec_rsc_0_5_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_9_64_512_512_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_5_i_qa,
      wea => vec_rsc_0_5_wea,
      da => vec_rsc_0_5_i_da,
      adra => vec_rsc_0_5_i_adra,
      adra_d => vec_rsc_0_5_i_adra_d,
      da_d => vec_rsc_0_5_i_da_d,
      qa_d => vec_rsc_0_5_i_qa_d_1,
      wea_d => vec_rsc_0_5_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_5_i_wea_d_iff
    );
  vec_rsc_0_5_i_qa <= vec_rsc_0_5_qa;
  vec_rsc_0_5_da <= vec_rsc_0_5_i_da;
  vec_rsc_0_5_adra <= vec_rsc_0_5_i_adra;
  vec_rsc_0_5_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_5_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_5_i_qa_d <= vec_rsc_0_5_i_qa_d_1;

  vec_rsc_0_6_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_9_64_512_512_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_6_i_qa,
      wea => vec_rsc_0_6_wea,
      da => vec_rsc_0_6_i_da,
      adra => vec_rsc_0_6_i_adra,
      adra_d => vec_rsc_0_6_i_adra_d,
      da_d => vec_rsc_0_6_i_da_d,
      qa_d => vec_rsc_0_6_i_qa_d_1,
      wea_d => vec_rsc_0_6_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_6_i_wea_d_iff
    );
  vec_rsc_0_6_i_qa <= vec_rsc_0_6_qa;
  vec_rsc_0_6_da <= vec_rsc_0_6_i_da;
  vec_rsc_0_6_adra <= vec_rsc_0_6_i_adra;
  vec_rsc_0_6_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_6_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_6_i_qa_d <= vec_rsc_0_6_i_qa_d_1;

  vec_rsc_0_7_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_9_64_512_512_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_7_i_qa,
      wea => vec_rsc_0_7_wea,
      da => vec_rsc_0_7_i_da,
      adra => vec_rsc_0_7_i_adra,
      adra_d => vec_rsc_0_7_i_adra_d,
      da_d => vec_rsc_0_7_i_da_d,
      qa_d => vec_rsc_0_7_i_qa_d_1,
      wea_d => vec_rsc_0_7_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_7_i_wea_d_iff
    );
  vec_rsc_0_7_i_qa <= vec_rsc_0_7_qa;
  vec_rsc_0_7_da <= vec_rsc_0_7_i_da;
  vec_rsc_0_7_adra <= vec_rsc_0_7_i_adra;
  vec_rsc_0_7_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_7_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_7_i_qa_d <= vec_rsc_0_7_i_qa_d_1;

  inPlaceNTT_DIT_core_inst : inPlaceNTT_DIT_core
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_triosy_0_0_lz => vec_rsc_triosy_0_0_lz,
      vec_rsc_triosy_0_1_lz => vec_rsc_triosy_0_1_lz,
      vec_rsc_triosy_0_2_lz => vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz => vec_rsc_triosy_0_3_lz,
      vec_rsc_triosy_0_4_lz => vec_rsc_triosy_0_4_lz,
      vec_rsc_triosy_0_5_lz => vec_rsc_triosy_0_5_lz,
      vec_rsc_triosy_0_6_lz => vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz => vec_rsc_triosy_0_7_lz,
      p_rsc_dat => inPlaceNTT_DIT_core_inst_p_rsc_dat,
      p_rsc_triosy_lz => p_rsc_triosy_lz,
      r_rsc_dat => inPlaceNTT_DIT_core_inst_r_rsc_dat,
      r_rsc_triosy_lz => r_rsc_triosy_lz,
      vec_rsc_0_0_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_qa_d,
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_1_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_1_i_qa_d,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_2_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_2_i_qa_d,
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_3_i_qa_d,
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_4_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_4_i_qa_d,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_5_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_5_i_qa_d,
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_6_i_qa_d,
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_7_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_7_i_qa_d,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_0_i_adra_d_pff => inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_adra_d_pff,
      vec_rsc_0_0_i_da_d_pff => inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_da_d_pff,
      vec_rsc_0_0_i_wea_d_pff => vec_rsc_0_0_i_wea_d_iff,
      vec_rsc_0_1_i_wea_d_pff => vec_rsc_0_1_i_wea_d_iff,
      vec_rsc_0_2_i_wea_d_pff => vec_rsc_0_2_i_wea_d_iff,
      vec_rsc_0_3_i_wea_d_pff => vec_rsc_0_3_i_wea_d_iff,
      vec_rsc_0_4_i_wea_d_pff => vec_rsc_0_4_i_wea_d_iff,
      vec_rsc_0_5_i_wea_d_pff => vec_rsc_0_5_i_wea_d_iff,
      vec_rsc_0_6_i_wea_d_pff => vec_rsc_0_6_i_wea_d_iff,
      vec_rsc_0_7_i_wea_d_pff => vec_rsc_0_7_i_wea_d_iff
    );
  inPlaceNTT_DIT_core_inst_p_rsc_dat <= p_rsc_dat;
  inPlaceNTT_DIT_core_inst_r_rsc_dat <= r_rsc_dat;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_qa_d <= vec_rsc_0_0_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_1_i_qa_d <= vec_rsc_0_1_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_2_i_qa_d <= vec_rsc_0_2_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_3_i_qa_d <= vec_rsc_0_3_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_4_i_qa_d <= vec_rsc_0_4_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_5_i_qa_d <= vec_rsc_0_5_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_6_i_qa_d <= vec_rsc_0_6_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_7_i_qa_d <= vec_rsc_0_7_i_qa_d;
  vec_rsc_0_0_i_adra_d_iff <= inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_adra_d_pff;
  vec_rsc_0_0_i_da_d_iff <= inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_da_d_pff;

END v40;



