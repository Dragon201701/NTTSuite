
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.v 
module mgc_rem(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_b-1:0] z;  
   reg  [width_b-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  rem_s(a,b,z);
	else
          rem_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.v 
module mgc_div(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_a-1:0] z;  
   reg  [width_a-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  div_s(a,b,z);
	else
          div_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Wed Jun 30 21:15:29 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_10_64_1024_1024_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_10_64_1024_1024_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [9:0] adra;
  input [9:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_10_64_1024_1024_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_10_64_1024_1024_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [9:0] adra;
  input [9:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_10_64_1024_1024_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_10_64_1024_1024_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [9:0] adra;
  input [9:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_10_64_1024_1024_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_10_64_1024_1024_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [9:0] adra;
  input [9:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core_core_fsm (
  clk, rst, fsm_output, STAGE_LOOP_C_9_tr0, modExp_while_C_42_tr0, COMP_LOOP_C_1_tr0,
      COMP_LOOP_1_modExp_1_while_C_42_tr0, COMP_LOOP_C_68_tr0, COMP_LOOP_2_modExp_1_while_C_42_tr0,
      COMP_LOOP_C_136_tr0, COMP_LOOP_3_modExp_1_while_C_42_tr0, COMP_LOOP_C_204_tr0,
      COMP_LOOP_4_modExp_1_while_C_42_tr0, COMP_LOOP_C_272_tr0, VEC_LOOP_C_0_tr0,
      STAGE_LOOP_C_10_tr0
);
  input clk;
  input rst;
  output [8:0] fsm_output;
  reg [8:0] fsm_output;
  input STAGE_LOOP_C_9_tr0;
  input modExp_while_C_42_tr0;
  input COMP_LOOP_C_1_tr0;
  input COMP_LOOP_1_modExp_1_while_C_42_tr0;
  input COMP_LOOP_C_68_tr0;
  input COMP_LOOP_2_modExp_1_while_C_42_tr0;
  input COMP_LOOP_C_136_tr0;
  input COMP_LOOP_3_modExp_1_while_C_42_tr0;
  input COMP_LOOP_C_204_tr0;
  input COMP_LOOP_4_modExp_1_while_C_42_tr0;
  input COMP_LOOP_C_272_tr0;
  input VEC_LOOP_C_0_tr0;
  input STAGE_LOOP_C_10_tr0;


  // FSM State Type Declaration for inPlaceNTT_DIT_core_core_fsm_1
  parameter
    main_C_0 = 9'd0,
    STAGE_LOOP_C_0 = 9'd1,
    STAGE_LOOP_C_1 = 9'd2,
    STAGE_LOOP_C_2 = 9'd3,
    STAGE_LOOP_C_3 = 9'd4,
    STAGE_LOOP_C_4 = 9'd5,
    STAGE_LOOP_C_5 = 9'd6,
    STAGE_LOOP_C_6 = 9'd7,
    STAGE_LOOP_C_7 = 9'd8,
    STAGE_LOOP_C_8 = 9'd9,
    STAGE_LOOP_C_9 = 9'd10,
    modExp_while_C_0 = 9'd11,
    modExp_while_C_1 = 9'd12,
    modExp_while_C_2 = 9'd13,
    modExp_while_C_3 = 9'd14,
    modExp_while_C_4 = 9'd15,
    modExp_while_C_5 = 9'd16,
    modExp_while_C_6 = 9'd17,
    modExp_while_C_7 = 9'd18,
    modExp_while_C_8 = 9'd19,
    modExp_while_C_9 = 9'd20,
    modExp_while_C_10 = 9'd21,
    modExp_while_C_11 = 9'd22,
    modExp_while_C_12 = 9'd23,
    modExp_while_C_13 = 9'd24,
    modExp_while_C_14 = 9'd25,
    modExp_while_C_15 = 9'd26,
    modExp_while_C_16 = 9'd27,
    modExp_while_C_17 = 9'd28,
    modExp_while_C_18 = 9'd29,
    modExp_while_C_19 = 9'd30,
    modExp_while_C_20 = 9'd31,
    modExp_while_C_21 = 9'd32,
    modExp_while_C_22 = 9'd33,
    modExp_while_C_23 = 9'd34,
    modExp_while_C_24 = 9'd35,
    modExp_while_C_25 = 9'd36,
    modExp_while_C_26 = 9'd37,
    modExp_while_C_27 = 9'd38,
    modExp_while_C_28 = 9'd39,
    modExp_while_C_29 = 9'd40,
    modExp_while_C_30 = 9'd41,
    modExp_while_C_31 = 9'd42,
    modExp_while_C_32 = 9'd43,
    modExp_while_C_33 = 9'd44,
    modExp_while_C_34 = 9'd45,
    modExp_while_C_35 = 9'd46,
    modExp_while_C_36 = 9'd47,
    modExp_while_C_37 = 9'd48,
    modExp_while_C_38 = 9'd49,
    modExp_while_C_39 = 9'd50,
    modExp_while_C_40 = 9'd51,
    modExp_while_C_41 = 9'd52,
    modExp_while_C_42 = 9'd53,
    COMP_LOOP_C_0 = 9'd54,
    COMP_LOOP_C_1 = 9'd55,
    COMP_LOOP_1_modExp_1_while_C_0 = 9'd56,
    COMP_LOOP_1_modExp_1_while_C_1 = 9'd57,
    COMP_LOOP_1_modExp_1_while_C_2 = 9'd58,
    COMP_LOOP_1_modExp_1_while_C_3 = 9'd59,
    COMP_LOOP_1_modExp_1_while_C_4 = 9'd60,
    COMP_LOOP_1_modExp_1_while_C_5 = 9'd61,
    COMP_LOOP_1_modExp_1_while_C_6 = 9'd62,
    COMP_LOOP_1_modExp_1_while_C_7 = 9'd63,
    COMP_LOOP_1_modExp_1_while_C_8 = 9'd64,
    COMP_LOOP_1_modExp_1_while_C_9 = 9'd65,
    COMP_LOOP_1_modExp_1_while_C_10 = 9'd66,
    COMP_LOOP_1_modExp_1_while_C_11 = 9'd67,
    COMP_LOOP_1_modExp_1_while_C_12 = 9'd68,
    COMP_LOOP_1_modExp_1_while_C_13 = 9'd69,
    COMP_LOOP_1_modExp_1_while_C_14 = 9'd70,
    COMP_LOOP_1_modExp_1_while_C_15 = 9'd71,
    COMP_LOOP_1_modExp_1_while_C_16 = 9'd72,
    COMP_LOOP_1_modExp_1_while_C_17 = 9'd73,
    COMP_LOOP_1_modExp_1_while_C_18 = 9'd74,
    COMP_LOOP_1_modExp_1_while_C_19 = 9'd75,
    COMP_LOOP_1_modExp_1_while_C_20 = 9'd76,
    COMP_LOOP_1_modExp_1_while_C_21 = 9'd77,
    COMP_LOOP_1_modExp_1_while_C_22 = 9'd78,
    COMP_LOOP_1_modExp_1_while_C_23 = 9'd79,
    COMP_LOOP_1_modExp_1_while_C_24 = 9'd80,
    COMP_LOOP_1_modExp_1_while_C_25 = 9'd81,
    COMP_LOOP_1_modExp_1_while_C_26 = 9'd82,
    COMP_LOOP_1_modExp_1_while_C_27 = 9'd83,
    COMP_LOOP_1_modExp_1_while_C_28 = 9'd84,
    COMP_LOOP_1_modExp_1_while_C_29 = 9'd85,
    COMP_LOOP_1_modExp_1_while_C_30 = 9'd86,
    COMP_LOOP_1_modExp_1_while_C_31 = 9'd87,
    COMP_LOOP_1_modExp_1_while_C_32 = 9'd88,
    COMP_LOOP_1_modExp_1_while_C_33 = 9'd89,
    COMP_LOOP_1_modExp_1_while_C_34 = 9'd90,
    COMP_LOOP_1_modExp_1_while_C_35 = 9'd91,
    COMP_LOOP_1_modExp_1_while_C_36 = 9'd92,
    COMP_LOOP_1_modExp_1_while_C_37 = 9'd93,
    COMP_LOOP_1_modExp_1_while_C_38 = 9'd94,
    COMP_LOOP_1_modExp_1_while_C_39 = 9'd95,
    COMP_LOOP_1_modExp_1_while_C_40 = 9'd96,
    COMP_LOOP_1_modExp_1_while_C_41 = 9'd97,
    COMP_LOOP_1_modExp_1_while_C_42 = 9'd98,
    COMP_LOOP_C_2 = 9'd99,
    COMP_LOOP_C_3 = 9'd100,
    COMP_LOOP_C_4 = 9'd101,
    COMP_LOOP_C_5 = 9'd102,
    COMP_LOOP_C_6 = 9'd103,
    COMP_LOOP_C_7 = 9'd104,
    COMP_LOOP_C_8 = 9'd105,
    COMP_LOOP_C_9 = 9'd106,
    COMP_LOOP_C_10 = 9'd107,
    COMP_LOOP_C_11 = 9'd108,
    COMP_LOOP_C_12 = 9'd109,
    COMP_LOOP_C_13 = 9'd110,
    COMP_LOOP_C_14 = 9'd111,
    COMP_LOOP_C_15 = 9'd112,
    COMP_LOOP_C_16 = 9'd113,
    COMP_LOOP_C_17 = 9'd114,
    COMP_LOOP_C_18 = 9'd115,
    COMP_LOOP_C_19 = 9'd116,
    COMP_LOOP_C_20 = 9'd117,
    COMP_LOOP_C_21 = 9'd118,
    COMP_LOOP_C_22 = 9'd119,
    COMP_LOOP_C_23 = 9'd120,
    COMP_LOOP_C_24 = 9'd121,
    COMP_LOOP_C_25 = 9'd122,
    COMP_LOOP_C_26 = 9'd123,
    COMP_LOOP_C_27 = 9'd124,
    COMP_LOOP_C_28 = 9'd125,
    COMP_LOOP_C_29 = 9'd126,
    COMP_LOOP_C_30 = 9'd127,
    COMP_LOOP_C_31 = 9'd128,
    COMP_LOOP_C_32 = 9'd129,
    COMP_LOOP_C_33 = 9'd130,
    COMP_LOOP_C_34 = 9'd131,
    COMP_LOOP_C_35 = 9'd132,
    COMP_LOOP_C_36 = 9'd133,
    COMP_LOOP_C_37 = 9'd134,
    COMP_LOOP_C_38 = 9'd135,
    COMP_LOOP_C_39 = 9'd136,
    COMP_LOOP_C_40 = 9'd137,
    COMP_LOOP_C_41 = 9'd138,
    COMP_LOOP_C_42 = 9'd139,
    COMP_LOOP_C_43 = 9'd140,
    COMP_LOOP_C_44 = 9'd141,
    COMP_LOOP_C_45 = 9'd142,
    COMP_LOOP_C_46 = 9'd143,
    COMP_LOOP_C_47 = 9'd144,
    COMP_LOOP_C_48 = 9'd145,
    COMP_LOOP_C_49 = 9'd146,
    COMP_LOOP_C_50 = 9'd147,
    COMP_LOOP_C_51 = 9'd148,
    COMP_LOOP_C_52 = 9'd149,
    COMP_LOOP_C_53 = 9'd150,
    COMP_LOOP_C_54 = 9'd151,
    COMP_LOOP_C_55 = 9'd152,
    COMP_LOOP_C_56 = 9'd153,
    COMP_LOOP_C_57 = 9'd154,
    COMP_LOOP_C_58 = 9'd155,
    COMP_LOOP_C_59 = 9'd156,
    COMP_LOOP_C_60 = 9'd157,
    COMP_LOOP_C_61 = 9'd158,
    COMP_LOOP_C_62 = 9'd159,
    COMP_LOOP_C_63 = 9'd160,
    COMP_LOOP_C_64 = 9'd161,
    COMP_LOOP_C_65 = 9'd162,
    COMP_LOOP_C_66 = 9'd163,
    COMP_LOOP_C_67 = 9'd164,
    COMP_LOOP_C_68 = 9'd165,
    COMP_LOOP_C_69 = 9'd166,
    COMP_LOOP_2_modExp_1_while_C_0 = 9'd167,
    COMP_LOOP_2_modExp_1_while_C_1 = 9'd168,
    COMP_LOOP_2_modExp_1_while_C_2 = 9'd169,
    COMP_LOOP_2_modExp_1_while_C_3 = 9'd170,
    COMP_LOOP_2_modExp_1_while_C_4 = 9'd171,
    COMP_LOOP_2_modExp_1_while_C_5 = 9'd172,
    COMP_LOOP_2_modExp_1_while_C_6 = 9'd173,
    COMP_LOOP_2_modExp_1_while_C_7 = 9'd174,
    COMP_LOOP_2_modExp_1_while_C_8 = 9'd175,
    COMP_LOOP_2_modExp_1_while_C_9 = 9'd176,
    COMP_LOOP_2_modExp_1_while_C_10 = 9'd177,
    COMP_LOOP_2_modExp_1_while_C_11 = 9'd178,
    COMP_LOOP_2_modExp_1_while_C_12 = 9'd179,
    COMP_LOOP_2_modExp_1_while_C_13 = 9'd180,
    COMP_LOOP_2_modExp_1_while_C_14 = 9'd181,
    COMP_LOOP_2_modExp_1_while_C_15 = 9'd182,
    COMP_LOOP_2_modExp_1_while_C_16 = 9'd183,
    COMP_LOOP_2_modExp_1_while_C_17 = 9'd184,
    COMP_LOOP_2_modExp_1_while_C_18 = 9'd185,
    COMP_LOOP_2_modExp_1_while_C_19 = 9'd186,
    COMP_LOOP_2_modExp_1_while_C_20 = 9'd187,
    COMP_LOOP_2_modExp_1_while_C_21 = 9'd188,
    COMP_LOOP_2_modExp_1_while_C_22 = 9'd189,
    COMP_LOOP_2_modExp_1_while_C_23 = 9'd190,
    COMP_LOOP_2_modExp_1_while_C_24 = 9'd191,
    COMP_LOOP_2_modExp_1_while_C_25 = 9'd192,
    COMP_LOOP_2_modExp_1_while_C_26 = 9'd193,
    COMP_LOOP_2_modExp_1_while_C_27 = 9'd194,
    COMP_LOOP_2_modExp_1_while_C_28 = 9'd195,
    COMP_LOOP_2_modExp_1_while_C_29 = 9'd196,
    COMP_LOOP_2_modExp_1_while_C_30 = 9'd197,
    COMP_LOOP_2_modExp_1_while_C_31 = 9'd198,
    COMP_LOOP_2_modExp_1_while_C_32 = 9'd199,
    COMP_LOOP_2_modExp_1_while_C_33 = 9'd200,
    COMP_LOOP_2_modExp_1_while_C_34 = 9'd201,
    COMP_LOOP_2_modExp_1_while_C_35 = 9'd202,
    COMP_LOOP_2_modExp_1_while_C_36 = 9'd203,
    COMP_LOOP_2_modExp_1_while_C_37 = 9'd204,
    COMP_LOOP_2_modExp_1_while_C_38 = 9'd205,
    COMP_LOOP_2_modExp_1_while_C_39 = 9'd206,
    COMP_LOOP_2_modExp_1_while_C_40 = 9'd207,
    COMP_LOOP_2_modExp_1_while_C_41 = 9'd208,
    COMP_LOOP_2_modExp_1_while_C_42 = 9'd209,
    COMP_LOOP_C_70 = 9'd210,
    COMP_LOOP_C_71 = 9'd211,
    COMP_LOOP_C_72 = 9'd212,
    COMP_LOOP_C_73 = 9'd213,
    COMP_LOOP_C_74 = 9'd214,
    COMP_LOOP_C_75 = 9'd215,
    COMP_LOOP_C_76 = 9'd216,
    COMP_LOOP_C_77 = 9'd217,
    COMP_LOOP_C_78 = 9'd218,
    COMP_LOOP_C_79 = 9'd219,
    COMP_LOOP_C_80 = 9'd220,
    COMP_LOOP_C_81 = 9'd221,
    COMP_LOOP_C_82 = 9'd222,
    COMP_LOOP_C_83 = 9'd223,
    COMP_LOOP_C_84 = 9'd224,
    COMP_LOOP_C_85 = 9'd225,
    COMP_LOOP_C_86 = 9'd226,
    COMP_LOOP_C_87 = 9'd227,
    COMP_LOOP_C_88 = 9'd228,
    COMP_LOOP_C_89 = 9'd229,
    COMP_LOOP_C_90 = 9'd230,
    COMP_LOOP_C_91 = 9'd231,
    COMP_LOOP_C_92 = 9'd232,
    COMP_LOOP_C_93 = 9'd233,
    COMP_LOOP_C_94 = 9'd234,
    COMP_LOOP_C_95 = 9'd235,
    COMP_LOOP_C_96 = 9'd236,
    COMP_LOOP_C_97 = 9'd237,
    COMP_LOOP_C_98 = 9'd238,
    COMP_LOOP_C_99 = 9'd239,
    COMP_LOOP_C_100 = 9'd240,
    COMP_LOOP_C_101 = 9'd241,
    COMP_LOOP_C_102 = 9'd242,
    COMP_LOOP_C_103 = 9'd243,
    COMP_LOOP_C_104 = 9'd244,
    COMP_LOOP_C_105 = 9'd245,
    COMP_LOOP_C_106 = 9'd246,
    COMP_LOOP_C_107 = 9'd247,
    COMP_LOOP_C_108 = 9'd248,
    COMP_LOOP_C_109 = 9'd249,
    COMP_LOOP_C_110 = 9'd250,
    COMP_LOOP_C_111 = 9'd251,
    COMP_LOOP_C_112 = 9'd252,
    COMP_LOOP_C_113 = 9'd253,
    COMP_LOOP_C_114 = 9'd254,
    COMP_LOOP_C_115 = 9'd255,
    COMP_LOOP_C_116 = 9'd256,
    COMP_LOOP_C_117 = 9'd257,
    COMP_LOOP_C_118 = 9'd258,
    COMP_LOOP_C_119 = 9'd259,
    COMP_LOOP_C_120 = 9'd260,
    COMP_LOOP_C_121 = 9'd261,
    COMP_LOOP_C_122 = 9'd262,
    COMP_LOOP_C_123 = 9'd263,
    COMP_LOOP_C_124 = 9'd264,
    COMP_LOOP_C_125 = 9'd265,
    COMP_LOOP_C_126 = 9'd266,
    COMP_LOOP_C_127 = 9'd267,
    COMP_LOOP_C_128 = 9'd268,
    COMP_LOOP_C_129 = 9'd269,
    COMP_LOOP_C_130 = 9'd270,
    COMP_LOOP_C_131 = 9'd271,
    COMP_LOOP_C_132 = 9'd272,
    COMP_LOOP_C_133 = 9'd273,
    COMP_LOOP_C_134 = 9'd274,
    COMP_LOOP_C_135 = 9'd275,
    COMP_LOOP_C_136 = 9'd276,
    COMP_LOOP_C_137 = 9'd277,
    COMP_LOOP_3_modExp_1_while_C_0 = 9'd278,
    COMP_LOOP_3_modExp_1_while_C_1 = 9'd279,
    COMP_LOOP_3_modExp_1_while_C_2 = 9'd280,
    COMP_LOOP_3_modExp_1_while_C_3 = 9'd281,
    COMP_LOOP_3_modExp_1_while_C_4 = 9'd282,
    COMP_LOOP_3_modExp_1_while_C_5 = 9'd283,
    COMP_LOOP_3_modExp_1_while_C_6 = 9'd284,
    COMP_LOOP_3_modExp_1_while_C_7 = 9'd285,
    COMP_LOOP_3_modExp_1_while_C_8 = 9'd286,
    COMP_LOOP_3_modExp_1_while_C_9 = 9'd287,
    COMP_LOOP_3_modExp_1_while_C_10 = 9'd288,
    COMP_LOOP_3_modExp_1_while_C_11 = 9'd289,
    COMP_LOOP_3_modExp_1_while_C_12 = 9'd290,
    COMP_LOOP_3_modExp_1_while_C_13 = 9'd291,
    COMP_LOOP_3_modExp_1_while_C_14 = 9'd292,
    COMP_LOOP_3_modExp_1_while_C_15 = 9'd293,
    COMP_LOOP_3_modExp_1_while_C_16 = 9'd294,
    COMP_LOOP_3_modExp_1_while_C_17 = 9'd295,
    COMP_LOOP_3_modExp_1_while_C_18 = 9'd296,
    COMP_LOOP_3_modExp_1_while_C_19 = 9'd297,
    COMP_LOOP_3_modExp_1_while_C_20 = 9'd298,
    COMP_LOOP_3_modExp_1_while_C_21 = 9'd299,
    COMP_LOOP_3_modExp_1_while_C_22 = 9'd300,
    COMP_LOOP_3_modExp_1_while_C_23 = 9'd301,
    COMP_LOOP_3_modExp_1_while_C_24 = 9'd302,
    COMP_LOOP_3_modExp_1_while_C_25 = 9'd303,
    COMP_LOOP_3_modExp_1_while_C_26 = 9'd304,
    COMP_LOOP_3_modExp_1_while_C_27 = 9'd305,
    COMP_LOOP_3_modExp_1_while_C_28 = 9'd306,
    COMP_LOOP_3_modExp_1_while_C_29 = 9'd307,
    COMP_LOOP_3_modExp_1_while_C_30 = 9'd308,
    COMP_LOOP_3_modExp_1_while_C_31 = 9'd309,
    COMP_LOOP_3_modExp_1_while_C_32 = 9'd310,
    COMP_LOOP_3_modExp_1_while_C_33 = 9'd311,
    COMP_LOOP_3_modExp_1_while_C_34 = 9'd312,
    COMP_LOOP_3_modExp_1_while_C_35 = 9'd313,
    COMP_LOOP_3_modExp_1_while_C_36 = 9'd314,
    COMP_LOOP_3_modExp_1_while_C_37 = 9'd315,
    COMP_LOOP_3_modExp_1_while_C_38 = 9'd316,
    COMP_LOOP_3_modExp_1_while_C_39 = 9'd317,
    COMP_LOOP_3_modExp_1_while_C_40 = 9'd318,
    COMP_LOOP_3_modExp_1_while_C_41 = 9'd319,
    COMP_LOOP_3_modExp_1_while_C_42 = 9'd320,
    COMP_LOOP_C_138 = 9'd321,
    COMP_LOOP_C_139 = 9'd322,
    COMP_LOOP_C_140 = 9'd323,
    COMP_LOOP_C_141 = 9'd324,
    COMP_LOOP_C_142 = 9'd325,
    COMP_LOOP_C_143 = 9'd326,
    COMP_LOOP_C_144 = 9'd327,
    COMP_LOOP_C_145 = 9'd328,
    COMP_LOOP_C_146 = 9'd329,
    COMP_LOOP_C_147 = 9'd330,
    COMP_LOOP_C_148 = 9'd331,
    COMP_LOOP_C_149 = 9'd332,
    COMP_LOOP_C_150 = 9'd333,
    COMP_LOOP_C_151 = 9'd334,
    COMP_LOOP_C_152 = 9'd335,
    COMP_LOOP_C_153 = 9'd336,
    COMP_LOOP_C_154 = 9'd337,
    COMP_LOOP_C_155 = 9'd338,
    COMP_LOOP_C_156 = 9'd339,
    COMP_LOOP_C_157 = 9'd340,
    COMP_LOOP_C_158 = 9'd341,
    COMP_LOOP_C_159 = 9'd342,
    COMP_LOOP_C_160 = 9'd343,
    COMP_LOOP_C_161 = 9'd344,
    COMP_LOOP_C_162 = 9'd345,
    COMP_LOOP_C_163 = 9'd346,
    COMP_LOOP_C_164 = 9'd347,
    COMP_LOOP_C_165 = 9'd348,
    COMP_LOOP_C_166 = 9'd349,
    COMP_LOOP_C_167 = 9'd350,
    COMP_LOOP_C_168 = 9'd351,
    COMP_LOOP_C_169 = 9'd352,
    COMP_LOOP_C_170 = 9'd353,
    COMP_LOOP_C_171 = 9'd354,
    COMP_LOOP_C_172 = 9'd355,
    COMP_LOOP_C_173 = 9'd356,
    COMP_LOOP_C_174 = 9'd357,
    COMP_LOOP_C_175 = 9'd358,
    COMP_LOOP_C_176 = 9'd359,
    COMP_LOOP_C_177 = 9'd360,
    COMP_LOOP_C_178 = 9'd361,
    COMP_LOOP_C_179 = 9'd362,
    COMP_LOOP_C_180 = 9'd363,
    COMP_LOOP_C_181 = 9'd364,
    COMP_LOOP_C_182 = 9'd365,
    COMP_LOOP_C_183 = 9'd366,
    COMP_LOOP_C_184 = 9'd367,
    COMP_LOOP_C_185 = 9'd368,
    COMP_LOOP_C_186 = 9'd369,
    COMP_LOOP_C_187 = 9'd370,
    COMP_LOOP_C_188 = 9'd371,
    COMP_LOOP_C_189 = 9'd372,
    COMP_LOOP_C_190 = 9'd373,
    COMP_LOOP_C_191 = 9'd374,
    COMP_LOOP_C_192 = 9'd375,
    COMP_LOOP_C_193 = 9'd376,
    COMP_LOOP_C_194 = 9'd377,
    COMP_LOOP_C_195 = 9'd378,
    COMP_LOOP_C_196 = 9'd379,
    COMP_LOOP_C_197 = 9'd380,
    COMP_LOOP_C_198 = 9'd381,
    COMP_LOOP_C_199 = 9'd382,
    COMP_LOOP_C_200 = 9'd383,
    COMP_LOOP_C_201 = 9'd384,
    COMP_LOOP_C_202 = 9'd385,
    COMP_LOOP_C_203 = 9'd386,
    COMP_LOOP_C_204 = 9'd387,
    COMP_LOOP_C_205 = 9'd388,
    COMP_LOOP_4_modExp_1_while_C_0 = 9'd389,
    COMP_LOOP_4_modExp_1_while_C_1 = 9'd390,
    COMP_LOOP_4_modExp_1_while_C_2 = 9'd391,
    COMP_LOOP_4_modExp_1_while_C_3 = 9'd392,
    COMP_LOOP_4_modExp_1_while_C_4 = 9'd393,
    COMP_LOOP_4_modExp_1_while_C_5 = 9'd394,
    COMP_LOOP_4_modExp_1_while_C_6 = 9'd395,
    COMP_LOOP_4_modExp_1_while_C_7 = 9'd396,
    COMP_LOOP_4_modExp_1_while_C_8 = 9'd397,
    COMP_LOOP_4_modExp_1_while_C_9 = 9'd398,
    COMP_LOOP_4_modExp_1_while_C_10 = 9'd399,
    COMP_LOOP_4_modExp_1_while_C_11 = 9'd400,
    COMP_LOOP_4_modExp_1_while_C_12 = 9'd401,
    COMP_LOOP_4_modExp_1_while_C_13 = 9'd402,
    COMP_LOOP_4_modExp_1_while_C_14 = 9'd403,
    COMP_LOOP_4_modExp_1_while_C_15 = 9'd404,
    COMP_LOOP_4_modExp_1_while_C_16 = 9'd405,
    COMP_LOOP_4_modExp_1_while_C_17 = 9'd406,
    COMP_LOOP_4_modExp_1_while_C_18 = 9'd407,
    COMP_LOOP_4_modExp_1_while_C_19 = 9'd408,
    COMP_LOOP_4_modExp_1_while_C_20 = 9'd409,
    COMP_LOOP_4_modExp_1_while_C_21 = 9'd410,
    COMP_LOOP_4_modExp_1_while_C_22 = 9'd411,
    COMP_LOOP_4_modExp_1_while_C_23 = 9'd412,
    COMP_LOOP_4_modExp_1_while_C_24 = 9'd413,
    COMP_LOOP_4_modExp_1_while_C_25 = 9'd414,
    COMP_LOOP_4_modExp_1_while_C_26 = 9'd415,
    COMP_LOOP_4_modExp_1_while_C_27 = 9'd416,
    COMP_LOOP_4_modExp_1_while_C_28 = 9'd417,
    COMP_LOOP_4_modExp_1_while_C_29 = 9'd418,
    COMP_LOOP_4_modExp_1_while_C_30 = 9'd419,
    COMP_LOOP_4_modExp_1_while_C_31 = 9'd420,
    COMP_LOOP_4_modExp_1_while_C_32 = 9'd421,
    COMP_LOOP_4_modExp_1_while_C_33 = 9'd422,
    COMP_LOOP_4_modExp_1_while_C_34 = 9'd423,
    COMP_LOOP_4_modExp_1_while_C_35 = 9'd424,
    COMP_LOOP_4_modExp_1_while_C_36 = 9'd425,
    COMP_LOOP_4_modExp_1_while_C_37 = 9'd426,
    COMP_LOOP_4_modExp_1_while_C_38 = 9'd427,
    COMP_LOOP_4_modExp_1_while_C_39 = 9'd428,
    COMP_LOOP_4_modExp_1_while_C_40 = 9'd429,
    COMP_LOOP_4_modExp_1_while_C_41 = 9'd430,
    COMP_LOOP_4_modExp_1_while_C_42 = 9'd431,
    COMP_LOOP_C_206 = 9'd432,
    COMP_LOOP_C_207 = 9'd433,
    COMP_LOOP_C_208 = 9'd434,
    COMP_LOOP_C_209 = 9'd435,
    COMP_LOOP_C_210 = 9'd436,
    COMP_LOOP_C_211 = 9'd437,
    COMP_LOOP_C_212 = 9'd438,
    COMP_LOOP_C_213 = 9'd439,
    COMP_LOOP_C_214 = 9'd440,
    COMP_LOOP_C_215 = 9'd441,
    COMP_LOOP_C_216 = 9'd442,
    COMP_LOOP_C_217 = 9'd443,
    COMP_LOOP_C_218 = 9'd444,
    COMP_LOOP_C_219 = 9'd445,
    COMP_LOOP_C_220 = 9'd446,
    COMP_LOOP_C_221 = 9'd447,
    COMP_LOOP_C_222 = 9'd448,
    COMP_LOOP_C_223 = 9'd449,
    COMP_LOOP_C_224 = 9'd450,
    COMP_LOOP_C_225 = 9'd451,
    COMP_LOOP_C_226 = 9'd452,
    COMP_LOOP_C_227 = 9'd453,
    COMP_LOOP_C_228 = 9'd454,
    COMP_LOOP_C_229 = 9'd455,
    COMP_LOOP_C_230 = 9'd456,
    COMP_LOOP_C_231 = 9'd457,
    COMP_LOOP_C_232 = 9'd458,
    COMP_LOOP_C_233 = 9'd459,
    COMP_LOOP_C_234 = 9'd460,
    COMP_LOOP_C_235 = 9'd461,
    COMP_LOOP_C_236 = 9'd462,
    COMP_LOOP_C_237 = 9'd463,
    COMP_LOOP_C_238 = 9'd464,
    COMP_LOOP_C_239 = 9'd465,
    COMP_LOOP_C_240 = 9'd466,
    COMP_LOOP_C_241 = 9'd467,
    COMP_LOOP_C_242 = 9'd468,
    COMP_LOOP_C_243 = 9'd469,
    COMP_LOOP_C_244 = 9'd470,
    COMP_LOOP_C_245 = 9'd471,
    COMP_LOOP_C_246 = 9'd472,
    COMP_LOOP_C_247 = 9'd473,
    COMP_LOOP_C_248 = 9'd474,
    COMP_LOOP_C_249 = 9'd475,
    COMP_LOOP_C_250 = 9'd476,
    COMP_LOOP_C_251 = 9'd477,
    COMP_LOOP_C_252 = 9'd478,
    COMP_LOOP_C_253 = 9'd479,
    COMP_LOOP_C_254 = 9'd480,
    COMP_LOOP_C_255 = 9'd481,
    COMP_LOOP_C_256 = 9'd482,
    COMP_LOOP_C_257 = 9'd483,
    COMP_LOOP_C_258 = 9'd484,
    COMP_LOOP_C_259 = 9'd485,
    COMP_LOOP_C_260 = 9'd486,
    COMP_LOOP_C_261 = 9'd487,
    COMP_LOOP_C_262 = 9'd488,
    COMP_LOOP_C_263 = 9'd489,
    COMP_LOOP_C_264 = 9'd490,
    COMP_LOOP_C_265 = 9'd491,
    COMP_LOOP_C_266 = 9'd492,
    COMP_LOOP_C_267 = 9'd493,
    COMP_LOOP_C_268 = 9'd494,
    COMP_LOOP_C_269 = 9'd495,
    COMP_LOOP_C_270 = 9'd496,
    COMP_LOOP_C_271 = 9'd497,
    COMP_LOOP_C_272 = 9'd498,
    VEC_LOOP_C_0 = 9'd499,
    STAGE_LOOP_C_10 = 9'd500,
    main_C_1 = 9'd501;

  reg [8:0] state_var;
  reg [8:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : inPlaceNTT_DIT_core_core_fsm_1
    case (state_var)
      STAGE_LOOP_C_0 : begin
        fsm_output = 9'b000000001;
        state_var_NS = STAGE_LOOP_C_1;
      end
      STAGE_LOOP_C_1 : begin
        fsm_output = 9'b000000010;
        state_var_NS = STAGE_LOOP_C_2;
      end
      STAGE_LOOP_C_2 : begin
        fsm_output = 9'b000000011;
        state_var_NS = STAGE_LOOP_C_3;
      end
      STAGE_LOOP_C_3 : begin
        fsm_output = 9'b000000100;
        state_var_NS = STAGE_LOOP_C_4;
      end
      STAGE_LOOP_C_4 : begin
        fsm_output = 9'b000000101;
        state_var_NS = STAGE_LOOP_C_5;
      end
      STAGE_LOOP_C_5 : begin
        fsm_output = 9'b000000110;
        state_var_NS = STAGE_LOOP_C_6;
      end
      STAGE_LOOP_C_6 : begin
        fsm_output = 9'b000000111;
        state_var_NS = STAGE_LOOP_C_7;
      end
      STAGE_LOOP_C_7 : begin
        fsm_output = 9'b000001000;
        state_var_NS = STAGE_LOOP_C_8;
      end
      STAGE_LOOP_C_8 : begin
        fsm_output = 9'b000001001;
        state_var_NS = STAGE_LOOP_C_9;
      end
      STAGE_LOOP_C_9 : begin
        fsm_output = 9'b000001010;
        if ( STAGE_LOOP_C_9_tr0 ) begin
          state_var_NS = COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_while_C_0;
        end
      end
      modExp_while_C_0 : begin
        fsm_output = 9'b000001011;
        state_var_NS = modExp_while_C_1;
      end
      modExp_while_C_1 : begin
        fsm_output = 9'b000001100;
        state_var_NS = modExp_while_C_2;
      end
      modExp_while_C_2 : begin
        fsm_output = 9'b000001101;
        state_var_NS = modExp_while_C_3;
      end
      modExp_while_C_3 : begin
        fsm_output = 9'b000001110;
        state_var_NS = modExp_while_C_4;
      end
      modExp_while_C_4 : begin
        fsm_output = 9'b000001111;
        state_var_NS = modExp_while_C_5;
      end
      modExp_while_C_5 : begin
        fsm_output = 9'b000010000;
        state_var_NS = modExp_while_C_6;
      end
      modExp_while_C_6 : begin
        fsm_output = 9'b000010001;
        state_var_NS = modExp_while_C_7;
      end
      modExp_while_C_7 : begin
        fsm_output = 9'b000010010;
        state_var_NS = modExp_while_C_8;
      end
      modExp_while_C_8 : begin
        fsm_output = 9'b000010011;
        state_var_NS = modExp_while_C_9;
      end
      modExp_while_C_9 : begin
        fsm_output = 9'b000010100;
        state_var_NS = modExp_while_C_10;
      end
      modExp_while_C_10 : begin
        fsm_output = 9'b000010101;
        state_var_NS = modExp_while_C_11;
      end
      modExp_while_C_11 : begin
        fsm_output = 9'b000010110;
        state_var_NS = modExp_while_C_12;
      end
      modExp_while_C_12 : begin
        fsm_output = 9'b000010111;
        state_var_NS = modExp_while_C_13;
      end
      modExp_while_C_13 : begin
        fsm_output = 9'b000011000;
        state_var_NS = modExp_while_C_14;
      end
      modExp_while_C_14 : begin
        fsm_output = 9'b000011001;
        state_var_NS = modExp_while_C_15;
      end
      modExp_while_C_15 : begin
        fsm_output = 9'b000011010;
        state_var_NS = modExp_while_C_16;
      end
      modExp_while_C_16 : begin
        fsm_output = 9'b000011011;
        state_var_NS = modExp_while_C_17;
      end
      modExp_while_C_17 : begin
        fsm_output = 9'b000011100;
        state_var_NS = modExp_while_C_18;
      end
      modExp_while_C_18 : begin
        fsm_output = 9'b000011101;
        state_var_NS = modExp_while_C_19;
      end
      modExp_while_C_19 : begin
        fsm_output = 9'b000011110;
        state_var_NS = modExp_while_C_20;
      end
      modExp_while_C_20 : begin
        fsm_output = 9'b000011111;
        state_var_NS = modExp_while_C_21;
      end
      modExp_while_C_21 : begin
        fsm_output = 9'b000100000;
        state_var_NS = modExp_while_C_22;
      end
      modExp_while_C_22 : begin
        fsm_output = 9'b000100001;
        state_var_NS = modExp_while_C_23;
      end
      modExp_while_C_23 : begin
        fsm_output = 9'b000100010;
        state_var_NS = modExp_while_C_24;
      end
      modExp_while_C_24 : begin
        fsm_output = 9'b000100011;
        state_var_NS = modExp_while_C_25;
      end
      modExp_while_C_25 : begin
        fsm_output = 9'b000100100;
        state_var_NS = modExp_while_C_26;
      end
      modExp_while_C_26 : begin
        fsm_output = 9'b000100101;
        state_var_NS = modExp_while_C_27;
      end
      modExp_while_C_27 : begin
        fsm_output = 9'b000100110;
        state_var_NS = modExp_while_C_28;
      end
      modExp_while_C_28 : begin
        fsm_output = 9'b000100111;
        state_var_NS = modExp_while_C_29;
      end
      modExp_while_C_29 : begin
        fsm_output = 9'b000101000;
        state_var_NS = modExp_while_C_30;
      end
      modExp_while_C_30 : begin
        fsm_output = 9'b000101001;
        state_var_NS = modExp_while_C_31;
      end
      modExp_while_C_31 : begin
        fsm_output = 9'b000101010;
        state_var_NS = modExp_while_C_32;
      end
      modExp_while_C_32 : begin
        fsm_output = 9'b000101011;
        state_var_NS = modExp_while_C_33;
      end
      modExp_while_C_33 : begin
        fsm_output = 9'b000101100;
        state_var_NS = modExp_while_C_34;
      end
      modExp_while_C_34 : begin
        fsm_output = 9'b000101101;
        state_var_NS = modExp_while_C_35;
      end
      modExp_while_C_35 : begin
        fsm_output = 9'b000101110;
        state_var_NS = modExp_while_C_36;
      end
      modExp_while_C_36 : begin
        fsm_output = 9'b000101111;
        state_var_NS = modExp_while_C_37;
      end
      modExp_while_C_37 : begin
        fsm_output = 9'b000110000;
        state_var_NS = modExp_while_C_38;
      end
      modExp_while_C_38 : begin
        fsm_output = 9'b000110001;
        state_var_NS = modExp_while_C_39;
      end
      modExp_while_C_39 : begin
        fsm_output = 9'b000110010;
        state_var_NS = modExp_while_C_40;
      end
      modExp_while_C_40 : begin
        fsm_output = 9'b000110011;
        state_var_NS = modExp_while_C_41;
      end
      modExp_while_C_41 : begin
        fsm_output = 9'b000110100;
        state_var_NS = modExp_while_C_42;
      end
      modExp_while_C_42 : begin
        fsm_output = 9'b000110101;
        if ( modExp_while_C_42_tr0 ) begin
          state_var_NS = COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_while_C_0;
        end
      end
      COMP_LOOP_C_0 : begin
        fsm_output = 9'b000110110;
        state_var_NS = COMP_LOOP_C_1;
      end
      COMP_LOOP_C_1 : begin
        fsm_output = 9'b000110111;
        if ( COMP_LOOP_C_1_tr0 ) begin
          state_var_NS = COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_1_modExp_1_while_C_0 : begin
        fsm_output = 9'b000111000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_1;
      end
      COMP_LOOP_1_modExp_1_while_C_1 : begin
        fsm_output = 9'b000111001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_2;
      end
      COMP_LOOP_1_modExp_1_while_C_2 : begin
        fsm_output = 9'b000111010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_3;
      end
      COMP_LOOP_1_modExp_1_while_C_3 : begin
        fsm_output = 9'b000111011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_4;
      end
      COMP_LOOP_1_modExp_1_while_C_4 : begin
        fsm_output = 9'b000111100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_5;
      end
      COMP_LOOP_1_modExp_1_while_C_5 : begin
        fsm_output = 9'b000111101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_6;
      end
      COMP_LOOP_1_modExp_1_while_C_6 : begin
        fsm_output = 9'b000111110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_7;
      end
      COMP_LOOP_1_modExp_1_while_C_7 : begin
        fsm_output = 9'b000111111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_8;
      end
      COMP_LOOP_1_modExp_1_while_C_8 : begin
        fsm_output = 9'b001000000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_9;
      end
      COMP_LOOP_1_modExp_1_while_C_9 : begin
        fsm_output = 9'b001000001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_10;
      end
      COMP_LOOP_1_modExp_1_while_C_10 : begin
        fsm_output = 9'b001000010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_11;
      end
      COMP_LOOP_1_modExp_1_while_C_11 : begin
        fsm_output = 9'b001000011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_12;
      end
      COMP_LOOP_1_modExp_1_while_C_12 : begin
        fsm_output = 9'b001000100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_13;
      end
      COMP_LOOP_1_modExp_1_while_C_13 : begin
        fsm_output = 9'b001000101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_14;
      end
      COMP_LOOP_1_modExp_1_while_C_14 : begin
        fsm_output = 9'b001000110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_15;
      end
      COMP_LOOP_1_modExp_1_while_C_15 : begin
        fsm_output = 9'b001000111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_16;
      end
      COMP_LOOP_1_modExp_1_while_C_16 : begin
        fsm_output = 9'b001001000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_17;
      end
      COMP_LOOP_1_modExp_1_while_C_17 : begin
        fsm_output = 9'b001001001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_18;
      end
      COMP_LOOP_1_modExp_1_while_C_18 : begin
        fsm_output = 9'b001001010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_19;
      end
      COMP_LOOP_1_modExp_1_while_C_19 : begin
        fsm_output = 9'b001001011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_20;
      end
      COMP_LOOP_1_modExp_1_while_C_20 : begin
        fsm_output = 9'b001001100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_21;
      end
      COMP_LOOP_1_modExp_1_while_C_21 : begin
        fsm_output = 9'b001001101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_22;
      end
      COMP_LOOP_1_modExp_1_while_C_22 : begin
        fsm_output = 9'b001001110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_23;
      end
      COMP_LOOP_1_modExp_1_while_C_23 : begin
        fsm_output = 9'b001001111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_24;
      end
      COMP_LOOP_1_modExp_1_while_C_24 : begin
        fsm_output = 9'b001010000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_25;
      end
      COMP_LOOP_1_modExp_1_while_C_25 : begin
        fsm_output = 9'b001010001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_26;
      end
      COMP_LOOP_1_modExp_1_while_C_26 : begin
        fsm_output = 9'b001010010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_27;
      end
      COMP_LOOP_1_modExp_1_while_C_27 : begin
        fsm_output = 9'b001010011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_28;
      end
      COMP_LOOP_1_modExp_1_while_C_28 : begin
        fsm_output = 9'b001010100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_29;
      end
      COMP_LOOP_1_modExp_1_while_C_29 : begin
        fsm_output = 9'b001010101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_30;
      end
      COMP_LOOP_1_modExp_1_while_C_30 : begin
        fsm_output = 9'b001010110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_31;
      end
      COMP_LOOP_1_modExp_1_while_C_31 : begin
        fsm_output = 9'b001010111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_32;
      end
      COMP_LOOP_1_modExp_1_while_C_32 : begin
        fsm_output = 9'b001011000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_33;
      end
      COMP_LOOP_1_modExp_1_while_C_33 : begin
        fsm_output = 9'b001011001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_34;
      end
      COMP_LOOP_1_modExp_1_while_C_34 : begin
        fsm_output = 9'b001011010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_35;
      end
      COMP_LOOP_1_modExp_1_while_C_35 : begin
        fsm_output = 9'b001011011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_36;
      end
      COMP_LOOP_1_modExp_1_while_C_36 : begin
        fsm_output = 9'b001011100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_37;
      end
      COMP_LOOP_1_modExp_1_while_C_37 : begin
        fsm_output = 9'b001011101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_38;
      end
      COMP_LOOP_1_modExp_1_while_C_38 : begin
        fsm_output = 9'b001011110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_39;
      end
      COMP_LOOP_1_modExp_1_while_C_39 : begin
        fsm_output = 9'b001011111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_40;
      end
      COMP_LOOP_1_modExp_1_while_C_40 : begin
        fsm_output = 9'b001100000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_41;
      end
      COMP_LOOP_1_modExp_1_while_C_41 : begin
        fsm_output = 9'b001100001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_42;
      end
      COMP_LOOP_1_modExp_1_while_C_42 : begin
        fsm_output = 9'b001100010;
        if ( COMP_LOOP_1_modExp_1_while_C_42_tr0 ) begin
          state_var_NS = COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_2 : begin
        fsm_output = 9'b001100011;
        state_var_NS = COMP_LOOP_C_3;
      end
      COMP_LOOP_C_3 : begin
        fsm_output = 9'b001100100;
        state_var_NS = COMP_LOOP_C_4;
      end
      COMP_LOOP_C_4 : begin
        fsm_output = 9'b001100101;
        state_var_NS = COMP_LOOP_C_5;
      end
      COMP_LOOP_C_5 : begin
        fsm_output = 9'b001100110;
        state_var_NS = COMP_LOOP_C_6;
      end
      COMP_LOOP_C_6 : begin
        fsm_output = 9'b001100111;
        state_var_NS = COMP_LOOP_C_7;
      end
      COMP_LOOP_C_7 : begin
        fsm_output = 9'b001101000;
        state_var_NS = COMP_LOOP_C_8;
      end
      COMP_LOOP_C_8 : begin
        fsm_output = 9'b001101001;
        state_var_NS = COMP_LOOP_C_9;
      end
      COMP_LOOP_C_9 : begin
        fsm_output = 9'b001101010;
        state_var_NS = COMP_LOOP_C_10;
      end
      COMP_LOOP_C_10 : begin
        fsm_output = 9'b001101011;
        state_var_NS = COMP_LOOP_C_11;
      end
      COMP_LOOP_C_11 : begin
        fsm_output = 9'b001101100;
        state_var_NS = COMP_LOOP_C_12;
      end
      COMP_LOOP_C_12 : begin
        fsm_output = 9'b001101101;
        state_var_NS = COMP_LOOP_C_13;
      end
      COMP_LOOP_C_13 : begin
        fsm_output = 9'b001101110;
        state_var_NS = COMP_LOOP_C_14;
      end
      COMP_LOOP_C_14 : begin
        fsm_output = 9'b001101111;
        state_var_NS = COMP_LOOP_C_15;
      end
      COMP_LOOP_C_15 : begin
        fsm_output = 9'b001110000;
        state_var_NS = COMP_LOOP_C_16;
      end
      COMP_LOOP_C_16 : begin
        fsm_output = 9'b001110001;
        state_var_NS = COMP_LOOP_C_17;
      end
      COMP_LOOP_C_17 : begin
        fsm_output = 9'b001110010;
        state_var_NS = COMP_LOOP_C_18;
      end
      COMP_LOOP_C_18 : begin
        fsm_output = 9'b001110011;
        state_var_NS = COMP_LOOP_C_19;
      end
      COMP_LOOP_C_19 : begin
        fsm_output = 9'b001110100;
        state_var_NS = COMP_LOOP_C_20;
      end
      COMP_LOOP_C_20 : begin
        fsm_output = 9'b001110101;
        state_var_NS = COMP_LOOP_C_21;
      end
      COMP_LOOP_C_21 : begin
        fsm_output = 9'b001110110;
        state_var_NS = COMP_LOOP_C_22;
      end
      COMP_LOOP_C_22 : begin
        fsm_output = 9'b001110111;
        state_var_NS = COMP_LOOP_C_23;
      end
      COMP_LOOP_C_23 : begin
        fsm_output = 9'b001111000;
        state_var_NS = COMP_LOOP_C_24;
      end
      COMP_LOOP_C_24 : begin
        fsm_output = 9'b001111001;
        state_var_NS = COMP_LOOP_C_25;
      end
      COMP_LOOP_C_25 : begin
        fsm_output = 9'b001111010;
        state_var_NS = COMP_LOOP_C_26;
      end
      COMP_LOOP_C_26 : begin
        fsm_output = 9'b001111011;
        state_var_NS = COMP_LOOP_C_27;
      end
      COMP_LOOP_C_27 : begin
        fsm_output = 9'b001111100;
        state_var_NS = COMP_LOOP_C_28;
      end
      COMP_LOOP_C_28 : begin
        fsm_output = 9'b001111101;
        state_var_NS = COMP_LOOP_C_29;
      end
      COMP_LOOP_C_29 : begin
        fsm_output = 9'b001111110;
        state_var_NS = COMP_LOOP_C_30;
      end
      COMP_LOOP_C_30 : begin
        fsm_output = 9'b001111111;
        state_var_NS = COMP_LOOP_C_31;
      end
      COMP_LOOP_C_31 : begin
        fsm_output = 9'b010000000;
        state_var_NS = COMP_LOOP_C_32;
      end
      COMP_LOOP_C_32 : begin
        fsm_output = 9'b010000001;
        state_var_NS = COMP_LOOP_C_33;
      end
      COMP_LOOP_C_33 : begin
        fsm_output = 9'b010000010;
        state_var_NS = COMP_LOOP_C_34;
      end
      COMP_LOOP_C_34 : begin
        fsm_output = 9'b010000011;
        state_var_NS = COMP_LOOP_C_35;
      end
      COMP_LOOP_C_35 : begin
        fsm_output = 9'b010000100;
        state_var_NS = COMP_LOOP_C_36;
      end
      COMP_LOOP_C_36 : begin
        fsm_output = 9'b010000101;
        state_var_NS = COMP_LOOP_C_37;
      end
      COMP_LOOP_C_37 : begin
        fsm_output = 9'b010000110;
        state_var_NS = COMP_LOOP_C_38;
      end
      COMP_LOOP_C_38 : begin
        fsm_output = 9'b010000111;
        state_var_NS = COMP_LOOP_C_39;
      end
      COMP_LOOP_C_39 : begin
        fsm_output = 9'b010001000;
        state_var_NS = COMP_LOOP_C_40;
      end
      COMP_LOOP_C_40 : begin
        fsm_output = 9'b010001001;
        state_var_NS = COMP_LOOP_C_41;
      end
      COMP_LOOP_C_41 : begin
        fsm_output = 9'b010001010;
        state_var_NS = COMP_LOOP_C_42;
      end
      COMP_LOOP_C_42 : begin
        fsm_output = 9'b010001011;
        state_var_NS = COMP_LOOP_C_43;
      end
      COMP_LOOP_C_43 : begin
        fsm_output = 9'b010001100;
        state_var_NS = COMP_LOOP_C_44;
      end
      COMP_LOOP_C_44 : begin
        fsm_output = 9'b010001101;
        state_var_NS = COMP_LOOP_C_45;
      end
      COMP_LOOP_C_45 : begin
        fsm_output = 9'b010001110;
        state_var_NS = COMP_LOOP_C_46;
      end
      COMP_LOOP_C_46 : begin
        fsm_output = 9'b010001111;
        state_var_NS = COMP_LOOP_C_47;
      end
      COMP_LOOP_C_47 : begin
        fsm_output = 9'b010010000;
        state_var_NS = COMP_LOOP_C_48;
      end
      COMP_LOOP_C_48 : begin
        fsm_output = 9'b010010001;
        state_var_NS = COMP_LOOP_C_49;
      end
      COMP_LOOP_C_49 : begin
        fsm_output = 9'b010010010;
        state_var_NS = COMP_LOOP_C_50;
      end
      COMP_LOOP_C_50 : begin
        fsm_output = 9'b010010011;
        state_var_NS = COMP_LOOP_C_51;
      end
      COMP_LOOP_C_51 : begin
        fsm_output = 9'b010010100;
        state_var_NS = COMP_LOOP_C_52;
      end
      COMP_LOOP_C_52 : begin
        fsm_output = 9'b010010101;
        state_var_NS = COMP_LOOP_C_53;
      end
      COMP_LOOP_C_53 : begin
        fsm_output = 9'b010010110;
        state_var_NS = COMP_LOOP_C_54;
      end
      COMP_LOOP_C_54 : begin
        fsm_output = 9'b010010111;
        state_var_NS = COMP_LOOP_C_55;
      end
      COMP_LOOP_C_55 : begin
        fsm_output = 9'b010011000;
        state_var_NS = COMP_LOOP_C_56;
      end
      COMP_LOOP_C_56 : begin
        fsm_output = 9'b010011001;
        state_var_NS = COMP_LOOP_C_57;
      end
      COMP_LOOP_C_57 : begin
        fsm_output = 9'b010011010;
        state_var_NS = COMP_LOOP_C_58;
      end
      COMP_LOOP_C_58 : begin
        fsm_output = 9'b010011011;
        state_var_NS = COMP_LOOP_C_59;
      end
      COMP_LOOP_C_59 : begin
        fsm_output = 9'b010011100;
        state_var_NS = COMP_LOOP_C_60;
      end
      COMP_LOOP_C_60 : begin
        fsm_output = 9'b010011101;
        state_var_NS = COMP_LOOP_C_61;
      end
      COMP_LOOP_C_61 : begin
        fsm_output = 9'b010011110;
        state_var_NS = COMP_LOOP_C_62;
      end
      COMP_LOOP_C_62 : begin
        fsm_output = 9'b010011111;
        state_var_NS = COMP_LOOP_C_63;
      end
      COMP_LOOP_C_63 : begin
        fsm_output = 9'b010100000;
        state_var_NS = COMP_LOOP_C_64;
      end
      COMP_LOOP_C_64 : begin
        fsm_output = 9'b010100001;
        state_var_NS = COMP_LOOP_C_65;
      end
      COMP_LOOP_C_65 : begin
        fsm_output = 9'b010100010;
        state_var_NS = COMP_LOOP_C_66;
      end
      COMP_LOOP_C_66 : begin
        fsm_output = 9'b010100011;
        state_var_NS = COMP_LOOP_C_67;
      end
      COMP_LOOP_C_67 : begin
        fsm_output = 9'b010100100;
        state_var_NS = COMP_LOOP_C_68;
      end
      COMP_LOOP_C_68 : begin
        fsm_output = 9'b010100101;
        if ( COMP_LOOP_C_68_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_69;
        end
      end
      COMP_LOOP_C_69 : begin
        fsm_output = 9'b010100110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_0;
      end
      COMP_LOOP_2_modExp_1_while_C_0 : begin
        fsm_output = 9'b010100111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_1;
      end
      COMP_LOOP_2_modExp_1_while_C_1 : begin
        fsm_output = 9'b010101000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_2;
      end
      COMP_LOOP_2_modExp_1_while_C_2 : begin
        fsm_output = 9'b010101001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_3;
      end
      COMP_LOOP_2_modExp_1_while_C_3 : begin
        fsm_output = 9'b010101010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_4;
      end
      COMP_LOOP_2_modExp_1_while_C_4 : begin
        fsm_output = 9'b010101011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_5;
      end
      COMP_LOOP_2_modExp_1_while_C_5 : begin
        fsm_output = 9'b010101100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_6;
      end
      COMP_LOOP_2_modExp_1_while_C_6 : begin
        fsm_output = 9'b010101101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_7;
      end
      COMP_LOOP_2_modExp_1_while_C_7 : begin
        fsm_output = 9'b010101110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_8;
      end
      COMP_LOOP_2_modExp_1_while_C_8 : begin
        fsm_output = 9'b010101111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_9;
      end
      COMP_LOOP_2_modExp_1_while_C_9 : begin
        fsm_output = 9'b010110000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_10;
      end
      COMP_LOOP_2_modExp_1_while_C_10 : begin
        fsm_output = 9'b010110001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_11;
      end
      COMP_LOOP_2_modExp_1_while_C_11 : begin
        fsm_output = 9'b010110010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_12;
      end
      COMP_LOOP_2_modExp_1_while_C_12 : begin
        fsm_output = 9'b010110011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_13;
      end
      COMP_LOOP_2_modExp_1_while_C_13 : begin
        fsm_output = 9'b010110100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_14;
      end
      COMP_LOOP_2_modExp_1_while_C_14 : begin
        fsm_output = 9'b010110101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_15;
      end
      COMP_LOOP_2_modExp_1_while_C_15 : begin
        fsm_output = 9'b010110110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_16;
      end
      COMP_LOOP_2_modExp_1_while_C_16 : begin
        fsm_output = 9'b010110111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_17;
      end
      COMP_LOOP_2_modExp_1_while_C_17 : begin
        fsm_output = 9'b010111000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_18;
      end
      COMP_LOOP_2_modExp_1_while_C_18 : begin
        fsm_output = 9'b010111001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_19;
      end
      COMP_LOOP_2_modExp_1_while_C_19 : begin
        fsm_output = 9'b010111010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_20;
      end
      COMP_LOOP_2_modExp_1_while_C_20 : begin
        fsm_output = 9'b010111011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_21;
      end
      COMP_LOOP_2_modExp_1_while_C_21 : begin
        fsm_output = 9'b010111100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_22;
      end
      COMP_LOOP_2_modExp_1_while_C_22 : begin
        fsm_output = 9'b010111101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_23;
      end
      COMP_LOOP_2_modExp_1_while_C_23 : begin
        fsm_output = 9'b010111110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_24;
      end
      COMP_LOOP_2_modExp_1_while_C_24 : begin
        fsm_output = 9'b010111111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_25;
      end
      COMP_LOOP_2_modExp_1_while_C_25 : begin
        fsm_output = 9'b011000000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_26;
      end
      COMP_LOOP_2_modExp_1_while_C_26 : begin
        fsm_output = 9'b011000001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_27;
      end
      COMP_LOOP_2_modExp_1_while_C_27 : begin
        fsm_output = 9'b011000010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_28;
      end
      COMP_LOOP_2_modExp_1_while_C_28 : begin
        fsm_output = 9'b011000011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_29;
      end
      COMP_LOOP_2_modExp_1_while_C_29 : begin
        fsm_output = 9'b011000100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_30;
      end
      COMP_LOOP_2_modExp_1_while_C_30 : begin
        fsm_output = 9'b011000101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_31;
      end
      COMP_LOOP_2_modExp_1_while_C_31 : begin
        fsm_output = 9'b011000110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_32;
      end
      COMP_LOOP_2_modExp_1_while_C_32 : begin
        fsm_output = 9'b011000111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_33;
      end
      COMP_LOOP_2_modExp_1_while_C_33 : begin
        fsm_output = 9'b011001000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_34;
      end
      COMP_LOOP_2_modExp_1_while_C_34 : begin
        fsm_output = 9'b011001001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_35;
      end
      COMP_LOOP_2_modExp_1_while_C_35 : begin
        fsm_output = 9'b011001010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_36;
      end
      COMP_LOOP_2_modExp_1_while_C_36 : begin
        fsm_output = 9'b011001011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_37;
      end
      COMP_LOOP_2_modExp_1_while_C_37 : begin
        fsm_output = 9'b011001100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_38;
      end
      COMP_LOOP_2_modExp_1_while_C_38 : begin
        fsm_output = 9'b011001101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_39;
      end
      COMP_LOOP_2_modExp_1_while_C_39 : begin
        fsm_output = 9'b011001110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_40;
      end
      COMP_LOOP_2_modExp_1_while_C_40 : begin
        fsm_output = 9'b011001111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_41;
      end
      COMP_LOOP_2_modExp_1_while_C_41 : begin
        fsm_output = 9'b011010000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_42;
      end
      COMP_LOOP_2_modExp_1_while_C_42 : begin
        fsm_output = 9'b011010001;
        if ( COMP_LOOP_2_modExp_1_while_C_42_tr0 ) begin
          state_var_NS = COMP_LOOP_C_70;
        end
        else begin
          state_var_NS = COMP_LOOP_2_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_70 : begin
        fsm_output = 9'b011010010;
        state_var_NS = COMP_LOOP_C_71;
      end
      COMP_LOOP_C_71 : begin
        fsm_output = 9'b011010011;
        state_var_NS = COMP_LOOP_C_72;
      end
      COMP_LOOP_C_72 : begin
        fsm_output = 9'b011010100;
        state_var_NS = COMP_LOOP_C_73;
      end
      COMP_LOOP_C_73 : begin
        fsm_output = 9'b011010101;
        state_var_NS = COMP_LOOP_C_74;
      end
      COMP_LOOP_C_74 : begin
        fsm_output = 9'b011010110;
        state_var_NS = COMP_LOOP_C_75;
      end
      COMP_LOOP_C_75 : begin
        fsm_output = 9'b011010111;
        state_var_NS = COMP_LOOP_C_76;
      end
      COMP_LOOP_C_76 : begin
        fsm_output = 9'b011011000;
        state_var_NS = COMP_LOOP_C_77;
      end
      COMP_LOOP_C_77 : begin
        fsm_output = 9'b011011001;
        state_var_NS = COMP_LOOP_C_78;
      end
      COMP_LOOP_C_78 : begin
        fsm_output = 9'b011011010;
        state_var_NS = COMP_LOOP_C_79;
      end
      COMP_LOOP_C_79 : begin
        fsm_output = 9'b011011011;
        state_var_NS = COMP_LOOP_C_80;
      end
      COMP_LOOP_C_80 : begin
        fsm_output = 9'b011011100;
        state_var_NS = COMP_LOOP_C_81;
      end
      COMP_LOOP_C_81 : begin
        fsm_output = 9'b011011101;
        state_var_NS = COMP_LOOP_C_82;
      end
      COMP_LOOP_C_82 : begin
        fsm_output = 9'b011011110;
        state_var_NS = COMP_LOOP_C_83;
      end
      COMP_LOOP_C_83 : begin
        fsm_output = 9'b011011111;
        state_var_NS = COMP_LOOP_C_84;
      end
      COMP_LOOP_C_84 : begin
        fsm_output = 9'b011100000;
        state_var_NS = COMP_LOOP_C_85;
      end
      COMP_LOOP_C_85 : begin
        fsm_output = 9'b011100001;
        state_var_NS = COMP_LOOP_C_86;
      end
      COMP_LOOP_C_86 : begin
        fsm_output = 9'b011100010;
        state_var_NS = COMP_LOOP_C_87;
      end
      COMP_LOOP_C_87 : begin
        fsm_output = 9'b011100011;
        state_var_NS = COMP_LOOP_C_88;
      end
      COMP_LOOP_C_88 : begin
        fsm_output = 9'b011100100;
        state_var_NS = COMP_LOOP_C_89;
      end
      COMP_LOOP_C_89 : begin
        fsm_output = 9'b011100101;
        state_var_NS = COMP_LOOP_C_90;
      end
      COMP_LOOP_C_90 : begin
        fsm_output = 9'b011100110;
        state_var_NS = COMP_LOOP_C_91;
      end
      COMP_LOOP_C_91 : begin
        fsm_output = 9'b011100111;
        state_var_NS = COMP_LOOP_C_92;
      end
      COMP_LOOP_C_92 : begin
        fsm_output = 9'b011101000;
        state_var_NS = COMP_LOOP_C_93;
      end
      COMP_LOOP_C_93 : begin
        fsm_output = 9'b011101001;
        state_var_NS = COMP_LOOP_C_94;
      end
      COMP_LOOP_C_94 : begin
        fsm_output = 9'b011101010;
        state_var_NS = COMP_LOOP_C_95;
      end
      COMP_LOOP_C_95 : begin
        fsm_output = 9'b011101011;
        state_var_NS = COMP_LOOP_C_96;
      end
      COMP_LOOP_C_96 : begin
        fsm_output = 9'b011101100;
        state_var_NS = COMP_LOOP_C_97;
      end
      COMP_LOOP_C_97 : begin
        fsm_output = 9'b011101101;
        state_var_NS = COMP_LOOP_C_98;
      end
      COMP_LOOP_C_98 : begin
        fsm_output = 9'b011101110;
        state_var_NS = COMP_LOOP_C_99;
      end
      COMP_LOOP_C_99 : begin
        fsm_output = 9'b011101111;
        state_var_NS = COMP_LOOP_C_100;
      end
      COMP_LOOP_C_100 : begin
        fsm_output = 9'b011110000;
        state_var_NS = COMP_LOOP_C_101;
      end
      COMP_LOOP_C_101 : begin
        fsm_output = 9'b011110001;
        state_var_NS = COMP_LOOP_C_102;
      end
      COMP_LOOP_C_102 : begin
        fsm_output = 9'b011110010;
        state_var_NS = COMP_LOOP_C_103;
      end
      COMP_LOOP_C_103 : begin
        fsm_output = 9'b011110011;
        state_var_NS = COMP_LOOP_C_104;
      end
      COMP_LOOP_C_104 : begin
        fsm_output = 9'b011110100;
        state_var_NS = COMP_LOOP_C_105;
      end
      COMP_LOOP_C_105 : begin
        fsm_output = 9'b011110101;
        state_var_NS = COMP_LOOP_C_106;
      end
      COMP_LOOP_C_106 : begin
        fsm_output = 9'b011110110;
        state_var_NS = COMP_LOOP_C_107;
      end
      COMP_LOOP_C_107 : begin
        fsm_output = 9'b011110111;
        state_var_NS = COMP_LOOP_C_108;
      end
      COMP_LOOP_C_108 : begin
        fsm_output = 9'b011111000;
        state_var_NS = COMP_LOOP_C_109;
      end
      COMP_LOOP_C_109 : begin
        fsm_output = 9'b011111001;
        state_var_NS = COMP_LOOP_C_110;
      end
      COMP_LOOP_C_110 : begin
        fsm_output = 9'b011111010;
        state_var_NS = COMP_LOOP_C_111;
      end
      COMP_LOOP_C_111 : begin
        fsm_output = 9'b011111011;
        state_var_NS = COMP_LOOP_C_112;
      end
      COMP_LOOP_C_112 : begin
        fsm_output = 9'b011111100;
        state_var_NS = COMP_LOOP_C_113;
      end
      COMP_LOOP_C_113 : begin
        fsm_output = 9'b011111101;
        state_var_NS = COMP_LOOP_C_114;
      end
      COMP_LOOP_C_114 : begin
        fsm_output = 9'b011111110;
        state_var_NS = COMP_LOOP_C_115;
      end
      COMP_LOOP_C_115 : begin
        fsm_output = 9'b011111111;
        state_var_NS = COMP_LOOP_C_116;
      end
      COMP_LOOP_C_116 : begin
        fsm_output = 9'b100000000;
        state_var_NS = COMP_LOOP_C_117;
      end
      COMP_LOOP_C_117 : begin
        fsm_output = 9'b100000001;
        state_var_NS = COMP_LOOP_C_118;
      end
      COMP_LOOP_C_118 : begin
        fsm_output = 9'b100000010;
        state_var_NS = COMP_LOOP_C_119;
      end
      COMP_LOOP_C_119 : begin
        fsm_output = 9'b100000011;
        state_var_NS = COMP_LOOP_C_120;
      end
      COMP_LOOP_C_120 : begin
        fsm_output = 9'b100000100;
        state_var_NS = COMP_LOOP_C_121;
      end
      COMP_LOOP_C_121 : begin
        fsm_output = 9'b100000101;
        state_var_NS = COMP_LOOP_C_122;
      end
      COMP_LOOP_C_122 : begin
        fsm_output = 9'b100000110;
        state_var_NS = COMP_LOOP_C_123;
      end
      COMP_LOOP_C_123 : begin
        fsm_output = 9'b100000111;
        state_var_NS = COMP_LOOP_C_124;
      end
      COMP_LOOP_C_124 : begin
        fsm_output = 9'b100001000;
        state_var_NS = COMP_LOOP_C_125;
      end
      COMP_LOOP_C_125 : begin
        fsm_output = 9'b100001001;
        state_var_NS = COMP_LOOP_C_126;
      end
      COMP_LOOP_C_126 : begin
        fsm_output = 9'b100001010;
        state_var_NS = COMP_LOOP_C_127;
      end
      COMP_LOOP_C_127 : begin
        fsm_output = 9'b100001011;
        state_var_NS = COMP_LOOP_C_128;
      end
      COMP_LOOP_C_128 : begin
        fsm_output = 9'b100001100;
        state_var_NS = COMP_LOOP_C_129;
      end
      COMP_LOOP_C_129 : begin
        fsm_output = 9'b100001101;
        state_var_NS = COMP_LOOP_C_130;
      end
      COMP_LOOP_C_130 : begin
        fsm_output = 9'b100001110;
        state_var_NS = COMP_LOOP_C_131;
      end
      COMP_LOOP_C_131 : begin
        fsm_output = 9'b100001111;
        state_var_NS = COMP_LOOP_C_132;
      end
      COMP_LOOP_C_132 : begin
        fsm_output = 9'b100010000;
        state_var_NS = COMP_LOOP_C_133;
      end
      COMP_LOOP_C_133 : begin
        fsm_output = 9'b100010001;
        state_var_NS = COMP_LOOP_C_134;
      end
      COMP_LOOP_C_134 : begin
        fsm_output = 9'b100010010;
        state_var_NS = COMP_LOOP_C_135;
      end
      COMP_LOOP_C_135 : begin
        fsm_output = 9'b100010011;
        state_var_NS = COMP_LOOP_C_136;
      end
      COMP_LOOP_C_136 : begin
        fsm_output = 9'b100010100;
        if ( COMP_LOOP_C_136_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_137;
        end
      end
      COMP_LOOP_C_137 : begin
        fsm_output = 9'b100010101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_0;
      end
      COMP_LOOP_3_modExp_1_while_C_0 : begin
        fsm_output = 9'b100010110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_1;
      end
      COMP_LOOP_3_modExp_1_while_C_1 : begin
        fsm_output = 9'b100010111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_2;
      end
      COMP_LOOP_3_modExp_1_while_C_2 : begin
        fsm_output = 9'b100011000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_3;
      end
      COMP_LOOP_3_modExp_1_while_C_3 : begin
        fsm_output = 9'b100011001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_4;
      end
      COMP_LOOP_3_modExp_1_while_C_4 : begin
        fsm_output = 9'b100011010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_5;
      end
      COMP_LOOP_3_modExp_1_while_C_5 : begin
        fsm_output = 9'b100011011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_6;
      end
      COMP_LOOP_3_modExp_1_while_C_6 : begin
        fsm_output = 9'b100011100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_7;
      end
      COMP_LOOP_3_modExp_1_while_C_7 : begin
        fsm_output = 9'b100011101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_8;
      end
      COMP_LOOP_3_modExp_1_while_C_8 : begin
        fsm_output = 9'b100011110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_9;
      end
      COMP_LOOP_3_modExp_1_while_C_9 : begin
        fsm_output = 9'b100011111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_10;
      end
      COMP_LOOP_3_modExp_1_while_C_10 : begin
        fsm_output = 9'b100100000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_11;
      end
      COMP_LOOP_3_modExp_1_while_C_11 : begin
        fsm_output = 9'b100100001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_12;
      end
      COMP_LOOP_3_modExp_1_while_C_12 : begin
        fsm_output = 9'b100100010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_13;
      end
      COMP_LOOP_3_modExp_1_while_C_13 : begin
        fsm_output = 9'b100100011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_14;
      end
      COMP_LOOP_3_modExp_1_while_C_14 : begin
        fsm_output = 9'b100100100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_15;
      end
      COMP_LOOP_3_modExp_1_while_C_15 : begin
        fsm_output = 9'b100100101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_16;
      end
      COMP_LOOP_3_modExp_1_while_C_16 : begin
        fsm_output = 9'b100100110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_17;
      end
      COMP_LOOP_3_modExp_1_while_C_17 : begin
        fsm_output = 9'b100100111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_18;
      end
      COMP_LOOP_3_modExp_1_while_C_18 : begin
        fsm_output = 9'b100101000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_19;
      end
      COMP_LOOP_3_modExp_1_while_C_19 : begin
        fsm_output = 9'b100101001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_20;
      end
      COMP_LOOP_3_modExp_1_while_C_20 : begin
        fsm_output = 9'b100101010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_21;
      end
      COMP_LOOP_3_modExp_1_while_C_21 : begin
        fsm_output = 9'b100101011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_22;
      end
      COMP_LOOP_3_modExp_1_while_C_22 : begin
        fsm_output = 9'b100101100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_23;
      end
      COMP_LOOP_3_modExp_1_while_C_23 : begin
        fsm_output = 9'b100101101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_24;
      end
      COMP_LOOP_3_modExp_1_while_C_24 : begin
        fsm_output = 9'b100101110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_25;
      end
      COMP_LOOP_3_modExp_1_while_C_25 : begin
        fsm_output = 9'b100101111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_26;
      end
      COMP_LOOP_3_modExp_1_while_C_26 : begin
        fsm_output = 9'b100110000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_27;
      end
      COMP_LOOP_3_modExp_1_while_C_27 : begin
        fsm_output = 9'b100110001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_28;
      end
      COMP_LOOP_3_modExp_1_while_C_28 : begin
        fsm_output = 9'b100110010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_29;
      end
      COMP_LOOP_3_modExp_1_while_C_29 : begin
        fsm_output = 9'b100110011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_30;
      end
      COMP_LOOP_3_modExp_1_while_C_30 : begin
        fsm_output = 9'b100110100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_31;
      end
      COMP_LOOP_3_modExp_1_while_C_31 : begin
        fsm_output = 9'b100110101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_32;
      end
      COMP_LOOP_3_modExp_1_while_C_32 : begin
        fsm_output = 9'b100110110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_33;
      end
      COMP_LOOP_3_modExp_1_while_C_33 : begin
        fsm_output = 9'b100110111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_34;
      end
      COMP_LOOP_3_modExp_1_while_C_34 : begin
        fsm_output = 9'b100111000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_35;
      end
      COMP_LOOP_3_modExp_1_while_C_35 : begin
        fsm_output = 9'b100111001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_36;
      end
      COMP_LOOP_3_modExp_1_while_C_36 : begin
        fsm_output = 9'b100111010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_37;
      end
      COMP_LOOP_3_modExp_1_while_C_37 : begin
        fsm_output = 9'b100111011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_38;
      end
      COMP_LOOP_3_modExp_1_while_C_38 : begin
        fsm_output = 9'b100111100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_39;
      end
      COMP_LOOP_3_modExp_1_while_C_39 : begin
        fsm_output = 9'b100111101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_40;
      end
      COMP_LOOP_3_modExp_1_while_C_40 : begin
        fsm_output = 9'b100111110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_41;
      end
      COMP_LOOP_3_modExp_1_while_C_41 : begin
        fsm_output = 9'b100111111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_42;
      end
      COMP_LOOP_3_modExp_1_while_C_42 : begin
        fsm_output = 9'b101000000;
        if ( COMP_LOOP_3_modExp_1_while_C_42_tr0 ) begin
          state_var_NS = COMP_LOOP_C_138;
        end
        else begin
          state_var_NS = COMP_LOOP_3_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_138 : begin
        fsm_output = 9'b101000001;
        state_var_NS = COMP_LOOP_C_139;
      end
      COMP_LOOP_C_139 : begin
        fsm_output = 9'b101000010;
        state_var_NS = COMP_LOOP_C_140;
      end
      COMP_LOOP_C_140 : begin
        fsm_output = 9'b101000011;
        state_var_NS = COMP_LOOP_C_141;
      end
      COMP_LOOP_C_141 : begin
        fsm_output = 9'b101000100;
        state_var_NS = COMP_LOOP_C_142;
      end
      COMP_LOOP_C_142 : begin
        fsm_output = 9'b101000101;
        state_var_NS = COMP_LOOP_C_143;
      end
      COMP_LOOP_C_143 : begin
        fsm_output = 9'b101000110;
        state_var_NS = COMP_LOOP_C_144;
      end
      COMP_LOOP_C_144 : begin
        fsm_output = 9'b101000111;
        state_var_NS = COMP_LOOP_C_145;
      end
      COMP_LOOP_C_145 : begin
        fsm_output = 9'b101001000;
        state_var_NS = COMP_LOOP_C_146;
      end
      COMP_LOOP_C_146 : begin
        fsm_output = 9'b101001001;
        state_var_NS = COMP_LOOP_C_147;
      end
      COMP_LOOP_C_147 : begin
        fsm_output = 9'b101001010;
        state_var_NS = COMP_LOOP_C_148;
      end
      COMP_LOOP_C_148 : begin
        fsm_output = 9'b101001011;
        state_var_NS = COMP_LOOP_C_149;
      end
      COMP_LOOP_C_149 : begin
        fsm_output = 9'b101001100;
        state_var_NS = COMP_LOOP_C_150;
      end
      COMP_LOOP_C_150 : begin
        fsm_output = 9'b101001101;
        state_var_NS = COMP_LOOP_C_151;
      end
      COMP_LOOP_C_151 : begin
        fsm_output = 9'b101001110;
        state_var_NS = COMP_LOOP_C_152;
      end
      COMP_LOOP_C_152 : begin
        fsm_output = 9'b101001111;
        state_var_NS = COMP_LOOP_C_153;
      end
      COMP_LOOP_C_153 : begin
        fsm_output = 9'b101010000;
        state_var_NS = COMP_LOOP_C_154;
      end
      COMP_LOOP_C_154 : begin
        fsm_output = 9'b101010001;
        state_var_NS = COMP_LOOP_C_155;
      end
      COMP_LOOP_C_155 : begin
        fsm_output = 9'b101010010;
        state_var_NS = COMP_LOOP_C_156;
      end
      COMP_LOOP_C_156 : begin
        fsm_output = 9'b101010011;
        state_var_NS = COMP_LOOP_C_157;
      end
      COMP_LOOP_C_157 : begin
        fsm_output = 9'b101010100;
        state_var_NS = COMP_LOOP_C_158;
      end
      COMP_LOOP_C_158 : begin
        fsm_output = 9'b101010101;
        state_var_NS = COMP_LOOP_C_159;
      end
      COMP_LOOP_C_159 : begin
        fsm_output = 9'b101010110;
        state_var_NS = COMP_LOOP_C_160;
      end
      COMP_LOOP_C_160 : begin
        fsm_output = 9'b101010111;
        state_var_NS = COMP_LOOP_C_161;
      end
      COMP_LOOP_C_161 : begin
        fsm_output = 9'b101011000;
        state_var_NS = COMP_LOOP_C_162;
      end
      COMP_LOOP_C_162 : begin
        fsm_output = 9'b101011001;
        state_var_NS = COMP_LOOP_C_163;
      end
      COMP_LOOP_C_163 : begin
        fsm_output = 9'b101011010;
        state_var_NS = COMP_LOOP_C_164;
      end
      COMP_LOOP_C_164 : begin
        fsm_output = 9'b101011011;
        state_var_NS = COMP_LOOP_C_165;
      end
      COMP_LOOP_C_165 : begin
        fsm_output = 9'b101011100;
        state_var_NS = COMP_LOOP_C_166;
      end
      COMP_LOOP_C_166 : begin
        fsm_output = 9'b101011101;
        state_var_NS = COMP_LOOP_C_167;
      end
      COMP_LOOP_C_167 : begin
        fsm_output = 9'b101011110;
        state_var_NS = COMP_LOOP_C_168;
      end
      COMP_LOOP_C_168 : begin
        fsm_output = 9'b101011111;
        state_var_NS = COMP_LOOP_C_169;
      end
      COMP_LOOP_C_169 : begin
        fsm_output = 9'b101100000;
        state_var_NS = COMP_LOOP_C_170;
      end
      COMP_LOOP_C_170 : begin
        fsm_output = 9'b101100001;
        state_var_NS = COMP_LOOP_C_171;
      end
      COMP_LOOP_C_171 : begin
        fsm_output = 9'b101100010;
        state_var_NS = COMP_LOOP_C_172;
      end
      COMP_LOOP_C_172 : begin
        fsm_output = 9'b101100011;
        state_var_NS = COMP_LOOP_C_173;
      end
      COMP_LOOP_C_173 : begin
        fsm_output = 9'b101100100;
        state_var_NS = COMP_LOOP_C_174;
      end
      COMP_LOOP_C_174 : begin
        fsm_output = 9'b101100101;
        state_var_NS = COMP_LOOP_C_175;
      end
      COMP_LOOP_C_175 : begin
        fsm_output = 9'b101100110;
        state_var_NS = COMP_LOOP_C_176;
      end
      COMP_LOOP_C_176 : begin
        fsm_output = 9'b101100111;
        state_var_NS = COMP_LOOP_C_177;
      end
      COMP_LOOP_C_177 : begin
        fsm_output = 9'b101101000;
        state_var_NS = COMP_LOOP_C_178;
      end
      COMP_LOOP_C_178 : begin
        fsm_output = 9'b101101001;
        state_var_NS = COMP_LOOP_C_179;
      end
      COMP_LOOP_C_179 : begin
        fsm_output = 9'b101101010;
        state_var_NS = COMP_LOOP_C_180;
      end
      COMP_LOOP_C_180 : begin
        fsm_output = 9'b101101011;
        state_var_NS = COMP_LOOP_C_181;
      end
      COMP_LOOP_C_181 : begin
        fsm_output = 9'b101101100;
        state_var_NS = COMP_LOOP_C_182;
      end
      COMP_LOOP_C_182 : begin
        fsm_output = 9'b101101101;
        state_var_NS = COMP_LOOP_C_183;
      end
      COMP_LOOP_C_183 : begin
        fsm_output = 9'b101101110;
        state_var_NS = COMP_LOOP_C_184;
      end
      COMP_LOOP_C_184 : begin
        fsm_output = 9'b101101111;
        state_var_NS = COMP_LOOP_C_185;
      end
      COMP_LOOP_C_185 : begin
        fsm_output = 9'b101110000;
        state_var_NS = COMP_LOOP_C_186;
      end
      COMP_LOOP_C_186 : begin
        fsm_output = 9'b101110001;
        state_var_NS = COMP_LOOP_C_187;
      end
      COMP_LOOP_C_187 : begin
        fsm_output = 9'b101110010;
        state_var_NS = COMP_LOOP_C_188;
      end
      COMP_LOOP_C_188 : begin
        fsm_output = 9'b101110011;
        state_var_NS = COMP_LOOP_C_189;
      end
      COMP_LOOP_C_189 : begin
        fsm_output = 9'b101110100;
        state_var_NS = COMP_LOOP_C_190;
      end
      COMP_LOOP_C_190 : begin
        fsm_output = 9'b101110101;
        state_var_NS = COMP_LOOP_C_191;
      end
      COMP_LOOP_C_191 : begin
        fsm_output = 9'b101110110;
        state_var_NS = COMP_LOOP_C_192;
      end
      COMP_LOOP_C_192 : begin
        fsm_output = 9'b101110111;
        state_var_NS = COMP_LOOP_C_193;
      end
      COMP_LOOP_C_193 : begin
        fsm_output = 9'b101111000;
        state_var_NS = COMP_LOOP_C_194;
      end
      COMP_LOOP_C_194 : begin
        fsm_output = 9'b101111001;
        state_var_NS = COMP_LOOP_C_195;
      end
      COMP_LOOP_C_195 : begin
        fsm_output = 9'b101111010;
        state_var_NS = COMP_LOOP_C_196;
      end
      COMP_LOOP_C_196 : begin
        fsm_output = 9'b101111011;
        state_var_NS = COMP_LOOP_C_197;
      end
      COMP_LOOP_C_197 : begin
        fsm_output = 9'b101111100;
        state_var_NS = COMP_LOOP_C_198;
      end
      COMP_LOOP_C_198 : begin
        fsm_output = 9'b101111101;
        state_var_NS = COMP_LOOP_C_199;
      end
      COMP_LOOP_C_199 : begin
        fsm_output = 9'b101111110;
        state_var_NS = COMP_LOOP_C_200;
      end
      COMP_LOOP_C_200 : begin
        fsm_output = 9'b101111111;
        state_var_NS = COMP_LOOP_C_201;
      end
      COMP_LOOP_C_201 : begin
        fsm_output = 9'b110000000;
        state_var_NS = COMP_LOOP_C_202;
      end
      COMP_LOOP_C_202 : begin
        fsm_output = 9'b110000001;
        state_var_NS = COMP_LOOP_C_203;
      end
      COMP_LOOP_C_203 : begin
        fsm_output = 9'b110000010;
        state_var_NS = COMP_LOOP_C_204;
      end
      COMP_LOOP_C_204 : begin
        fsm_output = 9'b110000011;
        if ( COMP_LOOP_C_204_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_205;
        end
      end
      COMP_LOOP_C_205 : begin
        fsm_output = 9'b110000100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_0;
      end
      COMP_LOOP_4_modExp_1_while_C_0 : begin
        fsm_output = 9'b110000101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_1;
      end
      COMP_LOOP_4_modExp_1_while_C_1 : begin
        fsm_output = 9'b110000110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_2;
      end
      COMP_LOOP_4_modExp_1_while_C_2 : begin
        fsm_output = 9'b110000111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_3;
      end
      COMP_LOOP_4_modExp_1_while_C_3 : begin
        fsm_output = 9'b110001000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_4;
      end
      COMP_LOOP_4_modExp_1_while_C_4 : begin
        fsm_output = 9'b110001001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_5;
      end
      COMP_LOOP_4_modExp_1_while_C_5 : begin
        fsm_output = 9'b110001010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_6;
      end
      COMP_LOOP_4_modExp_1_while_C_6 : begin
        fsm_output = 9'b110001011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_7;
      end
      COMP_LOOP_4_modExp_1_while_C_7 : begin
        fsm_output = 9'b110001100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_8;
      end
      COMP_LOOP_4_modExp_1_while_C_8 : begin
        fsm_output = 9'b110001101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_9;
      end
      COMP_LOOP_4_modExp_1_while_C_9 : begin
        fsm_output = 9'b110001110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_10;
      end
      COMP_LOOP_4_modExp_1_while_C_10 : begin
        fsm_output = 9'b110001111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_11;
      end
      COMP_LOOP_4_modExp_1_while_C_11 : begin
        fsm_output = 9'b110010000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_12;
      end
      COMP_LOOP_4_modExp_1_while_C_12 : begin
        fsm_output = 9'b110010001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_13;
      end
      COMP_LOOP_4_modExp_1_while_C_13 : begin
        fsm_output = 9'b110010010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_14;
      end
      COMP_LOOP_4_modExp_1_while_C_14 : begin
        fsm_output = 9'b110010011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_15;
      end
      COMP_LOOP_4_modExp_1_while_C_15 : begin
        fsm_output = 9'b110010100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_16;
      end
      COMP_LOOP_4_modExp_1_while_C_16 : begin
        fsm_output = 9'b110010101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_17;
      end
      COMP_LOOP_4_modExp_1_while_C_17 : begin
        fsm_output = 9'b110010110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_18;
      end
      COMP_LOOP_4_modExp_1_while_C_18 : begin
        fsm_output = 9'b110010111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_19;
      end
      COMP_LOOP_4_modExp_1_while_C_19 : begin
        fsm_output = 9'b110011000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_20;
      end
      COMP_LOOP_4_modExp_1_while_C_20 : begin
        fsm_output = 9'b110011001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_21;
      end
      COMP_LOOP_4_modExp_1_while_C_21 : begin
        fsm_output = 9'b110011010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_22;
      end
      COMP_LOOP_4_modExp_1_while_C_22 : begin
        fsm_output = 9'b110011011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_23;
      end
      COMP_LOOP_4_modExp_1_while_C_23 : begin
        fsm_output = 9'b110011100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_24;
      end
      COMP_LOOP_4_modExp_1_while_C_24 : begin
        fsm_output = 9'b110011101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_25;
      end
      COMP_LOOP_4_modExp_1_while_C_25 : begin
        fsm_output = 9'b110011110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_26;
      end
      COMP_LOOP_4_modExp_1_while_C_26 : begin
        fsm_output = 9'b110011111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_27;
      end
      COMP_LOOP_4_modExp_1_while_C_27 : begin
        fsm_output = 9'b110100000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_28;
      end
      COMP_LOOP_4_modExp_1_while_C_28 : begin
        fsm_output = 9'b110100001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_29;
      end
      COMP_LOOP_4_modExp_1_while_C_29 : begin
        fsm_output = 9'b110100010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_30;
      end
      COMP_LOOP_4_modExp_1_while_C_30 : begin
        fsm_output = 9'b110100011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_31;
      end
      COMP_LOOP_4_modExp_1_while_C_31 : begin
        fsm_output = 9'b110100100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_32;
      end
      COMP_LOOP_4_modExp_1_while_C_32 : begin
        fsm_output = 9'b110100101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_33;
      end
      COMP_LOOP_4_modExp_1_while_C_33 : begin
        fsm_output = 9'b110100110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_34;
      end
      COMP_LOOP_4_modExp_1_while_C_34 : begin
        fsm_output = 9'b110100111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_35;
      end
      COMP_LOOP_4_modExp_1_while_C_35 : begin
        fsm_output = 9'b110101000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_36;
      end
      COMP_LOOP_4_modExp_1_while_C_36 : begin
        fsm_output = 9'b110101001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_37;
      end
      COMP_LOOP_4_modExp_1_while_C_37 : begin
        fsm_output = 9'b110101010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_38;
      end
      COMP_LOOP_4_modExp_1_while_C_38 : begin
        fsm_output = 9'b110101011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_39;
      end
      COMP_LOOP_4_modExp_1_while_C_39 : begin
        fsm_output = 9'b110101100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_40;
      end
      COMP_LOOP_4_modExp_1_while_C_40 : begin
        fsm_output = 9'b110101101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_41;
      end
      COMP_LOOP_4_modExp_1_while_C_41 : begin
        fsm_output = 9'b110101110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_42;
      end
      COMP_LOOP_4_modExp_1_while_C_42 : begin
        fsm_output = 9'b110101111;
        if ( COMP_LOOP_4_modExp_1_while_C_42_tr0 ) begin
          state_var_NS = COMP_LOOP_C_206;
        end
        else begin
          state_var_NS = COMP_LOOP_4_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_206 : begin
        fsm_output = 9'b110110000;
        state_var_NS = COMP_LOOP_C_207;
      end
      COMP_LOOP_C_207 : begin
        fsm_output = 9'b110110001;
        state_var_NS = COMP_LOOP_C_208;
      end
      COMP_LOOP_C_208 : begin
        fsm_output = 9'b110110010;
        state_var_NS = COMP_LOOP_C_209;
      end
      COMP_LOOP_C_209 : begin
        fsm_output = 9'b110110011;
        state_var_NS = COMP_LOOP_C_210;
      end
      COMP_LOOP_C_210 : begin
        fsm_output = 9'b110110100;
        state_var_NS = COMP_LOOP_C_211;
      end
      COMP_LOOP_C_211 : begin
        fsm_output = 9'b110110101;
        state_var_NS = COMP_LOOP_C_212;
      end
      COMP_LOOP_C_212 : begin
        fsm_output = 9'b110110110;
        state_var_NS = COMP_LOOP_C_213;
      end
      COMP_LOOP_C_213 : begin
        fsm_output = 9'b110110111;
        state_var_NS = COMP_LOOP_C_214;
      end
      COMP_LOOP_C_214 : begin
        fsm_output = 9'b110111000;
        state_var_NS = COMP_LOOP_C_215;
      end
      COMP_LOOP_C_215 : begin
        fsm_output = 9'b110111001;
        state_var_NS = COMP_LOOP_C_216;
      end
      COMP_LOOP_C_216 : begin
        fsm_output = 9'b110111010;
        state_var_NS = COMP_LOOP_C_217;
      end
      COMP_LOOP_C_217 : begin
        fsm_output = 9'b110111011;
        state_var_NS = COMP_LOOP_C_218;
      end
      COMP_LOOP_C_218 : begin
        fsm_output = 9'b110111100;
        state_var_NS = COMP_LOOP_C_219;
      end
      COMP_LOOP_C_219 : begin
        fsm_output = 9'b110111101;
        state_var_NS = COMP_LOOP_C_220;
      end
      COMP_LOOP_C_220 : begin
        fsm_output = 9'b110111110;
        state_var_NS = COMP_LOOP_C_221;
      end
      COMP_LOOP_C_221 : begin
        fsm_output = 9'b110111111;
        state_var_NS = COMP_LOOP_C_222;
      end
      COMP_LOOP_C_222 : begin
        fsm_output = 9'b111000000;
        state_var_NS = COMP_LOOP_C_223;
      end
      COMP_LOOP_C_223 : begin
        fsm_output = 9'b111000001;
        state_var_NS = COMP_LOOP_C_224;
      end
      COMP_LOOP_C_224 : begin
        fsm_output = 9'b111000010;
        state_var_NS = COMP_LOOP_C_225;
      end
      COMP_LOOP_C_225 : begin
        fsm_output = 9'b111000011;
        state_var_NS = COMP_LOOP_C_226;
      end
      COMP_LOOP_C_226 : begin
        fsm_output = 9'b111000100;
        state_var_NS = COMP_LOOP_C_227;
      end
      COMP_LOOP_C_227 : begin
        fsm_output = 9'b111000101;
        state_var_NS = COMP_LOOP_C_228;
      end
      COMP_LOOP_C_228 : begin
        fsm_output = 9'b111000110;
        state_var_NS = COMP_LOOP_C_229;
      end
      COMP_LOOP_C_229 : begin
        fsm_output = 9'b111000111;
        state_var_NS = COMP_LOOP_C_230;
      end
      COMP_LOOP_C_230 : begin
        fsm_output = 9'b111001000;
        state_var_NS = COMP_LOOP_C_231;
      end
      COMP_LOOP_C_231 : begin
        fsm_output = 9'b111001001;
        state_var_NS = COMP_LOOP_C_232;
      end
      COMP_LOOP_C_232 : begin
        fsm_output = 9'b111001010;
        state_var_NS = COMP_LOOP_C_233;
      end
      COMP_LOOP_C_233 : begin
        fsm_output = 9'b111001011;
        state_var_NS = COMP_LOOP_C_234;
      end
      COMP_LOOP_C_234 : begin
        fsm_output = 9'b111001100;
        state_var_NS = COMP_LOOP_C_235;
      end
      COMP_LOOP_C_235 : begin
        fsm_output = 9'b111001101;
        state_var_NS = COMP_LOOP_C_236;
      end
      COMP_LOOP_C_236 : begin
        fsm_output = 9'b111001110;
        state_var_NS = COMP_LOOP_C_237;
      end
      COMP_LOOP_C_237 : begin
        fsm_output = 9'b111001111;
        state_var_NS = COMP_LOOP_C_238;
      end
      COMP_LOOP_C_238 : begin
        fsm_output = 9'b111010000;
        state_var_NS = COMP_LOOP_C_239;
      end
      COMP_LOOP_C_239 : begin
        fsm_output = 9'b111010001;
        state_var_NS = COMP_LOOP_C_240;
      end
      COMP_LOOP_C_240 : begin
        fsm_output = 9'b111010010;
        state_var_NS = COMP_LOOP_C_241;
      end
      COMP_LOOP_C_241 : begin
        fsm_output = 9'b111010011;
        state_var_NS = COMP_LOOP_C_242;
      end
      COMP_LOOP_C_242 : begin
        fsm_output = 9'b111010100;
        state_var_NS = COMP_LOOP_C_243;
      end
      COMP_LOOP_C_243 : begin
        fsm_output = 9'b111010101;
        state_var_NS = COMP_LOOP_C_244;
      end
      COMP_LOOP_C_244 : begin
        fsm_output = 9'b111010110;
        state_var_NS = COMP_LOOP_C_245;
      end
      COMP_LOOP_C_245 : begin
        fsm_output = 9'b111010111;
        state_var_NS = COMP_LOOP_C_246;
      end
      COMP_LOOP_C_246 : begin
        fsm_output = 9'b111011000;
        state_var_NS = COMP_LOOP_C_247;
      end
      COMP_LOOP_C_247 : begin
        fsm_output = 9'b111011001;
        state_var_NS = COMP_LOOP_C_248;
      end
      COMP_LOOP_C_248 : begin
        fsm_output = 9'b111011010;
        state_var_NS = COMP_LOOP_C_249;
      end
      COMP_LOOP_C_249 : begin
        fsm_output = 9'b111011011;
        state_var_NS = COMP_LOOP_C_250;
      end
      COMP_LOOP_C_250 : begin
        fsm_output = 9'b111011100;
        state_var_NS = COMP_LOOP_C_251;
      end
      COMP_LOOP_C_251 : begin
        fsm_output = 9'b111011101;
        state_var_NS = COMP_LOOP_C_252;
      end
      COMP_LOOP_C_252 : begin
        fsm_output = 9'b111011110;
        state_var_NS = COMP_LOOP_C_253;
      end
      COMP_LOOP_C_253 : begin
        fsm_output = 9'b111011111;
        state_var_NS = COMP_LOOP_C_254;
      end
      COMP_LOOP_C_254 : begin
        fsm_output = 9'b111100000;
        state_var_NS = COMP_LOOP_C_255;
      end
      COMP_LOOP_C_255 : begin
        fsm_output = 9'b111100001;
        state_var_NS = COMP_LOOP_C_256;
      end
      COMP_LOOP_C_256 : begin
        fsm_output = 9'b111100010;
        state_var_NS = COMP_LOOP_C_257;
      end
      COMP_LOOP_C_257 : begin
        fsm_output = 9'b111100011;
        state_var_NS = COMP_LOOP_C_258;
      end
      COMP_LOOP_C_258 : begin
        fsm_output = 9'b111100100;
        state_var_NS = COMP_LOOP_C_259;
      end
      COMP_LOOP_C_259 : begin
        fsm_output = 9'b111100101;
        state_var_NS = COMP_LOOP_C_260;
      end
      COMP_LOOP_C_260 : begin
        fsm_output = 9'b111100110;
        state_var_NS = COMP_LOOP_C_261;
      end
      COMP_LOOP_C_261 : begin
        fsm_output = 9'b111100111;
        state_var_NS = COMP_LOOP_C_262;
      end
      COMP_LOOP_C_262 : begin
        fsm_output = 9'b111101000;
        state_var_NS = COMP_LOOP_C_263;
      end
      COMP_LOOP_C_263 : begin
        fsm_output = 9'b111101001;
        state_var_NS = COMP_LOOP_C_264;
      end
      COMP_LOOP_C_264 : begin
        fsm_output = 9'b111101010;
        state_var_NS = COMP_LOOP_C_265;
      end
      COMP_LOOP_C_265 : begin
        fsm_output = 9'b111101011;
        state_var_NS = COMP_LOOP_C_266;
      end
      COMP_LOOP_C_266 : begin
        fsm_output = 9'b111101100;
        state_var_NS = COMP_LOOP_C_267;
      end
      COMP_LOOP_C_267 : begin
        fsm_output = 9'b111101101;
        state_var_NS = COMP_LOOP_C_268;
      end
      COMP_LOOP_C_268 : begin
        fsm_output = 9'b111101110;
        state_var_NS = COMP_LOOP_C_269;
      end
      COMP_LOOP_C_269 : begin
        fsm_output = 9'b111101111;
        state_var_NS = COMP_LOOP_C_270;
      end
      COMP_LOOP_C_270 : begin
        fsm_output = 9'b111110000;
        state_var_NS = COMP_LOOP_C_271;
      end
      COMP_LOOP_C_271 : begin
        fsm_output = 9'b111110001;
        state_var_NS = COMP_LOOP_C_272;
      end
      COMP_LOOP_C_272 : begin
        fsm_output = 9'b111110010;
        if ( COMP_LOOP_C_272_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_C_0 : begin
        fsm_output = 9'b111110011;
        if ( VEC_LOOP_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_10;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      STAGE_LOOP_C_10 : begin
        fsm_output = 9'b111110100;
        if ( STAGE_LOOP_C_10_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = STAGE_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 9'b111110101;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 9'b000000000;
        state_var_NS = STAGE_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core (
  clk, rst, vec_rsc_triosy_0_0_lz, vec_rsc_triosy_0_1_lz, vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz, p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz,
      vec_rsc_0_0_i_qa_d, vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_1_i_qa_d,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_qa_d, vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_0_i_adra_d_pff,
      vec_rsc_0_0_i_da_d_pff, vec_rsc_0_0_i_wea_d_pff, vec_rsc_0_1_i_wea_d_pff, vec_rsc_0_2_i_wea_d_pff,
      vec_rsc_0_3_i_wea_d_pff
);
  input clk;
  input rst;
  output vec_rsc_triosy_0_0_lz;
  output vec_rsc_triosy_0_1_lz;
  output vec_rsc_triosy_0_2_lz;
  output vec_rsc_triosy_0_3_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  input [63:0] vec_rsc_0_0_i_qa_d;
  output vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_1_i_qa_d;
  output vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_2_i_qa_d;
  output vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_3_i_qa_d;
  output vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [9:0] vec_rsc_0_0_i_adra_d_pff;
  output [63:0] vec_rsc_0_0_i_da_d_pff;
  output vec_rsc_0_0_i_wea_d_pff;
  output vec_rsc_0_1_i_wea_d_pff;
  output vec_rsc_0_2_i_wea_d_pff;
  output vec_rsc_0_3_i_wea_d_pff;


  // Interconnect Declarations
  wire [63:0] p_rsci_idat;
  wire [63:0] r_rsci_idat;
  reg [63:0] modulo_result_rem_cmp_a;
  reg [63:0] modulo_result_rem_cmp_b;
  wire [63:0] modulo_result_rem_cmp_z;
  reg [64:0] operator_66_true_div_cmp_a;
  wire [64:0] operator_66_true_div_cmp_z;
  reg [9:0] operator_66_true_div_cmp_b_9_0;
  wire [8:0] fsm_output;
  wire and_dcpl_1;
  wire nor_tmp_16;
  wire mux_tmp_41;
  wire nor_tmp_24;
  wire or_tmp_70;
  wire mux_tmp_86;
  wire nor_tmp_63;
  wire and_dcpl_25;
  wire and_dcpl_26;
  wire and_dcpl_27;
  wire and_dcpl_28;
  wire and_dcpl_29;
  wire and_dcpl_30;
  wire and_dcpl_31;
  wire and_dcpl_33;
  wire and_dcpl_34;
  wire and_dcpl_36;
  wire and_dcpl_38;
  wire and_dcpl_39;
  wire and_dcpl_42;
  wire and_dcpl_43;
  wire and_dcpl_44;
  wire and_dcpl_45;
  wire and_dcpl_46;
  wire and_dcpl_47;
  wire and_dcpl_48;
  wire and_dcpl_49;
  wire and_dcpl_50;
  wire and_dcpl_53;
  wire and_dcpl_54;
  wire and_dcpl_62;
  wire and_dcpl_65;
  wire and_dcpl_67;
  wire and_dcpl_72;
  wire and_dcpl_75;
  wire and_dcpl_85;
  wire and_dcpl_86;
  wire and_dcpl_88;
  wire and_dcpl_89;
  wire and_dcpl_91;
  wire not_tmp_154;
  wire or_tmp_254;
  wire or_tmp_256;
  wire mux_tmp_212;
  wire not_tmp_158;
  wire or_tmp_262;
  wire and_dcpl_102;
  wire mux_tmp_230;
  wire or_tmp_275;
  wire or_tmp_277;
  wire mux_tmp_239;
  wire or_tmp_288;
  wire and_dcpl_105;
  wire and_dcpl_111;
  wire and_dcpl_122;
  wire and_dcpl_128;
  wire and_dcpl_132;
  wire or_tmp_300;
  wire mux_tmp_272;
  wire mux_tmp_273;
  wire mux_tmp_274;
  wire mux_tmp_276;
  wire mux_tmp_278;
  wire mux_tmp_282;
  wire mux_tmp_283;
  wire nor_tmp_120;
  wire mux_tmp_303;
  wire mux_tmp_321;
  wire and_dcpl_137;
  wire and_dcpl_138;
  wire and_dcpl_139;
  wire mux_tmp_329;
  wire mux_tmp_330;
  wire and_tmp_8;
  wire and_tmp_9;
  wire mux_tmp_333;
  wire mux_tmp_336;
  wire mux_tmp_337;
  wire mux_tmp_339;
  wire not_tmp_221;
  wire mux_tmp_344;
  wire mux_tmp_352;
  wire or_tmp_331;
  wire mux_tmp_354;
  wire and_dcpl_140;
  wire not_tmp_235;
  wire and_dcpl_141;
  wire not_tmp_239;
  wire not_tmp_242;
  wire mux_tmp_392;
  wire mux_tmp_397;
  wire not_tmp_246;
  wire mux_tmp_404;
  wire mux_tmp_408;
  wire mux_tmp_409;
  wire mux_tmp_411;
  wire mux_tmp_412;
  wire mux_tmp_420;
  wire mux_tmp_427;
  wire mux_tmp_428;
  wire not_tmp_253;
  wire or_tmp_382;
  wire mux_tmp_462;
  wire mux_tmp_463;
  wire mux_tmp_466;
  wire mux_tmp_469;
  wire not_tmp_265;
  wire mux_tmp_471;
  wire mux_tmp_473;
  wire mux_tmp_474;
  wire mux_tmp_476;
  wire mux_tmp_481;
  wire and_dcpl_166;
  wire or_dcpl_35;
  wire or_dcpl_36;
  wire or_dcpl_38;
  wire or_dcpl_41;
  wire or_dcpl_42;
  wire or_dcpl_43;
  wire mux_tmp_495;
  wire nor_tmp_162;
  wire and_dcpl_168;
  wire not_tmp_279;
  wire and_dcpl_169;
  wire or_dcpl_47;
  wire or_dcpl_53;
  wire or_dcpl_54;
  wire or_dcpl_59;
  reg exit_COMP_LOOP_1_modExp_1_while_sva;
  reg modExp_exp_1_0_1_sva;
  reg COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  reg [11:0] VEC_LOOP_j_sva_11_0;
  reg [6:0] COMP_LOOP_k_9_2_sva_6_0;
  reg [11:0] COMP_LOOP_acc_1_cse_2_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_sva;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_sva;
  reg [10:0] COMP_LOOP_acc_11_psp_sva;
  reg [11:0] COMP_LOOP_acc_10_cse_12_1_1_sva;
  reg [63:0] COMP_LOOP_1_acc_5_mut;
  wire and_144_m1c;
  wire and_198_m1c;
  reg reg_vec_rsc_triosy_0_3_obj_ld_cse;
  wire or_644_cse;
  wire or_287_cse;
  wire and_289_cse;
  wire or_319_cse;
  wire and_281_cse;
  wire and_273_cse;
  wire and_93_cse;
  wire and_206_cse;
  wire nor_380_cse;
  wire and_333_cse;
  wire and_332_cse;
  wire or_604_cse;
  wire nor_92_cse;
  wire or_585_cse;
  wire [63:0] modulo_result_mux_1_cse;
  wire and_313_cse;
  wire nand_53_cse;
  wire or_641_cse;
  wire nand_79_cse;
  wire or_625_cse;
  wire or_92_cse;
  wire nor_246_cse;
  wire or_481_cse;
  wire mux_152_cse;
  wire mux_150_cse;
  wire and_365_cse;
  wire or_642_cse;
  wire mux_66_cse;
  wire or_589_cse;
  wire mux_93_cse;
  wire mux_180_cse;
  wire or_643_cse;
  wire mux_561_cse;
  wire mux_558_cse;
  wire [9:0] COMP_LOOP_acc_psp_sva_1;
  wire [10:0] nl_COMP_LOOP_acc_psp_sva_1;
  reg [9:0] COMP_LOOP_acc_psp_sva;
  wire mux_139_itm;
  wire mux_351_itm;
  wire mux_391_itm;
  wire mux_522_itm;
  wire and_dcpl_194;
  wire [64:0] z_out;
  wire [64:0] z_out_1;
  wire [65:0] nl_z_out_1;
  wire and_dcpl_225;
  wire [12:0] z_out_2;
  wire [13:0] nl_z_out_2;
  wire and_dcpl_250;
  wire and_dcpl_257;
  wire and_dcpl_273;
  wire and_dcpl_279;
  wire and_dcpl_281;
  wire and_dcpl_285;
  wire and_dcpl_292;
  wire and_dcpl_301;
  wire [63:0] z_out_5;
  wire [64:0] nl_z_out_5;
  wire and_dcpl_309;
  wire and_dcpl_312;
  wire and_dcpl_317;
  wire and_dcpl_320;
  wire and_dcpl_325;
  wire [11:0] z_out_6;
  wire not_tmp_390;
  wire [63:0] z_out_7;
  wire signed [128:0] nl_z_out_7;
  reg [63:0] p_sva;
  reg [63:0] r_sva;
  reg [3:0] STAGE_LOOP_i_3_0_sva;
  reg [9:0] STAGE_LOOP_lshift_psp_sva;
  reg [63:0] modExp_result_sva;
  reg modExp_exp_1_7_1_sva;
  reg modExp_exp_1_5_1_sva;
  reg modExp_exp_1_4_1_sva;
  reg modExp_exp_1_3_1_sva;
  reg modExp_exp_1_2_1_sva;
  reg modExp_exp_1_1_1_sva;
  reg modExp_exp_1_0_1_sva_1;
  reg modExp_exp_1_5_1_sva_1;
  reg [63:0] modExp_while_if_mul_mut;
  reg [63:0] COMP_LOOP_1_modExp_1_while_if_mul_mut;
  reg [63:0] COMP_LOOP_1_mul_mut;
  reg [63:0] COMP_LOOP_2_modExp_1_while_mul_mut;
  reg [63:0] COMP_LOOP_2_mul_mut;
  reg [63:0] COMP_LOOP_3_modExp_1_while_mul_mut;
  reg [63:0] COMP_LOOP_3_mul_mut;
  reg [63:0] COMP_LOOP_4_modExp_1_while_mul_mut;
  reg [63:0] COMP_LOOP_4_mul_mut;
  reg [63:0] modExp_while_mul_itm;
  reg [63:0] COMP_LOOP_1_modExp_1_while_mul_itm;
  reg [63:0] COMP_LOOP_2_modExp_1_while_if_mul_itm;
  reg [63:0] COMP_LOOP_3_modExp_1_while_if_mul_itm;
  reg [63:0] COMP_LOOP_4_modExp_1_while_if_mul_itm;
  reg [63:0] COMP_LOOP_1_acc_8_itm;
  wire STAGE_LOOP_i_3_0_sva_mx0c1;
  wire [3:0] STAGE_LOOP_i_3_0_sva_2;
  wire [4:0] nl_STAGE_LOOP_i_3_0_sva_2;
  wire [63:0] modulo_qr_sva_1_mx0w1;
  wire [64:0] nl_modulo_qr_sva_1_mx0w1;
  wire [63:0] COMP_LOOP_1_acc_5_mut_mx0w7;
  wire [64:0] nl_COMP_LOOP_1_acc_5_mut_mx0w7;
  wire [63:0] COMP_LOOP_1_modExp_1_while_if_mul_mut_1;
  wire signed [127:0] nl_COMP_LOOP_1_modExp_1_while_if_mul_mut_1;
  wire [9:0] STAGE_LOOP_lshift_psp_sva_mx0w0;
  wire VEC_LOOP_j_sva_11_0_mx0c1;
  wire modExp_result_sva_mx0c0;
  wire [62:0] operator_64_false_slc_modExp_exp_63_1_3;
  wire modExp_while_and_3;
  wire modExp_while_and_5;
  wire and_156_m1c;
  wire modExp_result_and_rgt;
  wire modExp_result_and_1_rgt;
  wire and_390_ssc;
  wire COMP_LOOP_or_2_cse;
  wire nor_353_cse;
  wire nor_399_cse;
  wire and_323_cse;
  wire and_441_cse;
  wire nor_tmp;
  wire mux_tmp;
  wire nor_tmp_210;
  wire mux_tmp_613;
  wire or_tmp;
  wire mux_tmp_616;
  wire not_tmp_397;
  wire [64:0] operator_64_false_mux1h_1_rgt;
  wire not_tmp_400;
  reg operator_64_false_acc_mut_64;
  reg [63:0] operator_64_false_acc_mut_63_0;
  wire COMP_LOOP_or_22_itm;
  wire COMP_LOOP_or_24_itm;
  wire STAGE_LOOP_acc_itm_2_1;

  wire[0:0] nor_323_nl;
  wire[0:0] nor_324_nl;
  wire[0:0] mux_151_nl;
  wire[0:0] or_164_nl;
  wire[0:0] nand_5_nl;
  wire[0:0] mux_179_nl;
  wire[0:0] nor_300_nl;
  wire[0:0] and_301_nl;
  wire[0:0] nor_303_nl;
  wire[0:0] modulo_result_or_nl;
  wire[0:0] and_96_nl;
  wire[0:0] and_101_nl;
  wire[0:0] mux_206_nl;
  wire[0:0] nor_279_nl;
  wire[0:0] mux_205_nl;
  wire[0:0] or_279_nl;
  wire[0:0] nand_20_nl;
  wire[0:0] mux_204_nl;
  wire[0:0] nor_280_nl;
  wire[0:0] nor_281_nl;
  wire[0:0] nor_282_nl;
  wire[0:0] mux_203_nl;
  wire[0:0] nand_104_nl;
  wire[0:0] or_271_nl;
  wire[0:0] and_102_nl;
  wire[0:0] mux_209_nl;
  wire[0:0] mux_208_nl;
  wire[0:0] mux_207_nl;
  wire[0:0] or_281_nl;
  wire[0:0] and_104_nl;
  wire[0:0] mux_214_nl;
  wire[0:0] mux_213_nl;
  wire[0:0] mux_211_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] and_107_nl;
  wire[0:0] mux_229_nl;
  wire[0:0] mux_228_nl;
  wire[0:0] nor_276_nl;
  wire[0:0] mux_227_nl;
  wire[0:0] nand_24_nl;
  wire[0:0] and_288_nl;
  wire[0:0] mux_226_nl;
  wire[0:0] and_366_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] mux_224_nl;
  wire[0:0] nand_121_nl;
  wire[0:0] and_291_nl;
  wire[0:0] mux_223_nl;
  wire[0:0] mux_222_nl;
  wire[0:0] and_362_nl;
  wire[0:0] mux_221_nl;
  wire[0:0] mux_220_nl;
  wire[0:0] nor_278_nl;
  wire[0:0] nor_382_nl;
  wire[0:0] mux_219_nl;
  wire[0:0] or_298_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] mux_246_nl;
  wire[0:0] mux_245_nl;
  wire[0:0] mux_244_nl;
  wire[0:0] mux_243_nl;
  wire[0:0] nand_100_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] or_312_nl;
  wire[0:0] nand_26_nl;
  wire[0:0] mux_241_nl;
  wire[0:0] nand_102_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] mux_236_nl;
  wire[0:0] or_308_nl;
  wire[0:0] mux_235_nl;
  wire[0:0] mux_234_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] nand_55_nl;
  wire[0:0] mux_232_nl;
  wire[0:0] nand_56_nl;
  wire[0:0] mux_231_nl;
  wire[0:0] and_114_nl;
  wire[0:0] mux_250_nl;
  wire[0:0] nand_107_nl;
  wire[0:0] and_115_nl;
  wire[0:0] mux_253_nl;
  wire[0:0] nand_27_nl;
  wire[0:0] mux_252_nl;
  wire[0:0] mux_251_nl;
  wire[0:0] nand_54_nl;
  wire[0:0] and_117_nl;
  wire[0:0] mux_257_nl;
  wire[0:0] mux_256_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] mux_254_nl;
  wire[0:0] and_119_nl;
  wire[0:0] mux_261_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] mux_259_nl;
  wire[0:0] mux_645_nl;
  wire[0:0] and_123_nl;
  wire[0:0] and_126_nl;
  wire[0:0] mux_262_nl;
  wire[0:0] nor_275_nl;
  wire[0:0] and_128_nl;
  wire[0:0] and_130_nl;
  wire[0:0] mux_265_nl;
  wire[0:0] mux_264_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] mux_614_nl;
  wire[0:0] and_131_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] mux_267_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] and_278_nl;
  wire[0:0] nor_273_nl;
  wire[0:0] nor_274_nl;
  wire[0:0] mux_132_nl;
  wire[0:0] nor_272_nl;
  wire[63:0] COMP_LOOP_mux1h_44_nl;
  wire[0:0] COMP_LOOP_or_6_nl;
  wire[0:0] mux_565_nl;
  wire[0:0] mux_564_nl;
  wire[0:0] nor_218_nl;
  wire[0:0] nor_219_nl;
  wire[0:0] nor_220_nl;
  wire[0:0] COMP_LOOP_or_7_nl;
  wire[0:0] mux_567_nl;
  wire[0:0] mux_566_nl;
  wire[0:0] nor_215_nl;
  wire[0:0] nor_216_nl;
  wire[0:0] nor_217_nl;
  wire[0:0] COMP_LOOP_or_8_nl;
  wire[0:0] mux_569_nl;
  wire[0:0] mux_568_nl;
  wire[0:0] nor_212_nl;
  wire[0:0] nor_213_nl;
  wire[0:0] nor_214_nl;
  wire[0:0] COMP_LOOP_or_9_nl;
  wire[0:0] mux_571_nl;
  wire[0:0] mux_570_nl;
  wire[0:0] nor_210_nl;
  wire[0:0] nor_211_nl;
  wire[0:0] and_213_nl;
  wire[0:0] and_137_nl;
  wire[0:0] mux_289_nl;
  wire[0:0] mux_288_nl;
  wire[0:0] mux_287_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] mux_285_nl;
  wire[0:0] mux_284_nl;
  wire[0:0] mux_281_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] mux_279_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] mux_635_nl;
  wire[0:0] mux_634_nl;
  wire[0:0] mux_633_nl;
  wire[0:0] mux_632_nl;
  wire[0:0] or_671_nl;
  wire[0:0] or_670_nl;
  wire[0:0] or_669_nl;
  wire[0:0] mux_631_nl;
  wire[0:0] mux_630_nl;
  wire[0:0] mux_629_nl;
  wire[0:0] mux_628_nl;
  wire[0:0] and_521_nl;
  wire[0:0] mux_627_nl;
  wire[0:0] mux_626_nl;
  wire[0:0] mux_625_nl;
  wire[0:0] mux_624_nl;
  wire[0:0] mux_623_nl;
  wire[0:0] mux_622_nl;
  wire[0:0] mux_621_nl;
  wire[0:0] mux_620_nl;
  wire[0:0] mux_618_nl;
  wire[0:0] mux_617_nl;
  wire[0:0] mux_615_nl;
  wire[0:0] mux_640_nl;
  wire[0:0] mux_639_nl;
  wire[0:0] mux_638_nl;
  wire[0:0] or_688_nl;
  wire[0:0] nand_138_nl;
  wire[0:0] or_689_nl;
  wire[0:0] mux_637_nl;
  wire[0:0] or_690_nl;
  wire[0:0] nand_139_nl;
  wire[0:0] mux_313_nl;
  wire[0:0] or_nl;
  wire[0:0] nand_134_nl;
  wire[0:0] mux_312_nl;
  wire[0:0] nor_268_nl;
  wire[0:0] nor_269_nl;
  wire[0:0] nor_420_nl;
  wire[0:0] mux_642_nl;
  wire[0:0] or_686_nl;
  wire[0:0] or_685_nl;
  wire[0:0] nor_421_nl;
  wire[0:0] mux_641_nl;
  wire[0:0] or_682_nl;
  wire[0:0] or_680_nl;
  wire[0:0] mux_325_nl;
  wire[0:0] mux_324_nl;
  wire[0:0] nor_261_nl;
  wire[0:0] COMP_LOOP_and_nl;
  wire[0:0] COMP_LOOP_and_1_nl;
  wire[0:0] mux_380_nl;
  wire[0:0] mux_379_nl;
  wire[0:0] mux_378_nl;
  wire[0:0] mux_377_nl;
  wire[0:0] mux_376_nl;
  wire[0:0] mux_375_nl;
  wire[0:0] mux_374_nl;
  wire[0:0] mux_373_nl;
  wire[0:0] mux_372_nl;
  wire[0:0] mux_371_nl;
  wire[0:0] mux_370_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] mux_368_nl;
  wire[0:0] mux_367_nl;
  wire[0:0] mux_366_nl;
  wire[0:0] mux_365_nl;
  wire[0:0] or_366_nl;
  wire[0:0] mux_364_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] mux_362_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] mux_360_nl;
  wire[0:0] mux_359_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] mux_357_nl;
  wire[0:0] mux_356_nl;
  wire[0:0] mux_355_nl;
  wire[0:0] mux_350_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] mux_348_nl;
  wire[0:0] mux_347_nl;
  wire[0:0] mux_346_nl;
  wire[0:0] and_150_nl;
  wire[0:0] mux_345_nl;
  wire[0:0] and_258_nl;
  wire[0:0] mux_343_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] mux_341_nl;
  wire[0:0] mux_338_nl;
  wire[0:0] mux_335_nl;
  wire[0:0] mux_334_nl;
  wire[0:0] mux_331_nl;
  wire[0:0] mux_386_nl;
  wire[0:0] and_364_nl;
  wire[0:0] nor_255_nl;
  wire[0:0] and_153_nl;
  wire[0:0] COMP_LOOP_or_12_nl;
  wire[0:0] COMP_LOOP_or_13_nl;
  wire[0:0] nor_388_nl;
  wire[0:0] and_162_nl;
  wire[0:0] and_165_nl;
  wire[0:0] and_168_nl;
  wire[0:0] mux_441_nl;
  wire[0:0] mux_440_nl;
  wire[0:0] mux_439_nl;
  wire[0:0] mux_438_nl;
  wire[0:0] mux_437_nl;
  wire[0:0] mux_436_nl;
  wire[0:0] mux_435_nl;
  wire[0:0] mux_434_nl;
  wire[0:0] mux_433_nl;
  wire[0:0] mux_432_nl;
  wire[0:0] mux_431_nl;
  wire[0:0] mux_430_nl;
  wire[0:0] mux_429_nl;
  wire[0:0] mux_426_nl;
  wire[0:0] mux_425_nl;
  wire[0:0] mux_424_nl;
  wire[0:0] mux_423_nl;
  wire[0:0] mux_422_nl;
  wire[0:0] mux_421_nl;
  wire[0:0] mux_418_nl;
  wire[0:0] mux_417_nl;
  wire[0:0] mux_416_nl;
  wire[0:0] mux_415_nl;
  wire[0:0] mux_414_nl;
  wire[0:0] mux_413_nl;
  wire[0:0] mux_410_nl;
  wire[0:0] mux_407_nl;
  wire[0:0] mux_406_nl;
  wire[0:0] mux_405_nl;
  wire[0:0] mux_402_nl;
  wire[0:0] mux_401_nl;
  wire[0:0] mux_400_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] nand_49_nl;
  wire[0:0] mux_398_nl;
  wire[0:0] mux_396_nl;
  wire[0:0] mux_395_nl;
  wire[0:0] and_337_nl;
  wire[0:0] COMP_LOOP_mux1h_18_nl;
  wire[0:0] COMP_LOOP_and_9_nl;
  wire[0:0] mux_460_nl;
  wire[0:0] mux_459_nl;
  wire[0:0] mux_458_nl;
  wire[0:0] mux_457_nl;
  wire[0:0] mux_75_nl;
  wire[0:0] and_335_nl;
  wire[0:0] nor_351_nl;
  wire[0:0] mux_455_nl;
  wire[0:0] or_75_nl;
  wire[0:0] or_409_nl;
  wire[0:0] or_408_nl;
  wire[0:0] mux_454_nl;
  wire[0:0] mux_453_nl;
  wire[0:0] or_405_nl;
  wire[0:0] or_403_nl;
  wire[0:0] or_402_nl;
  wire[0:0] mux_72_nl;
  wire[0:0] mux_71_nl;
  wire[0:0] mux_70_nl;
  wire[0:0] mux_69_nl;
  wire[0:0] nand_93_nl;
  wire[0:0] nand_94_nl;
  wire[0:0] mux_68_nl;
  wire[0:0] nor_378_nl;
  wire[0:0] mux_67_nl;
  wire[0:0] nor_379_nl;
  wire[0:0] mux_445_nl;
  wire[0:0] nor_245_nl;
  wire[0:0] mux_488_nl;
  wire[0:0] mux_487_nl;
  wire[0:0] mux_486_nl;
  wire[0:0] mux_485_nl;
  wire[0:0] mux_484_nl;
  wire[0:0] mux_483_nl;
  wire[0:0] mux_482_nl;
  wire[0:0] mux_480_nl;
  wire[0:0] mux_479_nl;
  wire[0:0] mux_478_nl;
  wire[0:0] mux_477_nl;
  wire[0:0] mux_472_nl;
  wire[0:0] mux_489_nl;
  wire[0:0] nand_106_nl;
  wire[9:0] COMP_LOOP_1_acc_nl;
  wire[10:0] nl_COMP_LOOP_1_acc_nl;
  wire[0:0] mux_493_nl;
  wire[0:0] nor_369_nl;
  wire[0:0] mux_492_nl;
  wire[0:0] nor_370_nl;
  wire[0:0] and_361_nl;
  wire[0:0] mux_501_nl;
  wire[0:0] mux_500_nl;
  wire[0:0] mux_499_nl;
  wire[0:0] mux_498_nl;
  wire[0:0] mux_497_nl;
  wire[0:0] mux_496_nl;
  wire[0:0] mux_494_nl;
  wire[0:0] mux_505_nl;
  wire[0:0] nor_239_nl;
  wire[0:0] mux_504_nl;
  wire[0:0] nor_240_nl;
  wire[0:0] mux_503_nl;
  wire[0:0] and_241_nl;
  wire[0:0] COMP_LOOP_mux_24_nl;
  wire[0:0] mux_538_nl;
  wire[0:0] and_226_nl;
  wire[0:0] mux_537_nl;
  wire[0:0] nor_228_nl;
  wire[0:0] mux_536_nl;
  wire[0:0] or_478_nl;
  wire[0:0] or_477_nl;
  wire[0:0] nor_229_nl;
  wire[0:0] nor_230_nl;
  wire[0:0] mux_524_nl;
  wire[0:0] nor_234_nl;
  wire[0:0] nor_235_nl;
  wire[0:0] mux_549_nl;
  wire[0:0] mux_548_nl;
  wire[0:0] mux_547_nl;
  wire[0:0] nand_34_nl;
  wire[0:0] mux_546_nl;
  wire[0:0] nand_39_nl;
  wire[0:0] nor_225_nl;
  wire[0:0] mux_545_nl;
  wire[0:0] or_490_nl;
  wire[0:0] mux_544_nl;
  wire[0:0] or_489_nl;
  wire[0:0] or_487_nl;
  wire[0:0] mux_543_nl;
  wire[0:0] mux_542_nl;
  wire[0:0] mux_541_nl;
  wire[0:0] nand_41_nl;
  wire[0:0] or_483_nl;
  wire[0:0] mux_540_nl;
  wire[0:0] mux_539_nl;
  wire[0:0] or_12_nl;
  wire[0:0] COMP_LOOP_mux1h_29_nl;
  wire[0:0] mux_551_nl;
  wire[0:0] nand_130_nl;
  wire[0:0] mux_550_nl;
  wire[0:0] nor_222_nl;
  wire[0:0] nor_223_nl;
  wire[0:0] nand_131_nl;
  wire[0:0] and_190_nl;
  wire[0:0] mux_560_nl;
  wire[0:0] or_506_nl;
  wire[0:0] mux_557_nl;
  wire[0:0] mux_556_nl;
  wire[0:0] mux_555_nl;
  wire[0:0] and_215_nl;
  wire[0:0] mux_529_nl;
  wire[0:0] or_500_nl;
  wire[0:0] mux_525_nl;
  wire[0:0] or_465_nl;
  wire[0:0] COMP_LOOP_mux1h_43_nl;
  wire[0:0] mux_563_nl;
  wire[0:0] mux_562_nl;
  wire[0:0] mux_559_nl;
  wire[0:0] or_504_nl;
  wire[0:0] mux_587_nl;
  wire[0:0] mux_586_nl;
  wire[0:0] or_533_nl;
  wire[10:0] acc_3_nl;
  wire[11:0] nl_acc_3_nl;
  wire[1:0] COMP_LOOP_mux_28_nl;
  wire[0:0] and_527_nl;
  wire[0:0] mux_598_nl;
  wire[0:0] mux_597_nl;
  wire[0:0] mux_596_nl;
  wire[0:0] mux_595_nl;
  wire[0:0] mux_600_nl;
  wire[0:0] mux_599_nl;
  wire[0:0] mux_603_nl;
  wire[0:0] mux_602_nl;
  wire[0:0] mux_601_nl;
  wire[0:0] or_40_nl;
  wire[0:0] or_38_nl;
  wire[0:0] mux_138_nl;
  wire[0:0] nor_338_nl;
  wire[0:0] and_30_nl;
  wire[0:0] or_611_nl;
  wire[0:0] nand_61_nl;
  wire[0:0] mux_218_nl;
  wire[0:0] nor_336_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] or_295_nl;
  wire[0:0] nor_337_nl;
  wire[0:0] mux_216_nl;
  wire[0:0] or_291_nl;
  wire[0:0] or_309_nl;
  wire[0:0] mux_238_nl;
  wire[0:0] nand_25_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] mux_249_nl;
  wire[0:0] mux_271_nl;
  wire[0:0] and_277_nl;
  wire[0:0] nor_271_nl;
  wire[0:0] mux_277_nl;
  wire[0:0] nor_263_nl;
  wire[0:0] and_358_nl;
  wire[0:0] mux_328_nl;
  wire[0:0] mux_326_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] mux_353_nl;
  wire[0:0] mux_43_nl;
  wire[0:0] mux_38_nl;
  wire[0:0] or_36_nl;
  wire[0:0] or_34_nl;
  wire[0:0] nor_256_nl;
  wire[0:0] mux_384_nl;
  wire[0:0] or_375_nl;
  wire[0:0] or_373_nl;
  wire[0:0] and_257_nl;
  wire[0:0] mux_383_nl;
  wire[0:0] nor_257_nl;
  wire[0:0] nor_258_nl;
  wire[0:0] and_255_nl;
  wire[0:0] mux_388_nl;
  wire[0:0] nor_250_nl;
  wire[0:0] nor_251_nl;
  wire[0:0] and_256_nl;
  wire[0:0] mux_387_nl;
  wire[0:0] nor_252_nl;
  wire[0:0] nor_253_nl;
  wire[0:0] mux_390_nl;
  wire[0:0] mux_419_nl;
  wire[0:0] mux_443_nl;
  wire[0:0] nor_247_nl;
  wire[0:0] nor_248_nl;
  wire[0:0] nor_249_nl;
  wire[0:0] and_176_nl;
  wire[0:0] mux_465_nl;
  wire[0:0] mux_464_nl;
  wire[0:0] mux_468_nl;
  wire[0:0] mux_467_nl;
  wire[0:0] mux_470_nl;
  wire[0:0] mux_475_nl;
  wire[0:0] and_177_nl;
  wire[0:0] nor_237_nl;
  wire[0:0] mux_508_nl;
  wire[0:0] or_450_nl;
  wire[0:0] or_449_nl;
  wire[0:0] nor_238_nl;
  wire[0:0] mux_507_nl;
  wire[0:0] or_446_nl;
  wire[0:0] or_445_nl;
  wire[0:0] mux_521_nl;
  wire[0:0] mux_518_nl;
  wire[0:0] or_459_nl;
  wire[0:0] mux_517_nl;
  wire[0:0] or_458_nl;
  wire[0:0] mux_42_nl;
  wire[0:0] or_32_nl;
  wire[0:0] mux_322_nl;
  wire[0:0] nor_262_nl;
  wire[2:0] STAGE_LOOP_acc_nl;
  wire[3:0] nl_STAGE_LOOP_acc_nl;
  wire[0:0] and_63_nl;
  wire[0:0] nor_377_nl;
  wire[0:0] mux_143_nl;
  wire[0:0] nand_112_nl;
  wire[0:0] mux_142_nl;
  wire[0:0] nor_332_nl;
  wire[0:0] mux_141_nl;
  wire[0:0] nand_82_nl;
  wire[0:0] or_137_nl;
  wire[0:0] nor_333_nl;
  wire[0:0] and_67_nl;
  wire[0:0] mux_144_nl;
  wire[0:0] nor_330_nl;
  wire[0:0] nor_331_nl;
  wire[0:0] and_75_nl;
  wire[0:0] mux_145_nl;
  wire[0:0] nor_329_nl;
  wire[0:0] and_308_nl;
  wire[0:0] and_80_nl;
  wire[0:0] mux_146_nl;
  wire[0:0] nor_327_nl;
  wire[0:0] nor_328_nl;
  wire[0:0] nor_322_nl;
  wire[0:0] and_307_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] nor_325_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] or_156_nl;
  wire[0:0] or_154_nl;
  wire[0:0] nor_326_nl;
  wire[0:0] mux_147_nl;
  wire[0:0] or_151_nl;
  wire[0:0] or_149_nl;
  wire[0:0] mux_160_nl;
  wire[0:0] nand_111_nl;
  wire[0:0] mux_159_nl;
  wire[0:0] mux_158_nl;
  wire[0:0] nor_317_nl;
  wire[0:0] nor_318_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] nor_319_nl;
  wire[0:0] nor_320_nl;
  wire[0:0] or_640_nl;
  wire[0:0] mux_156_nl;
  wire[0:0] or_172_nl;
  wire[0:0] mux_155_nl;
  wire[0:0] or_171_nl;
  wire[0:0] or_170_nl;
  wire[0:0] mux_154_nl;
  wire[0:0] or_168_nl;
  wire[0:0] or_167_nl;
  wire[0:0] nor_311_nl;
  wire[0:0] and_304_nl;
  wire[0:0] mux_163_nl;
  wire[0:0] and_305_nl;
  wire[0:0] mux_162_nl;
  wire[0:0] nor_314_nl;
  wire[0:0] nor_315_nl;
  wire[0:0] nor_316_nl;
  wire[0:0] mux_161_nl;
  wire[0:0] or_183_nl;
  wire[0:0] or_181_nl;
  wire[0:0] mux_174_nl;
  wire[0:0] nand_110_nl;
  wire[0:0] mux_173_nl;
  wire[0:0] mux_172_nl;
  wire[0:0] nor_306_nl;
  wire[0:0] nor_307_nl;
  wire[0:0] mux_171_nl;
  wire[0:0] nor_308_nl;
  wire[0:0] nor_309_nl;
  wire[0:0] or_639_nl;
  wire[0:0] mux_170_nl;
  wire[0:0] or_202_nl;
  wire[0:0] mux_169_nl;
  wire[0:0] or_201_nl;
  wire[0:0] or_200_nl;
  wire[0:0] mux_168_nl;
  wire[0:0] or_198_nl;
  wire[0:0] or_197_nl;
  wire[0:0] and_300_nl;
  wire[0:0] and_302_nl;
  wire[0:0] mux_177_nl;
  wire[0:0] nor_304_nl;
  wire[0:0] mux_176_nl;
  wire[0:0] or_218_nl;
  wire[0:0] or_216_nl;
  wire[0:0] nor_305_nl;
  wire[0:0] mux_175_nl;
  wire[0:0] or_213_nl;
  wire[0:0] or_211_nl;
  wire[0:0] mux_188_nl;
  wire[0:0] nand_109_nl;
  wire[0:0] mux_187_nl;
  wire[0:0] mux_186_nl;
  wire[0:0] nor_295_nl;
  wire[0:0] nor_296_nl;
  wire[0:0] mux_185_nl;
  wire[0:0] nor_297_nl;
  wire[0:0] nor_298_nl;
  wire[0:0] or_638_nl;
  wire[0:0] mux_184_nl;
  wire[0:0] or_232_nl;
  wire[0:0] mux_183_nl;
  wire[0:0] or_231_nl;
  wire[0:0] or_230_nl;
  wire[0:0] mux_182_nl;
  wire[0:0] or_228_nl;
  wire[0:0] or_227_nl;
  wire[0:0] and_295_nl;
  wire[0:0] and_297_nl;
  wire[0:0] mux_191_nl;
  wire[0:0] and_298_nl;
  wire[0:0] mux_190_nl;
  wire[0:0] nor_292_nl;
  wire[0:0] nor_293_nl;
  wire[0:0] nor_294_nl;
  wire[0:0] mux_189_nl;
  wire[0:0] or_242_nl;
  wire[0:0] nand_105_nl;
  wire[0:0] mux_202_nl;
  wire[0:0] nand_108_nl;
  wire[0:0] mux_201_nl;
  wire[0:0] mux_200_nl;
  wire[0:0] and_363_nl;
  wire[0:0] nor_284_nl;
  wire[0:0] mux_199_nl;
  wire[0:0] nor_285_nl;
  wire[0:0] nor_286_nl;
  wire[0:0] or_637_nl;
  wire[0:0] mux_198_nl;
  wire[0:0] or_259_nl;
  wire[0:0] mux_197_nl;
  wire[0:0] nand_64_nl;
  wire[0:0] or_257_nl;
  wire[0:0] mux_196_nl;
  wire[0:0] or_255_nl;
  wire[0:0] or_254_nl;
  wire[0:0] mux_608_nl;
  wire[0:0] and_nl;
  wire[0:0] mux_607_nl;
  wire[0:0] nor_nl;
  wire[0:0] nor_392_nl;
  wire[0:0] nor_393_nl;
  wire[0:0] nor_423_nl;
  wire[0:0] nor_424_nl;
  wire[65:0] acc_nl;
  wire[66:0] nl_acc_nl;
  wire[63:0] COMP_LOOP_mux_26_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_nand_2_nl;
  wire[0:0] mux_646_nl;
  wire[0:0] and_525_nl;
  wire[0:0] mux_647_nl;
  wire[0:0] and_526_nl;
  wire[0:0] mux_648_nl;
  wire[0:0] nor_425_nl;
  wire[0:0] nor_426_nl;
  wire[0:0] nor_427_nl;
  wire[0:0] nor_428_nl;
  wire[63:0] COMP_LOOP_COMP_LOOP_nand_3_nl;
  wire[0:0] COMP_LOOP_not_101_nl;
  wire[56:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_52_nl;
  wire[0:0] COMP_LOOP_not_102_nl;
  wire[6:0] COMP_LOOP_mux_27_nl;
  wire[11:0] operator_64_false_1_mux_2_nl;
  wire[9:0] operator_64_false_1_mux_3_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_4_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_53_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_54_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_55_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_56_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_57_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_58_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_59_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_60_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_61_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_62_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_63_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_64_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_65_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_66_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_67_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_68_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_69_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_70_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_71_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_72_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_73_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_74_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_75_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_76_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_77_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_78_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_79_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_80_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_81_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_82_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_83_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_84_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_85_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_86_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_87_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_88_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_89_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_90_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_91_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_92_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_93_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_94_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_95_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_96_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_97_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_98_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_99_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_100_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_101_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_102_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_103_nl;
  wire[11:0] COMP_LOOP_mux1h_89_nl;
  wire[9:0] COMP_LOOP_mux1h_90_nl;
  wire[9:0] COMP_LOOP_acc_35_nl;
  wire[10:0] nl_COMP_LOOP_acc_35_nl;
  wire[1:0] COMP_LOOP_COMP_LOOP_or_3_nl;
  wire[1:0] COMP_LOOP_COMP_LOOP_nor_2_nl;
  wire[1:0] COMP_LOOP_mux_29_nl;
  wire[0:0] and_528_nl;
  wire[0:0] and_529_nl;
  wire[12:0] acc_6_nl;
  wire[13:0] nl_acc_6_nl;
  wire[3:0] COMP_LOOP_COMP_LOOP_or_5_nl;
  wire[3:0] COMP_LOOP_and_16_nl;
  wire[0:0] not_1471_nl;
  wire[0:0] COMP_LOOP_or_30_nl;
  wire[0:0] COMP_LOOP_mux1h_91_nl;
  wire[0:0] COMP_LOOP_mux1h_92_nl;
  wire[0:0] COMP_LOOP_mux1h_93_nl;
  wire[0:0] COMP_LOOP_mux1h_94_nl;
  wire[0:0] COMP_LOOP_mux1h_95_nl;
  wire[0:0] COMP_LOOP_mux1h_96_nl;
  wire[0:0] COMP_LOOP_mux1h_97_nl;
  wire[0:0] COMP_LOOP_mux1h_98_nl;
  wire[0:0] COMP_LOOP_or_31_nl;
  wire[8:0] COMP_LOOP_mux1h_99_nl;
  wire[63:0] modExp_while_if_mux_1_nl;
  wire[0:0] nor_429_nl;
  wire[0:0] mux_649_nl;
  wire[0:0] mux_650_nl;
  wire[0:0] or_694_nl;
  wire[0:0] mux_651_nl;
  wire[0:0] or_695_nl;
  wire[0:0] or_696_nl;
  wire[0:0] or_697_nl;
  wire[0:0] mux_652_nl;
  wire[0:0] or_698_nl;
  wire[0:0] or_699_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [10:0] nl_operator_66_true_div_cmp_b;
  assign nl_operator_66_true_div_cmp_b = {1'b0, operator_66_true_div_cmp_b_9_0};
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0 = ~ (z_out_1[64]);
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0 = ~ modExp_exp_1_0_1_sva;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_68_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_68_tr0 = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_42_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_42_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_136_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_136_tr0 = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_42_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_42_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_204_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_204_tr0 = ~ modExp_exp_1_0_1_sva;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_42_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_42_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 = z_out_2[12];
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_10_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_10_tr0 = ~ STAGE_LOOP_acc_itm_2_1;
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd64)) r_rsci (
      .dat(r_rsc_dat),
      .idat(r_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_3_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(vec_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_2_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(vec_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_1_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(vec_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(vec_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd1)) modulo_result_rem_cmp (
      .a(modulo_result_rem_cmp_a),
      .b(modulo_result_rem_cmp_b),
      .z(modulo_result_rem_cmp_z)
    );
  mgc_div #(.width_a(32'sd65),
  .width_b(32'sd11),
  .signd(32'sd1)) operator_66_true_div_cmp (
      .a(operator_66_true_div_cmp_a),
      .b(nl_operator_66_true_div_cmp_b[10:0]),
      .z(operator_66_true_div_cmp_z)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd10)) STAGE_LOOP_lshift_rg (
      .a(1'b1),
      .s(STAGE_LOOP_i_3_0_sva),
      .z(STAGE_LOOP_lshift_psp_sva_mx0w0)
    );
  inPlaceNTT_DIT_core_core_fsm inPlaceNTT_DIT_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .STAGE_LOOP_C_9_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0[0:0]),
      .modExp_while_C_42_tr0(exit_COMP_LOOP_1_modExp_1_while_sva),
      .COMP_LOOP_C_1_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0[0:0]),
      .COMP_LOOP_1_modExp_1_while_C_42_tr0(exit_COMP_LOOP_1_modExp_1_while_sva),
      .COMP_LOOP_C_68_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_68_tr0[0:0]),
      .COMP_LOOP_2_modExp_1_while_C_42_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_42_tr0[0:0]),
      .COMP_LOOP_C_136_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_136_tr0[0:0]),
      .COMP_LOOP_3_modExp_1_while_C_42_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_42_tr0[0:0]),
      .COMP_LOOP_C_204_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_204_tr0[0:0]),
      .COMP_LOOP_4_modExp_1_while_C_42_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_42_tr0[0:0]),
      .COMP_LOOP_C_272_tr0(exit_COMP_LOOP_1_modExp_1_while_sva),
      .VEC_LOOP_C_0_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0[0:0]),
      .STAGE_LOOP_C_10_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_10_tr0[0:0])
    );
  assign nor_323_nl = ~((~ (fsm_output[1])) | (fsm_output[6]) | (~ (fsm_output[8]))
      | (fsm_output[7]));
  assign nor_324_nl = ~((fsm_output[1]) | nand_53_cse);
  assign mux_150_cse = MUX_s_1_2_2(nor_323_nl, nor_324_nl, fsm_output[5]);
  assign or_164_nl = (fsm_output[0]) | (fsm_output[5]) | (~ (fsm_output[1])) | (fsm_output[6])
      | nand_79_cse;
  assign nand_5_nl = ~((fsm_output[0]) & mux_150_cse);
  assign mux_151_nl = MUX_s_1_2_2(or_164_nl, nand_5_nl, fsm_output[4]);
  assign mux_152_cse = MUX_s_1_2_2(mux_151_nl, or_641_cse, fsm_output[2]);
  assign nor_300_nl = ~((fsm_output[0]) | (fsm_output[5]) | (~ (fsm_output[1])) |
      (fsm_output[6]) | nand_79_cse);
  assign and_301_nl = (fsm_output[0]) & mux_150_cse;
  assign mux_179_nl = MUX_s_1_2_2(nor_300_nl, and_301_nl, fsm_output[4]);
  assign nor_303_nl = ~((fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[5])) |
      (fsm_output[1]) | (fsm_output[6]) | (fsm_output[8]) | (~ (fsm_output[7])));
  assign mux_180_cse = MUX_s_1_2_2(mux_179_nl, nor_303_nl, fsm_output[2]);
  assign or_644_cse = (fsm_output[1:0]!=2'b00);
  assign or_287_cse = (fsm_output[2:1]!=2'b00);
  assign and_289_cse = (fsm_output[1:0]==2'b11);
  assign or_319_cse = (fsm_output[2:0]!=3'b000);
  assign and_281_cse = (fsm_output[2:0]==3'b111);
  assign and_93_cse = (fsm_output[3:2]==2'b11);
  assign nor_92_cse = ~((fsm_output[3]) | (~ (fsm_output[6])));
  assign and_365_cse = or_644_cse & (fsm_output[2]);
  assign or_642_cse = and_289_cse | (fsm_output[2]);
  assign or_643_cse = and_365_cse | (fsm_output[3]);
  assign and_313_cse = (fsm_output[2]) & (fsm_output[5]) & (fsm_output[4]) & (fsm_output[7])
      & (fsm_output[8]);
  assign and_273_cse = (fsm_output[5:4]==2'b11);
  assign and_206_cse = (fsm_output[2:1]==2'b11);
  assign or_604_cse = (fsm_output[5:4]!=2'b00);
  assign nor_218_nl = ~((COMP_LOOP_acc_1_cse_sva[1:0]!=2'b00) | (fsm_output[5:4]!=2'b00)
      | (~ nor_tmp_16));
  assign nor_219_nl = ~((COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b00) | (~ (fsm_output[5]))
      | (fsm_output[4]) | (fsm_output[8]) | (~ (fsm_output[7])));
  assign mux_564_nl = MUX_s_1_2_2(nor_218_nl, nor_219_nl, fsm_output[1]);
  assign nor_220_nl = ~((VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (~ (fsm_output[1])) |
      (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[8]) | (fsm_output[7]));
  assign mux_565_nl = MUX_s_1_2_2(mux_564_nl, nor_220_nl, fsm_output[0]);
  assign COMP_LOOP_or_6_nl = (mux_565_nl & and_dcpl_1) | ((~((VEC_LOOP_j_sva_11_0[0])
      | (COMP_LOOP_acc_11_psp_sva[0]))) & and_198_m1c);
  assign nor_215_nl = ~((COMP_LOOP_acc_1_cse_sva[1:0]!=2'b01) | (fsm_output[5:4]!=2'b00)
      | (~ nor_tmp_16));
  assign nor_216_nl = ~((COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b01) | (~ (fsm_output[5]))
      | (fsm_output[4]) | (fsm_output[8]) | (~ (fsm_output[7])));
  assign mux_566_nl = MUX_s_1_2_2(nor_215_nl, nor_216_nl, fsm_output[1]);
  assign nor_217_nl = ~((VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (~ (fsm_output[1])) |
      (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[8]) | (fsm_output[7]));
  assign mux_567_nl = MUX_s_1_2_2(mux_566_nl, nor_217_nl, fsm_output[0]);
  assign COMP_LOOP_or_7_nl = (mux_567_nl & and_dcpl_1) | ((VEC_LOOP_j_sva_11_0[0])
      & (~ (COMP_LOOP_acc_11_psp_sva[0])) & and_198_m1c);
  assign nor_212_nl = ~((COMP_LOOP_acc_1_cse_sva[1:0]!=2'b10) | (fsm_output[5:4]!=2'b00)
      | (~ nor_tmp_16));
  assign nor_213_nl = ~((COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b10) | (~ (fsm_output[5]))
      | (fsm_output[4]) | (fsm_output[8]) | (~ (fsm_output[7])));
  assign mux_568_nl = MUX_s_1_2_2(nor_212_nl, nor_213_nl, fsm_output[1]);
  assign nor_214_nl = ~((VEC_LOOP_j_sva_11_0[1:0]!=2'b10) | (~ (fsm_output[1])) |
      (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[8]) | (fsm_output[7]));
  assign mux_569_nl = MUX_s_1_2_2(mux_568_nl, nor_214_nl, fsm_output[0]);
  assign COMP_LOOP_or_8_nl = (mux_569_nl & and_dcpl_1) | ((COMP_LOOP_acc_11_psp_sva[0])
      & (~ (VEC_LOOP_j_sva_11_0[0])) & and_198_m1c);
  assign nor_210_nl = ~((COMP_LOOP_acc_1_cse_sva[1:0]!=2'b11) | (fsm_output[5:4]!=2'b00)
      | (~ nor_tmp_16));
  assign nor_211_nl = ~((COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b11) | (~ (fsm_output[5]))
      | (fsm_output[4]) | (fsm_output[8]) | (~ (fsm_output[7])));
  assign mux_570_nl = MUX_s_1_2_2(nor_210_nl, nor_211_nl, fsm_output[1]);
  assign and_213_nl = (VEC_LOOP_j_sva_11_0[1:0]==2'b11) & (fsm_output[1]) & (fsm_output[5])
      & (fsm_output[4]) & (~ (fsm_output[8])) & (~ (fsm_output[7]));
  assign mux_571_nl = MUX_s_1_2_2(mux_570_nl, and_213_nl, fsm_output[0]);
  assign COMP_LOOP_or_9_nl = (mux_571_nl & and_dcpl_1) | ((VEC_LOOP_j_sva_11_0[0])
      & (COMP_LOOP_acc_11_psp_sva[0]) & and_198_m1c);
  assign COMP_LOOP_mux1h_44_nl = MUX1HOT_v_64_4_2(vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d,
      vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d, {COMP_LOOP_or_6_nl , COMP_LOOP_or_7_nl
      , COMP_LOOP_or_8_nl , COMP_LOOP_or_9_nl});
  assign and_137_nl = and_dcpl_31 & and_dcpl_46 & and_dcpl_25;
  assign mux_285_nl = MUX_s_1_2_2(mux_tmp_282, mux_tmp_274, fsm_output[1]);
  assign mux_286_nl = MUX_s_1_2_2(mux_285_nl, mux_tmp_278, fsm_output[0]);
  assign mux_287_nl = MUX_s_1_2_2(mux_tmp_283, mux_286_nl, fsm_output[2]);
  assign mux_284_nl = MUX_s_1_2_2(mux_tmp_283, mux_tmp_282, and_281_cse);
  assign mux_288_nl = MUX_s_1_2_2((~ mux_287_nl), mux_284_nl, fsm_output[6]);
  assign mux_275_nl = MUX_s_1_2_2(mux_tmp_274, mux_tmp_273, fsm_output[1]);
  assign mux_279_nl = MUX_s_1_2_2(mux_tmp_278, mux_275_nl, fsm_output[0]);
  assign mux_280_nl = MUX_s_1_2_2(mux_279_nl, mux_tmp_273, fsm_output[2]);
  assign mux_281_nl = MUX_s_1_2_2((~ mux_tmp_273), mux_280_nl, fsm_output[6]);
  assign mux_289_nl = MUX_s_1_2_2(mux_288_nl, mux_281_nl, fsm_output[3]);
  assign operator_64_false_mux1h_1_rgt = MUX1HOT_v_65_3_2(z_out, ({2'b00 , operator_64_false_slc_modExp_exp_63_1_3}),
      ({1'b0 , COMP_LOOP_mux1h_44_nl}), {and_137_nl , and_dcpl_132 , (~ mux_289_nl)});
  assign nand_53_cse = ~((fsm_output[8:6]==3'b111));
  assign mux_93_cse = MUX_s_1_2_2((~ (fsm_output[8])), mux_tmp_86, fsm_output[4]);
  assign and_144_m1c = and_dcpl_30 & and_dcpl_36 & and_dcpl_27;
  assign modExp_result_and_rgt = (~ modExp_while_and_5) & and_144_m1c;
  assign modExp_result_and_1_rgt = modExp_while_and_5 & and_144_m1c;
  assign modulo_result_mux_1_cse = MUX_v_64_2_2(modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w1,
      modulo_result_rem_cmp_z[63]);
  assign and_364_nl = (fsm_output[2]) & (fsm_output[0]) & (~ (fsm_output[1])) & (fsm_output[4]);
  assign nor_255_nl = ~((fsm_output[2]) | (fsm_output[0]) | (~ (fsm_output[1])) |
      (fsm_output[4]));
  assign mux_386_nl = MUX_s_1_2_2(and_364_nl, nor_255_nl, fsm_output[6]);
  assign and_156_m1c = mux_386_nl & and_dcpl_29 & (fsm_output[5]) & (~ (fsm_output[3]));
  assign nor_380_cse = ~((fsm_output[6]) | (fsm_output[8]));
  assign nor_246_cse = ~((~ (fsm_output[5])) | (fsm_output[8]));
  assign nor_353_cse = ~((fsm_output[3]) | (fsm_output[8]));
  assign and_337_nl = (fsm_output[3]) & (fsm_output[8]);
  assign mux_66_cse = MUX_s_1_2_2(nor_353_cse, and_337_nl, and_281_cse);
  assign and_333_cse = (fsm_output[2]) & (fsm_output[0]) & (fsm_output[1]) & (fsm_output[5])
      & (fsm_output[4]);
  assign and_332_cse = (fsm_output[2]) & (fsm_output[0]);
  assign or_625_cse = (fsm_output[5:4]!=2'b10);
  assign or_92_cse = (fsm_output[5]) | (fsm_output[8]);
  assign or_585_cse = (fsm_output[3:2]!=2'b00);
  assign or_481_cse = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[8]);
  assign or_589_cse = and_206_cse | (fsm_output[3]);
  assign and_190_nl = (fsm_output[4]) & nor_tmp_24;
  assign or_506_nl = (or_319_cse & (fsm_output[3])) | (fsm_output[8]);
  assign mux_560_nl = MUX_s_1_2_2((fsm_output[8]), or_506_nl, fsm_output[4]);
  assign mux_561_cse = MUX_s_1_2_2(and_190_nl, mux_560_nl, fsm_output[5]);
  assign and_215_nl = or_585_cse & (fsm_output[8]);
  assign mux_555_nl = MUX_s_1_2_2(nor_tmp_24, and_215_nl, fsm_output[0]);
  assign mux_556_nl = MUX_s_1_2_2(mux_555_nl, (fsm_output[8]), fsm_output[4]);
  assign mux_529_nl = MUX_s_1_2_2(mux_66_cse, (fsm_output[8]), fsm_output[4]);
  assign mux_557_nl = MUX_s_1_2_2((~ mux_556_nl), mux_529_nl, fsm_output[5]);
  assign or_465_nl = (fsm_output[2]) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[3])
      | (fsm_output[8]);
  assign mux_525_nl = MUX_s_1_2_2((fsm_output[8]), or_465_nl, fsm_output[4]);
  assign or_500_nl = (fsm_output[5]) | mux_525_nl;
  assign mux_558_cse = MUX_s_1_2_2(mux_557_nl, or_500_nl, fsm_output[6]);
  assign COMP_LOOP_or_2_cse = and_dcpl_49 | and_dcpl_65 | and_dcpl_72 | and_dcpl_75;
  assign nl_STAGE_LOOP_i_3_0_sva_2 = STAGE_LOOP_i_3_0_sva + 4'b0001;
  assign STAGE_LOOP_i_3_0_sva_2 = nl_STAGE_LOOP_i_3_0_sva_2[3:0];
  assign nl_COMP_LOOP_acc_psp_sva_1 = (VEC_LOOP_j_sva_11_0[11:2]) + conv_u2u_7_10(COMP_LOOP_k_9_2_sva_6_0);
  assign COMP_LOOP_acc_psp_sva_1 = nl_COMP_LOOP_acc_psp_sva_1[9:0];
  assign or_641_cse = (fsm_output[8]) | (fsm_output[6]) | (fsm_output[1]) | (~ (fsm_output[5]))
      | (~ (fsm_output[7])) | (fsm_output[0]) | (fsm_output[4]);
  assign nl_modulo_qr_sva_1_mx0w1 = modulo_result_rem_cmp_z + p_sva;
  assign modulo_qr_sva_1_mx0w1 = nl_modulo_qr_sva_1_mx0w1[63:0];
  assign nl_COMP_LOOP_1_acc_5_mut_mx0w7 = operator_64_false_acc_mut_63_0 + modulo_result_mux_1_cse;
  assign COMP_LOOP_1_acc_5_mut_mx0w7 = nl_COMP_LOOP_1_acc_5_mut_mx0w7[63:0];
  assign nl_COMP_LOOP_1_modExp_1_while_if_mul_mut_1 = $signed(COMP_LOOP_1_acc_5_mut)
      * $signed(COMP_LOOP_1_acc_8_itm);
  assign COMP_LOOP_1_modExp_1_while_if_mul_mut_1 = nl_COMP_LOOP_1_modExp_1_while_if_mul_mut_1[63:0];
  assign operator_64_false_slc_modExp_exp_63_1_3 = MUX_v_63_2_2((operator_66_true_div_cmp_z[63:1]),
      (COMP_LOOP_1_acc_5_mut[63:1]), and_dcpl_139);
  assign modExp_while_and_3 = (~ (modulo_result_rem_cmp_z[63])) & modExp_exp_1_0_1_sva;
  assign modExp_while_and_5 = (modulo_result_rem_cmp_z[63]) & modExp_exp_1_0_1_sva;
  assign and_dcpl_1 = (fsm_output[2]) & (~ (fsm_output[6])) & (~ (fsm_output[3]));
  assign nor_tmp_16 = (fsm_output[8:7]==2'b11);
  assign or_40_nl = (fsm_output[5:4]!=2'b00) | (~ nor_tmp_16);
  assign or_38_nl = (~ (fsm_output[5])) | (fsm_output[4]) | (~ (fsm_output[7])) |
      (fsm_output[8]);
  assign mux_tmp_41 = MUX_s_1_2_2(or_40_nl, or_38_nl, fsm_output[1]);
  assign nor_tmp_24 = or_589_cse & (fsm_output[8]);
  assign or_tmp_70 = (fsm_output[8:7]!=2'b00);
  assign mux_tmp_86 = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[8]);
  assign nor_tmp_63 = (fsm_output[8:4]==5'b11111);
  assign nor_338_nl = ~((fsm_output[2]) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[5])
      | (fsm_output[4]) | (fsm_output[8]) | (fsm_output[7]));
  assign and_30_nl = (fsm_output[2]) & or_644_cse & (fsm_output[5]) & (fsm_output[4])
      & (fsm_output[8]) & (fsm_output[7]);
  assign mux_138_nl = MUX_s_1_2_2(nor_338_nl, and_30_nl, fsm_output[6]);
  assign mux_139_itm = MUX_s_1_2_2(mux_138_nl, nor_tmp_63, fsm_output[3]);
  assign and_dcpl_25 = ~((fsm_output[6]) | (fsm_output[3]));
  assign and_dcpl_26 = ~((fsm_output[0]) | (fsm_output[2]));
  assign and_dcpl_27 = and_dcpl_26 & and_dcpl_25;
  assign and_dcpl_28 = ~((fsm_output[5]) | (fsm_output[1]));
  assign and_dcpl_29 = ~((fsm_output[8:7]!=2'b00));
  assign and_dcpl_30 = and_dcpl_29 & (~ (fsm_output[4]));
  assign and_dcpl_31 = and_dcpl_30 & and_dcpl_28;
  assign and_dcpl_33 = (fsm_output[6]) & (~ (fsm_output[3]));
  assign and_dcpl_34 = (~ (fsm_output[0])) & (fsm_output[2]);
  assign and_dcpl_36 = (fsm_output[5]) & (~ (fsm_output[1]));
  assign and_dcpl_38 = nor_tmp_16 & (fsm_output[4]);
  assign and_dcpl_39 = and_dcpl_38 & and_dcpl_36;
  assign and_dcpl_42 = (fsm_output[5]) & (fsm_output[1]);
  assign and_dcpl_43 = and_dcpl_29 & (fsm_output[4]);
  assign and_dcpl_44 = and_dcpl_43 & and_dcpl_42;
  assign and_dcpl_45 = and_dcpl_44 & and_dcpl_34 & and_dcpl_25;
  assign and_dcpl_46 = (fsm_output[0]) & (~ (fsm_output[2]));
  assign and_dcpl_47 = and_dcpl_46 & and_dcpl_33;
  assign and_dcpl_48 = and_dcpl_30 & and_dcpl_42;
  assign and_dcpl_49 = and_dcpl_48 & and_dcpl_47;
  assign and_dcpl_50 = (~ (fsm_output[6])) & (fsm_output[3]);
  assign and_dcpl_53 = (~ (fsm_output[5])) & (fsm_output[1]);
  assign and_dcpl_54 = (fsm_output[8:7]==2'b01);
  assign and_dcpl_62 = and_dcpl_26 & and_dcpl_33;
  assign and_dcpl_65 = and_dcpl_54 & (fsm_output[4]) & and_dcpl_53 & and_dcpl_62;
  assign and_dcpl_67 = (fsm_output[8:7]==2'b10);
  assign and_dcpl_72 = and_dcpl_67 & (~ (fsm_output[4])) & and_dcpl_28 & and_dcpl_47;
  assign and_dcpl_75 = and_dcpl_39 & and_dcpl_27;
  assign nand_79_cse = ~((fsm_output[8:7]==2'b11));
  assign and_dcpl_85 = and_dcpl_30 & and_dcpl_53;
  assign and_dcpl_86 = and_dcpl_85 & and_dcpl_46 & and_dcpl_50;
  assign and_dcpl_88 = ~((fsm_output[6:5]!=2'b00));
  assign and_dcpl_89 = and_dcpl_29 & and_dcpl_88;
  assign and_dcpl_91 = (fsm_output[6:5]==2'b01);
  assign not_tmp_154 = ~(or_319_cse & (fsm_output[5:4]==2'b11));
  assign or_tmp_254 = (fsm_output[6:4]!=3'b100);
  assign or_tmp_256 = (fsm_output[5:4]!=2'b01);
  assign mux_tmp_212 = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), fsm_output[5]);
  assign or_611_nl = and_206_cse | (fsm_output[4]);
  assign nand_61_nl = ~(or_287_cse & (fsm_output[4]));
  assign not_tmp_158 = MUX_s_1_2_2(or_611_nl, nand_61_nl, fsm_output[3]);
  assign or_tmp_262 = (fsm_output[2]) | (~ (fsm_output[3])) | (~ (fsm_output[5]))
      | (fsm_output[8]);
  assign or_295_nl = (fsm_output[2]) | (~ (fsm_output[3])) | (fsm_output[5]) | (~
      (fsm_output[8]));
  assign mux_217_nl = MUX_s_1_2_2(or_295_nl, or_tmp_262, fsm_output[1]);
  assign nor_336_nl = ~((~ (fsm_output[4])) | (fsm_output[7]) | mux_217_nl);
  assign or_291_nl = (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[5]) | (~
      (fsm_output[8]));
  assign mux_216_nl = MUX_s_1_2_2(or_tmp_262, or_291_nl, fsm_output[1]);
  assign nor_337_nl = ~((fsm_output[4]) | (~ (fsm_output[7])) | mux_216_nl);
  assign mux_218_nl = MUX_s_1_2_2(nor_336_nl, nor_337_nl, fsm_output[0]);
  assign and_dcpl_102 = mux_218_nl & (fsm_output[6]);
  assign mux_tmp_230 = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), fsm_output[7]);
  assign or_tmp_275 = (fsm_output[8:7]!=2'b10);
  assign or_tmp_277 = (fsm_output[8:7]!=2'b01);
  assign mux_238_nl = MUX_s_1_2_2(or_tmp_275, or_tmp_277, fsm_output[4]);
  assign or_309_nl = (fsm_output[5]) | mux_238_nl;
  assign mux_237_nl = MUX_s_1_2_2(nand_79_cse, or_tmp_275, fsm_output[4]);
  assign nand_25_nl = ~((fsm_output[5]) & (~ mux_237_nl));
  assign mux_tmp_239 = MUX_s_1_2_2(or_309_nl, nand_25_nl, fsm_output[6]);
  assign or_tmp_288 = (~ (fsm_output[1])) | (fsm_output[5]) | (~ (fsm_output[4]))
      | (~ (fsm_output[8])) | (fsm_output[7]);
  assign mux_249_nl = MUX_s_1_2_2(or_tmp_288, mux_tmp_41, fsm_output[0]);
  assign and_dcpl_105 = (~ mux_249_nl) & and_dcpl_1;
  assign and_dcpl_111 = and_dcpl_67 & (~ (fsm_output[6]));
  assign and_dcpl_122 = nor_tmp_16 & (~ (fsm_output[6]));
  assign and_dcpl_128 = ~((~(or_287_cse ^ (fsm_output[3]))) | (fsm_output[7]) | (fsm_output[8])
      | (fsm_output[4]) | (~ and_dcpl_88));
  assign and_277_nl = (fsm_output[2:0]==3'b101) & and_273_cse;
  assign nor_271_nl = ~((fsm_output[2]) | (fsm_output[0]) | (~ (fsm_output[1])) |
      (fsm_output[5]) | (fsm_output[4]));
  assign mux_271_nl = MUX_s_1_2_2(and_277_nl, nor_271_nl, fsm_output[3]);
  assign and_dcpl_132 = mux_271_nl & and_dcpl_29 & (~ (fsm_output[6]));
  assign or_tmp_300 = (fsm_output[4]) | (fsm_output[8]) | (fsm_output[7]);
  assign mux_tmp_272 = MUX_s_1_2_2(nor_tmp_16, (fsm_output[8]), fsm_output[4]);
  assign mux_tmp_273 = MUX_s_1_2_2(mux_tmp_272, or_tmp_300, fsm_output[5]);
  assign mux_tmp_274 = MUX_s_1_2_2(mux_tmp_272, or_tmp_70, fsm_output[5]);
  assign mux_tmp_276 = MUX_s_1_2_2((fsm_output[8]), or_tmp_70, fsm_output[4]);
  assign mux_277_nl = MUX_s_1_2_2(mux_tmp_272, mux_tmp_276, fsm_output[5]);
  assign mux_tmp_278 = MUX_s_1_2_2(mux_277_nl, mux_tmp_273, fsm_output[1]);
  assign mux_tmp_282 = MUX_s_1_2_2(nor_tmp_16, mux_tmp_276, fsm_output[5]);
  assign mux_tmp_283 = MUX_s_1_2_2(and_dcpl_38, mux_tmp_276, fsm_output[5]);
  assign nor_tmp_120 = (fsm_output[5]) & (fsm_output[8]);
  assign mux_tmp_303 = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), fsm_output[5]);
  assign nor_263_nl = ~((fsm_output[2]) | and_289_cse | (fsm_output[5]) | (fsm_output[4])
      | (fsm_output[8]) | (fsm_output[7]));
  assign and_358_nl = (fsm_output[5]) & (fsm_output[4]) & (fsm_output[7]) & (fsm_output[8]);
  assign mux_tmp_321 = MUX_s_1_2_2(nor_263_nl, and_358_nl, fsm_output[6]);
  assign and_dcpl_137 = and_332_cse & and_dcpl_25;
  assign and_dcpl_138 = and_dcpl_43 & and_dcpl_36;
  assign and_dcpl_139 = and_dcpl_138 & and_dcpl_137;
  assign mux_328_nl = MUX_s_1_2_2(mux_tmp_86, or_tmp_277, fsm_output[6]);
  assign mux_326_nl = MUX_s_1_2_2(nor_tmp_16, or_tmp_70, fsm_output[6]);
  assign mux_tmp_329 = MUX_s_1_2_2(mux_328_nl, mux_326_nl, fsm_output[3]);
  assign mux_tmp_330 = MUX_s_1_2_2(nor_tmp_16, or_tmp_277, fsm_output[6]);
  assign and_tmp_8 = (fsm_output[6]) & or_tmp_275;
  assign and_tmp_9 = (fsm_output[6]) & or_tmp_277;
  assign mux_332_nl = MUX_s_1_2_2((~ or_tmp_277), or_tmp_275, fsm_output[6]);
  assign mux_tmp_333 = MUX_s_1_2_2(mux_332_nl, and_tmp_9, fsm_output[3]);
  assign mux_tmp_336 = MUX_s_1_2_2((~ or_tmp_277), (fsm_output[7]), fsm_output[6]);
  assign mux_tmp_337 = MUX_s_1_2_2(or_tmp_277, mux_tmp_86, fsm_output[6]);
  assign mux_tmp_339 = MUX_s_1_2_2(mux_tmp_86, or_tmp_275, fsm_output[6]);
  assign not_tmp_221 = MUX_s_1_2_2((fsm_output[7]), (~ (fsm_output[8])), fsm_output[6]);
  assign mux_tmp_344 = MUX_s_1_2_2(nor_tmp_16, (fsm_output[8]), fsm_output[6]);
  assign mux_351_itm = MUX_s_1_2_2(or_tmp_277, (fsm_output[8]), fsm_output[6]);
  assign mux_tmp_352 = MUX_s_1_2_2((~ mux_351_itm), or_tmp_275, fsm_output[3]);
  assign or_tmp_331 = (~((~ (fsm_output[6])) | (fsm_output[8]))) | (fsm_output[7]);
  assign mux_353_nl = MUX_s_1_2_2(or_tmp_277, nor_tmp_16, fsm_output[6]);
  assign mux_tmp_354 = MUX_s_1_2_2((~ mux_353_nl), or_tmp_331, fsm_output[3]);
  assign or_36_nl = (fsm_output[5]) | (~ (fsm_output[4])) | (fsm_output[7]) | (~
      (fsm_output[8]));
  assign or_34_nl = (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[7]) |
      (fsm_output[8]);
  assign mux_38_nl = MUX_s_1_2_2(or_36_nl, or_34_nl, fsm_output[1]);
  assign mux_43_nl = MUX_s_1_2_2(mux_tmp_41, mux_38_nl, fsm_output[0]);
  assign and_dcpl_140 = (~ mux_43_nl) & and_dcpl_1;
  assign or_375_nl = (~ (fsm_output[8])) | (fsm_output[4]) | (fsm_output[7]) | (fsm_output[1])
      | (fsm_output[5]) | (~ (fsm_output[6]));
  assign or_373_nl = (fsm_output[8]) | (~ (fsm_output[4])) | (~ (fsm_output[7]))
      | (fsm_output[1]) | (fsm_output[5]) | (~ (fsm_output[6]));
  assign mux_384_nl = MUX_s_1_2_2(or_375_nl, or_373_nl, fsm_output[0]);
  assign nor_256_nl = ~((fsm_output[3]) | mux_384_nl);
  assign nor_257_nl = ~((fsm_output[4]) | (fsm_output[7]) | (fsm_output[1]) | (fsm_output[5])
      | (~ (fsm_output[6])));
  assign nor_258_nl = ~((fsm_output[4]) | (~ (fsm_output[7])) | (~ (fsm_output[1]))
      | (~ (fsm_output[5])) | (fsm_output[6]));
  assign mux_383_nl = MUX_s_1_2_2(nor_257_nl, nor_258_nl, fsm_output[8]);
  assign and_257_nl = (fsm_output[3]) & (fsm_output[0]) & mux_383_nl;
  assign not_tmp_235 = MUX_s_1_2_2(nor_256_nl, and_257_nl, fsm_output[2]);
  assign and_dcpl_141 = and_dcpl_26 & and_dcpl_50;
  assign not_tmp_239 = ~((fsm_output[0]) & (fsm_output[4]) & (fsm_output[7]));
  assign nor_250_nl = ~((~ (fsm_output[8])) | (fsm_output[2]) | not_tmp_239);
  assign nor_251_nl = ~((fsm_output[8]) | (~ (fsm_output[2])) | (fsm_output[0]) |
      (fsm_output[4]) | (fsm_output[7]));
  assign mux_388_nl = MUX_s_1_2_2(nor_250_nl, nor_251_nl, fsm_output[6]);
  assign and_255_nl = (fsm_output[5]) & mux_388_nl;
  assign nor_252_nl = ~((fsm_output[2]) | not_tmp_239);
  assign nor_253_nl = ~((fsm_output[2]) | (fsm_output[0]) | (fsm_output[4]) | (fsm_output[7]));
  assign mux_387_nl = MUX_s_1_2_2(nor_252_nl, nor_253_nl, fsm_output[8]);
  assign and_256_nl = (~((fsm_output[6:5]!=2'b10))) & mux_387_nl;
  assign not_tmp_242 = MUX_s_1_2_2(and_255_nl, and_256_nl, fsm_output[1]);
  assign mux_391_itm = MUX_s_1_2_2((fsm_output[7]), (fsm_output[8]), fsm_output[4]);
  assign mux_390_nl = MUX_s_1_2_2(and_dcpl_29, nor_tmp_16, fsm_output[4]);
  assign mux_tmp_392 = MUX_s_1_2_2((~ mux_391_itm), mux_390_nl, fsm_output[5]);
  assign mux_tmp_397 = MUX_s_1_2_2(and_dcpl_29, mux_tmp_86, fsm_output[4]);
  assign not_tmp_246 = MUX_s_1_2_2(mux_tmp_86, (~ (fsm_output[7])), fsm_output[4]);
  assign mux_tmp_404 = MUX_s_1_2_2(not_tmp_246, mux_93_cse, fsm_output[5]);
  assign mux_tmp_408 = MUX_s_1_2_2((~ nor_tmp_16), or_tmp_275, fsm_output[4]);
  assign mux_tmp_409 = MUX_s_1_2_2((~ nor_tmp_16), (fsm_output[7]), fsm_output[4]);
  assign mux_tmp_411 = MUX_s_1_2_2(mux_tmp_86, or_tmp_277, fsm_output[4]);
  assign mux_tmp_412 = MUX_s_1_2_2(mux_tmp_411, mux_tmp_408, fsm_output[5]);
  assign mux_419_nl = MUX_s_1_2_2(and_dcpl_54, nor_tmp_16, fsm_output[4]);
  assign mux_tmp_420 = MUX_s_1_2_2((~ mux_419_nl), mux_93_cse, fsm_output[5]);
  assign mux_tmp_427 = MUX_s_1_2_2((~ (fsm_output[7])), or_tmp_275, fsm_output[4]);
  assign mux_tmp_428 = MUX_s_1_2_2(mux_tmp_411, mux_tmp_427, fsm_output[5]);
  assign nor_247_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (~ and_dcpl_38));
  assign nor_248_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[5])) | (fsm_output[4])
      | (~ (fsm_output[8])) | (fsm_output[7]));
  assign mux_443_nl = MUX_s_1_2_2(nor_247_nl, nor_248_nl, fsm_output[0]);
  assign nor_249_nl = ~((fsm_output[0]) | (fsm_output[1]) | (~ (fsm_output[5])) |
      (~ (fsm_output[4])) | (fsm_output[8]) | (~ (fsm_output[7])));
  assign not_tmp_253 = MUX_s_1_2_2(mux_443_nl, nor_249_nl, fsm_output[2]);
  assign or_tmp_382 = (fsm_output[7]) | nor_246_cse;
  assign and_176_nl = (fsm_output[7]) & mux_tmp_303;
  assign mux_tmp_462 = MUX_s_1_2_2(and_176_nl, or_tmp_382, fsm_output[6]);
  assign mux_tmp_463 = MUX_s_1_2_2(nor_246_cse, or_92_cse, fsm_output[7]);
  assign mux_464_nl = MUX_s_1_2_2(mux_tmp_303, or_92_cse, fsm_output[7]);
  assign mux_465_nl = MUX_s_1_2_2((~ mux_464_nl), mux_tmp_463, fsm_output[6]);
  assign mux_tmp_466 = MUX_s_1_2_2(mux_465_nl, mux_tmp_462, fsm_output[4]);
  assign mux_467_nl = MUX_s_1_2_2(nor_tmp_120, or_92_cse, fsm_output[7]);
  assign mux_468_nl = MUX_s_1_2_2((~ mux_467_nl), mux_tmp_463, fsm_output[6]);
  assign mux_tmp_469 = MUX_s_1_2_2(mux_468_nl, mux_tmp_462, fsm_output[4]);
  assign not_tmp_265 = ~(((fsm_output[7]) | (fsm_output[5])) & (fsm_output[8]));
  assign mux_470_nl = MUX_s_1_2_2(not_tmp_265, mux_tmp_463, fsm_output[6]);
  assign mux_tmp_471 = MUX_s_1_2_2(mux_470_nl, mux_tmp_462, fsm_output[4]);
  assign mux_tmp_473 = MUX_s_1_2_2((~ mux_tmp_303), mux_tmp_303, fsm_output[7]);
  assign mux_tmp_474 = MUX_s_1_2_2(mux_tmp_473, or_tmp_382, fsm_output[6]);
  assign mux_475_nl = MUX_s_1_2_2((~ nor_tmp_120), mux_tmp_463, fsm_output[6]);
  assign mux_tmp_476 = MUX_s_1_2_2(mux_475_nl, mux_tmp_474, fsm_output[4]);
  assign and_177_nl = (fsm_output[7]) & or_92_cse;
  assign mux_tmp_481 = MUX_s_1_2_2(not_tmp_265, and_177_nl, fsm_output[6]);
  assign and_dcpl_166 = and_dcpl_138 & and_dcpl_141;
  assign or_dcpl_35 = (fsm_output[6]) | (~ (fsm_output[3]));
  assign or_dcpl_36 = (fsm_output[0]) | (~ (fsm_output[2]));
  assign or_dcpl_38 = (fsm_output[5]) | (fsm_output[1]);
  assign or_dcpl_41 = (fsm_output[6]) | (fsm_output[3]);
  assign or_dcpl_42 = or_dcpl_36 | or_dcpl_41;
  assign or_dcpl_43 = ~((fsm_output[5]) & (fsm_output[1]));
  assign mux_tmp_495 = MUX_s_1_2_2(nor_tmp_16, (fsm_output[8]), and_273_cse);
  assign nor_tmp_162 = (fsm_output[5]) & (fsm_output[8]) & (fsm_output[7]);
  assign and_dcpl_168 = and_dcpl_44 & and_dcpl_137;
  assign or_450_nl = (~ (fsm_output[8])) | (fsm_output[0]) | (fsm_output[7]);
  assign or_449_nl = (fsm_output[8]) | (~((fsm_output[0]) & (fsm_output[7])));
  assign mux_508_nl = MUX_s_1_2_2(or_450_nl, or_449_nl, fsm_output[4]);
  assign nor_237_nl = ~((fsm_output[5]) | (~ (fsm_output[6])) | (fsm_output[1]) |
      (fsm_output[2]) | mux_508_nl);
  assign or_446_nl = (fsm_output[2]) | (~ (fsm_output[4])) | (fsm_output[8]) | (fsm_output[0])
      | (fsm_output[7]);
  assign or_445_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (~((fsm_output[8]) &
      (fsm_output[0]) & (fsm_output[7])));
  assign mux_507_nl = MUX_s_1_2_2(or_446_nl, or_445_nl, fsm_output[1]);
  assign nor_238_nl = ~((fsm_output[6:5]!=2'b01) | mux_507_nl);
  assign not_tmp_279 = MUX_s_1_2_2(nor_237_nl, nor_238_nl, fsm_output[3]);
  assign or_458_nl = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[8]);
  assign mux_517_nl = MUX_s_1_2_2(or_458_nl, or_481_cse, fsm_output[0]);
  assign or_459_nl = (fsm_output[4]) | mux_517_nl;
  assign mux_518_nl = MUX_s_1_2_2((fsm_output[8]), or_459_nl, fsm_output[5]);
  assign mux_521_nl = MUX_s_1_2_2((~ mux_561_cse), mux_518_nl, fsm_output[6]);
  assign mux_522_itm = MUX_s_1_2_2(mux_521_nl, mux_558_cse, fsm_output[7]);
  assign or_32_nl = (fsm_output[1]) | (fsm_output[5]) | (~ (fsm_output[4])) | (fsm_output[7])
      | (~ (fsm_output[8]));
  assign mux_42_nl = MUX_s_1_2_2(mux_tmp_41, or_32_nl, fsm_output[0]);
  assign and_dcpl_169 = (~ mux_42_nl) & and_dcpl_1;
  assign and_323_cse = (fsm_output[4]) & (fsm_output[7]);
  assign or_dcpl_47 = (~ (fsm_output[0])) | (fsm_output[2]);
  assign or_dcpl_53 = (~ (fsm_output[6])) | (fsm_output[3]);
  assign or_dcpl_54 = ~((fsm_output[0]) & (fsm_output[2]));
  assign or_dcpl_59 = or_dcpl_54 | or_dcpl_41;
  assign STAGE_LOOP_i_3_0_sva_mx0c1 = and_dcpl_39 & and_dcpl_34 & and_dcpl_33;
  assign VEC_LOOP_j_sva_11_0_mx0c1 = and_dcpl_38 & and_dcpl_42 & and_dcpl_47;
  assign nor_262_nl = ~((fsm_output[5]) | (fsm_output[4]) | (fsm_output[8]) | (fsm_output[7]));
  assign mux_322_nl = MUX_s_1_2_2(nor_262_nl, and_313_cse, fsm_output[6]);
  assign modExp_result_sva_mx0c0 = MUX_s_1_2_2(mux_322_nl, mux_tmp_321, fsm_output[3]);
  assign nl_STAGE_LOOP_acc_nl = (STAGE_LOOP_i_3_0_sva_2[3:1]) + 3'b011;
  assign STAGE_LOOP_acc_nl = nl_STAGE_LOOP_acc_nl[2:0];
  assign STAGE_LOOP_acc_itm_2_1 = readslicef_3_1_2(STAGE_LOOP_acc_nl);
  assign and_198_m1c = and_dcpl_67 & (fsm_output[4]) & and_dcpl_28 & and_dcpl_137;
  assign and_63_nl = and_dcpl_54 & (~ (fsm_output[4])) & and_dcpl_53 & and_332_cse
      & and_dcpl_50;
  assign nand_82_nl = ~((fsm_output[0]) & (fsm_output[4]));
  assign or_137_nl = (fsm_output[0]) | (fsm_output[4]);
  assign mux_141_nl = MUX_s_1_2_2(nand_82_nl, or_137_nl, fsm_output[7]);
  assign nor_332_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | mux_141_nl);
  assign nor_333_nl = ~((fsm_output[1]) | (~((fsm_output[5]) & (fsm_output[7]) &
      (fsm_output[0]) & (fsm_output[4]))));
  assign mux_142_nl = MUX_s_1_2_2(nor_332_nl, nor_333_nl, fsm_output[6]);
  assign nand_112_nl = ~((fsm_output[8]) & mux_142_nl);
  assign mux_143_nl = MUX_s_1_2_2(nand_112_nl, or_641_cse, fsm_output[2]);
  assign nor_377_nl = ~(mux_143_nl | (fsm_output[3]));
  assign nor_330_nl = ~((fsm_output[6]) | (~ (fsm_output[0])) | (fsm_output[1]) |
      (fsm_output[4]));
  assign nor_331_nl = ~((~ (fsm_output[6])) | (fsm_output[0]) | (~((fsm_output[1])
      & (fsm_output[4]))));
  assign mux_144_nl = MUX_s_1_2_2(nor_330_nl, nor_331_nl, fsm_output[3]);
  assign and_67_nl = mux_144_nl & and_dcpl_54 & (fsm_output[5]) & (fsm_output[2]);
  assign nor_329_nl = ~((fsm_output[6]) | (fsm_output[0]) | (fsm_output[5]) | (~
      (fsm_output[4])));
  assign and_308_nl = (fsm_output[6]) & (fsm_output[0]) & (fsm_output[5]) & (~ (fsm_output[4]));
  assign mux_145_nl = MUX_s_1_2_2(nor_329_nl, and_308_nl, fsm_output[3]);
  assign and_75_nl = mux_145_nl & and_dcpl_67 & (fsm_output[2:1]==2'b10);
  assign nor_327_nl = ~((fsm_output[6]) | (fsm_output[2]) | (~ (fsm_output[0])) |
      (~ (fsm_output[1])) | (fsm_output[4]));
  assign nor_328_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[2])) | (fsm_output[0])
      | (fsm_output[1]) | (~ (fsm_output[4])));
  assign mux_146_nl = MUX_s_1_2_2(nor_327_nl, nor_328_nl, fsm_output[3]);
  assign and_80_nl = mux_146_nl & nor_tmp_16 & (~ (fsm_output[5]));
  assign vec_rsc_0_0_i_adra_d_pff = MUX1HOT_v_10_7_2(COMP_LOOP_acc_psp_sva_1, (z_out_5[12:3]),
      COMP_LOOP_acc_psp_sva, (COMP_LOOP_acc_10_cse_12_1_1_sva[11:2]), (COMP_LOOP_acc_1_cse_2_sva[11:2]),
      (COMP_LOOP_acc_11_psp_sva[10:1]), (COMP_LOOP_acc_1_cse_sva[11:2]), {and_dcpl_45
      , COMP_LOOP_or_2_cse , and_63_nl , nor_377_nl , and_67_nl , and_75_nl , and_80_nl});
  assign vec_rsc_0_0_i_da_d_pff = modulo_result_mux_1_cse;
  assign nor_322_nl = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b00) | mux_152_cse);
  assign or_156_nl = (~ (fsm_output[1])) | (VEC_LOOP_j_sva_11_0[1]) | (fsm_output[8:6]!=3'b010);
  assign or_154_nl = (fsm_output[1]) | (~ (fsm_output[6])) | (COMP_LOOP_acc_11_psp_sva[0])
      | (fsm_output[8:7]!=2'b10);
  assign mux_148_nl = MUX_s_1_2_2(or_156_nl, or_154_nl, fsm_output[5]);
  assign nor_325_nl = ~((~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0]) | mux_148_nl);
  assign or_151_nl = (fsm_output[1]) | (COMP_LOOP_acc_1_cse_sva[1:0]!=2'b00) | nand_53_cse;
  assign or_149_nl = (~ (fsm_output[1])) | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b00)
      | (fsm_output[8:7]!=2'b01);
  assign mux_147_nl = MUX_s_1_2_2(or_151_nl, or_149_nl, fsm_output[5]);
  assign nor_326_nl = ~((fsm_output[0]) | mux_147_nl);
  assign mux_149_nl = MUX_s_1_2_2(nor_325_nl, nor_326_nl, fsm_output[4]);
  assign and_307_nl = (fsm_output[2]) & mux_149_nl;
  assign vec_rsc_0_0_i_wea_d_pff = MUX_s_1_2_2(nor_322_nl, and_307_nl, fsm_output[3]);
  assign nor_317_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[6])) | (z_out_5[2:1]!=2'b00)
      | (fsm_output[8:7]!=2'b01));
  assign nor_318_nl = ~((fsm_output[1]) | (fsm_output[6]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_11_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[8:7]!=2'b10));
  assign mux_158_nl = MUX_s_1_2_2(nor_317_nl, nor_318_nl, fsm_output[2]);
  assign nor_319_nl = ~((fsm_output[1]) | (z_out_5[2:1]!=2'b00) | (fsm_output[6])
      | nand_79_cse);
  assign nor_320_nl = ~((~ (fsm_output[1])) | (fsm_output[6]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (fsm_output[8:7]!=2'b00));
  assign mux_157_nl = MUX_s_1_2_2(nor_319_nl, nor_320_nl, fsm_output[2]);
  assign mux_159_nl = MUX_s_1_2_2(mux_158_nl, mux_157_nl, fsm_output[5]);
  assign nand_111_nl = ~((fsm_output[4]) & mux_159_nl);
  assign or_171_nl = (~ (fsm_output[6])) | (z_out_5[2:1]!=2'b00) | (fsm_output[8:7]!=2'b10);
  assign or_170_nl = (~ modExp_exp_1_0_1_sva) | (COMP_LOOP_acc_1_cse_sva[1:0]!=2'b00)
      | (fsm_output[6]) | nand_79_cse;
  assign mux_155_nl = MUX_s_1_2_2(or_171_nl, or_170_nl, fsm_output[1]);
  assign or_172_nl = (fsm_output[2]) | mux_155_nl;
  assign or_168_nl = (~ (fsm_output[1])) | (~ (fsm_output[6])) | (z_out_5[2:1]!=2'b00)
      | (fsm_output[8:7]!=2'b00);
  assign or_167_nl = (fsm_output[1]) | (fsm_output[6]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b00) | (fsm_output[8:7]!=2'b01);
  assign mux_154_nl = MUX_s_1_2_2(or_168_nl, or_167_nl, fsm_output[2]);
  assign mux_156_nl = MUX_s_1_2_2(or_172_nl, mux_154_nl, fsm_output[5]);
  assign or_640_nl = (fsm_output[4]) | mux_156_nl;
  assign mux_160_nl = MUX_s_1_2_2(nand_111_nl, or_640_nl, fsm_output[0]);
  assign vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~(mux_160_nl | (fsm_output[3]));
  assign nor_311_nl = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b01) | mux_152_cse);
  assign nor_314_nl = ~((~ (fsm_output[1])) | (VEC_LOOP_j_sva_11_0[1]) | (fsm_output[8:6]!=3'b010));
  assign nor_315_nl = ~((fsm_output[1]) | (~ (fsm_output[6])) | (COMP_LOOP_acc_11_psp_sva[0])
      | (fsm_output[8:7]!=2'b10));
  assign mux_162_nl = MUX_s_1_2_2(nor_314_nl, nor_315_nl, fsm_output[5]);
  assign and_305_nl = (fsm_output[0]) & (VEC_LOOP_j_sva_11_0[0]) & mux_162_nl;
  assign or_183_nl = (fsm_output[1]) | (COMP_LOOP_acc_1_cse_sva[1:0]!=2'b01) | nand_53_cse;
  assign or_181_nl = (~ (fsm_output[1])) | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b01)
      | (fsm_output[8:7]!=2'b01);
  assign mux_161_nl = MUX_s_1_2_2(or_183_nl, or_181_nl, fsm_output[5]);
  assign nor_316_nl = ~((fsm_output[0]) | mux_161_nl);
  assign mux_163_nl = MUX_s_1_2_2(and_305_nl, nor_316_nl, fsm_output[4]);
  assign and_304_nl = (fsm_output[2]) & mux_163_nl;
  assign vec_rsc_0_1_i_wea_d_pff = MUX_s_1_2_2(nor_311_nl, and_304_nl, fsm_output[3]);
  assign nor_306_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[6])) | (z_out_5[2:1]!=2'b01)
      | (fsm_output[8:7]!=2'b01));
  assign nor_307_nl = ~((fsm_output[1]) | (fsm_output[6]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_11_psp_sva[0]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[8:7]!=2'b10));
  assign mux_172_nl = MUX_s_1_2_2(nor_306_nl, nor_307_nl, fsm_output[2]);
  assign nor_308_nl = ~((fsm_output[1]) | (z_out_5[2:1]!=2'b01) | (fsm_output[6])
      | nand_79_cse);
  assign nor_309_nl = ~((~ (fsm_output[1])) | (fsm_output[6]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (fsm_output[8:7]!=2'b00));
  assign mux_171_nl = MUX_s_1_2_2(nor_308_nl, nor_309_nl, fsm_output[2]);
  assign mux_173_nl = MUX_s_1_2_2(mux_172_nl, mux_171_nl, fsm_output[5]);
  assign nand_110_nl = ~((fsm_output[4]) & mux_173_nl);
  assign or_201_nl = (~ (fsm_output[6])) | (z_out_5[2:1]!=2'b01) | (fsm_output[8:7]!=2'b10);
  assign or_200_nl = (~ modExp_exp_1_0_1_sva) | (COMP_LOOP_acc_1_cse_sva[1:0]!=2'b01)
      | (fsm_output[6]) | nand_79_cse;
  assign mux_169_nl = MUX_s_1_2_2(or_201_nl, or_200_nl, fsm_output[1]);
  assign or_202_nl = (fsm_output[2]) | mux_169_nl;
  assign or_198_nl = (~ (fsm_output[1])) | (~ (fsm_output[6])) | (z_out_5[2:1]!=2'b01)
      | (fsm_output[8:7]!=2'b00);
  assign or_197_nl = (fsm_output[1]) | (fsm_output[6]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b01) | (fsm_output[8:7]!=2'b01);
  assign mux_168_nl = MUX_s_1_2_2(or_198_nl, or_197_nl, fsm_output[2]);
  assign mux_170_nl = MUX_s_1_2_2(or_202_nl, mux_168_nl, fsm_output[5]);
  assign or_639_nl = (fsm_output[4]) | mux_170_nl;
  assign mux_174_nl = MUX_s_1_2_2(nand_110_nl, or_639_nl, fsm_output[0]);
  assign vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~(mux_174_nl | (fsm_output[3]));
  assign and_300_nl = (~((COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b10))) & mux_180_cse;
  assign or_218_nl = (~ (fsm_output[1])) | (~ (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[8:6]!=3'b010);
  assign or_216_nl = (fsm_output[1]) | (~ (fsm_output[6])) | (~ (COMP_LOOP_acc_11_psp_sva[0]))
      | (fsm_output[8:7]!=2'b10);
  assign mux_176_nl = MUX_s_1_2_2(or_218_nl, or_216_nl, fsm_output[5]);
  assign nor_304_nl = ~((~ (fsm_output[0])) | (VEC_LOOP_j_sva_11_0[0]) | mux_176_nl);
  assign or_213_nl = (fsm_output[1]) | (COMP_LOOP_acc_1_cse_sva[0]) | (~((COMP_LOOP_acc_1_cse_sva[1])
      & (fsm_output[8:6]==3'b111)));
  assign or_211_nl = (~ (fsm_output[1])) | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b10)
      | (fsm_output[8:7]!=2'b01);
  assign mux_175_nl = MUX_s_1_2_2(or_213_nl, or_211_nl, fsm_output[5]);
  assign nor_305_nl = ~((fsm_output[0]) | mux_175_nl);
  assign mux_177_nl = MUX_s_1_2_2(nor_304_nl, nor_305_nl, fsm_output[4]);
  assign and_302_nl = (fsm_output[2]) & mux_177_nl;
  assign vec_rsc_0_2_i_wea_d_pff = MUX_s_1_2_2(and_300_nl, and_302_nl, fsm_output[3]);
  assign nor_295_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[6])) | (z_out_5[2:1]!=2'b10)
      | (fsm_output[8:7]!=2'b01));
  assign nor_296_nl = ~((fsm_output[1]) | (fsm_output[6]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (~ (COMP_LOOP_acc_11_psp_sva[0])) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[8:7]!=2'b10));
  assign mux_186_nl = MUX_s_1_2_2(nor_295_nl, nor_296_nl, fsm_output[2]);
  assign nor_297_nl = ~((fsm_output[1]) | (z_out_5[2:1]!=2'b10) | (fsm_output[6])
      | nand_79_cse);
  assign nor_298_nl = ~((~ (fsm_output[1])) | (fsm_output[6]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10)
      | (fsm_output[8:7]!=2'b00));
  assign mux_185_nl = MUX_s_1_2_2(nor_297_nl, nor_298_nl, fsm_output[2]);
  assign mux_187_nl = MUX_s_1_2_2(mux_186_nl, mux_185_nl, fsm_output[5]);
  assign nand_109_nl = ~((fsm_output[4]) & mux_187_nl);
  assign or_231_nl = (~ (fsm_output[6])) | (z_out_5[2:1]!=2'b10) | (fsm_output[8:7]!=2'b10);
  assign or_230_nl = (~ modExp_exp_1_0_1_sva) | (COMP_LOOP_acc_1_cse_sva[1:0]!=2'b10)
      | (fsm_output[6]) | nand_79_cse;
  assign mux_183_nl = MUX_s_1_2_2(or_231_nl, or_230_nl, fsm_output[1]);
  assign or_232_nl = (fsm_output[2]) | mux_183_nl;
  assign or_228_nl = (~ (fsm_output[1])) | (~ (fsm_output[6])) | (z_out_5[2:1]!=2'b10)
      | (fsm_output[8:7]!=2'b00);
  assign or_227_nl = (fsm_output[1]) | (fsm_output[6]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b10) | (fsm_output[8:7]!=2'b01);
  assign mux_182_nl = MUX_s_1_2_2(or_228_nl, or_227_nl, fsm_output[2]);
  assign mux_184_nl = MUX_s_1_2_2(or_232_nl, mux_182_nl, fsm_output[5]);
  assign or_638_nl = (fsm_output[4]) | mux_184_nl;
  assign mux_188_nl = MUX_s_1_2_2(nand_109_nl, or_638_nl, fsm_output[0]);
  assign vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~(mux_188_nl | (fsm_output[3]));
  assign and_295_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]==2'b11) & mux_180_cse;
  assign nor_292_nl = ~((~ (fsm_output[1])) | (~ (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[8:6]!=3'b010));
  assign nor_293_nl = ~((fsm_output[1]) | (~ (fsm_output[6])) | (~ (COMP_LOOP_acc_11_psp_sva[0]))
      | (fsm_output[8:7]!=2'b10));
  assign mux_190_nl = MUX_s_1_2_2(nor_292_nl, nor_293_nl, fsm_output[5]);
  assign and_298_nl = (fsm_output[0]) & (VEC_LOOP_j_sva_11_0[0]) & mux_190_nl;
  assign or_242_nl = (fsm_output[1]) | (~((COMP_LOOP_acc_1_cse_sva[1:0]==2'b11) &
      (fsm_output[8:6]==3'b111)));
  assign nand_105_nl = ~((fsm_output[1]) & (fsm_output[6]) & (COMP_LOOP_acc_1_cse_2_sva[1:0]==2'b11)
      & (fsm_output[8:7]==2'b01));
  assign mux_189_nl = MUX_s_1_2_2(or_242_nl, nand_105_nl, fsm_output[5]);
  assign nor_294_nl = ~((fsm_output[0]) | mux_189_nl);
  assign mux_191_nl = MUX_s_1_2_2(and_298_nl, nor_294_nl, fsm_output[4]);
  assign and_297_nl = (fsm_output[2]) & mux_191_nl;
  assign vec_rsc_0_3_i_wea_d_pff = MUX_s_1_2_2(and_295_nl, and_297_nl, fsm_output[3]);
  assign and_363_nl = (fsm_output[1]) & (fsm_output[6]) & (z_out_5[2:1]==2'b11) &
      (fsm_output[8:7]==2'b01);
  assign nor_284_nl = ~((fsm_output[1]) | (fsm_output[6]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (~ (COMP_LOOP_acc_11_psp_sva[0])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[8:7]!=2'b10));
  assign mux_200_nl = MUX_s_1_2_2(and_363_nl, nor_284_nl, fsm_output[2]);
  assign nor_285_nl = ~((fsm_output[1]) | (z_out_5[2:1]!=2'b11) | (fsm_output[6])
      | nand_79_cse);
  assign nor_286_nl = ~((~ (fsm_output[1])) | (fsm_output[6]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11)
      | (fsm_output[8:7]!=2'b00));
  assign mux_199_nl = MUX_s_1_2_2(nor_285_nl, nor_286_nl, fsm_output[2]);
  assign mux_201_nl = MUX_s_1_2_2(mux_200_nl, mux_199_nl, fsm_output[5]);
  assign nand_108_nl = ~((fsm_output[4]) & mux_201_nl);
  assign nand_64_nl = ~((fsm_output[6]) & (z_out_5[2:1]==2'b11) & (fsm_output[8:7]==2'b10));
  assign or_257_nl = (~(modExp_exp_1_0_1_sva & (COMP_LOOP_acc_1_cse_sva[1:0]==2'b11)
      & (~ (fsm_output[6])))) | nand_79_cse;
  assign mux_197_nl = MUX_s_1_2_2(nand_64_nl, or_257_nl, fsm_output[1]);
  assign or_259_nl = (fsm_output[2]) | mux_197_nl;
  assign or_255_nl = (~ (fsm_output[1])) | (~ (fsm_output[6])) | (z_out_5[2:1]!=2'b11)
      | (fsm_output[8:7]!=2'b00);
  assign or_254_nl = (fsm_output[1]) | (fsm_output[6]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b11) | (fsm_output[8:7]!=2'b01);
  assign mux_196_nl = MUX_s_1_2_2(or_255_nl, or_254_nl, fsm_output[2]);
  assign mux_198_nl = MUX_s_1_2_2(or_259_nl, mux_196_nl, fsm_output[5]);
  assign or_637_nl = (fsm_output[4]) | mux_198_nl;
  assign mux_202_nl = MUX_s_1_2_2(nand_108_nl, or_637_nl, fsm_output[0]);
  assign vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d = ~(mux_202_nl | (fsm_output[3]));
  assign nor_399_cse = ~((fsm_output[7]) | (fsm_output[4]));
  assign and_dcpl_194 = (~ (fsm_output[2])) & (fsm_output[0]) & (~ (fsm_output[1]))
      & (~((fsm_output[3]) | (fsm_output[5]))) & nor_380_cse & nor_399_cse;
  assign and_dcpl_225 = (fsm_output==9'b111110011);
  assign and_dcpl_250 = (fsm_output[6:5]==2'b10);
  assign and_dcpl_257 = (~ (fsm_output[3])) & (fsm_output[8]);
  assign and_441_cse = and_dcpl_46 & (~ (fsm_output[1])) & and_dcpl_257 & and_dcpl_250
      & nor_399_cse;
  assign and_dcpl_273 = (fsm_output[2:0]==3'b110) & nor_353_cse & and_dcpl_91 & (~
      (fsm_output[7])) & (fsm_output[4]);
  assign and_dcpl_279 = and_dcpl_46 & (fsm_output[1]);
  assign and_dcpl_281 = and_dcpl_279 & (fsm_output[3]) & (~ (fsm_output[8])) & (~
      (fsm_output[5])) & (~ (fsm_output[6])) & nor_399_cse;
  assign and_dcpl_285 = and_dcpl_279 & nor_353_cse & (fsm_output[6:5]==2'b11) & nor_399_cse;
  assign and_dcpl_292 = and_dcpl_26 & (fsm_output[1]) & nor_353_cse & and_dcpl_250
      & and_323_cse;
  assign and_dcpl_301 = and_dcpl_26 & (~ (fsm_output[1])) & and_dcpl_257 & and_dcpl_91
      & and_323_cse;
  assign and_dcpl_309 = (fsm_output==9'b101000001);
  assign and_dcpl_312 = (fsm_output[7:4]==4'b0011);
  assign and_dcpl_317 = (fsm_output[2]) & (~ (fsm_output[0])) & (fsm_output[1]) &
      (~ (fsm_output[3])) & (~ (fsm_output[8])) & and_dcpl_312;
  assign nor_nl = ~((~ (fsm_output[8])) | (fsm_output[1]) | (~ (fsm_output[0])));
  assign nor_392_nl = ~((fsm_output[8]) | (~((fsm_output[1:0]==2'b11))));
  assign mux_607_nl = MUX_s_1_2_2(nor_nl, nor_392_nl, fsm_output[5]);
  assign and_nl = (fsm_output[7]) & mux_607_nl;
  assign nor_393_nl = ~((fsm_output[7]) | (fsm_output[5]) | (~ (fsm_output[8])) |
      (~ (fsm_output[1])) | (fsm_output[0]));
  assign mux_608_nl = MUX_s_1_2_2(and_nl, nor_393_nl, fsm_output[4]);
  assign and_dcpl_320 = mux_608_nl & (fsm_output[2]) & (~ (fsm_output[3])) & (~ (fsm_output[6]));
  assign and_dcpl_325 = (~ (fsm_output[2])) & (~ (fsm_output[0])) & (~ (fsm_output[1]))
      & (fsm_output[3]) & (~ (fsm_output[8])) & and_dcpl_312;
  assign not_tmp_390 = ~((fsm_output[0]) & (fsm_output[2]) & (fsm_output[7]));
  assign and_390_ssc = and_dcpl_26 & (fsm_output[1]) & (fsm_output[3]) & (~ (fsm_output[8]))
      & and_dcpl_88 & nor_399_cse;
  assign nor_tmp = (fsm_output[6]) & (fsm_output[3]);
  assign mux_tmp = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), fsm_output[6]);
  assign nor_tmp_210 = (fsm_output[1]) & (fsm_output[3]);
  assign mux_tmp_613 = MUX_s_1_2_2((~ (fsm_output[3])), nor_tmp_210, fsm_output[6]);
  assign or_tmp = (fsm_output[1]) | (fsm_output[3]);
  assign mux_tmp_616 = MUX_s_1_2_2((~ or_tmp), (fsm_output[3]), fsm_output[6]);
  assign nor_423_nl = ~((fsm_output[0]) | (~ (fsm_output[7])) | (fsm_output[3]));
  assign nor_424_nl = ~((~ (fsm_output[0])) | (fsm_output[7]) | (fsm_output[3]));
  assign not_tmp_397 = MUX_s_1_2_2(nor_423_nl, nor_424_nl, fsm_output[4]);
  assign not_tmp_400 = ~((fsm_output[5:4]==2'b11));
  assign COMP_LOOP_or_22_itm = and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301;
  assign COMP_LOOP_or_24_itm = and_dcpl_320 | and_dcpl_325;
  always @(posedge clk) begin
    if ( mux_139_itm ) begin
      p_sva <= p_rsci_idat;
      r_sva <= r_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( (and_dcpl_31 & and_dcpl_27) | STAGE_LOOP_i_3_0_sva_mx0c1 ) begin
      STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(4'b0001, STAGE_LOOP_i_3_0_sva_2, STAGE_LOOP_i_3_0_sva_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_vec_rsc_triosy_0_3_obj_ld_cse <= 1'b0;
      modExp_exp_1_0_1_sva <= 1'b0;
      modExp_exp_1_0_1_sva_1 <= 1'b0;
      modExp_exp_1_7_1_sva <= 1'b0;
      modExp_exp_1_1_1_sva <= 1'b0;
    end
    else begin
      reg_vec_rsc_triosy_0_3_obj_ld_cse <= and_dcpl_39 & and_dcpl_34 & (fsm_output[6])
          & (~ (fsm_output[3])) & (~ STAGE_LOOP_acc_itm_2_1);
      modExp_exp_1_0_1_sva <= (COMP_LOOP_mux1h_18_nl & (~(mux_445_nl & (~ (fsm_output[7]))
          & (fsm_output[4]) & and_dcpl_137))) | mux_488_nl;
      modExp_exp_1_0_1_sva_1 <= (COMP_LOOP_mux_24_nl & (~(mux_524_nl & (~ (fsm_output[8]))
          & (fsm_output[5]) & (fsm_output[1]) & (fsm_output[2]) & and_dcpl_25)))
          | mux_549_nl;
      modExp_exp_1_7_1_sva <= COMP_LOOP_mux1h_29_nl & mux_551_nl;
      modExp_exp_1_1_1_sva <= COMP_LOOP_mux1h_43_nl & (~(and_dcpl_48 & and_dcpl_62));
    end
  end
  always @(posedge clk) begin
    modulo_result_rem_cmp_a <= MUX1HOT_v_64_19_2(z_out_7, modExp_while_if_mul_mut,
        modExp_while_mul_itm, COMP_LOOP_1_modExp_1_while_if_mul_mut_1, COMP_LOOP_1_modExp_1_while_if_mul_mut,
        COMP_LOOP_1_modExp_1_while_mul_itm, COMP_LOOP_1_mul_mut, COMP_LOOP_1_acc_5_mut_mx0w7,
        COMP_LOOP_1_acc_5_mut, COMP_LOOP_1_acc_8_itm, COMP_LOOP_2_modExp_1_while_mul_mut,
        COMP_LOOP_2_modExp_1_while_if_mul_itm, COMP_LOOP_2_mul_mut, COMP_LOOP_3_modExp_1_while_mul_mut,
        COMP_LOOP_3_modExp_1_while_if_mul_itm, COMP_LOOP_3_mul_mut, COMP_LOOP_4_modExp_1_while_mul_mut,
        COMP_LOOP_4_modExp_1_while_if_mul_itm, COMP_LOOP_4_mul_mut, {modulo_result_or_nl
        , and_96_nl , and_101_nl , mux_206_nl , and_102_nl , and_104_nl , and_107_nl
        , and_dcpl_102 , mux_229_nl , (~ mux_247_nl) , and_114_nl , and_115_nl ,
        and_117_nl , and_119_nl , and_123_nl , and_126_nl , and_128_nl , and_130_nl
        , and_131_nl});
    modulo_result_rem_cmp_b <= p_sva;
    operator_66_true_div_cmp_a <= MUX_v_65_2_2(z_out, ({operator_64_false_acc_mut_64
        , operator_64_false_acc_mut_63_0}), and_dcpl_128);
    operator_66_true_div_cmp_b_9_0 <= MUX_v_10_2_2(STAGE_LOOP_lshift_psp_sva_mx0w0,
        STAGE_LOOP_lshift_psp_sva, and_dcpl_128);
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_132_nl, nor_tmp_63, fsm_output[3]) ) begin
      STAGE_LOOP_lshift_psp_sva <= STAGE_LOOP_lshift_psp_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ mux_635_nl ) begin
      operator_64_false_acc_mut_64 <= operator_64_false_mux1h_1_rgt[64];
    end
  end
  always @(posedge clk) begin
    if ( ~(mux_640_nl | (fsm_output[6])) ) begin
      operator_64_false_acc_mut_63_0 <= operator_64_false_mux1h_1_rgt[63:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      VEC_LOOP_j_sva_11_0 <= 12'b000000000000;
    end
    else if ( and_dcpl_132 | VEC_LOOP_j_sva_11_0_mx0c1 ) begin
      VEC_LOOP_j_sva_11_0 <= MUX_v_12_2_2(12'b000000000000, (z_out_2[11:0]), VEC_LOOP_j_sva_11_0_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_k_9_2_sva_6_0 <= 7'b0000000;
    end
    else if ( MUX_s_1_2_2(nor_420_nl, nor_421_nl, fsm_output[7]) ) begin
      COMP_LOOP_k_9_2_sva_6_0 <= MUX_v_7_2_2(7'b0000000, (z_out_1[6:0]), mux_313_nl);
    end
  end
  always @(posedge clk) begin
    if ( (modExp_while_and_3 | modExp_while_and_5 | modExp_result_sva_mx0c0 | (~
        mux_325_nl)) & (modExp_result_sva_mx0c0 | modExp_result_and_rgt | modExp_result_and_1_rgt)
        ) begin
      modExp_result_sva <= MUX1HOT_v_64_3_2(64'b0000000000000000000000000000000000000000000000000000000000000001,
          modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w1, {modExp_result_sva_mx0c0
          , modExp_result_and_rgt , modExp_result_and_1_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_1_acc_5_mut <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( (modExp_while_and_3 | modExp_while_and_5 | and_dcpl_132 | and_dcpl_140
        | and_dcpl_102) & mux_380_nl ) begin
      COMP_LOOP_1_acc_5_mut <= MUX1HOT_v_64_5_2(({1'b0 , operator_64_false_slc_modExp_exp_63_1_3}),
          64'b0000000000000000000000000000000000000000000000000000000000000001, modulo_result_rem_cmp_z,
          modulo_qr_sva_1_mx0w1, COMP_LOOP_1_acc_5_mut_mx0w7, {and_dcpl_132 , and_dcpl_140
          , COMP_LOOP_and_nl , COMP_LOOP_and_1_nl , and_dcpl_102});
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_441_nl, mux_418_nl, fsm_output[3]) ) begin
      COMP_LOOP_1_acc_8_itm <= MUX1HOT_v_64_9_2(r_sva, modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w1,
          modExp_result_sva, vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d,
          vec_rsc_0_3_i_qa_d, (z_out[63:0]), {and_153_nl , COMP_LOOP_or_12_nl , COMP_LOOP_or_13_nl
          , and_dcpl_140 , nor_388_nl , and_162_nl , and_165_nl , and_168_nl , and_dcpl_102});
    end
  end
  always @(posedge clk) begin
    if ( ~(mux_489_nl & and_dcpl_89) ) begin
      modExp_while_if_mul_mut <= z_out_7;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      exit_COMP_LOOP_1_modExp_1_while_sva <= 1'b0;
    end
    else if ( and_dcpl_86 | and_dcpl_166 | and_dcpl_75 ) begin
      exit_COMP_LOOP_1_modExp_1_while_sva <= MUX1HOT_s_1_3_2((~ (z_out_5[63])), (~
          (z_out_6[8])), (~ (readslicef_10_1_9(COMP_LOOP_1_acc_nl))), {and_dcpl_86
          , and_dcpl_166 , and_dcpl_75});
    end
  end
  always @(posedge clk) begin
    if ( ~(or_tmp_300 | or_dcpl_38 | or_dcpl_36 | or_dcpl_35) ) begin
      modExp_while_mul_itm <= z_out_7;
    end
  end
  always @(posedge clk) begin
    if ( ~(or_tmp_70 | (~ (fsm_output[4])) | or_dcpl_43 | or_dcpl_42) ) begin
      COMP_LOOP_acc_psp_sva <= COMP_LOOP_acc_psp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_2_sva <= 12'b000000000000;
    end
    else if ( mux_493_nl | (fsm_output[8]) ) begin
      COMP_LOOP_acc_1_cse_2_sva <= z_out_6;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_11_psp_sva <= 11'b00000000000;
    end
    else if ( MUX_s_1_2_2(mux_501_nl, mux_499_nl, fsm_output[3]) ) begin
      COMP_LOOP_acc_11_psp_sva <= z_out_5[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_sva <= 12'b000000000000;
    end
    else if ( MUX_s_1_2_2(mux_505_nl, mux_504_nl, fsm_output[3]) ) begin
      COMP_LOOP_acc_1_cse_sva <= nl_COMP_LOOP_acc_1_cse_sva[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_5_1_sva_1 <= 1'b0;
      modExp_exp_1_5_1_sva <= 1'b0;
      modExp_exp_1_4_1_sva <= 1'b0;
      modExp_exp_1_3_1_sva <= 1'b0;
      modExp_exp_1_2_1_sva <= 1'b0;
    end
    else if ( mux_522_itm ) begin
      modExp_exp_1_5_1_sva_1 <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_2_sva_6_0[4]), modExp_exp_1_7_1_sva,
          (COMP_LOOP_k_9_2_sva_6_0[5]), {and_dcpl_168 , not_tmp_279 , and_dcpl_169});
      modExp_exp_1_5_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_2_sva_6_0[3]), modExp_exp_1_5_1_sva_1,
          (COMP_LOOP_k_9_2_sva_6_0[4]), {and_dcpl_168 , not_tmp_279 , and_dcpl_169});
      modExp_exp_1_4_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_2_sva_6_0[2]), modExp_exp_1_5_1_sva,
          (COMP_LOOP_k_9_2_sva_6_0[3]), {and_dcpl_168 , not_tmp_279 , and_dcpl_169});
      modExp_exp_1_3_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_2_sva_6_0[1]), modExp_exp_1_4_1_sva,
          (COMP_LOOP_k_9_2_sva_6_0[2]), {and_dcpl_168 , not_tmp_279 , and_dcpl_169});
      modExp_exp_1_2_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_2_sva_6_0[0]), modExp_exp_1_3_1_sva,
          (COMP_LOOP_k_9_2_sva_6_0[1]), {and_dcpl_168 , not_tmp_279 , and_dcpl_169});
    end
  end
  always @(posedge clk) begin
    if ( ~((~ mux_587_nl) & and_dcpl_29) ) begin
      COMP_LOOP_1_modExp_1_while_if_mul_mut <= COMP_LOOP_1_modExp_1_while_if_mul_mut_1;
    end
  end
  always @(posedge clk) begin
    if ( ~((fsm_output[1]) | (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[8])
        | (fsm_output[7]) | or_dcpl_47 | or_dcpl_35) ) begin
      COMP_LOOP_1_modExp_1_while_mul_itm <= z_out_7;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_12_1_1_sva <= 12'b000000000000;
    end
    else if ( COMP_LOOP_or_2_cse ) begin
      COMP_LOOP_acc_10_cse_12_1_1_sva <= z_out_5[12:1];
    end
  end
  always @(posedge clk) begin
    if ( and_dcpl_49 | and_dcpl_105 | and_dcpl_65 ) begin
      COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm <= MUX_s_1_2_2((readslicef_11_1_10(acc_3_nl)),
          (z_out_6[8]), and_dcpl_105);
    end
  end
  always @(posedge clk) begin
    if ( ~(or_tmp_300 | (~ (fsm_output[5])) | (fsm_output[1]) | or_dcpl_54 | or_dcpl_53)
        ) begin
      COMP_LOOP_1_mul_mut <= COMP_LOOP_1_modExp_1_while_if_mul_mut_1;
    end
  end
  always @(posedge clk) begin
    if ( ~(or_tmp_277 | (fsm_output[4]) | or_dcpl_43 | or_dcpl_59) ) begin
      COMP_LOOP_2_modExp_1_while_mul_mut <= z_out_7;
    end
  end
  always @(posedge clk) begin
    if ( ~((~ mux_598_nl) & and_dcpl_54) ) begin
      COMP_LOOP_2_modExp_1_while_if_mul_itm <= COMP_LOOP_1_modExp_1_while_if_mul_mut_1;
    end
  end
  always @(posedge clk) begin
    if ( ~(or_tmp_277 | (~ (fsm_output[4])) | or_dcpl_38 | or_dcpl_36 | or_dcpl_53)
        ) begin
      COMP_LOOP_2_mul_mut <= COMP_LOOP_1_modExp_1_while_if_mul_mut_1;
    end
  end
  always @(posedge clk) begin
    if ( ~(or_tmp_288 | or_dcpl_42) ) begin
      COMP_LOOP_3_modExp_1_while_mul_mut <= z_out_7;
    end
  end
  always @(posedge clk) begin
    if ( ~(mux_600_nl & and_dcpl_111) ) begin
      COMP_LOOP_3_modExp_1_while_if_mul_itm <= COMP_LOOP_1_modExp_1_while_if_mul_mut_1;
    end
  end
  always @(posedge clk) begin
    if ( ~(or_tmp_275 | (fsm_output[4]) | (fsm_output[5]) | (~ (fsm_output[1])) |
        or_dcpl_47 | or_dcpl_53) ) begin
      COMP_LOOP_3_mul_mut <= COMP_LOOP_1_modExp_1_while_if_mul_mut_1;
    end
  end
  always @(posedge clk) begin
    if ( ~((~ nor_tmp_16) | (fsm_output[4]) | or_dcpl_38 | or_dcpl_59) ) begin
      COMP_LOOP_4_modExp_1_while_mul_mut <= z_out_7;
    end
  end
  always @(posedge clk) begin
    if ( ~((~ mux_603_nl) & and_dcpl_122) ) begin
      COMP_LOOP_4_modExp_1_while_if_mul_itm <= COMP_LOOP_1_modExp_1_while_if_mul_mut_1;
    end
  end
  always @(posedge clk) begin
    if ( ~((~ and_dcpl_38) | or_dcpl_43 | (fsm_output[0]) | (fsm_output[2]) | or_dcpl_41)
        ) begin
      COMP_LOOP_4_mul_mut <= COMP_LOOP_1_modExp_1_while_if_mul_mut_1;
    end
  end
  assign modulo_result_or_nl = and_dcpl_86 | and_dcpl_105;
  assign and_96_nl = and_dcpl_89 & (and_93_cse | (fsm_output[4]));
  assign and_101_nl = (~(or_643_cse & (fsm_output[4]))) & and_dcpl_29 & and_dcpl_91;
  assign or_279_nl = (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[0]) | (~ (fsm_output[4]));
  assign nor_280_nl = ~((~ (fsm_output[7])) | (fsm_output[0]) | (~ (fsm_output[4])));
  assign nor_281_nl = ~((fsm_output[7]) | (~ (fsm_output[0])) | (fsm_output[4]));
  assign mux_204_nl = MUX_s_1_2_2(nor_280_nl, nor_281_nl, fsm_output[5]);
  assign nand_20_nl = ~(nor_92_cse & mux_204_nl);
  assign mux_205_nl = MUX_s_1_2_2(or_279_nl, nand_20_nl, fsm_output[2]);
  assign nor_279_nl = ~((fsm_output[8]) | mux_205_nl);
  assign nand_104_nl = ~((fsm_output[5]) & (fsm_output[7]) & (~ (fsm_output[0]))
      & (fsm_output[4]));
  assign or_271_nl = (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[0])) | (fsm_output[4]);
  assign mux_203_nl = MUX_s_1_2_2(nand_104_nl, or_271_nl, fsm_output[6]);
  assign nor_282_nl = ~((~ (fsm_output[8])) | (fsm_output[2]) | (fsm_output[3]) |
      mux_203_nl);
  assign mux_206_nl = MUX_s_1_2_2(nor_279_nl, nor_282_nl, fsm_output[1]);
  assign or_281_nl = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[5]) | (fsm_output[4]);
  assign mux_207_nl = MUX_s_1_2_2(or_604_cse, or_281_nl, fsm_output[2]);
  assign mux_208_nl = MUX_s_1_2_2(not_tmp_154, mux_207_nl, fsm_output[6]);
  assign mux_209_nl = MUX_s_1_2_2(or_tmp_254, mux_208_nl, fsm_output[3]);
  assign and_102_nl = (~ mux_209_nl) & and_dcpl_29;
  assign mux_213_nl = MUX_s_1_2_2(mux_tmp_212, or_tmp_256, or_287_cse);
  assign mux_210_nl = MUX_s_1_2_2(or_tmp_256, (fsm_output[5]), or_644_cse);
  assign mux_211_nl = MUX_s_1_2_2(or_tmp_256, mux_210_nl, fsm_output[2]);
  assign mux_214_nl = MUX_s_1_2_2(mux_213_nl, mux_211_nl, fsm_output[3]);
  assign and_104_nl = (~ mux_214_nl) & and_dcpl_29 & (fsm_output[6]);
  assign and_107_nl = not_tmp_158 & and_dcpl_29 & (fsm_output[6:5]==2'b11);
  assign nand_24_nl = ~((fsm_output[7]) & (~((fsm_output[2:0]==3'b111))));
  assign mux_227_nl = MUX_s_1_2_2((~ (fsm_output[7])), nand_24_nl, fsm_output[3]);
  assign nor_276_nl = ~((fsm_output[5:4]!=2'b00) | mux_227_nl);
  assign and_366_nl = (fsm_output[3]) & (fsm_output[7]) & or_287_cse;
  assign nand_121_nl = ~((fsm_output[2:1]==2'b11));
  assign mux_224_nl = MUX_s_1_2_2(or_642_cse, nand_121_nl, fsm_output[7]);
  assign mux_225_nl = MUX_s_1_2_2((fsm_output[7]), mux_224_nl, fsm_output[3]);
  assign mux_226_nl = MUX_s_1_2_2(and_366_nl, mux_225_nl, fsm_output[4]);
  assign and_288_nl = (fsm_output[5]) & mux_226_nl;
  assign mux_228_nl = MUX_s_1_2_2(nor_276_nl, and_288_nl, fsm_output[6]);
  assign and_362_nl = (fsm_output[3]) & (fsm_output[7]);
  assign nor_278_nl = ~((fsm_output[2:0]!=3'b000));
  assign mux_220_nl = MUX_s_1_2_2(nor_278_nl, (fsm_output[2]), fsm_output[7]);
  assign mux_221_nl = MUX_s_1_2_2((fsm_output[7]), (~ mux_220_nl), fsm_output[3]);
  assign mux_222_nl = MUX_s_1_2_2(and_362_nl, mux_221_nl, fsm_output[4]);
  assign or_298_nl = (fsm_output[7]) | and_365_cse;
  assign mux_219_nl = MUX_s_1_2_2((fsm_output[7]), or_298_nl, fsm_output[3]);
  assign nor_382_nl = ~((fsm_output[4]) | mux_219_nl);
  assign mux_223_nl = MUX_s_1_2_2(mux_222_nl, nor_382_nl, fsm_output[5]);
  assign and_291_nl = (fsm_output[6]) & mux_223_nl;
  assign mux_229_nl = MUX_s_1_2_2(mux_228_nl, and_291_nl, fsm_output[8]);
  assign nand_100_nl = ~((~((fsm_output[1]) & (fsm_output[7]))) & (fsm_output[8]));
  assign mux_242_nl = MUX_s_1_2_2(mux_tmp_230, or_tmp_277, and_289_cse);
  assign mux_243_nl = MUX_s_1_2_2(nand_100_nl, mux_242_nl, fsm_output[4]);
  assign or_312_nl = (fsm_output[4]) | (~ (fsm_output[7])) | (fsm_output[8]);
  assign mux_244_nl = MUX_s_1_2_2(mux_243_nl, or_312_nl, fsm_output[5]);
  assign nand_102_nl = ~((~(or_644_cse & (fsm_output[7]))) & (fsm_output[8]));
  assign mux_241_nl = MUX_s_1_2_2(nand_79_cse, nand_102_nl, fsm_output[4]);
  assign nand_26_nl = ~((fsm_output[5]) & (~ mux_241_nl));
  assign mux_245_nl = MUX_s_1_2_2(mux_244_nl, nand_26_nl, fsm_output[6]);
  assign mux_246_nl = MUX_s_1_2_2(mux_245_nl, mux_tmp_239, fsm_output[3]);
  assign mux_234_nl = MUX_s_1_2_2(or_tmp_275, mux_tmp_230, and_289_cse);
  assign mux_235_nl = MUX_s_1_2_2(mux_234_nl, or_tmp_277, fsm_output[4]);
  assign or_308_nl = (fsm_output[5]) | mux_235_nl;
  assign nand_55_nl = ~((fsm_output[4]) & (fsm_output[7]) & (fsm_output[8]));
  assign nand_56_nl = ~(((fsm_output[0]) | (fsm_output[1]) | (fsm_output[7])) & (fsm_output[8]));
  assign mux_231_nl = MUX_s_1_2_2(or_tmp_275, mux_tmp_230, fsm_output[1]);
  assign mux_232_nl = MUX_s_1_2_2(nand_56_nl, mux_231_nl, fsm_output[4]);
  assign mux_233_nl = MUX_s_1_2_2(nand_55_nl, mux_232_nl, fsm_output[5]);
  assign mux_236_nl = MUX_s_1_2_2(or_308_nl, mux_233_nl, fsm_output[6]);
  assign mux_240_nl = MUX_s_1_2_2(mux_tmp_239, mux_236_nl, fsm_output[3]);
  assign mux_247_nl = MUX_s_1_2_2(mux_246_nl, mux_240_nl, fsm_output[2]);
  assign nand_107_nl = ~((fsm_output[2]) & (fsm_output[4]));
  assign mux_250_nl = MUX_s_1_2_2((fsm_output[4]), nand_107_nl, fsm_output[3]);
  assign and_114_nl = and_dcpl_54 & and_dcpl_91 & mux_250_nl;
  assign mux_252_nl = MUX_s_1_2_2((fsm_output[5]), or_604_cse, or_319_cse);
  assign nand_27_nl = ~((fsm_output[6]) & (~ mux_252_nl));
  assign nand_54_nl = ~((fsm_output[2]) & (fsm_output[5]) & (fsm_output[4]));
  assign mux_251_nl = MUX_s_1_2_2(nand_54_nl, or_604_cse, fsm_output[6]);
  assign mux_253_nl = MUX_s_1_2_2(nand_27_nl, mux_251_nl, fsm_output[3]);
  assign and_115_nl = (~ mux_253_nl) & and_dcpl_54;
  assign mux_255_nl = MUX_s_1_2_2(or_625_cse, mux_tmp_212, or_644_cse);
  assign mux_256_nl = MUX_s_1_2_2(or_625_cse, mux_255_nl, fsm_output[2]);
  assign mux_254_nl = MUX_s_1_2_2(mux_tmp_212, or_tmp_256, or_319_cse);
  assign mux_257_nl = MUX_s_1_2_2(mux_256_nl, mux_254_nl, fsm_output[3]);
  assign and_117_nl = (~ mux_257_nl) & and_dcpl_54 & (fsm_output[6]);
  assign mux_260_nl = MUX_s_1_2_2(or_625_cse, mux_tmp_212, and_281_cse);
  assign mux_645_nl = MUX_s_1_2_2(mux_tmp_212, or_tmp_256, and_289_cse);
  assign mux_259_nl = MUX_s_1_2_2(mux_645_nl, or_tmp_256, fsm_output[2]);
  assign mux_261_nl = MUX_s_1_2_2(mux_260_nl, mux_259_nl, fsm_output[3]);
  assign and_119_nl = (~ mux_261_nl) & and_dcpl_111;
  assign and_123_nl = ((or_642_cse & (fsm_output[3])) | (fsm_output[4])) & and_dcpl_67
      & and_dcpl_91;
  assign nor_275_nl = ~((fsm_output[2]) | (fsm_output[4]));
  assign mux_262_nl = MUX_s_1_2_2(nor_275_nl, (fsm_output[4]), fsm_output[3]);
  assign and_126_nl = and_dcpl_67 & (fsm_output[6:5]==2'b10) & (~ mux_262_nl);
  assign and_128_nl = not_tmp_158 & nor_tmp_16 & and_dcpl_88;
  assign mux_263_nl = MUX_s_1_2_2(or_625_cse, mux_tmp_212, fsm_output[1]);
  assign mux_614_nl = MUX_s_1_2_2(mux_tmp_212, or_tmp_256, and_289_cse);
  assign mux_264_nl = MUX_s_1_2_2(mux_263_nl, mux_614_nl, fsm_output[2]);
  assign mux_265_nl = MUX_s_1_2_2(or_625_cse, mux_264_nl, fsm_output[3]);
  assign and_130_nl = (~ mux_265_nl) & and_dcpl_122;
  assign and_278_nl = (fsm_output[0]) & (fsm_output[1]) & (fsm_output[5]) & (fsm_output[4]);
  assign mux_266_nl = MUX_s_1_2_2(and_278_nl, and_273_cse, fsm_output[2]);
  assign nor_273_nl = ~(and_281_cse | (fsm_output[5:4]!=2'b00));
  assign mux_267_nl = MUX_s_1_2_2(mux_266_nl, nor_273_nl, fsm_output[6]);
  assign nor_274_nl = ~((fsm_output[6]) | (~ and_273_cse));
  assign mux_268_nl = MUX_s_1_2_2(mux_267_nl, nor_274_nl, fsm_output[3]);
  assign and_131_nl = mux_268_nl & nor_tmp_16;
  assign COMP_LOOP_and_9_nl = (~ and_dcpl_139) & and_dcpl_132;
  assign and_335_nl = (fsm_output[0]) & (fsm_output[1]) & (fsm_output[3]) & (~ (fsm_output[8]));
  assign nor_351_nl = ~((~ (fsm_output[3])) | (fsm_output[8]));
  assign mux_75_nl = MUX_s_1_2_2(and_335_nl, nor_351_nl, fsm_output[2]);
  assign or_75_nl = (fsm_output[1]) | (fsm_output[3]) | (~ (fsm_output[8]));
  assign or_409_nl = (fsm_output[1]) | (~ (fsm_output[0])) | (~ (fsm_output[3]))
      | (fsm_output[8]);
  assign mux_455_nl = MUX_s_1_2_2(or_75_nl, or_409_nl, fsm_output[2]);
  assign mux_457_nl = MUX_s_1_2_2(mux_75_nl, mux_455_nl, fsm_output[6]);
  assign or_408_nl = (fsm_output[6]) | and_206_cse | (fsm_output[3]) | (~ (fsm_output[8]));
  assign mux_458_nl = MUX_s_1_2_2(mux_457_nl, or_408_nl, fsm_output[4]);
  assign or_405_nl = (~(and_289_cse | (fsm_output[3]))) | (fsm_output[8]);
  assign or_403_nl = (~ (fsm_output[6])) | (fsm_output[2]);
  assign mux_453_nl = MUX_s_1_2_2(or_405_nl, (fsm_output[8]), or_403_nl);
  assign or_402_nl = (~((fsm_output[6]) | (~ (fsm_output[3])))) | (fsm_output[8]);
  assign mux_454_nl = MUX_s_1_2_2(mux_453_nl, or_402_nl, fsm_output[4]);
  assign mux_459_nl = MUX_s_1_2_2(mux_458_nl, mux_454_nl, fsm_output[5]);
  assign nand_93_nl = ~(((~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[3]))
      & (fsm_output[8]));
  assign nand_94_nl = ~(((fsm_output[0]) | (fsm_output[1]) | (fsm_output[3])) & (fsm_output[8]));
  assign mux_69_nl = MUX_s_1_2_2(nand_93_nl, nand_94_nl, fsm_output[2]);
  assign mux_70_nl = MUX_s_1_2_2(mux_69_nl, (fsm_output[8]), fsm_output[6]);
  assign nor_378_nl = ~((fsm_output[2]) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[3])
      | (fsm_output[8]));
  assign mux_68_nl = MUX_s_1_2_2((fsm_output[8]), nor_378_nl, fsm_output[6]);
  assign mux_71_nl = MUX_s_1_2_2((~ mux_70_nl), mux_68_nl, fsm_output[4]);
  assign nor_379_nl = ~((fsm_output[6]) | mux_66_cse);
  assign mux_67_nl = MUX_s_1_2_2(nor_379_nl, nor_380_cse, fsm_output[4]);
  assign mux_72_nl = MUX_s_1_2_2(mux_71_nl, mux_67_nl, fsm_output[5]);
  assign mux_460_nl = MUX_s_1_2_2(mux_459_nl, mux_72_nl, fsm_output[7]);
  assign COMP_LOOP_mux1h_18_nl = MUX1HOT_s_1_6_2((operator_66_true_div_cmp_z[0]),
      (COMP_LOOP_1_acc_5_mut[0]), (z_out_2[7]), modExp_exp_1_0_1_sva_1, modExp_exp_1_0_1_sva,
      (z_out_6[7]), {COMP_LOOP_and_9_nl , and_dcpl_139 , and_dcpl_45 , not_tmp_235
      , mux_460_nl , and_dcpl_72});
  assign nor_245_nl = ~((fsm_output[5]) | (~ (fsm_output[8])));
  assign mux_445_nl = MUX_s_1_2_2(nor_245_nl, nor_246_cse, fsm_output[1]);
  assign mux_484_nl = MUX_s_1_2_2(mux_tmp_473, mux_tmp_463, fsm_output[6]);
  assign mux_485_nl = MUX_s_1_2_2(mux_tmp_481, mux_484_nl, fsm_output[4]);
  assign mux_482_nl = MUX_s_1_2_2(mux_tmp_481, mux_tmp_474, fsm_output[4]);
  assign mux_483_nl = MUX_s_1_2_2(mux_482_nl, mux_tmp_476, fsm_output[0]);
  assign mux_486_nl = MUX_s_1_2_2(mux_485_nl, mux_483_nl, fsm_output[1]);
  assign mux_480_nl = MUX_s_1_2_2(mux_tmp_469, mux_tmp_466, fsm_output[1]);
  assign mux_487_nl = MUX_s_1_2_2(mux_486_nl, mux_480_nl, fsm_output[3]);
  assign mux_477_nl = MUX_s_1_2_2(mux_tmp_476, mux_tmp_471, fsm_output[0]);
  assign mux_472_nl = MUX_s_1_2_2(mux_tmp_471, mux_tmp_469, fsm_output[0]);
  assign mux_478_nl = MUX_s_1_2_2(mux_477_nl, mux_472_nl, fsm_output[1]);
  assign mux_479_nl = MUX_s_1_2_2(mux_478_nl, mux_tmp_466, fsm_output[3]);
  assign mux_488_nl = MUX_s_1_2_2(mux_487_nl, mux_479_nl, fsm_output[2]);
  assign or_478_nl = (fsm_output[4]) | or_dcpl_43;
  assign or_477_nl = (fsm_output[4]) | (fsm_output[1]) | (fsm_output[5]);
  assign mux_536_nl = MUX_s_1_2_2(or_478_nl, or_477_nl, fsm_output[8]);
  assign nor_228_nl = ~((fsm_output[7]) | mux_536_nl);
  assign nor_229_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[4]))
      | (fsm_output[1]) | (fsm_output[5]));
  assign mux_537_nl = MUX_s_1_2_2(nor_228_nl, nor_229_nl, fsm_output[0]);
  assign and_226_nl = nor_92_cse & mux_537_nl;
  assign nor_230_nl = ~((~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[0]))
      | (~ (fsm_output[7])) | (~ (fsm_output[8])) | (fsm_output[4]) | or_dcpl_43);
  assign mux_538_nl = MUX_s_1_2_2(and_226_nl, nor_230_nl, fsm_output[2]);
  assign COMP_LOOP_mux_24_nl = MUX_s_1_2_2(modExp_exp_1_0_1_sva_1, modExp_exp_1_1_1_sva,
      mux_538_nl);
  assign nor_234_nl = ~((fsm_output[4]) | (~ (fsm_output[7])));
  assign nor_235_nl = ~((~ (fsm_output[4])) | (fsm_output[7]));
  assign mux_524_nl = MUX_s_1_2_2(nor_234_nl, nor_235_nl, fsm_output[0]);
  assign nand_39_nl = ~(or_585_cse & (fsm_output[8]));
  assign nor_225_nl = ~(and_93_cse | (fsm_output[8]));
  assign mux_546_nl = MUX_s_1_2_2(nand_39_nl, nor_225_nl, or_644_cse);
  assign nand_34_nl = ~((fsm_output[6]) & mux_546_nl);
  assign or_490_nl = (fsm_output[0]) | (~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[3])
      | (fsm_output[8]);
  assign mux_545_nl = MUX_s_1_2_2((~ (fsm_output[8])), or_490_nl, fsm_output[6]);
  assign mux_547_nl = MUX_s_1_2_2(nand_34_nl, mux_545_nl, fsm_output[5]);
  assign or_489_nl = (fsm_output[6]) | (~(or_589_cse & (fsm_output[8])));
  assign or_487_nl = (fsm_output[6]) | (~(and_281_cse | (fsm_output[3]) | (fsm_output[8])));
  assign mux_544_nl = MUX_s_1_2_2(or_489_nl, or_487_nl, fsm_output[5]);
  assign mux_548_nl = MUX_s_1_2_2(mux_547_nl, mux_544_nl, fsm_output[4]);
  assign nand_41_nl = ~(or_643_cse & (fsm_output[8]));
  assign mux_541_nl = MUX_s_1_2_2(nand_41_nl, (fsm_output[8]), fsm_output[6]);
  assign or_483_nl = (fsm_output[6]) | (~(and_206_cse | (fsm_output[3]) | (fsm_output[8])));
  assign mux_542_nl = MUX_s_1_2_2(mux_541_nl, or_483_nl, fsm_output[5]);
  assign mux_539_nl = MUX_s_1_2_2((~ (fsm_output[8])), or_481_cse, fsm_output[6]);
  assign or_12_nl = (fsm_output[8]) | (fsm_output[6]);
  assign mux_540_nl = MUX_s_1_2_2(mux_539_nl, or_12_nl, fsm_output[5]);
  assign mux_543_nl = MUX_s_1_2_2(mux_542_nl, mux_540_nl, fsm_output[4]);
  assign mux_549_nl = MUX_s_1_2_2(mux_548_nl, mux_543_nl, fsm_output[7]);
  assign COMP_LOOP_mux1h_29_nl = MUX1HOT_s_1_4_2((COMP_LOOP_k_9_2_sva_6_0[5]), modExp_exp_1_1_1_sva,
      modExp_exp_1_7_1_sva, (COMP_LOOP_k_9_2_sva_6_0[6]), {and_dcpl_168 , and_dcpl_166
      , (~ mux_522_itm) , and_dcpl_169});
  assign nor_222_nl = ~((fsm_output[7]) | (fsm_output[4]) | (~ (fsm_output[8])));
  assign nor_223_nl = ~((~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_550_nl = MUX_s_1_2_2(nor_222_nl, nor_223_nl, fsm_output[0]);
  assign nand_130_nl = ~((~((fsm_output[2]) | (fsm_output[3]) | (fsm_output[5]) |
      (~ (fsm_output[6])))) & mux_550_nl);
  assign nand_131_nl = ~((fsm_output[2]) & (fsm_output[3]) & (fsm_output[5]) & (~
      (fsm_output[6])) & (fsm_output[0]) & (fsm_output[7]) & (~ (fsm_output[4]))
      & (fsm_output[8]));
  assign mux_551_nl = MUX_s_1_2_2(nand_130_nl, nand_131_nl, fsm_output[1]);
  assign or_504_nl = (fsm_output[4]) | (fsm_output[2]) | (fsm_output[1]) | (fsm_output[3])
      | (fsm_output[8]);
  assign mux_559_nl = MUX_s_1_2_2((fsm_output[8]), or_504_nl, fsm_output[5]);
  assign mux_562_nl = MUX_s_1_2_2((~ mux_561_cse), mux_559_nl, fsm_output[6]);
  assign mux_563_nl = MUX_s_1_2_2(mux_562_nl, mux_558_cse, fsm_output[7]);
  assign COMP_LOOP_mux1h_43_nl = MUX1HOT_s_1_4_2((COMP_LOOP_k_9_2_sva_6_0[6]), modExp_exp_1_2_1_sva,
      modExp_exp_1_1_1_sva, (COMP_LOOP_k_9_2_sva_6_0[0]), {and_dcpl_168 , not_tmp_279
      , (~ mux_563_nl) , and_dcpl_169});
  assign nor_272_nl = ~((fsm_output[2]) | (fsm_output[1]) | (fsm_output[5]) | (fsm_output[4])
      | (fsm_output[8]) | (fsm_output[7]));
  assign mux_132_nl = MUX_s_1_2_2(nor_272_nl, and_313_cse, fsm_output[6]);
  assign or_671_nl = (fsm_output[6]) | nor_tmp_210;
  assign or_670_nl = (fsm_output[6]) | (~ or_tmp);
  assign mux_632_nl = MUX_s_1_2_2(or_671_nl, or_670_nl, fsm_output[0]);
  assign or_669_nl = (fsm_output[4]) | (fsm_output[7]) | (fsm_output[2]);
  assign mux_633_nl = MUX_s_1_2_2(mux_632_nl, (fsm_output[6]), or_669_nl);
  assign and_521_nl = (fsm_output[6]) & or_tmp;
  assign mux_628_nl = MUX_s_1_2_2(nor_tmp, and_521_nl, fsm_output[0]);
  assign mux_629_nl = MUX_s_1_2_2(mux_tmp, mux_628_nl, fsm_output[2]);
  assign mux_630_nl = MUX_s_1_2_2((~ (fsm_output[6])), mux_629_nl, fsm_output[7]);
  assign mux_625_nl = MUX_s_1_2_2(mux_tmp_616, nor_tmp, fsm_output[0]);
  assign mux_626_nl = MUX_s_1_2_2(mux_tmp, mux_625_nl, fsm_output[2]);
  assign mux_627_nl = MUX_s_1_2_2(mux_626_nl, (fsm_output[6]), fsm_output[7]);
  assign mux_631_nl = MUX_s_1_2_2(mux_630_nl, mux_627_nl, fsm_output[4]);
  assign mux_634_nl = MUX_s_1_2_2((~ mux_633_nl), mux_631_nl, fsm_output[8]);
  assign mux_620_nl = MUX_s_1_2_2(mux_tmp_613, mux_tmp, fsm_output[0]);
  assign mux_621_nl = MUX_s_1_2_2(mux_620_nl, mux_tmp_616, fsm_output[2]);
  assign mux_622_nl = MUX_s_1_2_2((~ (fsm_output[6])), mux_621_nl, fsm_output[7]);
  assign mux_615_nl = MUX_s_1_2_2(mux_tmp, nor_tmp, fsm_output[0]);
  assign mux_617_nl = MUX_s_1_2_2(mux_tmp_613, mux_615_nl, fsm_output[2]);
  assign mux_618_nl = MUX_s_1_2_2(mux_617_nl, (fsm_output[6]), fsm_output[7]);
  assign mux_623_nl = MUX_s_1_2_2(mux_622_nl, mux_618_nl, fsm_output[4]);
  assign mux_624_nl = MUX_s_1_2_2(mux_623_nl, (fsm_output[6]), fsm_output[8]);
  assign mux_635_nl = MUX_s_1_2_2(mux_634_nl, mux_624_nl, fsm_output[5]);
  assign or_688_nl = (fsm_output[2]) | (fsm_output[4]) | (~ (fsm_output[0])) | (fsm_output[7])
      | (fsm_output[3]);
  assign nand_138_nl = ~((fsm_output[2]) & not_tmp_397);
  assign mux_638_nl = MUX_s_1_2_2(or_688_nl, nand_138_nl, fsm_output[8]);
  assign or_689_nl = (fsm_output[8]) | (fsm_output[2]) | (fsm_output[4]) | (fsm_output[0])
      | (fsm_output[7]) | (~ (fsm_output[3]));
  assign mux_639_nl = MUX_s_1_2_2(mux_638_nl, or_689_nl, fsm_output[1]);
  assign or_690_nl = (fsm_output[8]) | (~ (fsm_output[2])) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (fsm_output[7]) | (fsm_output[3]);
  assign nand_139_nl = ~((~((fsm_output[8]) | (~ (fsm_output[2])))) & not_tmp_397);
  assign mux_637_nl = MUX_s_1_2_2(or_690_nl, nand_139_nl, fsm_output[1]);
  assign mux_640_nl = MUX_s_1_2_2(mux_639_nl, mux_637_nl, fsm_output[5]);
  assign or_nl = (fsm_output[8:1]!=8'b00000101);
  assign nor_268_nl = ~((~ (fsm_output[2])) | (fsm_output[6]) | (fsm_output[7]) |
      (fsm_output[8]));
  assign nor_269_nl = ~((fsm_output[2]) | nand_53_cse);
  assign mux_312_nl = MUX_s_1_2_2(nor_268_nl, nor_269_nl, fsm_output[1]);
  assign nand_134_nl = ~((~((fsm_output[5:3]!=3'b110))) & mux_312_nl);
  assign mux_313_nl = MUX_s_1_2_2(or_nl, nand_134_nl, fsm_output[0]);
  assign or_686_nl = (fsm_output[0]) | (fsm_output[6]) | (~ (fsm_output[1])) | (~
      (fsm_output[3])) | (fsm_output[4]) | (fsm_output[5]);
  assign or_685_nl = (~ (fsm_output[0])) | (fsm_output[6]) | (fsm_output[1]) | (fsm_output[3])
      | not_tmp_400;
  assign mux_642_nl = MUX_s_1_2_2(or_686_nl, or_685_nl, fsm_output[2]);
  assign nor_420_nl = ~((fsm_output[8]) | mux_642_nl);
  assign or_682_nl = (fsm_output[6]) | (fsm_output[1]) | (fsm_output[3]) | not_tmp_400;
  assign or_680_nl = (~ (fsm_output[6])) | (~ (fsm_output[1])) | (fsm_output[3])
      | not_tmp_400;
  assign mux_641_nl = MUX_s_1_2_2(or_682_nl, or_680_nl, fsm_output[0]);
  assign nor_421_nl = ~((~ (fsm_output[8])) | (fsm_output[2]) | mux_641_nl);
  assign nor_261_nl = ~((or_319_cse & (fsm_output[5])) | (fsm_output[4]) | (fsm_output[8])
      | (fsm_output[7]));
  assign mux_324_nl = MUX_s_1_2_2(nor_261_nl, and_313_cse, fsm_output[6]);
  assign mux_325_nl = MUX_s_1_2_2(mux_324_nl, mux_tmp_321, fsm_output[3]);
  assign COMP_LOOP_and_nl = (~ modExp_while_and_5) & not_tmp_235;
  assign COMP_LOOP_and_1_nl = modExp_while_and_5 & not_tmp_235;
  assign mux_375_nl = MUX_s_1_2_2((~ mux_351_itm), or_tmp_331, fsm_output[3]);
  assign mux_376_nl = MUX_s_1_2_2(mux_375_nl, mux_tmp_354, fsm_output[0]);
  assign mux_373_nl = MUX_s_1_2_2(mux_tmp_339, mux_tmp_337, fsm_output[3]);
  assign mux_372_nl = MUX_s_1_2_2(mux_tmp_86, or_tmp_277, fsm_output[3]);
  assign mux_374_nl = MUX_s_1_2_2(mux_373_nl, mux_372_nl, fsm_output[0]);
  assign mux_377_nl = MUX_s_1_2_2(mux_376_nl, mux_374_nl, fsm_output[4]);
  assign mux_370_nl = MUX_s_1_2_2(mux_tmp_336, and_tmp_8, fsm_output[3]);
  assign mux_369_nl = MUX_s_1_2_2(and_tmp_9, mux_tmp_330, fsm_output[3]);
  assign mux_371_nl = MUX_s_1_2_2(mux_370_nl, mux_369_nl, fsm_output[4]);
  assign mux_378_nl = MUX_s_1_2_2((~ mux_377_nl), mux_371_nl, fsm_output[5]);
  assign or_366_nl = nor_380_cse | (fsm_output[7]);
  assign mux_365_nl = MUX_s_1_2_2(not_tmp_221, or_366_nl, fsm_output[3]);
  assign mux_366_nl = MUX_s_1_2_2(mux_tmp_352, mux_365_nl, fsm_output[0]);
  assign mux_364_nl = MUX_s_1_2_2((~ mux_tmp_86), mux_tmp_336, fsm_output[3]);
  assign mux_367_nl = MUX_s_1_2_2((~ mux_366_nl), mux_364_nl, fsm_output[4]);
  assign mux_361_nl = MUX_s_1_2_2(mux_tmp_336, and_tmp_9, fsm_output[3]);
  assign mux_362_nl = MUX_s_1_2_2(mux_361_nl, mux_tmp_333, fsm_output[0]);
  assign mux_359_nl = MUX_s_1_2_2(mux_tmp_330, mux_tmp_344, fsm_output[3]);
  assign mux_360_nl = MUX_s_1_2_2(mux_359_nl, mux_tmp_329, fsm_output[0]);
  assign mux_363_nl = MUX_s_1_2_2(mux_362_nl, mux_360_nl, fsm_output[4]);
  assign mux_368_nl = MUX_s_1_2_2(mux_367_nl, mux_363_nl, fsm_output[5]);
  assign mux_379_nl = MUX_s_1_2_2(mux_378_nl, mux_368_nl, fsm_output[2]);
  assign mux_355_nl = MUX_s_1_2_2(mux_tmp_354, mux_tmp_352, fsm_output[0]);
  assign mux_349_nl = MUX_s_1_2_2(mux_tmp_339, or_tmp_277, fsm_output[3]);
  assign mux_348_nl = MUX_s_1_2_2((~ mux_tmp_339), mux_tmp_336, fsm_output[3]);
  assign mux_350_nl = MUX_s_1_2_2((~ mux_349_nl), mux_348_nl, fsm_output[0]);
  assign mux_356_nl = MUX_s_1_2_2((~ mux_355_nl), mux_350_nl, fsm_output[4]);
  assign and_150_nl = (fsm_output[6]) & mux_tmp_86;
  assign mux_346_nl = MUX_s_1_2_2(mux_tmp_336, and_150_nl, fsm_output[3]);
  assign and_258_nl = (fsm_output[0]) & (fsm_output[3]);
  assign mux_345_nl = MUX_s_1_2_2(mux_tmp_330, mux_tmp_344, and_258_nl);
  assign mux_347_nl = MUX_s_1_2_2(mux_346_nl, mux_345_nl, fsm_output[4]);
  assign mux_357_nl = MUX_s_1_2_2(mux_356_nl, mux_347_nl, fsm_output[5]);
  assign mux_341_nl = MUX_s_1_2_2(not_tmp_221, mux_tmp_339, fsm_output[3]);
  assign mux_338_nl = MUX_s_1_2_2((~ mux_tmp_337), mux_tmp_336, fsm_output[3]);
  assign mux_342_nl = MUX_s_1_2_2((~ mux_341_nl), mux_338_nl, fsm_output[4]);
  assign mux_331_nl = MUX_s_1_2_2(and_tmp_8, mux_tmp_330, fsm_output[3]);
  assign mux_334_nl = MUX_s_1_2_2(mux_tmp_333, mux_331_nl, fsm_output[0]);
  assign mux_335_nl = MUX_s_1_2_2(mux_334_nl, mux_tmp_329, fsm_output[4]);
  assign mux_343_nl = MUX_s_1_2_2(mux_342_nl, mux_335_nl, fsm_output[5]);
  assign mux_358_nl = MUX_s_1_2_2(mux_357_nl, mux_343_nl, fsm_output[2]);
  assign mux_380_nl = MUX_s_1_2_2(mux_379_nl, mux_358_nl, fsm_output[1]);
  assign and_153_nl = and_dcpl_85 & and_dcpl_141;
  assign COMP_LOOP_or_12_nl = ((~ (modulo_result_rem_cmp_z[63])) & and_156_m1c) |
      (not_tmp_253 & and_dcpl_50 & (~ (modulo_result_rem_cmp_z[63])));
  assign COMP_LOOP_or_13_nl = ((modulo_result_rem_cmp_z[63]) & and_156_m1c) | (not_tmp_253
      & and_dcpl_50 & (modulo_result_rem_cmp_z[63]));
  assign nor_388_nl = ~((~ not_tmp_242) | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b00)
      | (fsm_output[3]));
  assign and_162_nl = not_tmp_242 & (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]==2'b01)
      & (~ (fsm_output[3]));
  assign and_165_nl = not_tmp_242 & (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]==2'b10)
      & (~ (fsm_output[3]));
  assign and_168_nl = not_tmp_242 & (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]==2'b11)
      & (~ (fsm_output[3]));
  assign mux_437_nl = MUX_s_1_2_2(mux_tmp_397, mux_tmp_427, fsm_output[5]);
  assign mux_438_nl = MUX_s_1_2_2(mux_437_nl, mux_tmp_428, fsm_output[1]);
  assign mux_435_nl = MUX_s_1_2_2(mux_tmp_86, mux_tmp_427, fsm_output[5]);
  assign mux_436_nl = MUX_s_1_2_2(mux_435_nl, mux_tmp_412, fsm_output[1]);
  assign mux_439_nl = MUX_s_1_2_2(mux_438_nl, mux_436_nl, fsm_output[0]);
  assign mux_432_nl = MUX_s_1_2_2(mux_tmp_86, mux_tmp_408, fsm_output[5]);
  assign mux_433_nl = MUX_s_1_2_2(mux_tmp_412, mux_432_nl, fsm_output[1]);
  assign mux_429_nl = MUX_s_1_2_2(and_dcpl_29, or_tmp_277, fsm_output[4]);
  assign mux_430_nl = MUX_s_1_2_2(mux_429_nl, mux_tmp_408, fsm_output[5]);
  assign mux_431_nl = MUX_s_1_2_2(mux_430_nl, mux_tmp_428, fsm_output[1]);
  assign mux_434_nl = MUX_s_1_2_2(mux_433_nl, mux_431_nl, fsm_output[0]);
  assign mux_440_nl = MUX_s_1_2_2(mux_439_nl, mux_434_nl, fsm_output[2]);
  assign mux_424_nl = MUX_s_1_2_2(mux_tmp_404, mux_tmp_420, fsm_output[1]);
  assign mux_421_nl = MUX_s_1_2_2(and_dcpl_54, (fsm_output[7]), fsm_output[4]);
  assign mux_422_nl = MUX_s_1_2_2((~ mux_421_nl), mux_93_cse, fsm_output[5]);
  assign mux_423_nl = MUX_s_1_2_2(mux_422_nl, mux_tmp_420, fsm_output[1]);
  assign mux_425_nl = MUX_s_1_2_2(mux_424_nl, mux_423_nl, fsm_output[0]);
  assign mux_426_nl = MUX_s_1_2_2(mux_425_nl, mux_tmp_420, fsm_output[2]);
  assign mux_441_nl = MUX_s_1_2_2(mux_440_nl, mux_426_nl, fsm_output[6]);
  assign mux_414_nl = MUX_s_1_2_2(mux_tmp_411, mux_tmp_409, fsm_output[5]);
  assign mux_415_nl = MUX_s_1_2_2(mux_414_nl, mux_tmp_412, fsm_output[1]);
  assign mux_410_nl = MUX_s_1_2_2((~ mux_tmp_409), mux_tmp_408, fsm_output[5]);
  assign mux_413_nl = MUX_s_1_2_2(mux_tmp_412, mux_410_nl, fsm_output[1]);
  assign mux_416_nl = MUX_s_1_2_2(mux_415_nl, mux_413_nl, fsm_output[0]);
  assign mux_405_nl = MUX_s_1_2_2((~ (fsm_output[8])), or_tmp_275, fsm_output[4]);
  assign mux_406_nl = MUX_s_1_2_2(not_tmp_246, mux_405_nl, fsm_output[5]);
  assign mux_407_nl = MUX_s_1_2_2(mux_406_nl, mux_tmp_404, or_644_cse);
  assign mux_417_nl = MUX_s_1_2_2(mux_416_nl, mux_407_nl, fsm_output[2]);
  assign nand_49_nl = ~(((~ (fsm_output[4])) | (fsm_output[8])) & (fsm_output[7]));
  assign mux_399_nl = MUX_s_1_2_2(nand_49_nl, mux_93_cse, fsm_output[5]);
  assign mux_398_nl = MUX_s_1_2_2((~ mux_391_itm), mux_tmp_397, fsm_output[5]);
  assign mux_400_nl = MUX_s_1_2_2(mux_399_nl, mux_398_nl, fsm_output[1]);
  assign mux_395_nl = MUX_s_1_2_2((~ mux_391_itm), mux_93_cse, fsm_output[5]);
  assign mux_396_nl = MUX_s_1_2_2(mux_395_nl, mux_tmp_392, fsm_output[1]);
  assign mux_401_nl = MUX_s_1_2_2(mux_400_nl, mux_396_nl, fsm_output[0]);
  assign mux_402_nl = MUX_s_1_2_2(mux_401_nl, mux_tmp_392, fsm_output[2]);
  assign mux_418_nl = MUX_s_1_2_2(mux_417_nl, mux_402_nl, fsm_output[6]);
  assign nand_106_nl = ~((fsm_output[0]) & (fsm_output[1]) & (fsm_output[4]));
  assign mux_489_nl = MUX_s_1_2_2((fsm_output[4]), nand_106_nl, and_93_cse);
  assign nl_COMP_LOOP_1_acc_nl = ({(z_out_1[7:0]) , 2'b00}) + ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[9:1]))})
      + 10'b0000000001;
  assign COMP_LOOP_1_acc_nl = nl_COMP_LOOP_1_acc_nl[9:0];
  assign nor_369_nl = ~((fsm_output[6]) | and_333_cse | (fsm_output[7]));
  assign nor_370_nl = ~(and_273_cse | (fsm_output[7]));
  assign and_361_nl = (fsm_output[2]) & (fsm_output[1]) & (fsm_output[5]) & (fsm_output[4])
      & (fsm_output[7]);
  assign mux_492_nl = MUX_s_1_2_2(nor_370_nl, and_361_nl, fsm_output[6]);
  assign mux_493_nl = MUX_s_1_2_2(nor_369_nl, mux_492_nl, fsm_output[3]);
  assign mux_500_nl = MUX_s_1_2_2(mux_tmp_86, nor_tmp_16, and_333_cse);
  assign mux_501_nl = MUX_s_1_2_2(mux_500_nl, mux_tmp_495, fsm_output[6]);
  assign mux_498_nl = MUX_s_1_2_2(mux_tmp_86, nor_tmp_16, and_273_cse);
  assign mux_494_nl = MUX_s_1_2_2(nor_tmp_16, (fsm_output[8]), fsm_output[5]);
  assign mux_496_nl = MUX_s_1_2_2(mux_tmp_495, mux_494_nl, or_644_cse);
  assign mux_497_nl = MUX_s_1_2_2(mux_tmp_495, mux_496_nl, fsm_output[2]);
  assign mux_499_nl = MUX_s_1_2_2(mux_498_nl, mux_497_nl, fsm_output[6]);
  assign nl_COMP_LOOP_acc_1_cse_sva  = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_2_sva_6_0
      , 2'b11});
  assign nor_239_nl = ~(and_333_cse | (fsm_output[8:7]!=2'b00));
  assign mux_505_nl = MUX_s_1_2_2(nor_239_nl, nor_tmp_162, fsm_output[6]);
  assign nor_240_nl = ~(and_273_cse | (fsm_output[8:7]!=2'b00));
  assign and_241_nl = or_604_cse & (fsm_output[8:7]==2'b11);
  assign mux_503_nl = MUX_s_1_2_2(nor_tmp_162, and_241_nl, fsm_output[2]);
  assign mux_504_nl = MUX_s_1_2_2(nor_240_nl, mux_503_nl, fsm_output[6]);
  assign or_533_nl = (fsm_output[2]) | (fsm_output[5]) | (fsm_output[4]);
  assign mux_586_nl = MUX_s_1_2_2(not_tmp_154, or_533_nl, fsm_output[6]);
  assign mux_587_nl = MUX_s_1_2_2(or_tmp_254, mux_586_nl, fsm_output[3]);
  assign and_527_nl = (fsm_output[2:0]==3'b010) & nor_353_cse & (fsm_output[7:4]==4'b1101);
  assign COMP_LOOP_mux_28_nl = MUX_v_2_2_2(2'b01, 2'b10, and_527_nl);
  assign nl_acc_3_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[9:1])) , 1'b1}) + conv_u2u_10_11({COMP_LOOP_k_9_2_sva_6_0
      , COMP_LOOP_mux_28_nl , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[10:0];
  assign mux_597_nl = MUX_s_1_2_2((~ and_273_cse), or_604_cse, fsm_output[6]);
  assign mux_595_nl = MUX_s_1_2_2(and_273_cse, (fsm_output[5]), or_319_cse);
  assign mux_596_nl = MUX_s_1_2_2((~ mux_595_nl), or_604_cse, fsm_output[6]);
  assign mux_598_nl = MUX_s_1_2_2(mux_597_nl, mux_596_nl, fsm_output[3]);
  assign mux_599_nl = MUX_s_1_2_2(or_604_cse, (~ mux_tmp_212), and_281_cse);
  assign mux_600_nl = MUX_s_1_2_2((fsm_output[5]), mux_599_nl, fsm_output[3]);
  assign mux_602_nl = MUX_s_1_2_2(mux_tmp_212, and_273_cse, and_281_cse);
  assign mux_601_nl = MUX_s_1_2_2(and_273_cse, (fsm_output[5]), and_206_cse);
  assign mux_603_nl = MUX_s_1_2_2(mux_602_nl, mux_601_nl, fsm_output[3]);
  assign COMP_LOOP_mux_26_nl = MUX_v_64_2_2(operator_64_false_acc_mut_63_0, p_sva,
      and_dcpl_194);
  assign nor_425_nl = ~((~ (fsm_output[7])) | (fsm_output[4]) | (~ (fsm_output[0])));
  assign nor_426_nl = ~((fsm_output[7]) | (~ (fsm_output[4])) | (fsm_output[0]));
  assign mux_648_nl = MUX_s_1_2_2(nor_425_nl, nor_426_nl, fsm_output[1]);
  assign and_526_nl = (fsm_output[5]) & mux_648_nl;
  assign nor_427_nl = ~((fsm_output[5]) | (fsm_output[1]) | (fsm_output[7]) | (~
      (fsm_output[4])) | (fsm_output[0]));
  assign mux_647_nl = MUX_s_1_2_2(and_526_nl, nor_427_nl, fsm_output[8]);
  assign and_525_nl = (fsm_output[3]) & mux_647_nl;
  assign nor_428_nl = ~((fsm_output[3]) | (~ (fsm_output[8])) | (fsm_output[5]) |
      (~ (fsm_output[1])) | (~ (fsm_output[7])) | (fsm_output[4]) | (~ (fsm_output[0])));
  assign mux_646_nl = MUX_s_1_2_2(and_525_nl, nor_428_nl, fsm_output[2]);
  assign COMP_LOOP_COMP_LOOP_nand_2_nl = ~(and_dcpl_194 & (~(mux_646_nl & (fsm_output[6]))));
  assign COMP_LOOP_not_101_nl = ~ and_dcpl_194;
  assign COMP_LOOP_COMP_LOOP_nand_3_nl = ~(MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
      modulo_result_mux_1_cse, COMP_LOOP_not_101_nl));
  assign nl_acc_nl = conv_u2u_65_66({COMP_LOOP_mux_26_nl , COMP_LOOP_COMP_LOOP_nand_2_nl})
      + conv_s2u_65_66({COMP_LOOP_COMP_LOOP_nand_3_nl , 1'b1});
  assign acc_nl = nl_acc_nl[65:0];
  assign z_out = readslicef_66_65_1(acc_nl);
  assign COMP_LOOP_not_102_nl = ~ and_390_ssc;
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_52_nl = ~(MUX_v_57_2_2((operator_66_true_div_cmp_z[63:7]),
      57'b111111111111111111111111111111111111111111111111111111111, COMP_LOOP_not_102_nl));
  assign COMP_LOOP_mux_27_nl = MUX_v_7_2_2(COMP_LOOP_k_9_2_sva_6_0, (~ (operator_66_true_div_cmp_z[6:0])),
      and_390_ssc);
  assign nl_z_out_1 = ({and_390_ssc , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_52_nl , COMP_LOOP_mux_27_nl})
      + 65'b00000000000000000000000000000000000000000000000000000000000000001;
  assign z_out_1 = nl_z_out_1[64:0];
  assign operator_64_false_1_mux_2_nl = MUX_v_12_2_2(({5'b00001 , (~ COMP_LOOP_k_9_2_sva_6_0)}),
      VEC_LOOP_j_sva_11_0, and_dcpl_225);
  assign operator_64_false_1_mux_3_nl = MUX_v_10_2_2(10'b0000000001, STAGE_LOOP_lshift_psp_sva,
      and_dcpl_225);
  assign nl_z_out_2 = conv_u2u_12_13(operator_64_false_1_mux_2_nl) + conv_u2u_10_13(operator_64_false_1_mux_3_nl);
  assign z_out_2 = nl_z_out_2[12:0];
  assign COMP_LOOP_COMP_LOOP_or_4_nl = (~(and_dcpl_273 | and_dcpl_285 | and_dcpl_292
      | and_441_cse | and_dcpl_301)) | and_dcpl_281;
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_53_nl = ~((operator_64_false_acc_mut_63_0[62])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_54_nl = ~((operator_64_false_acc_mut_63_0[61])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_55_nl = ~((operator_64_false_acc_mut_63_0[60])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_56_nl = ~((operator_64_false_acc_mut_63_0[59])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_57_nl = ~((operator_64_false_acc_mut_63_0[58])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_58_nl = ~((operator_64_false_acc_mut_63_0[57])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_59_nl = ~((operator_64_false_acc_mut_63_0[56])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_60_nl = ~((operator_64_false_acc_mut_63_0[55])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_61_nl = ~((operator_64_false_acc_mut_63_0[54])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_62_nl = ~((operator_64_false_acc_mut_63_0[53])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_63_nl = ~((operator_64_false_acc_mut_63_0[52])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_64_nl = ~((operator_64_false_acc_mut_63_0[51])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_65_nl = ~((operator_64_false_acc_mut_63_0[50])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_66_nl = ~((operator_64_false_acc_mut_63_0[49])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_67_nl = ~((operator_64_false_acc_mut_63_0[48])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_68_nl = ~((operator_64_false_acc_mut_63_0[47])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_69_nl = ~((operator_64_false_acc_mut_63_0[46])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_70_nl = ~((operator_64_false_acc_mut_63_0[45])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_71_nl = ~((operator_64_false_acc_mut_63_0[44])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_72_nl = ~((operator_64_false_acc_mut_63_0[43])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_73_nl = ~((operator_64_false_acc_mut_63_0[42])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_74_nl = ~((operator_64_false_acc_mut_63_0[41])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_75_nl = ~((operator_64_false_acc_mut_63_0[40])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_76_nl = ~((operator_64_false_acc_mut_63_0[39])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_77_nl = ~((operator_64_false_acc_mut_63_0[38])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_78_nl = ~((operator_64_false_acc_mut_63_0[37])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_79_nl = ~((operator_64_false_acc_mut_63_0[36])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_80_nl = ~((operator_64_false_acc_mut_63_0[35])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_81_nl = ~((operator_64_false_acc_mut_63_0[34])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_82_nl = ~((operator_64_false_acc_mut_63_0[33])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_83_nl = ~((operator_64_false_acc_mut_63_0[32])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_84_nl = ~((operator_64_false_acc_mut_63_0[31])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_85_nl = ~((operator_64_false_acc_mut_63_0[30])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_86_nl = ~((operator_64_false_acc_mut_63_0[29])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_87_nl = ~((operator_64_false_acc_mut_63_0[28])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_88_nl = ~((operator_64_false_acc_mut_63_0[27])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_89_nl = ~((operator_64_false_acc_mut_63_0[26])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_90_nl = ~((operator_64_false_acc_mut_63_0[25])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_91_nl = ~((operator_64_false_acc_mut_63_0[24])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_92_nl = ~((operator_64_false_acc_mut_63_0[23])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_93_nl = ~((operator_64_false_acc_mut_63_0[22])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_94_nl = ~((operator_64_false_acc_mut_63_0[21])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_95_nl = ~((operator_64_false_acc_mut_63_0[20])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_96_nl = ~((operator_64_false_acc_mut_63_0[19])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_97_nl = ~((operator_64_false_acc_mut_63_0[18])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_98_nl = ~((operator_64_false_acc_mut_63_0[17])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_99_nl = ~((operator_64_false_acc_mut_63_0[16])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_100_nl = ~((operator_64_false_acc_mut_63_0[15])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_101_nl = ~((operator_64_false_acc_mut_63_0[14])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_102_nl = ~((operator_64_false_acc_mut_63_0[13])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_103_nl = ~((operator_64_false_acc_mut_63_0[12])
      | and_dcpl_273 | and_dcpl_285 | and_dcpl_292 | and_441_cse | and_dcpl_301);
  assign COMP_LOOP_mux1h_89_nl = MUX1HOT_v_12_3_2(({1'b0 , (VEC_LOOP_j_sva_11_0[11:1])}),
      (~ (operator_64_false_acc_mut_63_0[11:0])), VEC_LOOP_j_sva_11_0, {and_dcpl_273
      , and_dcpl_281 , COMP_LOOP_or_22_itm});
  assign COMP_LOOP_mux_29_nl = MUX_v_2_2_2(2'b10, 2'b01, and_441_cse);
  assign and_528_nl = and_dcpl_46 & (fsm_output[1]) & nor_353_cse & (fsm_output[6:5]==2'b11)
      & nor_399_cse;
  assign COMP_LOOP_COMP_LOOP_nor_2_nl = ~(MUX_v_2_2_2(COMP_LOOP_mux_29_nl, 2'b11,
      and_528_nl));
  assign and_529_nl = and_dcpl_26 & (~ (fsm_output[1])) & and_dcpl_257 & (fsm_output[6:5]==2'b01)
      & and_323_cse;
  assign COMP_LOOP_COMP_LOOP_or_3_nl = MUX_v_2_2_2(COMP_LOOP_COMP_LOOP_nor_2_nl,
      2'b11, and_529_nl);
  assign nl_COMP_LOOP_acc_35_nl = STAGE_LOOP_lshift_psp_sva + conv_u2u_9_10({COMP_LOOP_k_9_2_sva_6_0
      , COMP_LOOP_COMP_LOOP_or_3_nl});
  assign COMP_LOOP_acc_35_nl = nl_COMP_LOOP_acc_35_nl[9:0];
  assign COMP_LOOP_mux1h_90_nl = MUX1HOT_v_10_3_2(({2'b00 , COMP_LOOP_k_9_2_sva_6_0
      , 1'b1}), 10'b0000000001, COMP_LOOP_acc_35_nl, {and_dcpl_273 , and_dcpl_281
      , COMP_LOOP_or_22_itm});
  assign nl_z_out_5 = ({COMP_LOOP_COMP_LOOP_or_4_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_53_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_54_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_55_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_56_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_57_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_58_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_59_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_60_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_61_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_62_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_63_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_64_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_65_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_66_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_67_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_68_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_69_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_70_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_71_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_72_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_73_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_74_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_75_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_76_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_77_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_78_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_79_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_80_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_81_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_82_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_83_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_84_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_85_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_86_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_87_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_88_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_89_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_90_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_91_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_92_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_93_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_94_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_95_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_96_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_97_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_98_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_99_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_100_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_101_nl
      , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_102_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_103_nl
      , COMP_LOOP_mux1h_89_nl}) + conv_u2u_10_64(COMP_LOOP_mux1h_90_nl);
  assign z_out_5 = nl_z_out_5[63:0];
  assign not_1471_nl = ~ and_dcpl_309;
  assign COMP_LOOP_and_16_nl = MUX_v_4_2_2(4'b0000, (VEC_LOOP_j_sva_11_0[11:8]),
      not_1471_nl);
  assign COMP_LOOP_COMP_LOOP_or_5_nl = MUX_v_4_2_2(COMP_LOOP_and_16_nl, 4'b1111,
      COMP_LOOP_or_24_itm);
  assign COMP_LOOP_mux1h_91_nl = MUX1HOT_s_1_3_2((VEC_LOOP_j_sva_11_0[7]), (~ modExp_exp_1_7_1_sva),
      (~ modExp_exp_1_1_1_sva), {and_dcpl_317 , and_dcpl_320 , and_dcpl_325});
  assign COMP_LOOP_or_30_nl = COMP_LOOP_mux1h_91_nl | and_dcpl_309;
  assign COMP_LOOP_mux1h_92_nl = MUX1HOT_s_1_4_2((~ (STAGE_LOOP_lshift_psp_sva[9])),
      (VEC_LOOP_j_sva_11_0[6]), (~ modExp_exp_1_5_1_sva_1), (~ modExp_exp_1_7_1_sva),
      {and_dcpl_309 , and_dcpl_317 , and_dcpl_320 , and_dcpl_325});
  assign COMP_LOOP_mux1h_93_nl = MUX1HOT_s_1_4_2((~ (STAGE_LOOP_lshift_psp_sva[8])),
      (VEC_LOOP_j_sva_11_0[5]), (~ modExp_exp_1_5_1_sva), (~ modExp_exp_1_5_1_sva_1),
      {and_dcpl_309 , and_dcpl_317 , and_dcpl_320 , and_dcpl_325});
  assign COMP_LOOP_mux1h_94_nl = MUX1HOT_s_1_4_2((~ (STAGE_LOOP_lshift_psp_sva[7])),
      (VEC_LOOP_j_sva_11_0[4]), (~ modExp_exp_1_4_1_sva), (~ modExp_exp_1_5_1_sva),
      {and_dcpl_309 , and_dcpl_317 , and_dcpl_320 , and_dcpl_325});
  assign COMP_LOOP_mux1h_95_nl = MUX1HOT_s_1_4_2((~ (STAGE_LOOP_lshift_psp_sva[6])),
      (VEC_LOOP_j_sva_11_0[3]), (~ modExp_exp_1_3_1_sva), (~ modExp_exp_1_4_1_sva),
      {and_dcpl_309 , and_dcpl_317 , and_dcpl_320 , and_dcpl_325});
  assign COMP_LOOP_mux1h_96_nl = MUX1HOT_s_1_4_2((~ (STAGE_LOOP_lshift_psp_sva[5])),
      (VEC_LOOP_j_sva_11_0[2]), (~ modExp_exp_1_2_1_sva), (~ modExp_exp_1_3_1_sva),
      {and_dcpl_309 , and_dcpl_317 , and_dcpl_320 , and_dcpl_325});
  assign COMP_LOOP_mux1h_97_nl = MUX1HOT_s_1_4_2((~ (STAGE_LOOP_lshift_psp_sva[4])),
      (VEC_LOOP_j_sva_11_0[1]), (~ modExp_exp_1_1_1_sva), (~ modExp_exp_1_2_1_sva),
      {and_dcpl_309 , and_dcpl_317 , and_dcpl_320 , and_dcpl_325});
  assign COMP_LOOP_mux1h_98_nl = MUX1HOT_s_1_3_2((~ (STAGE_LOOP_lshift_psp_sva[3])),
      (VEC_LOOP_j_sva_11_0[0]), (~ modExp_exp_1_0_1_sva_1), {and_dcpl_309 , and_dcpl_317
      , COMP_LOOP_or_24_itm});
  assign COMP_LOOP_or_31_nl = (~(and_dcpl_317 | and_dcpl_320 | and_dcpl_325)) | and_dcpl_309;
  assign COMP_LOOP_mux1h_99_nl = MUX1HOT_v_9_3_2(({2'b00 , COMP_LOOP_k_9_2_sva_6_0}),
      ({COMP_LOOP_k_9_2_sva_6_0 , 2'b01}), 9'b000000001, {and_dcpl_309 , and_dcpl_317
      , COMP_LOOP_or_24_itm});
  assign nl_acc_6_nl = ({COMP_LOOP_COMP_LOOP_or_5_nl , COMP_LOOP_or_30_nl , COMP_LOOP_mux1h_92_nl
      , COMP_LOOP_mux1h_93_nl , COMP_LOOP_mux1h_94_nl , COMP_LOOP_mux1h_95_nl , COMP_LOOP_mux1h_96_nl
      , COMP_LOOP_mux1h_97_nl , COMP_LOOP_mux1h_98_nl , COMP_LOOP_or_31_nl}) + conv_u2u_10_13({COMP_LOOP_mux1h_99_nl
      , 1'b1});
  assign acc_6_nl = nl_acc_6_nl[12:0];
  assign z_out_6 = readslicef_13_12_1(acc_6_nl);
  assign or_694_nl = (~ (fsm_output[8])) | (fsm_output[5]) | (fsm_output[4]) | not_tmp_390;
  assign or_695_nl = (fsm_output[5:4]!=2'b10) | not_tmp_390;
  assign or_696_nl = (fsm_output[5]) | (~ (fsm_output[4])) | (fsm_output[0]) | (~
      (fsm_output[2])) | (fsm_output[7]);
  assign mux_651_nl = MUX_s_1_2_2(or_695_nl, or_696_nl, fsm_output[8]);
  assign mux_650_nl = MUX_s_1_2_2(or_694_nl, mux_651_nl, fsm_output[1]);
  assign or_698_nl = (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[2])) | (fsm_output[7]);
  assign or_699_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (fsm_output[2])
      | (fsm_output[7]);
  assign mux_652_nl = MUX_s_1_2_2(or_698_nl, or_699_nl, fsm_output[5]);
  assign or_697_nl = (fsm_output[1]) | (fsm_output[8]) | mux_652_nl;
  assign mux_649_nl = MUX_s_1_2_2(mux_650_nl, or_697_nl, fsm_output[3]);
  assign nor_429_nl = ~(mux_649_nl | (fsm_output[6]));
  assign modExp_while_if_mux_1_nl = MUX_v_64_2_2(modExp_result_sva, COMP_LOOP_1_acc_8_itm,
      nor_429_nl);
  assign nl_z_out_7 = $signed(conv_u2s_64_65(modExp_while_if_mux_1_nl)) * $signed(COMP_LOOP_1_acc_8_itm);
  assign z_out_7 = nl_z_out_7[63:0];

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_6_2;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [5:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    MUX1HOT_s_1_6_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_3_2;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [2:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    MUX1HOT_v_10_3_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_7_2;
    input [9:0] input_6;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [6:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    result = result | ( input_4 & {10{sel[4]}});
    result = result | ( input_5 & {10{sel[5]}});
    result = result | ( input_6 & {10{sel[6]}});
    MUX1HOT_v_10_7_2 = result;
  end
  endfunction


  function automatic [11:0] MUX1HOT_v_12_3_2;
    input [11:0] input_2;
    input [11:0] input_1;
    input [11:0] input_0;
    input [2:0] sel;
    reg [11:0] result;
  begin
    result = input_0 & {12{sel[0]}};
    result = result | ( input_1 & {12{sel[1]}});
    result = result | ( input_2 & {12{sel[2]}});
    MUX1HOT_v_12_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_19_2;
    input [63:0] input_18;
    input [63:0] input_17;
    input [63:0] input_16;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [18:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    result = result | ( input_16 & {64{sel[16]}});
    result = result | ( input_17 & {64{sel[17]}});
    result = result | ( input_18 & {64{sel[18]}});
    MUX1HOT_v_64_19_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_4_2;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [3:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    MUX1HOT_v_64_4_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_5_2;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [4:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    MUX1HOT_v_64_5_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_9_2;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [8:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    MUX1HOT_v_64_9_2 = result;
  end
  endfunction


  function automatic [64:0] MUX1HOT_v_65_3_2;
    input [64:0] input_2;
    input [64:0] input_1;
    input [64:0] input_0;
    input [2:0] sel;
    reg [64:0] result;
  begin
    result = input_0 & {65{sel[0]}};
    result = result | ( input_1 & {65{sel[1]}});
    result = result | ( input_2 & {65{sel[2]}});
    MUX1HOT_v_65_3_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_3_2;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [2:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    MUX1HOT_v_9_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [0:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [56:0] MUX_v_57_2_2;
    input [56:0] input_0;
    input [56:0] input_1;
    input [0:0] sel;
    reg [56:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_57_2_2 = result;
  end
  endfunction


  function automatic [62:0] MUX_v_63_2_2;
    input [62:0] input_0;
    input [62:0] input_1;
    input [0:0] sel;
    reg [62:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_63_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [64:0] MUX_v_65_2_2;
    input [64:0] input_0;
    input [64:0] input_1;
    input [0:0] sel;
    reg [64:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_65_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function automatic [11:0] readslicef_13_12_1;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_13_12_1 = tmp[11:0];
  end
  endfunction


  function automatic [0:0] readslicef_3_1_2;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_3_1_2 = tmp[0:0];
  end
  endfunction


  function automatic [64:0] readslicef_66_65_1;
    input [65:0] vector;
    reg [65:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_66_65_1 = tmp[64:0];
  end
  endfunction


  function automatic [65:0] conv_s2u_65_66 ;
    input [64:0]  vector ;
  begin
    conv_s2u_65_66 = {vector[64], vector};
  end
  endfunction


  function automatic [64:0] conv_u2s_64_65 ;
    input [63:0]  vector ;
  begin
    conv_u2s_64_65 =  {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_7_10 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_10 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_9_12 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_12 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_10_13 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_13 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [63:0] conv_u2u_10_64 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_64 = {{54{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_12_13 ;
    input [11:0]  vector ;
  begin
    conv_u2u_12_13 = {1'b0, vector};
  end
  endfunction


  function automatic [65:0] conv_u2u_65_66 ;
    input [64:0]  vector ;
  begin
    conv_u2u_65_66 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT
// ------------------------------------------------------------------


module inPlaceNTT_DIT (
  clk, rst, vec_rsc_0_0_adra, vec_rsc_0_0_da, vec_rsc_0_0_wea, vec_rsc_0_0_qa, vec_rsc_triosy_0_0_lz,
      vec_rsc_0_1_adra, vec_rsc_0_1_da, vec_rsc_0_1_wea, vec_rsc_0_1_qa, vec_rsc_triosy_0_1_lz,
      vec_rsc_0_2_adra, vec_rsc_0_2_da, vec_rsc_0_2_wea, vec_rsc_0_2_qa, vec_rsc_triosy_0_2_lz,
      vec_rsc_0_3_adra, vec_rsc_0_3_da, vec_rsc_0_3_wea, vec_rsc_0_3_qa, vec_rsc_triosy_0_3_lz,
      p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz
);
  input clk;
  input rst;
  output [9:0] vec_rsc_0_0_adra;
  output [63:0] vec_rsc_0_0_da;
  output vec_rsc_0_0_wea;
  input [63:0] vec_rsc_0_0_qa;
  output vec_rsc_triosy_0_0_lz;
  output [9:0] vec_rsc_0_1_adra;
  output [63:0] vec_rsc_0_1_da;
  output vec_rsc_0_1_wea;
  input [63:0] vec_rsc_0_1_qa;
  output vec_rsc_triosy_0_1_lz;
  output [9:0] vec_rsc_0_2_adra;
  output [63:0] vec_rsc_0_2_da;
  output vec_rsc_0_2_wea;
  input [63:0] vec_rsc_0_2_qa;
  output vec_rsc_triosy_0_2_lz;
  output [9:0] vec_rsc_0_3_adra;
  output [63:0] vec_rsc_0_3_da;
  output vec_rsc_0_3_wea;
  input [63:0] vec_rsc_0_3_qa;
  output vec_rsc_triosy_0_3_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;


  // Interconnect Declarations
  wire [63:0] vec_rsc_0_0_i_qa_d;
  wire vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_1_i_qa_d;
  wire vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_2_i_qa_d;
  wire vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_3_i_qa_d;
  wire vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [9:0] vec_rsc_0_0_i_adra_d_iff;
  wire [63:0] vec_rsc_0_0_i_da_d_iff;
  wire vec_rsc_0_0_i_wea_d_iff;
  wire vec_rsc_0_1_i_wea_d_iff;
  wire vec_rsc_0_2_i_wea_d_iff;
  wire vec_rsc_0_3_i_wea_d_iff;


  // Interconnect Declarations for Component Instantiations 
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_10_64_1024_1024_64_1_gen
      vec_rsc_0_0_i (
      .qa(vec_rsc_0_0_qa),
      .wea(vec_rsc_0_0_wea),
      .da(vec_rsc_0_0_da),
      .adra(vec_rsc_0_0_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_0_i_qa_d),
      .wea_d(vec_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_0_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_10_64_1024_1024_64_1_gen
      vec_rsc_0_1_i (
      .qa(vec_rsc_0_1_qa),
      .wea(vec_rsc_0_1_wea),
      .da(vec_rsc_0_1_da),
      .adra(vec_rsc_0_1_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_1_i_qa_d),
      .wea_d(vec_rsc_0_1_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_1_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_10_64_1024_1024_64_1_gen
      vec_rsc_0_2_i (
      .qa(vec_rsc_0_2_qa),
      .wea(vec_rsc_0_2_wea),
      .da(vec_rsc_0_2_da),
      .adra(vec_rsc_0_2_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_2_i_qa_d),
      .wea_d(vec_rsc_0_2_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_2_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_10_64_1024_1024_64_1_gen
      vec_rsc_0_3_i (
      .qa(vec_rsc_0_3_qa),
      .wea(vec_rsc_0_3_wea),
      .da(vec_rsc_0_3_da),
      .adra(vec_rsc_0_3_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_3_i_qa_d),
      .wea_d(vec_rsc_0_3_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_3_i_wea_d_iff)
    );
  inPlaceNTT_DIT_core inPlaceNTT_DIT_core_inst (
      .clk(clk),
      .rst(rst),
      .vec_rsc_triosy_0_0_lz(vec_rsc_triosy_0_0_lz),
      .vec_rsc_triosy_0_1_lz(vec_rsc_triosy_0_1_lz),
      .vec_rsc_triosy_0_2_lz(vec_rsc_triosy_0_2_lz),
      .vec_rsc_triosy_0_3_lz(vec_rsc_triosy_0_3_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_dat(r_rsc_dat),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .vec_rsc_0_0_i_qa_d(vec_rsc_0_0_i_qa_d),
      .vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_1_i_qa_d(vec_rsc_0_1_i_qa_d),
      .vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_2_i_qa_d(vec_rsc_0_2_i_qa_d),
      .vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_3_i_qa_d(vec_rsc_0_3_i_qa_d),
      .vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_0_i_adra_d_pff(vec_rsc_0_0_i_adra_d_iff),
      .vec_rsc_0_0_i_da_d_pff(vec_rsc_0_0_i_da_d_iff),
      .vec_rsc_0_0_i_wea_d_pff(vec_rsc_0_0_i_wea_d_iff),
      .vec_rsc_0_1_i_wea_d_pff(vec_rsc_0_1_i_wea_d_iff),
      .vec_rsc_0_2_i_wea_d_pff(vec_rsc_0_2_i_wea_d_iff),
      .vec_rsc_0_3_i_wea_d_pff(vec_rsc_0_3_i_wea_d_iff)
    );
endmodule



