
--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_pkg_v1 IS

COMPONENT ccs_in_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    dat    : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_in_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    dat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_in_v1;

ARCHITECTURE beh OF ccs_in_v1 IS
BEGIN

  idat <= dat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_out_dreg_pkg_v2 IS

COMPONENT mgc_out_dreg_v2
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    d        : IN  std_logic_vector(width-1 DOWNTO 0);
    z        : OUT std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_out_dreg_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_out_dreg_v2 IS
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    d        : IN  std_logic_vector(width-1 DOWNTO 0);
    z        : OUT std_logic_vector(width-1 DOWNTO 0)
  );
END mgc_out_dreg_v2;

ARCHITECTURE beh OF mgc_out_dreg_v2 IS
BEGIN

  z <= d;

END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/src/funcs.vhd 

-- a package of attributes that give verification tools a hint about
-- the function being implemented
PACKAGE attributes IS
  ATTRIBUTE CALYPTO_FUNC : string;
  ATTRIBUTE CALYPTO_DATA_ORDER : string;
end attributes;

-----------------------------------------------------------------------
-- Package that declares synthesizable functions needed for RTL output
-----------------------------------------------------------------------

LIBRARY ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

PACKAGE funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

   FUNCTION maximum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION minimum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2 : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;
   
-----------------------------------------------------------------
-- logic functions
-----------------------------------------------------------------

   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION or_v (inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- mux functions
-----------------------------------------------------------------

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC_VECTOR;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- latch functions
-----------------------------------------------------------------
   FUNCTION lat_s(dinput: STD_LOGIC       ; clk: STD_LOGIC; doutput: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- tristate functions
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC       ; control: STD_LOGIC) RETURN STD_LOGIC;
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: SIGNED  ) RETURN STD_LOGIC;

   -- RETURN 2 bits (left => lt, right => eq)
   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED;
 
   FUNCTION fabs(arg1: SIGNED  ) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "**" (l, r: UNSIGNED) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "**" (l, r: SIGNED  ) RETURN SIGNED  ;

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-- *_stdar functions use shift functions from std_logic_arith
-----------------------------------------------------------------

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;

   -----------------------------------------------------------------
   -- *_stdar functions use shift functions from std_logic_arith
   -----------------------------------------------------------------
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC;
   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE;
   --FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR ;

   FUNCTION ceil_log2(size : NATURAL) return NATURAL;
   FUNCTION bits(size : NATURAL) return NATURAL;    

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   
END funcs;


--------------------------- B O D Y ----------------------------


PACKAGE BODY funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC IS
     BEGIN IF arg1 THEN RETURN '1'; ELSE RETURN '0'; END IF; END;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
--     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;

   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
     VARIABLE result: STD_LOGIC_VECTOR(0 DOWNTO 0);
   BEGIN
     result := (0 => arg1);
     RETURN result;
   END;

   FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 > arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION minimum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 < arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;

   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := input1'LENGTH;
     ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
     ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     --synopsys translate_off
     FOR i IN len-1 DOWNTO 0 LOOP
       result(i) := resolved(input1a(i) & input2a(i));
     END LOOP;
     --synopsys translate_on
     RETURN result;
   END;

   FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED) RETURN UNSIGNED IS
   BEGIN RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

   FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED) RETURN SIGNED IS
   BEGIN RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

-----------------------------------------------------------------
-- Logic Functions
-----------------------------------------------------------------

   FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;
   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(and_v(inputs, 1)); END;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(or_v(inputs, 1)); END;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(xor_v(inputs, 1)); END;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result AND inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

   FUNCTION or_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     -- this if is added as a quick fix for a bug in catapult evaluating the loop even if inputs'LENGTH==1
     -- see dts0100971279
     IF icnt2 > 1 THEN
       FOR i IN icnt2-1 DOWNTO 1 LOOP
         inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
         result := result OR inputsx(olenM1 DOWNTO 0);
       END LOOP;
     END IF;
     RETURN result;
   END;

   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result XOR inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

-----------------------------------------------------------------
-- Muxes
-----------------------------------------------------------------
   
   FUNCTION mux_sel2_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(1 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 4;
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector( size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "01" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "10" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "11" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel3_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(2 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 8;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "001" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "010" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "011" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN "100" =>
       result := inputs0(5*size-1 DOWNTO 4*size);
     WHEN "101" =>
       result := inputs0(6*size-1 DOWNTO 5*size);
     WHEN "110" =>
       result := inputs0(7*size-1 DOWNTO 6*size);
     WHEN "111" =>
       result := inputs0(8*size-1 DOWNTO 7*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel4_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(3 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 16;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "0000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "0001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "0010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "0011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "0100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "0101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "0110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "0111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "1000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "1001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "1010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "1011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "1100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "1101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "1110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "1111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel5_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(4 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 32;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0 );
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "00001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "00010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "00011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "00100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "00101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "00110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "00111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "01000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "01001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "01010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "01011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "01100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "01101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "01110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "01111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "10000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "10001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "10010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "10011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "10100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "10101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "10110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "10111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "11000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "11001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "11010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "11011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "11100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "11101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "11110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "11111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel6_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(5 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 64;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "000001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "000010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "000011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "000100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "000101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "000110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "000111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "001000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "001001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "001010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "001011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "001100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "001101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "001110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "001111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "010000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "010001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "010010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "010011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "010100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "010101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "010110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "010111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "011000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "011001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "011010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "011011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "011100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "011101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "011110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "011111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN "100000" =>
       result := inputs0( 33*size-1 DOWNTO 32*size);
     WHEN "100001" =>
       result := inputs0( 34*size-1 DOWNTO 33*size);
     WHEN "100010" =>
       result := inputs0( 35*size-1 DOWNTO 34*size);
     WHEN "100011" =>
       result := inputs0( 36*size-1 DOWNTO 35*size);
     WHEN "100100" =>
       result := inputs0( 37*size-1 DOWNTO 36*size);
     WHEN "100101" =>
       result := inputs0( 38*size-1 DOWNTO 37*size);
     WHEN "100110" =>
       result := inputs0( 39*size-1 DOWNTO 38*size);
     WHEN "100111" =>
       result := inputs0( 40*size-1 DOWNTO 39*size);
     WHEN "101000" =>
       result := inputs0( 41*size-1 DOWNTO 40*size);
     WHEN "101001" =>
       result := inputs0( 42*size-1 DOWNTO 41*size);
     WHEN "101010" =>
       result := inputs0( 43*size-1 DOWNTO 42*size);
     WHEN "101011" =>
       result := inputs0( 44*size-1 DOWNTO 43*size);
     WHEN "101100" =>
       result := inputs0( 45*size-1 DOWNTO 44*size);
     WHEN "101101" =>
       result := inputs0( 46*size-1 DOWNTO 45*size);
     WHEN "101110" =>
       result := inputs0( 47*size-1 DOWNTO 46*size);
     WHEN "101111" =>
       result := inputs0( 48*size-1 DOWNTO 47*size);
     WHEN "110000" =>
       result := inputs0( 49*size-1 DOWNTO 48*size);
     WHEN "110001" =>
       result := inputs0( 50*size-1 DOWNTO 49*size);
     WHEN "110010" =>
       result := inputs0( 51*size-1 DOWNTO 50*size);
     WHEN "110011" =>
       result := inputs0( 52*size-1 DOWNTO 51*size);
     WHEN "110100" =>
       result := inputs0( 53*size-1 DOWNTO 52*size);
     WHEN "110101" =>
       result := inputs0( 54*size-1 DOWNTO 53*size);
     WHEN "110110" =>
       result := inputs0( 55*size-1 DOWNTO 54*size);
     WHEN "110111" =>
       result := inputs0( 56*size-1 DOWNTO 55*size);
     WHEN "111000" =>
       result := inputs0( 57*size-1 DOWNTO 56*size);
     WHEN "111001" =>
       result := inputs0( 58*size-1 DOWNTO 57*size);
     WHEN "111010" =>
       result := inputs0( 59*size-1 DOWNTO 58*size);
     WHEN "111011" =>
       result := inputs0( 60*size-1 DOWNTO 59*size);
     WHEN "111100" =>
       result := inputs0( 61*size-1 DOWNTO 60*size);
     WHEN "111101" =>
       result := inputs0( 62*size-1 DOWNTO 61*size);
     WHEN "111110" =>
       result := inputs0( 63*size-1 DOWNTO 62*size);
     WHEN "111111" =>
       result := inputs0( 64*size-1 DOWNTO 63*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS  --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2 SEVERITY FAILURE;
     --synopsys translate_on
       CASE sel IS
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0( size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1  DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0(size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
       RETURN result;
   END;
--   BEGIN RETURN mux_v(inputs, TO_STDLOGICVECTOR(sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     ALIAS    sel0   : STD_LOGIC_VECTOR( sel'LENGTH-1 DOWNTO 0 ) IS sel;

     VARIABLE sellen : INTEGER RANGE 2-sel'LENGTH TO sel'LENGTH;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2**sel'LENGTH;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
     TYPE inputs_array_type is array(natural range <>) of std_logic_vector( olen - 1 DOWNTO 0);
     VARIABLE inputs_array : inputs_array_type( 2**sel'LENGTH - 1 DOWNTO 0);
   BEGIN
     sellen := sel'LENGTH;
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2**sellen SEVERITY FAILURE;
     sellen := 2-sellen;
     --synopsys translate_on
     CASE sellen IS
     WHEN 1 =>
       CASE sel0(0) IS

       WHEN '1' 
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0(  size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1 DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0( size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
     WHEN 2 =>
       result := mux_sel2_v(inputs, not sel);
     WHEN 3 =>
       result := mux_sel3_v(inputs, not sel);
     WHEN 4 =>
       result := mux_sel4_v(inputs, not sel);
     WHEN 5 =>
       result := mux_sel5_v(inputs, not sel);
     WHEN 6 =>
       result := mux_sel6_v(inputs, not sel);
     WHEN others =>
       -- synopsys translate_off
       IF(Is_X(sel0)) THEN
         result := (others => 'X');
       ELSE
       -- synopsys translate_on
         FOR i in 0 to 2**sel'LENGTH - 1 LOOP
           inputs_array(i) := inputs0( ((i + 1) * olen) - 1  DOWNTO i*olen);
         END LOOP;
         result := inputs_array(CONV_INTEGER( (UNSIGNED(NOT sel0)) ));
       -- synopsys translate_off
       END IF;
       -- synopsys translate_on
     END CASE;
     RETURN result;
   END;

 
-----------------------------------------------------------------
-- Latches
-----------------------------------------------------------------

   FUNCTION lat_s(dinput: STD_LOGIC; clk: STD_LOGIC; doutput: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN mux_s(STD_LOGIC_VECTOR'(doutput & dinput), clk); END;

   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR ; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR ) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     --synopsys translate_off
     ASSERT dinput'LENGTH = doutput'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN mux_v(doutput & dinput, clk);
   END;

-----------------------------------------------------------------
-- Tri-States
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC; control: STD_LOGIC) RETURN STD_LOGIC IS
--   BEGIN RETURN TO_STDLOGIC(tri_v(TO_STDLOGICVECTOR(dinput), control)); END;
--
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR ; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
--     VARIABLE result: STD_LOGIC_VECTOR(dinput'range);
--   BEGIN
--     CASE control IS
--     WHEN '0' | 'L' =>
--       result := (others => 'Z');
--     WHEN '1' | 'H' =>
--       FOR i IN dinput'range LOOP
--         result(i) := to_UX01(dinput(i));
--       END LOOP;
--     WHEN others =>
--       -- synopsys translate_off
--       result := (others => 'X');
--       -- synopsys translate_on
--     END CASE;
--     RETURN result;
--   END;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;

   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     VARIABLE diff: UNSIGNED(l'LENGTH DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     diff := ('0'&l) - ('0'&r);
     RETURN diff(l'LENGTH);
   END;
   FUNCTION "<"(l, r: SIGNED  ) RETURN STD_LOGIC IS
   BEGIN
     RETURN (UNSIGNED(l) < UNSIGNED(r)) xor (l(l'LEFT) xor r(r'LEFT));
   END;

   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION "<=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">"(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;
   FUNCTION ">=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;

   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN not or_s(l xor r);
   END;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   --some functions to placate spyglass
   FUNCTION mult_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a*b;
   END mult_natural;

   FUNCTION div_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a/b;
   END div_natural;

   FUNCTION mod_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a mod b;
   END mod_natural;

   FUNCTION add_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a+b;
   END add_unsigned;

   FUNCTION sub_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a-b;
   END sub_unsigned;

   FUNCTION sub_int(a,b : INTEGER) RETURN INTEGER IS
   BEGIN
     return a-b;
   END sub_int;

   FUNCTION concat_0(b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return '0' & b;
   END concat_0;

   FUNCTION concat_uns(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a&b;
   END concat_uns;

   FUNCTION concat_vect(a,b : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     return a&b;
   END concat_vect;





   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED IS
     CONSTANT ninps : NATURAL := arg'LENGTH / width;
     ALIAS    arg0  : UNSIGNED(arg'LENGTH-1 DOWNTO 0) IS arg;
     VARIABLE result: UNSIGNED(width-1 DOWNTO 0);
     VARIABLE from  : INTEGER;
     VARIABLE dto   : INTEGER;
   BEGIN
     --synopsys translate_off
     ASSERT arg'LENGTH = width * ninps SEVERITY FAILURE;
     --synopsys translate_on
     result := (OTHERS => '0');
     FOR i IN ninps-1 DOWNTO 0 LOOP
       --result := result + arg0((i+1)*width-1 DOWNTO i*width);
       from := mult_natural((i+1), width)-1; --2.1.6.3
       dto  := mult_natural(i,width); --2.1.6.3
       result := add_unsigned(result , arg0(from DOWNTO dto) );
     END LOOP;
     RETURN result;
   END faccu;

   FUNCTION  fabs (arg1: SIGNED) RETURN UNSIGNED IS
   BEGIN
     CASE arg1(arg1'LEFT) IS
     WHEN '1'
     --synopsys translate_off
          | 'H'
     --synopsys translate_on
       =>
       RETURN UNSIGNED'("0") - UNSIGNED(arg1);
     WHEN '0'
     --synopsys translate_off
          | 'L'
     --synopsys translate_on
       =>
       RETURN UNSIGNED(arg1);
     WHEN others =>
       RETURN resolve_unsigned(UNSIGNED(arg1), UNSIGNED'("0") - UNSIGNED(arg1));
     END CASE;
   END;

   PROCEDURE divmod(l, r: UNSIGNED; rdiv, rmod: OUT UNSIGNED) IS
     CONSTANT llen: INTEGER := l'LENGTH;
     CONSTANT rlen: INTEGER := r'LENGTH;
     CONSTANT llen_plus_rlen: INTEGER := llen + rlen;
     VARIABLE lbuf: UNSIGNED(llen+rlen-1 DOWNTO 0);
     VARIABLE diff: UNSIGNED(rlen DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT rdiv'LENGTH = llen AND rmod'LENGTH = rlen SEVERITY FAILURE;
     --synopsys translate_on
     lbuf := (others => '0');
     lbuf(llen-1 DOWNTO 0) := l;
     FOR i IN rdiv'range LOOP
       diff := sub_unsigned(lbuf(llen_plus_rlen-1 DOWNTO llen-1) ,(concat_0(r)));
       rdiv(i) := not diff(rlen);
       IF diff(rlen) = '0' THEN
         lbuf(llen_plus_rlen-1 DOWNTO llen-1) := diff;
       END IF;
       lbuf(llen_plus_rlen-1 DOWNTO 1) := lbuf(llen_plus_rlen-2 DOWNTO 0);
     END LOOP;
     rmod := lbuf(llen_plus_rlen-1 DOWNTO llen);
   END divmod;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rdiv;
   END "/";

   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rmod;
   END;

   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN l MOD r; END;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rdiv := UNSIGNED'("0") - rdiv;
     END IF;
     RETURN SIGNED(rdiv); -- overflow problem "1000" / "11"
   END "/";

   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
     CONSTANT rnul: UNSIGNED(r'LENGTH-1 DOWNTO 0) := (others => '0');
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     IF rmod /= rnul AND to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rmod := UNSIGNED(r) + rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "MOD";

   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "REM";

   FUNCTION mult_unsigned(l,r : UNSIGNED) return UNSIGNED is
   BEGIN
     return l*r; 
   END mult_unsigned;

   FUNCTION "**" (l, r : UNSIGNED) RETURN UNSIGNED IS
     CONSTANT llen  : NATURAL := l'LENGTH;
     VARIABLE result: UNSIGNED(llen-1 DOWNTO 0);
     VARIABLE fak   : UNSIGNED(llen-1 DOWNTO 0);
   BEGIN
     fak := l;
     result := (others => '0'); result(0) := '1';
     FOR i IN r'reverse_range LOOP
       --was:result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(result & (result*fak)), r(i)));
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR( concat_uns(result , mult_unsigned(result,fak) )), r(i)));

       fak := mult_unsigned(fak , fak);
     END LOOP;
     RETURN result;
   END "**";

   FUNCTION "**" (l, r : SIGNED) RETURN SIGNED IS
     CONSTANT rlen  : NATURAL := r'LENGTH;
     ALIAS    r0    : SIGNED(0 TO r'LENGTH-1) IS r;
     VARIABLE result: SIGNED(l'range);
   BEGIN
     CASE r(r'LEFT) IS
     WHEN '0'
   --synopsys translate_off
          | 'L'
   --synopsys translate_on
     =>
       result := SIGNED(UNSIGNED(l) ** UNSIGNED(r0(1 TO r'LENGTH-1)));
     WHEN '1'
   --synopsys translate_off
          | 'H'
   --synopsys translate_on
     =>
       result := (others => '0');
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END "**";

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-----------------------------------------------------------------

   FUNCTION add_nat(arg1 : NATURAL; arg2 : NATURAL ) RETURN NATURAL IS
   BEGIN
     return (arg1 + arg2);
   END;
   
--   FUNCTION UNSIGNED_2_BIT_VECTOR(arg1 : NATURAL; arg2 : NATURAL ) RETURN BIT_VECTOR IS
--   BEGIN
--     return (arg1 + arg2);
--   END;
   
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(SIGNED(result), arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
        =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
        =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;


   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     --SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: NATURAL range 1 TO len;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => '0');
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         --was:temp(i2+sw) := result(i2);
         temp_idx := add_nat(i2,sw);
         temp(temp_idx) := result(i2);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: sw_range;
     VARIABLE result_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => sbit);
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         -- was: temp(i2) := result(i2+sw);
         result_idx := add_nat(i2,sw);
         temp(i2) := result(result_idx);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;


   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := arg1'LENGTH;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     VARIABLE temp: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     SUBTYPE sw_range IS NATURAL range 0 TO len-1;
     VARIABLE sw: sw_range;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     result := (others=>'0');
     result := arg1;
     sw := sdir MOD len;
     FOR i IN arg2'reverse_range LOOP
       EXIT WHEN sw = 0;
       IF signd2 AND i = arg2'LEFT THEN 
         sw := sub_int(len,sw); 
       END IF;
       -- temp := result(len-sw-1 DOWNTO 0) & result(len-1 DOWNTO len-sw)
       FOR i2 IN len-1 DOWNTO 0 LOOP
         --was: temp((i2+sw) MOD len) := result(i2);
         temp_idx := add_nat(i2,sw) MOD len;
         temp(temp_idx) := result(i2);
       END LOOP;
       result := mux_v(STD_LOGIC_VECTOR(concat_vect(result,temp)), arg2(i));
       sw := mod_natural(mult_natural(sw,2), len);
     END LOOP;
     RETURN result;
   END frot;

   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, -1); END;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, -1); END;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC IS
     CONSTANT len : INTEGER := vec'LENGTH;
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
   BEGIN
     IF index >= len OR index < 0 THEN
       RETURN 'X';
     END IF;
     RETURN vec0(index);
   END;

   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     CONSTANT indexPwidthM1 : INTEGER := index+width-1; --2.1.6.3
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
     CONSTANT xxx : STD_LOGIC_VECTOR(width-1 DOWNTO 0) := (others => 'X');
   BEGIN
     IF index+width > len OR index < 0 THEN
       RETURN xxx;
     END IF;
     RETURN vec0(indexPwidthM1 DOWNTO index);
   END;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     VARIABLE vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     CONSTANT xxx : STD_LOGIC_VECTOR(len-1 DOWNTO 0) := (others => 'X');
   BEGIN
     vec0 := vec;
     IF index >= len OR index < 0 THEN
       RETURN xxx;
     END IF;
     vec0(index) := dinput;
     RETURN vec0;
   END;

   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE IS
     VARIABLE n_b : POSITIVE;
     VARIABLE p_v : NATURAL;
   BEGIN
     p_v := p;
     FOR i IN 1 TO 32 LOOP
       p_v := div_natural(p_v,2);
       n_b := i;
       EXIT WHEN (p_v = 0);
     END LOOP;
     RETURN n_b;
   END;


--   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
--
--     CONSTANT vlen: INTEGER := vec'LENGTH;
--     CONSTANT ilen: INTEGER := dinput'LENGTH;
--     CONSTANT max_shift: INTEGER := vlen-ilen;
--     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
--     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
--     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
--     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
--     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
--     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
--   BEGIN
--     inp := (others => '0');
--     mask := (others => '0');
--
--     IF index > max_shift OR index < 0 THEN
--       RETURN xxx;
--     END IF;
--
--     shift := CONV_UNSIGNED(index, shift'LENGTH);
--     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
--     mask(ilen-1 DOWNTO 0) := ones;
--     inp := fshl(inp, shift, vlen);
--     mask := fshl(mask, shift, vlen);
--     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
--     RETURN vec0;
--   END;

   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR IS

     type enable_matrix is array (0 to enable'LENGTH-1 ) of std_logic_vector(byte_width-1 downto 0);
     CONSTANT vlen: INTEGER := vec'LENGTH;
     CONSTANT ilen: INTEGER := dinput'LENGTH;
     CONSTANT max_shift: INTEGER := vlen-ilen;
     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask2: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE enables: enable_matrix;
     VARIABLE cat_enables: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0 );
     VARIABLE lsbi : INTEGER;
     VARIABLE msbi : INTEGER;

   BEGIN
     cat_enables := (others => '0');
     lsbi := 0;
     msbi := byte_width-1;
     inp := (others => '0');
     mask := (others => '0');

     IF index > max_shift OR index < 0 THEN
       RETURN xxx;
     END IF;

     --initialize enables
     for i in 0 TO (enable'LENGTH-1) loop
       enables(i)  := (others => enable(i));
       cat_enables(msbi downto lsbi) := enables(i) ;
       lsbi := msbi+1;
       msbi := msbi+byte_width;
     end loop;


     shift := CONV_UNSIGNED(index, shift'LENGTH);
     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
     mask(ilen-1 DOWNTO 0) := UNSIGNED((STD_LOGIC_VECTOR(ones) AND cat_enables));
     inp := fshl(inp, shift, vlen);
     mask := fshl(mask, shift, vlen);
     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
     RETURN vec0;
   END;


   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;
   
   FUNCTION bits(size : NATURAL) return NATURAL is
   begin
     return ceil_log2(size);
   END;

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH) xor conv_std_logic_vector(c, s'LENGTH);
     cout := ( (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH)) or (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) or (conv_std_logic_vector(b, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) );
   END PROCEDURE csa;

   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH);
     cout := (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH));
   END PROCEDURE csha;

END funcs;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_comps.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_comps IS
 
FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
FUNCTION ceil_log2(size : NATURAL) return NATURAL;
 

COMPONENT mgc_not
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_and
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nand
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_or
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xnor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux
  GENERIC (
    width  :  NATURAL;
    ctrlw  :  NATURAL;
    p2ctrlw : NATURAL := 0
  );
  PORT (
    a: in  std_logic_vector(width*(2**ctrlw) - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw            - 1 DOWNTO 0);
    z: out std_logic_vector(width            - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux1hot
  GENERIC (
    width  : NATURAL;
    ctrlw  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ctrlw - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw       - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_reg_pos
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;  -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL  -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_reg_neg
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;   -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_generic_reg
  GENERIC(
   width: natural := 8;
   ph_clk: integer range 0 to 1 := 1; -- clock polarity, 1=rising_edge
   ph_en: integer range 0 to 1 := 1;
   ph_a_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   ph_s_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   a_rst_used: integer range 0 to 1 := 1;
   s_rst_used: integer range 0 to 1 := 0;
   en_used: integer range 0 to 1 := 1
  );
  PORT(
   d: std_logic_vector(width-1 downto 0);
   clk: in std_logic;
   en: in std_logic;
   a_rst: in std_logic;
   s_rst: in std_logic;
   q: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_equal
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a : in  std_logic_vector(width-1 DOWNTO 0);
    b : in  std_logic_vector(width-1 DOWNTO 0);
    eq: out std_logic;
    ne: out std_logic
  );
END COMPONENT;

COMPONENT mgc_shift_l
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rot
  GENERIC (
    width  : NATURAL;
    width_s: NATURAL;
    signd_s: NATURAL;      -- 0:unsigned 1:signed
    sleft  : NATURAL;      -- 0:right 1:left;
    log2w  : NATURAL := 0; -- LOG2(width)
    l2wp2  : NATURAL := 0  --2**LOG2(width)
  );
  PORT (
    a : in  std_logic_vector(width  -1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width  -1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_sub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_ci
  GENERIC (
    width_a : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width_a, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width_a, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width_a,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width_a,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_addc
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add3
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_c : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_c : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(ifeqsel(width_c,0,width,width_c)-1 DOWNTO 0);
    d: in  std_logic_vector(0 DOWNTO 0);
    e: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_sub_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addc_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     c: in std_logic_vector(0 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addsub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    add: in  std_logic;
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_accu
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_abs
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_fast
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_pipe
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2  : NATURAL;
    add_d2  : NATURAL
  );
  PORT (
    a   : in  std_logic_vector(width_a-1 DOWNTO 0);
    b   : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2  : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c   : in  std_logic_vector(width_c-1 DOWNTO 0);
    d   : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2  : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst : in  std_logic_vector(width_e-1 DOWNTO 0);
    z   : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1_pipe
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2   : NATURAL;
    add_d2   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2     : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2     : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_e-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL
  );
  PORT (
    a:   in  std_logic_vector(width_a-1 DOWNTO 0);
    b:   in  std_logic_vector(width_b-1 DOWNTO 0);
    c:   in  std_logic_vector(width_c-1 DOWNTO 0);
    cst: in  std_logic_vector(width_cst-1 DOWNTO 0);
    d:   in  std_logic_vector(width_d-1 DOWNTO 0);
    z:   out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1_pipe
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_cst-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mulacc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2acc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    add_cxd : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    d         : in  std_logic_vector(width_d-1 DOWNTO 0);
    e         : in  std_logic_vector(width_e-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_div
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mod
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rem
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_csa
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     c: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_csha
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_rom
    GENERIC (
      rom_id : natural := 1;
      size : natural := 33;
      width : natural := 32
      );
    PORT (
      data_in : std_logic_vector((size*width)-1 downto 0);
      addr : std_logic_vector(ceil_log2(size)-1 downto 0);
      data_out : out std_logic_vector(width-1 downto 0)
    );
END COMPONENT;

END mgc_comps;

PACKAGE BODY mgc_comps IS
 
   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;
 
END mgc_comps;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_rem IS
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END mgc_rem;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

USE work.funcs.all;

ARCHITECTURE beh OF mgc_rem IS
BEGIN
  z <= std_logic_vector(unsigned(a) rem unsigned(b)) WHEN signd = 0 ELSE
       std_logic_vector(  signed(a) rem   signed(b));
END beh;

--------> ../td_ccore_solutions/modulo_dev_bb61c76201db0c9669a47462bb7d006361ff_0/rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Tue Jul 20 15:24:30 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    modulo_dev_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;
USE work.mgc_comps.ALL;


ENTITY modulo_dev_core IS
  PORT(
    base_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    m_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    return_rsc_z : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    ccs_ccore_start_rsc_dat : IN STD_LOGIC;
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_srst : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC
  );
END modulo_dev_core;

ARCHITECTURE v1 OF modulo_dev_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL base_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL return_rsci_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL ccs_ccore_start_rsci_idat : STD_LOGIC;
  SIGNAL rem_13_cmp_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_1_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_2_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_3_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_4_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_5_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_6_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_7_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_8_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_9_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_10_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_11_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_1_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_2_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_3_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_4_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_5_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_6_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_7_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_8_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_9_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_10_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_11_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_1_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_2_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_3_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_4_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_5_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_6_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_7_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_8_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_9_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_10_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_11_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL acc_tmp : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL acc_1_tmp : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL and_dcpl_1 : STD_LOGIC;
  SIGNAL and_dcpl_2 : STD_LOGIC;
  SIGNAL and_dcpl_3 : STD_LOGIC;
  SIGNAL and_dcpl_4 : STD_LOGIC;
  SIGNAL and_dcpl_6 : STD_LOGIC;
  SIGNAL and_dcpl_8 : STD_LOGIC;
  SIGNAL and_dcpl_9 : STD_LOGIC;
  SIGNAL and_dcpl_11 : STD_LOGIC;
  SIGNAL and_dcpl_13 : STD_LOGIC;
  SIGNAL and_dcpl_18 : STD_LOGIC;
  SIGNAL and_dcpl_23 : STD_LOGIC;
  SIGNAL and_dcpl_28 : STD_LOGIC;
  SIGNAL and_dcpl_29 : STD_LOGIC;
  SIGNAL and_dcpl_30 : STD_LOGIC;
  SIGNAL and_dcpl_31 : STD_LOGIC;
  SIGNAL and_dcpl_33 : STD_LOGIC;
  SIGNAL and_dcpl_35 : STD_LOGIC;
  SIGNAL and_dcpl_36 : STD_LOGIC;
  SIGNAL and_dcpl_38 : STD_LOGIC;
  SIGNAL and_dcpl_40 : STD_LOGIC;
  SIGNAL and_dcpl_45 : STD_LOGIC;
  SIGNAL and_dcpl_50 : STD_LOGIC;
  SIGNAL and_dcpl_55 : STD_LOGIC;
  SIGNAL and_dcpl_56 : STD_LOGIC;
  SIGNAL and_dcpl_57 : STD_LOGIC;
  SIGNAL and_dcpl_58 : STD_LOGIC;
  SIGNAL and_dcpl_60 : STD_LOGIC;
  SIGNAL and_dcpl_62 : STD_LOGIC;
  SIGNAL and_dcpl_63 : STD_LOGIC;
  SIGNAL and_dcpl_65 : STD_LOGIC;
  SIGNAL and_dcpl_67 : STD_LOGIC;
  SIGNAL and_dcpl_72 : STD_LOGIC;
  SIGNAL and_dcpl_77 : STD_LOGIC;
  SIGNAL and_dcpl_82 : STD_LOGIC;
  SIGNAL and_dcpl_83 : STD_LOGIC;
  SIGNAL and_dcpl_84 : STD_LOGIC;
  SIGNAL and_dcpl_85 : STD_LOGIC;
  SIGNAL and_dcpl_87 : STD_LOGIC;
  SIGNAL and_dcpl_89 : STD_LOGIC;
  SIGNAL and_dcpl_90 : STD_LOGIC;
  SIGNAL and_dcpl_92 : STD_LOGIC;
  SIGNAL and_dcpl_94 : STD_LOGIC;
  SIGNAL and_dcpl_99 : STD_LOGIC;
  SIGNAL and_dcpl_104 : STD_LOGIC;
  SIGNAL and_dcpl_109 : STD_LOGIC;
  SIGNAL and_dcpl_110 : STD_LOGIC;
  SIGNAL and_dcpl_111 : STD_LOGIC;
  SIGNAL and_dcpl_112 : STD_LOGIC;
  SIGNAL and_dcpl_114 : STD_LOGIC;
  SIGNAL and_dcpl_115 : STD_LOGIC;
  SIGNAL and_dcpl_117 : STD_LOGIC;
  SIGNAL and_dcpl_119 : STD_LOGIC;
  SIGNAL and_dcpl_121 : STD_LOGIC;
  SIGNAL and_dcpl_126 : STD_LOGIC;
  SIGNAL and_dcpl_129 : STD_LOGIC;
  SIGNAL and_dcpl_136 : STD_LOGIC;
  SIGNAL and_dcpl_137 : STD_LOGIC;
  SIGNAL and_dcpl_138 : STD_LOGIC;
  SIGNAL and_dcpl_139 : STD_LOGIC;
  SIGNAL and_dcpl_141 : STD_LOGIC;
  SIGNAL and_dcpl_143 : STD_LOGIC;
  SIGNAL and_dcpl_144 : STD_LOGIC;
  SIGNAL and_dcpl_146 : STD_LOGIC;
  SIGNAL and_dcpl_148 : STD_LOGIC;
  SIGNAL and_dcpl_153 : STD_LOGIC;
  SIGNAL and_dcpl_158 : STD_LOGIC;
  SIGNAL and_dcpl_163 : STD_LOGIC;
  SIGNAL and_dcpl_164 : STD_LOGIC;
  SIGNAL and_dcpl_165 : STD_LOGIC;
  SIGNAL and_dcpl_166 : STD_LOGIC;
  SIGNAL and_dcpl_168 : STD_LOGIC;
  SIGNAL and_dcpl_170 : STD_LOGIC;
  SIGNAL and_dcpl_171 : STD_LOGIC;
  SIGNAL and_dcpl_173 : STD_LOGIC;
  SIGNAL and_dcpl_175 : STD_LOGIC;
  SIGNAL and_dcpl_180 : STD_LOGIC;
  SIGNAL and_dcpl_185 : STD_LOGIC;
  SIGNAL and_dcpl_190 : STD_LOGIC;
  SIGNAL and_dcpl_191 : STD_LOGIC;
  SIGNAL and_dcpl_192 : STD_LOGIC;
  SIGNAL and_dcpl_193 : STD_LOGIC;
  SIGNAL and_dcpl_195 : STD_LOGIC;
  SIGNAL and_dcpl_197 : STD_LOGIC;
  SIGNAL and_dcpl_198 : STD_LOGIC;
  SIGNAL and_dcpl_200 : STD_LOGIC;
  SIGNAL and_dcpl_202 : STD_LOGIC;
  SIGNAL and_dcpl_207 : STD_LOGIC;
  SIGNAL and_dcpl_212 : STD_LOGIC;
  SIGNAL and_dcpl_217 : STD_LOGIC;
  SIGNAL and_dcpl_218 : STD_LOGIC;
  SIGNAL and_dcpl_219 : STD_LOGIC;
  SIGNAL and_dcpl_220 : STD_LOGIC;
  SIGNAL and_dcpl_222 : STD_LOGIC;
  SIGNAL and_dcpl_224 : STD_LOGIC;
  SIGNAL and_dcpl_225 : STD_LOGIC;
  SIGNAL and_dcpl_227 : STD_LOGIC;
  SIGNAL and_dcpl_229 : STD_LOGIC;
  SIGNAL and_dcpl_234 : STD_LOGIC;
  SIGNAL and_dcpl_239 : STD_LOGIC;
  SIGNAL and_dcpl_244 : STD_LOGIC;
  SIGNAL and_dcpl_245 : STD_LOGIC;
  SIGNAL and_dcpl_246 : STD_LOGIC;
  SIGNAL and_dcpl_247 : STD_LOGIC;
  SIGNAL and_dcpl_249 : STD_LOGIC;
  SIGNAL and_dcpl_251 : STD_LOGIC;
  SIGNAL and_dcpl_252 : STD_LOGIC;
  SIGNAL and_dcpl_254 : STD_LOGIC;
  SIGNAL and_dcpl_256 : STD_LOGIC;
  SIGNAL and_dcpl_261 : STD_LOGIC;
  SIGNAL and_dcpl_266 : STD_LOGIC;
  SIGNAL and_dcpl_271 : STD_LOGIC;
  SIGNAL and_dcpl_272 : STD_LOGIC;
  SIGNAL and_dcpl_274 : STD_LOGIC;
  SIGNAL and_dcpl_276 : STD_LOGIC;
  SIGNAL and_dcpl_278 : STD_LOGIC;
  SIGNAL and_dcpl_280 : STD_LOGIC;
  SIGNAL and_dcpl_285 : STD_LOGIC;
  SIGNAL and_dcpl_291 : STD_LOGIC;
  SIGNAL and_dcpl_292 : STD_LOGIC;
  SIGNAL and_dcpl_293 : STD_LOGIC;
  SIGNAL and_dcpl_294 : STD_LOGIC;
  SIGNAL and_dcpl_295 : STD_LOGIC;
  SIGNAL and_dcpl_296 : STD_LOGIC;
  SIGNAL and_dcpl_298 : STD_LOGIC;
  SIGNAL not_tmp_54 : STD_LOGIC;
  SIGNAL or_tmp_2 : STD_LOGIC;
  SIGNAL and_dcpl_300 : STD_LOGIC;
  SIGNAL and_dcpl_301 : STD_LOGIC;
  SIGNAL and_dcpl_302 : STD_LOGIC;
  SIGNAL and_dcpl_304 : STD_LOGIC;
  SIGNAL and_tmp : STD_LOGIC;
  SIGNAL and_dcpl_306 : STD_LOGIC;
  SIGNAL and_dcpl_307 : STD_LOGIC;
  SIGNAL and_dcpl_308 : STD_LOGIC;
  SIGNAL and_dcpl_310 : STD_LOGIC;
  SIGNAL and_tmp_2 : STD_LOGIC;
  SIGNAL and_dcpl_312 : STD_LOGIC;
  SIGNAL and_dcpl_313 : STD_LOGIC;
  SIGNAL and_dcpl_314 : STD_LOGIC;
  SIGNAL and_dcpl_316 : STD_LOGIC;
  SIGNAL and_tmp_5 : STD_LOGIC;
  SIGNAL and_dcpl_318 : STD_LOGIC;
  SIGNAL and_tmp_9 : STD_LOGIC;
  SIGNAL and_dcpl_324 : STD_LOGIC;
  SIGNAL and_tmp_13 : STD_LOGIC;
  SIGNAL and_dcpl_330 : STD_LOGIC;
  SIGNAL mux_tmp_19 : STD_LOGIC;
  SIGNAL and_tmp_17 : STD_LOGIC;
  SIGNAL and_dcpl_336 : STD_LOGIC;
  SIGNAL mux_tmp_22 : STD_LOGIC;
  SIGNAL mux_tmp_23 : STD_LOGIC;
  SIGNAL and_tmp_21 : STD_LOGIC;
  SIGNAL and_dcpl_342 : STD_LOGIC;
  SIGNAL mux_tmp_26 : STD_LOGIC;
  SIGNAL mux_tmp_27 : STD_LOGIC;
  SIGNAL mux_tmp_28 : STD_LOGIC;
  SIGNAL and_tmp_25 : STD_LOGIC;
  SIGNAL and_dcpl_348 : STD_LOGIC;
  SIGNAL and_tmp_35 : STD_LOGIC;
  SIGNAL and_dcpl_355 : STD_LOGIC;
  SIGNAL and_dcpl_356 : STD_LOGIC;
  SIGNAL and_dcpl_358 : STD_LOGIC;
  SIGNAL or_tmp_80 : STD_LOGIC;
  SIGNAL and_dcpl_360 : STD_LOGIC;
  SIGNAL and_dcpl_362 : STD_LOGIC;
  SIGNAL mux_tmp_32 : STD_LOGIC;
  SIGNAL and_dcpl_364 : STD_LOGIC;
  SIGNAL and_dcpl_366 : STD_LOGIC;
  SIGNAL mux_tmp_34 : STD_LOGIC;
  SIGNAL mux_tmp_35 : STD_LOGIC;
  SIGNAL and_dcpl_368 : STD_LOGIC;
  SIGNAL and_dcpl_370 : STD_LOGIC;
  SIGNAL mux_tmp_37 : STD_LOGIC;
  SIGNAL mux_tmp_38 : STD_LOGIC;
  SIGNAL mux_tmp_39 : STD_LOGIC;
  SIGNAL and_dcpl_372 : STD_LOGIC;
  SIGNAL mux_tmp_41 : STD_LOGIC;
  SIGNAL mux_tmp_42 : STD_LOGIC;
  SIGNAL mux_tmp_43 : STD_LOGIC;
  SIGNAL mux_tmp_44 : STD_LOGIC;
  SIGNAL and_dcpl_376 : STD_LOGIC;
  SIGNAL mux_tmp_46 : STD_LOGIC;
  SIGNAL mux_tmp_47 : STD_LOGIC;
  SIGNAL mux_tmp_48 : STD_LOGIC;
  SIGNAL mux_tmp_49 : STD_LOGIC;
  SIGNAL mux_tmp_50 : STD_LOGIC;
  SIGNAL and_dcpl_379 : STD_LOGIC;
  SIGNAL mux_tmp_52 : STD_LOGIC;
  SIGNAL mux_tmp_53 : STD_LOGIC;
  SIGNAL mux_tmp_54 : STD_LOGIC;
  SIGNAL mux_tmp_55 : STD_LOGIC;
  SIGNAL mux_tmp_56 : STD_LOGIC;
  SIGNAL mux_tmp_57 : STD_LOGIC;
  SIGNAL and_dcpl_382 : STD_LOGIC;
  SIGNAL mux_tmp_59 : STD_LOGIC;
  SIGNAL mux_tmp_60 : STD_LOGIC;
  SIGNAL mux_tmp_61 : STD_LOGIC;
  SIGNAL mux_tmp_62 : STD_LOGIC;
  SIGNAL mux_tmp_63 : STD_LOGIC;
  SIGNAL mux_tmp_64 : STD_LOGIC;
  SIGNAL mux_tmp_65 : STD_LOGIC;
  SIGNAL and_dcpl_385 : STD_LOGIC;
  SIGNAL mux_tmp_67 : STD_LOGIC;
  SIGNAL mux_tmp_68 : STD_LOGIC;
  SIGNAL mux_tmp_69 : STD_LOGIC;
  SIGNAL mux_tmp_70 : STD_LOGIC;
  SIGNAL mux_tmp_71 : STD_LOGIC;
  SIGNAL mux_tmp_72 : STD_LOGIC;
  SIGNAL mux_tmp_73 : STD_LOGIC;
  SIGNAL mux_tmp_74 : STD_LOGIC;
  SIGNAL and_dcpl_388 : STD_LOGIC;
  SIGNAL and_tmp_44 : STD_LOGIC;
  SIGNAL mux_tmp_76 : STD_LOGIC;
  SIGNAL and_dcpl_393 : STD_LOGIC;
  SIGNAL and_dcpl_394 : STD_LOGIC;
  SIGNAL and_dcpl_395 : STD_LOGIC;
  SIGNAL or_tmp_185 : STD_LOGIC;
  SIGNAL and_dcpl_397 : STD_LOGIC;
  SIGNAL and_dcpl_398 : STD_LOGIC;
  SIGNAL and_tmp_45 : STD_LOGIC;
  SIGNAL and_dcpl_400 : STD_LOGIC;
  SIGNAL and_dcpl_401 : STD_LOGIC;
  SIGNAL and_tmp_47 : STD_LOGIC;
  SIGNAL and_dcpl_403 : STD_LOGIC;
  SIGNAL and_dcpl_404 : STD_LOGIC;
  SIGNAL and_tmp_50 : STD_LOGIC;
  SIGNAL and_dcpl_406 : STD_LOGIC;
  SIGNAL and_tmp_54 : STD_LOGIC;
  SIGNAL and_dcpl_409 : STD_LOGIC;
  SIGNAL and_tmp_58 : STD_LOGIC;
  SIGNAL and_dcpl_413 : STD_LOGIC;
  SIGNAL mux_tmp_84 : STD_LOGIC;
  SIGNAL and_tmp_62 : STD_LOGIC;
  SIGNAL and_dcpl_417 : STD_LOGIC;
  SIGNAL mux_tmp_87 : STD_LOGIC;
  SIGNAL mux_tmp_88 : STD_LOGIC;
  SIGNAL and_tmp_66 : STD_LOGIC;
  SIGNAL and_dcpl_421 : STD_LOGIC;
  SIGNAL mux_tmp_91 : STD_LOGIC;
  SIGNAL mux_tmp_92 : STD_LOGIC;
  SIGNAL mux_tmp_93 : STD_LOGIC;
  SIGNAL and_tmp_70 : STD_LOGIC;
  SIGNAL and_dcpl_425 : STD_LOGIC;
  SIGNAL and_tmp_80 : STD_LOGIC;
  SIGNAL and_dcpl_430 : STD_LOGIC;
  SIGNAL and_dcpl_431 : STD_LOGIC;
  SIGNAL or_tmp_263 : STD_LOGIC;
  SIGNAL and_dcpl_433 : STD_LOGIC;
  SIGNAL mux_tmp_97 : STD_LOGIC;
  SIGNAL and_dcpl_435 : STD_LOGIC;
  SIGNAL mux_tmp_99 : STD_LOGIC;
  SIGNAL mux_tmp_100 : STD_LOGIC;
  SIGNAL and_dcpl_437 : STD_LOGIC;
  SIGNAL mux_tmp_102 : STD_LOGIC;
  SIGNAL mux_tmp_103 : STD_LOGIC;
  SIGNAL mux_tmp_104 : STD_LOGIC;
  SIGNAL and_dcpl_439 : STD_LOGIC;
  SIGNAL mux_tmp_106 : STD_LOGIC;
  SIGNAL mux_tmp_107 : STD_LOGIC;
  SIGNAL mux_tmp_108 : STD_LOGIC;
  SIGNAL mux_tmp_109 : STD_LOGIC;
  SIGNAL and_dcpl_442 : STD_LOGIC;
  SIGNAL mux_tmp_111 : STD_LOGIC;
  SIGNAL mux_tmp_112 : STD_LOGIC;
  SIGNAL mux_tmp_113 : STD_LOGIC;
  SIGNAL mux_tmp_114 : STD_LOGIC;
  SIGNAL mux_tmp_115 : STD_LOGIC;
  SIGNAL and_dcpl_445 : STD_LOGIC;
  SIGNAL mux_tmp_117 : STD_LOGIC;
  SIGNAL mux_tmp_118 : STD_LOGIC;
  SIGNAL mux_tmp_119 : STD_LOGIC;
  SIGNAL mux_tmp_120 : STD_LOGIC;
  SIGNAL mux_tmp_121 : STD_LOGIC;
  SIGNAL mux_tmp_122 : STD_LOGIC;
  SIGNAL and_dcpl_448 : STD_LOGIC;
  SIGNAL mux_tmp_124 : STD_LOGIC;
  SIGNAL mux_tmp_125 : STD_LOGIC;
  SIGNAL mux_tmp_126 : STD_LOGIC;
  SIGNAL mux_tmp_127 : STD_LOGIC;
  SIGNAL mux_tmp_128 : STD_LOGIC;
  SIGNAL mux_tmp_129 : STD_LOGIC;
  SIGNAL mux_tmp_130 : STD_LOGIC;
  SIGNAL and_dcpl_451 : STD_LOGIC;
  SIGNAL mux_tmp_132 : STD_LOGIC;
  SIGNAL mux_tmp_133 : STD_LOGIC;
  SIGNAL mux_tmp_134 : STD_LOGIC;
  SIGNAL mux_tmp_135 : STD_LOGIC;
  SIGNAL mux_tmp_136 : STD_LOGIC;
  SIGNAL mux_tmp_137 : STD_LOGIC;
  SIGNAL mux_tmp_138 : STD_LOGIC;
  SIGNAL mux_tmp_139 : STD_LOGIC;
  SIGNAL and_dcpl_454 : STD_LOGIC;
  SIGNAL and_tmp_89 : STD_LOGIC;
  SIGNAL mux_tmp_141 : STD_LOGIC;
  SIGNAL and_dcpl_460 : STD_LOGIC;
  SIGNAL and_dcpl_461 : STD_LOGIC;
  SIGNAL and_dcpl_462 : STD_LOGIC;
  SIGNAL and_dcpl_463 : STD_LOGIC;
  SIGNAL not_tmp_332 : STD_LOGIC;
  SIGNAL or_tmp_368 : STD_LOGIC;
  SIGNAL and_dcpl_465 : STD_LOGIC;
  SIGNAL and_dcpl_466 : STD_LOGIC;
  SIGNAL and_dcpl_467 : STD_LOGIC;
  SIGNAL and_tmp_90 : STD_LOGIC;
  SIGNAL and_dcpl_469 : STD_LOGIC;
  SIGNAL and_dcpl_470 : STD_LOGIC;
  SIGNAL and_dcpl_471 : STD_LOGIC;
  SIGNAL and_tmp_92 : STD_LOGIC;
  SIGNAL and_dcpl_473 : STD_LOGIC;
  SIGNAL and_dcpl_474 : STD_LOGIC;
  SIGNAL and_dcpl_475 : STD_LOGIC;
  SIGNAL and_tmp_95 : STD_LOGIC;
  SIGNAL and_dcpl_477 : STD_LOGIC;
  SIGNAL and_tmp_99 : STD_LOGIC;
  SIGNAL and_dcpl_480 : STD_LOGIC;
  SIGNAL and_tmp_103 : STD_LOGIC;
  SIGNAL and_dcpl_483 : STD_LOGIC;
  SIGNAL mux_tmp_149 : STD_LOGIC;
  SIGNAL and_tmp_107 : STD_LOGIC;
  SIGNAL and_dcpl_486 : STD_LOGIC;
  SIGNAL mux_tmp_152 : STD_LOGIC;
  SIGNAL mux_tmp_153 : STD_LOGIC;
  SIGNAL and_tmp_111 : STD_LOGIC;
  SIGNAL and_dcpl_489 : STD_LOGIC;
  SIGNAL mux_tmp_156 : STD_LOGIC;
  SIGNAL mux_tmp_157 : STD_LOGIC;
  SIGNAL mux_tmp_158 : STD_LOGIC;
  SIGNAL and_tmp_115 : STD_LOGIC;
  SIGNAL and_dcpl_492 : STD_LOGIC;
  SIGNAL and_tmp_125 : STD_LOGIC;
  SIGNAL and_dcpl_498 : STD_LOGIC;
  SIGNAL or_tmp_446 : STD_LOGIC;
  SIGNAL and_dcpl_500 : STD_LOGIC;
  SIGNAL mux_tmp_162 : STD_LOGIC;
  SIGNAL and_dcpl_502 : STD_LOGIC;
  SIGNAL mux_tmp_164 : STD_LOGIC;
  SIGNAL mux_tmp_165 : STD_LOGIC;
  SIGNAL and_dcpl_504 : STD_LOGIC;
  SIGNAL mux_tmp_167 : STD_LOGIC;
  SIGNAL mux_tmp_168 : STD_LOGIC;
  SIGNAL mux_tmp_169 : STD_LOGIC;
  SIGNAL and_dcpl_506 : STD_LOGIC;
  SIGNAL mux_tmp_171 : STD_LOGIC;
  SIGNAL mux_tmp_172 : STD_LOGIC;
  SIGNAL mux_tmp_173 : STD_LOGIC;
  SIGNAL mux_tmp_174 : STD_LOGIC;
  SIGNAL and_dcpl_508 : STD_LOGIC;
  SIGNAL mux_tmp_176 : STD_LOGIC;
  SIGNAL mux_tmp_177 : STD_LOGIC;
  SIGNAL mux_tmp_178 : STD_LOGIC;
  SIGNAL mux_tmp_179 : STD_LOGIC;
  SIGNAL mux_tmp_180 : STD_LOGIC;
  SIGNAL and_dcpl_510 : STD_LOGIC;
  SIGNAL mux_tmp_182 : STD_LOGIC;
  SIGNAL mux_tmp_183 : STD_LOGIC;
  SIGNAL mux_tmp_184 : STD_LOGIC;
  SIGNAL mux_tmp_185 : STD_LOGIC;
  SIGNAL mux_tmp_186 : STD_LOGIC;
  SIGNAL mux_tmp_187 : STD_LOGIC;
  SIGNAL and_dcpl_512 : STD_LOGIC;
  SIGNAL mux_tmp_189 : STD_LOGIC;
  SIGNAL mux_tmp_190 : STD_LOGIC;
  SIGNAL mux_tmp_191 : STD_LOGIC;
  SIGNAL mux_tmp_192 : STD_LOGIC;
  SIGNAL mux_tmp_193 : STD_LOGIC;
  SIGNAL mux_tmp_194 : STD_LOGIC;
  SIGNAL mux_tmp_195 : STD_LOGIC;
  SIGNAL and_dcpl_514 : STD_LOGIC;
  SIGNAL mux_tmp_197 : STD_LOGIC;
  SIGNAL mux_tmp_198 : STD_LOGIC;
  SIGNAL mux_tmp_199 : STD_LOGIC;
  SIGNAL mux_tmp_200 : STD_LOGIC;
  SIGNAL mux_tmp_201 : STD_LOGIC;
  SIGNAL mux_tmp_202 : STD_LOGIC;
  SIGNAL mux_tmp_203 : STD_LOGIC;
  SIGNAL mux_tmp_204 : STD_LOGIC;
  SIGNAL and_dcpl_516 : STD_LOGIC;
  SIGNAL and_tmp_134 : STD_LOGIC;
  SIGNAL mux_tmp_206 : STD_LOGIC;
  SIGNAL and_dcpl_520 : STD_LOGIC;
  SIGNAL and_dcpl_521 : STD_LOGIC;
  SIGNAL or_tmp_551 : STD_LOGIC;
  SIGNAL and_dcpl_523 : STD_LOGIC;
  SIGNAL and_dcpl_524 : STD_LOGIC;
  SIGNAL and_tmp_135 : STD_LOGIC;
  SIGNAL and_dcpl_526 : STD_LOGIC;
  SIGNAL and_dcpl_527 : STD_LOGIC;
  SIGNAL and_tmp_137 : STD_LOGIC;
  SIGNAL and_dcpl_529 : STD_LOGIC;
  SIGNAL and_dcpl_530 : STD_LOGIC;
  SIGNAL and_tmp_140 : STD_LOGIC;
  SIGNAL and_dcpl_532 : STD_LOGIC;
  SIGNAL and_tmp_144 : STD_LOGIC;
  SIGNAL and_dcpl_534 : STD_LOGIC;
  SIGNAL and_tmp_148 : STD_LOGIC;
  SIGNAL and_dcpl_536 : STD_LOGIC;
  SIGNAL mux_tmp_214 : STD_LOGIC;
  SIGNAL and_tmp_152 : STD_LOGIC;
  SIGNAL and_dcpl_538 : STD_LOGIC;
  SIGNAL mux_tmp_217 : STD_LOGIC;
  SIGNAL mux_tmp_218 : STD_LOGIC;
  SIGNAL and_tmp_156 : STD_LOGIC;
  SIGNAL and_dcpl_540 : STD_LOGIC;
  SIGNAL mux_tmp_221 : STD_LOGIC;
  SIGNAL mux_tmp_222 : STD_LOGIC;
  SIGNAL mux_tmp_223 : STD_LOGIC;
  SIGNAL and_tmp_160 : STD_LOGIC;
  SIGNAL and_dcpl_542 : STD_LOGIC;
  SIGNAL and_tmp_170 : STD_LOGIC;
  SIGNAL and_dcpl_546 : STD_LOGIC;
  SIGNAL or_tmp_629 : STD_LOGIC;
  SIGNAL and_dcpl_548 : STD_LOGIC;
  SIGNAL mux_tmp_227 : STD_LOGIC;
  SIGNAL and_dcpl_550 : STD_LOGIC;
  SIGNAL mux_tmp_229 : STD_LOGIC;
  SIGNAL mux_tmp_230 : STD_LOGIC;
  SIGNAL and_dcpl_552 : STD_LOGIC;
  SIGNAL mux_tmp_232 : STD_LOGIC;
  SIGNAL mux_tmp_233 : STD_LOGIC;
  SIGNAL mux_tmp_234 : STD_LOGIC;
  SIGNAL and_dcpl_554 : STD_LOGIC;
  SIGNAL mux_tmp_236 : STD_LOGIC;
  SIGNAL mux_tmp_237 : STD_LOGIC;
  SIGNAL mux_tmp_238 : STD_LOGIC;
  SIGNAL mux_tmp_239 : STD_LOGIC;
  SIGNAL and_dcpl_556 : STD_LOGIC;
  SIGNAL mux_tmp_241 : STD_LOGIC;
  SIGNAL mux_tmp_242 : STD_LOGIC;
  SIGNAL mux_tmp_243 : STD_LOGIC;
  SIGNAL mux_tmp_244 : STD_LOGIC;
  SIGNAL mux_tmp_245 : STD_LOGIC;
  SIGNAL and_dcpl_558 : STD_LOGIC;
  SIGNAL mux_tmp_247 : STD_LOGIC;
  SIGNAL mux_tmp_248 : STD_LOGIC;
  SIGNAL mux_tmp_249 : STD_LOGIC;
  SIGNAL mux_tmp_250 : STD_LOGIC;
  SIGNAL mux_tmp_251 : STD_LOGIC;
  SIGNAL mux_tmp_252 : STD_LOGIC;
  SIGNAL and_dcpl_560 : STD_LOGIC;
  SIGNAL mux_tmp_254 : STD_LOGIC;
  SIGNAL mux_tmp_255 : STD_LOGIC;
  SIGNAL mux_tmp_256 : STD_LOGIC;
  SIGNAL mux_tmp_257 : STD_LOGIC;
  SIGNAL mux_tmp_258 : STD_LOGIC;
  SIGNAL mux_tmp_259 : STD_LOGIC;
  SIGNAL mux_tmp_260 : STD_LOGIC;
  SIGNAL and_dcpl_562 : STD_LOGIC;
  SIGNAL mux_tmp_262 : STD_LOGIC;
  SIGNAL mux_tmp_263 : STD_LOGIC;
  SIGNAL mux_tmp_264 : STD_LOGIC;
  SIGNAL mux_tmp_265 : STD_LOGIC;
  SIGNAL mux_tmp_266 : STD_LOGIC;
  SIGNAL mux_tmp_267 : STD_LOGIC;
  SIGNAL mux_tmp_268 : STD_LOGIC;
  SIGNAL mux_tmp_269 : STD_LOGIC;
  SIGNAL and_dcpl_564 : STD_LOGIC;
  SIGNAL and_tmp_179 : STD_LOGIC;
  SIGNAL mux_tmp_271 : STD_LOGIC;
  SIGNAL and_dcpl_568 : STD_LOGIC;
  SIGNAL and_dcpl_569 : STD_LOGIC;
  SIGNAL and_dcpl_570 : STD_LOGIC;
  SIGNAL and_dcpl_571 : STD_LOGIC;
  SIGNAL or_tmp_733 : STD_LOGIC;
  SIGNAL and_dcpl_573 : STD_LOGIC;
  SIGNAL and_dcpl_574 : STD_LOGIC;
  SIGNAL and_dcpl_575 : STD_LOGIC;
  SIGNAL and_tmp_180 : STD_LOGIC;
  SIGNAL and_dcpl_577 : STD_LOGIC;
  SIGNAL and_dcpl_578 : STD_LOGIC;
  SIGNAL and_dcpl_579 : STD_LOGIC;
  SIGNAL and_tmp_182 : STD_LOGIC;
  SIGNAL and_dcpl_581 : STD_LOGIC;
  SIGNAL and_dcpl_582 : STD_LOGIC;
  SIGNAL and_dcpl_583 : STD_LOGIC;
  SIGNAL and_tmp_185 : STD_LOGIC;
  SIGNAL and_dcpl_585 : STD_LOGIC;
  SIGNAL and_tmp_189 : STD_LOGIC;
  SIGNAL and_dcpl_589 : STD_LOGIC;
  SIGNAL and_tmp_193 : STD_LOGIC;
  SIGNAL and_dcpl_593 : STD_LOGIC;
  SIGNAL mux_tmp_279 : STD_LOGIC;
  SIGNAL and_tmp_197 : STD_LOGIC;
  SIGNAL and_dcpl_597 : STD_LOGIC;
  SIGNAL mux_tmp_282 : STD_LOGIC;
  SIGNAL mux_tmp_283 : STD_LOGIC;
  SIGNAL and_tmp_201 : STD_LOGIC;
  SIGNAL and_dcpl_601 : STD_LOGIC;
  SIGNAL mux_tmp_286 : STD_LOGIC;
  SIGNAL mux_tmp_287 : STD_LOGIC;
  SIGNAL mux_tmp_288 : STD_LOGIC;
  SIGNAL and_tmp_205 : STD_LOGIC;
  SIGNAL and_dcpl_605 : STD_LOGIC;
  SIGNAL or_tmp_808 : STD_LOGIC;
  SIGNAL mux_tmp_291 : STD_LOGIC;
  SIGNAL mux_tmp_292 : STD_LOGIC;
  SIGNAL mux_tmp_293 : STD_LOGIC;
  SIGNAL mux_tmp_294 : STD_LOGIC;
  SIGNAL mux_tmp_295 : STD_LOGIC;
  SIGNAL mux_tmp_296 : STD_LOGIC;
  SIGNAL mux_tmp_297 : STD_LOGIC;
  SIGNAL mux_tmp_298 : STD_LOGIC;
  SIGNAL and_tmp_206 : STD_LOGIC;
  SIGNAL and_dcpl_610 : STD_LOGIC;
  SIGNAL or_tmp_820 : STD_LOGIC;
  SIGNAL and_dcpl_612 : STD_LOGIC;
  SIGNAL mux_tmp_301 : STD_LOGIC;
  SIGNAL and_dcpl_614 : STD_LOGIC;
  SIGNAL mux_tmp_303 : STD_LOGIC;
  SIGNAL mux_tmp_304 : STD_LOGIC;
  SIGNAL and_dcpl_616 : STD_LOGIC;
  SIGNAL mux_tmp_306 : STD_LOGIC;
  SIGNAL mux_tmp_307 : STD_LOGIC;
  SIGNAL mux_tmp_308 : STD_LOGIC;
  SIGNAL and_dcpl_618 : STD_LOGIC;
  SIGNAL mux_tmp_310 : STD_LOGIC;
  SIGNAL mux_tmp_311 : STD_LOGIC;
  SIGNAL mux_tmp_312 : STD_LOGIC;
  SIGNAL mux_tmp_313 : STD_LOGIC;
  SIGNAL and_dcpl_622 : STD_LOGIC;
  SIGNAL mux_tmp_315 : STD_LOGIC;
  SIGNAL mux_tmp_316 : STD_LOGIC;
  SIGNAL mux_tmp_317 : STD_LOGIC;
  SIGNAL mux_tmp_318 : STD_LOGIC;
  SIGNAL mux_tmp_319 : STD_LOGIC;
  SIGNAL and_dcpl_625 : STD_LOGIC;
  SIGNAL mux_tmp_321 : STD_LOGIC;
  SIGNAL mux_tmp_322 : STD_LOGIC;
  SIGNAL mux_tmp_323 : STD_LOGIC;
  SIGNAL mux_tmp_324 : STD_LOGIC;
  SIGNAL mux_tmp_325 : STD_LOGIC;
  SIGNAL mux_tmp_326 : STD_LOGIC;
  SIGNAL and_dcpl_628 : STD_LOGIC;
  SIGNAL mux_tmp_328 : STD_LOGIC;
  SIGNAL mux_tmp_329 : STD_LOGIC;
  SIGNAL mux_tmp_330 : STD_LOGIC;
  SIGNAL mux_tmp_331 : STD_LOGIC;
  SIGNAL mux_tmp_332 : STD_LOGIC;
  SIGNAL mux_tmp_333 : STD_LOGIC;
  SIGNAL mux_tmp_334 : STD_LOGIC;
  SIGNAL and_dcpl_631 : STD_LOGIC;
  SIGNAL mux_tmp_336 : STD_LOGIC;
  SIGNAL mux_tmp_337 : STD_LOGIC;
  SIGNAL mux_tmp_338 : STD_LOGIC;
  SIGNAL mux_tmp_339 : STD_LOGIC;
  SIGNAL mux_tmp_340 : STD_LOGIC;
  SIGNAL mux_tmp_341 : STD_LOGIC;
  SIGNAL mux_tmp_342 : STD_LOGIC;
  SIGNAL mux_tmp_343 : STD_LOGIC;
  SIGNAL and_dcpl_634 : STD_LOGIC;
  SIGNAL or_tmp_921 : STD_LOGIC;
  SIGNAL mux_tmp_345 : STD_LOGIC;
  SIGNAL mux_tmp_346 : STD_LOGIC;
  SIGNAL mux_tmp_347 : STD_LOGIC;
  SIGNAL mux_tmp_348 : STD_LOGIC;
  SIGNAL mux_tmp_349 : STD_LOGIC;
  SIGNAL mux_tmp_350 : STD_LOGIC;
  SIGNAL mux_tmp_351 : STD_LOGIC;
  SIGNAL mux_tmp_352 : STD_LOGIC;
  SIGNAL mux_tmp_353 : STD_LOGIC;
  SIGNAL mux_tmp_354 : STD_LOGIC;
  SIGNAL and_dcpl_638 : STD_LOGIC;
  SIGNAL and_dcpl_639 : STD_LOGIC;
  SIGNAL or_tmp_934 : STD_LOGIC;
  SIGNAL and_dcpl_641 : STD_LOGIC;
  SIGNAL and_dcpl_642 : STD_LOGIC;
  SIGNAL and_tmp_207 : STD_LOGIC;
  SIGNAL and_dcpl_644 : STD_LOGIC;
  SIGNAL and_dcpl_645 : STD_LOGIC;
  SIGNAL and_tmp_209 : STD_LOGIC;
  SIGNAL and_dcpl_647 : STD_LOGIC;
  SIGNAL and_dcpl_648 : STD_LOGIC;
  SIGNAL and_tmp_212 : STD_LOGIC;
  SIGNAL and_dcpl_650 : STD_LOGIC;
  SIGNAL and_tmp_216 : STD_LOGIC;
  SIGNAL and_dcpl_653 : STD_LOGIC;
  SIGNAL and_tmp_220 : STD_LOGIC;
  SIGNAL and_dcpl_657 : STD_LOGIC;
  SIGNAL mux_tmp_362 : STD_LOGIC;
  SIGNAL and_tmp_224 : STD_LOGIC;
  SIGNAL and_dcpl_661 : STD_LOGIC;
  SIGNAL mux_tmp_365 : STD_LOGIC;
  SIGNAL mux_tmp_366 : STD_LOGIC;
  SIGNAL and_tmp_228 : STD_LOGIC;
  SIGNAL and_dcpl_665 : STD_LOGIC;
  SIGNAL mux_tmp_369 : STD_LOGIC;
  SIGNAL mux_tmp_370 : STD_LOGIC;
  SIGNAL mux_tmp_371 : STD_LOGIC;
  SIGNAL and_tmp_232 : STD_LOGIC;
  SIGNAL and_dcpl_669 : STD_LOGIC;
  SIGNAL or_tmp_1009 : STD_LOGIC;
  SIGNAL mux_tmp_374 : STD_LOGIC;
  SIGNAL mux_tmp_375 : STD_LOGIC;
  SIGNAL mux_tmp_376 : STD_LOGIC;
  SIGNAL mux_tmp_377 : STD_LOGIC;
  SIGNAL mux_tmp_378 : STD_LOGIC;
  SIGNAL mux_tmp_379 : STD_LOGIC;
  SIGNAL mux_tmp_380 : STD_LOGIC;
  SIGNAL mux_tmp_381 : STD_LOGIC;
  SIGNAL and_tmp_233 : STD_LOGIC;
  SIGNAL and_dcpl_673 : STD_LOGIC;
  SIGNAL or_tmp_1021 : STD_LOGIC;
  SIGNAL and_dcpl_675 : STD_LOGIC;
  SIGNAL mux_tmp_384 : STD_LOGIC;
  SIGNAL and_dcpl_677 : STD_LOGIC;
  SIGNAL mux_tmp_386 : STD_LOGIC;
  SIGNAL mux_tmp_387 : STD_LOGIC;
  SIGNAL and_dcpl_679 : STD_LOGIC;
  SIGNAL mux_tmp_389 : STD_LOGIC;
  SIGNAL mux_tmp_390 : STD_LOGIC;
  SIGNAL mux_tmp_391 : STD_LOGIC;
  SIGNAL and_dcpl_681 : STD_LOGIC;
  SIGNAL mux_tmp_393 : STD_LOGIC;
  SIGNAL mux_tmp_394 : STD_LOGIC;
  SIGNAL mux_tmp_395 : STD_LOGIC;
  SIGNAL mux_tmp_396 : STD_LOGIC;
  SIGNAL and_dcpl_684 : STD_LOGIC;
  SIGNAL mux_tmp_398 : STD_LOGIC;
  SIGNAL mux_tmp_399 : STD_LOGIC;
  SIGNAL mux_tmp_400 : STD_LOGIC;
  SIGNAL mux_tmp_401 : STD_LOGIC;
  SIGNAL mux_tmp_402 : STD_LOGIC;
  SIGNAL and_dcpl_687 : STD_LOGIC;
  SIGNAL mux_tmp_404 : STD_LOGIC;
  SIGNAL mux_tmp_405 : STD_LOGIC;
  SIGNAL mux_tmp_406 : STD_LOGIC;
  SIGNAL mux_tmp_407 : STD_LOGIC;
  SIGNAL mux_tmp_408 : STD_LOGIC;
  SIGNAL mux_tmp_409 : STD_LOGIC;
  SIGNAL and_dcpl_690 : STD_LOGIC;
  SIGNAL mux_tmp_411 : STD_LOGIC;
  SIGNAL mux_tmp_412 : STD_LOGIC;
  SIGNAL mux_tmp_413 : STD_LOGIC;
  SIGNAL mux_tmp_414 : STD_LOGIC;
  SIGNAL mux_tmp_415 : STD_LOGIC;
  SIGNAL mux_tmp_416 : STD_LOGIC;
  SIGNAL mux_tmp_417 : STD_LOGIC;
  SIGNAL and_dcpl_693 : STD_LOGIC;
  SIGNAL mux_tmp_419 : STD_LOGIC;
  SIGNAL mux_tmp_420 : STD_LOGIC;
  SIGNAL mux_tmp_421 : STD_LOGIC;
  SIGNAL mux_tmp_422 : STD_LOGIC;
  SIGNAL mux_tmp_423 : STD_LOGIC;
  SIGNAL mux_tmp_424 : STD_LOGIC;
  SIGNAL mux_tmp_425 : STD_LOGIC;
  SIGNAL mux_tmp_426 : STD_LOGIC;
  SIGNAL and_dcpl_696 : STD_LOGIC;
  SIGNAL or_tmp_1122 : STD_LOGIC;
  SIGNAL mux_tmp_428 : STD_LOGIC;
  SIGNAL mux_tmp_429 : STD_LOGIC;
  SIGNAL mux_tmp_430 : STD_LOGIC;
  SIGNAL mux_tmp_431 : STD_LOGIC;
  SIGNAL mux_tmp_432 : STD_LOGIC;
  SIGNAL mux_tmp_433 : STD_LOGIC;
  SIGNAL mux_tmp_434 : STD_LOGIC;
  SIGNAL mux_tmp_435 : STD_LOGIC;
  SIGNAL mux_tmp_436 : STD_LOGIC;
  SIGNAL mux_tmp_437 : STD_LOGIC;
  SIGNAL rem_12cyc_st_10_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_10_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_9_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_9_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_8_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_8_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_7_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_7_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_6_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_6_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_5_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_5_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_4_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_4_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_3_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_3_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_2_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_2_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_12_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL result_sva_duc : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12cyc_st_12_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL asn_itm_12 : STD_LOGIC;
  SIGNAL main_stage_0_13 : STD_LOGIC;
  SIGNAL main_stage_0_3 : STD_LOGIC;
  SIGNAL asn_itm_1 : STD_LOGIC;
  SIGNAL main_stage_0_2 : STD_LOGIC;
  SIGNAL main_stage_0_4 : STD_LOGIC;
  SIGNAL asn_itm_2 : STD_LOGIC;
  SIGNAL main_stage_0_5 : STD_LOGIC;
  SIGNAL asn_itm_3 : STD_LOGIC;
  SIGNAL main_stage_0_6 : STD_LOGIC;
  SIGNAL asn_itm_4 : STD_LOGIC;
  SIGNAL asn_itm_5 : STD_LOGIC;
  SIGNAL main_stage_0_8 : STD_LOGIC;
  SIGNAL asn_itm_7 : STD_LOGIC;
  SIGNAL main_stage_0_9 : STD_LOGIC;
  SIGNAL asn_itm_8 : STD_LOGIC;
  SIGNAL main_stage_0_10 : STD_LOGIC;
  SIGNAL asn_itm_9 : STD_LOGIC;
  SIGNAL main_stage_0_7 : STD_LOGIC;
  SIGNAL asn_itm_6 : STD_LOGIC;
  SIGNAL main_stage_0_11 : STD_LOGIC;
  SIGNAL asn_itm_10 : STD_LOGIC;
  SIGNAL and_1173_cse : STD_LOGIC;
  SIGNAL and_1175_cse : STD_LOGIC;
  SIGNAL and_1177_cse : STD_LOGIC;
  SIGNAL and_1179_cse : STD_LOGIC;
  SIGNAL and_1181_cse : STD_LOGIC;
  SIGNAL and_1183_cse : STD_LOGIC;
  SIGNAL and_1185_cse : STD_LOGIC;
  SIGNAL and_1187_cse : STD_LOGIC;
  SIGNAL and_1189_cse : STD_LOGIC;
  SIGNAL and_1191_cse : STD_LOGIC;
  SIGNAL and_1193_cse : STD_LOGIC;
  SIGNAL and_1195_cse : STD_LOGIC;
  SIGNAL and_1197_cse : STD_LOGIC;
  SIGNAL or_1_cse : STD_LOGIC;
  SIGNAL or_6_cse : STD_LOGIC;
  SIGNAL or_10_cse : STD_LOGIC;
  SIGNAL or_15_cse : STD_LOGIC;
  SIGNAL or_21_cse : STD_LOGIC;
  SIGNAL or_28_cse : STD_LOGIC;
  SIGNAL or_37_cse : STD_LOGIC;
  SIGNAL or_48_cse : STD_LOGIC;
  SIGNAL or_83_cse : STD_LOGIC;
  SIGNAL nand_276_cse : STD_LOGIC;
  SIGNAL or_88_cse : STD_LOGIC;
  SIGNAL nand_274_cse : STD_LOGIC;
  SIGNAL or_93_cse : STD_LOGIC;
  SIGNAL nand_271_cse : STD_LOGIC;
  SIGNAL or_100_cse : STD_LOGIC;
  SIGNAL nand_267_cse : STD_LOGIC;
  SIGNAL or_109_cse : STD_LOGIC;
  SIGNAL or_120_cse : STD_LOGIC;
  SIGNAL or_133_cse : STD_LOGIC;
  SIGNAL or_148_cse : STD_LOGIC;
  SIGNAL or_190_cse : STD_LOGIC;
  SIGNAL or_195_cse : STD_LOGIC;
  SIGNAL or_199_cse : STD_LOGIC;
  SIGNAL or_204_cse : STD_LOGIC;
  SIGNAL or_210_cse : STD_LOGIC;
  SIGNAL or_217_cse : STD_LOGIC;
  SIGNAL or_226_cse : STD_LOGIC;
  SIGNAL or_237_cse : STD_LOGIC;
  SIGNAL or_270_cse : STD_LOGIC;
  SIGNAL or_275_cse : STD_LOGIC;
  SIGNAL or_280_cse : STD_LOGIC;
  SIGNAL or_287_cse : STD_LOGIC;
  SIGNAL or_296_cse : STD_LOGIC;
  SIGNAL or_307_cse : STD_LOGIC;
  SIGNAL or_320_cse : STD_LOGIC;
  SIGNAL or_335_cse : STD_LOGIC;
  SIGNAL nand_281_cse : STD_LOGIC;
  SIGNAL or_377_cse : STD_LOGIC;
  SIGNAL or_382_cse : STD_LOGIC;
  SIGNAL or_386_cse : STD_LOGIC;
  SIGNAL or_391_cse : STD_LOGIC;
  SIGNAL or_397_cse : STD_LOGIC;
  SIGNAL nand_215_cse : STD_LOGIC;
  SIGNAL or_404_cse : STD_LOGIC;
  SIGNAL nand_212_cse : STD_LOGIC;
  SIGNAL or_413_cse : STD_LOGIC;
  SIGNAL nand_208_cse : STD_LOGIC;
  SIGNAL or_424_cse : STD_LOGIC;
  SIGNAL or_458_cse : STD_LOGIC;
  SIGNAL or_463_cse : STD_LOGIC;
  SIGNAL nand_198_cse : STD_LOGIC;
  SIGNAL or_468_cse : STD_LOGIC;
  SIGNAL or_475_cse : STD_LOGIC;
  SIGNAL nand_189_cse : STD_LOGIC;
  SIGNAL or_484_cse : STD_LOGIC;
  SIGNAL or_495_cse : STD_LOGIC;
  SIGNAL or_508_cse : STD_LOGIC;
  SIGNAL nand_203_cse : STD_LOGIC;
  SIGNAL or_523_cse : STD_LOGIC;
  SIGNAL nand_250_cse : STD_LOGIC;
  SIGNAL or_564_cse : STD_LOGIC;
  SIGNAL or_569_cse : STD_LOGIC;
  SIGNAL or_573_cse : STD_LOGIC;
  SIGNAL or_578_cse : STD_LOGIC;
  SIGNAL or_584_cse : STD_LOGIC;
  SIGNAL or_591_cse : STD_LOGIC;
  SIGNAL or_600_cse : STD_LOGIC;
  SIGNAL or_611_cse : STD_LOGIC;
  SIGNAL or_643_cse : STD_LOGIC;
  SIGNAL or_648_cse : STD_LOGIC;
  SIGNAL or_653_cse : STD_LOGIC;
  SIGNAL or_660_cse : STD_LOGIC;
  SIGNAL or_669_cse : STD_LOGIC;
  SIGNAL or_680_cse : STD_LOGIC;
  SIGNAL or_693_cse : STD_LOGIC;
  SIGNAL or_708_cse : STD_LOGIC;
  SIGNAL or_748_cse : STD_LOGIC;
  SIGNAL or_753_cse : STD_LOGIC;
  SIGNAL or_757_cse : STD_LOGIC;
  SIGNAL or_762_cse : STD_LOGIC;
  SIGNAL or_768_cse : STD_LOGIC;
  SIGNAL or_775_cse : STD_LOGIC;
  SIGNAL or_784_cse : STD_LOGIC;
  SIGNAL or_795_cse : STD_LOGIC;
  SIGNAL or_837_cse : STD_LOGIC;
  SIGNAL nand_84_cse : STD_LOGIC;
  SIGNAL or_842_cse : STD_LOGIC;
  SIGNAL or_847_cse : STD_LOGIC;
  SIGNAL nand_79_cse : STD_LOGIC;
  SIGNAL or_854_cse : STD_LOGIC;
  SIGNAL or_863_cse : STD_LOGIC;
  SIGNAL or_874_cse : STD_LOGIC;
  SIGNAL or_887_cse : STD_LOGIC;
  SIGNAL or_902_cse : STD_LOGIC;
  SIGNAL or_952_cse : STD_LOGIC;
  SIGNAL or_957_cse : STD_LOGIC;
  SIGNAL or_961_cse : STD_LOGIC;
  SIGNAL or_966_cse : STD_LOGIC;
  SIGNAL or_972_cse : STD_LOGIC;
  SIGNAL or_979_cse : STD_LOGIC;
  SIGNAL or_988_cse : STD_LOGIC;
  SIGNAL or_999_cse : STD_LOGIC;
  SIGNAL nand_57_cse : STD_LOGIC;
  SIGNAL or_1045_cse : STD_LOGIC;
  SIGNAL or_1050_cse : STD_LOGIC;
  SIGNAL or_1057_cse : STD_LOGIC;
  SIGNAL or_1066_cse : STD_LOGIC;
  SIGNAL nand_36_cse : STD_LOGIC;
  SIGNAL nand_29_cse : STD_LOGIC;
  SIGNAL nand_21_cse : STD_LOGIC;
  SIGNAL nand_222_cse : STD_LOGIC;
  SIGNAL nand_223_cse : STD_LOGIC;
  SIGNAL main_stage_0_12 : STD_LOGIC;
  SIGNAL m_buf_sva_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_11 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_12 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL asn_itm_11 : STD_LOGIC;
  SIGNAL mut_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12cyc_st_11_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_11_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL result_sva_duc_mx0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL and_1203_cse : STD_LOGIC;
  SIGNAL and_1205_cse : STD_LOGIC;
  SIGNAL and_1207_cse : STD_LOGIC;
  SIGNAL and_1209_cse : STD_LOGIC;
  SIGNAL and_1211_cse : STD_LOGIC;
  SIGNAL and_1213_cse : STD_LOGIC;
  SIGNAL and_1215_cse : STD_LOGIC;
  SIGNAL and_1217_cse : STD_LOGIC;
  SIGNAL and_1219_cse : STD_LOGIC;
  SIGNAL and_1221_cse : STD_LOGIC;
  SIGNAL and_1223_cse : STD_LOGIC;
  SIGNAL and_1225_cse : STD_LOGIC;
  SIGNAL and_1227_cse : STD_LOGIC;
  SIGNAL and_1229_cse : STD_LOGIC;
  SIGNAL and_1231_cse : STD_LOGIC;
  SIGNAL and_1233_cse : STD_LOGIC;
  SIGNAL and_1235_cse : STD_LOGIC;
  SIGNAL and_1237_cse : STD_LOGIC;
  SIGNAL and_1239_cse : STD_LOGIC;
  SIGNAL and_1241_cse : STD_LOGIC;
  SIGNAL and_1243_cse : STD_LOGIC;
  SIGNAL and_1245_cse : STD_LOGIC;
  SIGNAL and_1247_cse : STD_LOGIC;
  SIGNAL and_1249_cse : STD_LOGIC;
  SIGNAL and_1251_cse : STD_LOGIC;
  SIGNAL and_1253_cse : STD_LOGIC;
  SIGNAL and_1255_cse : STD_LOGIC;
  SIGNAL and_1257_cse : STD_LOGIC;
  SIGNAL and_1259_cse : STD_LOGIC;
  SIGNAL and_1261_cse : STD_LOGIC;
  SIGNAL and_1263_cse : STD_LOGIC;
  SIGNAL and_1265_cse : STD_LOGIC;
  SIGNAL and_1267_cse : STD_LOGIC;
  SIGNAL and_1269_cse : STD_LOGIC;
  SIGNAL and_1271_cse : STD_LOGIC;
  SIGNAL and_1273_cse : STD_LOGIC;
  SIGNAL and_1275_cse : STD_LOGIC;
  SIGNAL and_1277_cse : STD_LOGIC;
  SIGNAL and_1279_cse : STD_LOGIC;
  SIGNAL and_1281_cse : STD_LOGIC;
  SIGNAL and_1283_cse : STD_LOGIC;
  SIGNAL and_1285_cse : STD_LOGIC;
  SIGNAL and_1287_cse : STD_LOGIC;
  SIGNAL and_1289_cse : STD_LOGIC;
  SIGNAL and_1291_cse : STD_LOGIC;
  SIGNAL and_1293_cse : STD_LOGIC;
  SIGNAL and_1295_cse : STD_LOGIC;
  SIGNAL and_1297_cse : STD_LOGIC;
  SIGNAL and_1299_cse : STD_LOGIC;
  SIGNAL and_1301_cse : STD_LOGIC;
  SIGNAL and_1303_cse : STD_LOGIC;
  SIGNAL and_1305_cse : STD_LOGIC;
  SIGNAL and_1307_cse : STD_LOGIC;
  SIGNAL and_1309_cse : STD_LOGIC;
  SIGNAL and_1311_cse : STD_LOGIC;
  SIGNAL and_1313_cse : STD_LOGIC;
  SIGNAL and_1315_cse : STD_LOGIC;
  SIGNAL and_1317_cse : STD_LOGIC;
  SIGNAL and_1319_cse : STD_LOGIC;
  SIGNAL and_1321_cse : STD_LOGIC;
  SIGNAL and_1323_cse : STD_LOGIC;
  SIGNAL and_1325_cse : STD_LOGIC;
  SIGNAL and_1327_cse : STD_LOGIC;
  SIGNAL and_1329_cse : STD_LOGIC;
  SIGNAL and_1331_cse : STD_LOGIC;
  SIGNAL and_1333_cse : STD_LOGIC;
  SIGNAL and_1335_cse : STD_LOGIC;
  SIGNAL and_1337_cse : STD_LOGIC;
  SIGNAL and_1339_cse : STD_LOGIC;
  SIGNAL and_1341_cse : STD_LOGIC;
  SIGNAL and_1343_cse : STD_LOGIC;
  SIGNAL and_1345_cse : STD_LOGIC;
  SIGNAL and_1347_cse : STD_LOGIC;
  SIGNAL and_1349_cse : STD_LOGIC;
  SIGNAL and_1351_cse : STD_LOGIC;
  SIGNAL and_1353_cse : STD_LOGIC;
  SIGNAL and_1355_cse : STD_LOGIC;
  SIGNAL and_1357_cse : STD_LOGIC;
  SIGNAL and_1359_cse : STD_LOGIC;
  SIGNAL and_1361_cse : STD_LOGIC;
  SIGNAL and_1363_cse : STD_LOGIC;
  SIGNAL and_1365_cse : STD_LOGIC;
  SIGNAL and_1367_cse : STD_LOGIC;
  SIGNAL and_1369_cse : STD_LOGIC;
  SIGNAL and_1371_cse : STD_LOGIC;
  SIGNAL and_1373_cse : STD_LOGIC;
  SIGNAL and_1375_cse : STD_LOGIC;
  SIGNAL and_1377_cse : STD_LOGIC;
  SIGNAL and_1379_cse : STD_LOGIC;
  SIGNAL and_1381_cse : STD_LOGIC;
  SIGNAL and_1383_cse : STD_LOGIC;
  SIGNAL and_1385_cse : STD_LOGIC;
  SIGNAL and_1387_cse : STD_LOGIC;
  SIGNAL and_1389_cse : STD_LOGIC;
  SIGNAL and_1391_cse : STD_LOGIC;
  SIGNAL and_1393_cse : STD_LOGIC;
  SIGNAL and_1395_cse : STD_LOGIC;
  SIGNAL and_1397_cse : STD_LOGIC;
  SIGNAL and_1399_cse : STD_LOGIC;
  SIGNAL and_1401_cse : STD_LOGIC;
  SIGNAL and_1403_cse : STD_LOGIC;
  SIGNAL and_1405_cse : STD_LOGIC;
  SIGNAL and_1407_cse : STD_LOGIC;
  SIGNAL and_1409_cse : STD_LOGIC;
  SIGNAL and_1411_cse : STD_LOGIC;
  SIGNAL and_1413_cse : STD_LOGIC;
  SIGNAL and_1415_cse : STD_LOGIC;
  SIGNAL and_1417_cse : STD_LOGIC;
  SIGNAL and_1419_cse : STD_LOGIC;
  SIGNAL and_1421_cse : STD_LOGIC;
  SIGNAL and_1423_cse : STD_LOGIC;
  SIGNAL and_1425_cse : STD_LOGIC;
  SIGNAL and_1427_cse : STD_LOGIC;
  SIGNAL and_1429_cse : STD_LOGIC;
  SIGNAL and_1431_cse : STD_LOGIC;
  SIGNAL and_1433_cse : STD_LOGIC;
  SIGNAL and_1435_cse : STD_LOGIC;
  SIGNAL and_1437_cse : STD_LOGIC;
  SIGNAL and_1439_cse : STD_LOGIC;
  SIGNAL and_1441_cse : STD_LOGIC;
  SIGNAL and_1443_cse : STD_LOGIC;
  SIGNAL and_1445_cse : STD_LOGIC;
  SIGNAL and_1447_cse : STD_LOGIC;
  SIGNAL and_1449_cse : STD_LOGIC;
  SIGNAL and_1451_cse : STD_LOGIC;
  SIGNAL and_1453_cse : STD_LOGIC;
  SIGNAL and_1455_cse : STD_LOGIC;
  SIGNAL and_1457_cse : STD_LOGIC;
  SIGNAL and_1459_cse : STD_LOGIC;
  SIGNAL and_1461_cse : STD_LOGIC;
  SIGNAL and_1463_cse : STD_LOGIC;

  SIGNAL qelse_acc_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mux_13_nl : STD_LOGIC;
  SIGNAL mux_12_nl : STD_LOGIC;
  SIGNAL mux_11_nl : STD_LOGIC;
  SIGNAL mux_10_nl : STD_LOGIC;
  SIGNAL mux_9_nl : STD_LOGIC;
  SIGNAL mux_8_nl : STD_LOGIC;
  SIGNAL mux_7_nl : STD_LOGIC;
  SIGNAL mux_6_nl : STD_LOGIC;
  SIGNAL mux_5_nl : STD_LOGIC;
  SIGNAL mux_4_nl : STD_LOGIC;
  SIGNAL mux_3_nl : STD_LOGIC;
  SIGNAL mux_2_nl : STD_LOGIC;
  SIGNAL and_273_nl : STD_LOGIC;
  SIGNAL and_275_nl : STD_LOGIC;
  SIGNAL and_277_nl : STD_LOGIC;
  SIGNAL and_279_nl : STD_LOGIC;
  SIGNAL and_281_nl : STD_LOGIC;
  SIGNAL and_282_nl : STD_LOGIC;
  SIGNAL and_283_nl : STD_LOGIC;
  SIGNAL and_284_nl : STD_LOGIC;
  SIGNAL and_286_nl : STD_LOGIC;
  SIGNAL and_287_nl : STD_LOGIC;
  SIGNAL and_288_nl : STD_LOGIC;
  SIGNAL and_289_nl : STD_LOGIC;
  SIGNAL and_290_nl : STD_LOGIC;
  SIGNAL xor_nl : STD_LOGIC;
  SIGNAL nor_nl : STD_LOGIC;
  SIGNAL mux_14_nl : STD_LOGIC;
  SIGNAL nor_518_nl : STD_LOGIC;
  SIGNAL mux_15_nl : STD_LOGIC;
  SIGNAL nor_517_nl : STD_LOGIC;
  SIGNAL mux_16_nl : STD_LOGIC;
  SIGNAL nor_516_nl : STD_LOGIC;
  SIGNAL mux_17_nl : STD_LOGIC;
  SIGNAL nor_515_nl : STD_LOGIC;
  SIGNAL mux_18_nl : STD_LOGIC;
  SIGNAL nor_514_nl : STD_LOGIC;
  SIGNAL mux_19_nl : STD_LOGIC;
  SIGNAL nor_512_nl : STD_LOGIC;
  SIGNAL mux_20_nl : STD_LOGIC;
  SIGNAL nor_513_nl : STD_LOGIC;
  SIGNAL nor_509_nl : STD_LOGIC;
  SIGNAL mux_22_nl : STD_LOGIC;
  SIGNAL nor_510_nl : STD_LOGIC;
  SIGNAL mux_23_nl : STD_LOGIC;
  SIGNAL nor_511_nl : STD_LOGIC;
  SIGNAL nor_505_nl : STD_LOGIC;
  SIGNAL nor_506_nl : STD_LOGIC;
  SIGNAL mux_26_nl : STD_LOGIC;
  SIGNAL nor_507_nl : STD_LOGIC;
  SIGNAL mux_27_nl : STD_LOGIC;
  SIGNAL nor_508_nl : STD_LOGIC;
  SIGNAL nor_500_nl : STD_LOGIC;
  SIGNAL or_61_nl : STD_LOGIC;
  SIGNAL nor_501_nl : STD_LOGIC;
  SIGNAL nor_502_nl : STD_LOGIC;
  SIGNAL mux_31_nl : STD_LOGIC;
  SIGNAL nor_503_nl : STD_LOGIC;
  SIGNAL mux_32_nl : STD_LOGIC;
  SIGNAL nor_504_nl : STD_LOGIC;
  SIGNAL mux_33_nl : STD_LOGIC;
  SIGNAL nor_499_nl : STD_LOGIC;
  SIGNAL and_1168_nl : STD_LOGIC;
  SIGNAL mux_35_nl : STD_LOGIC;
  SIGNAL nor_498_nl : STD_LOGIC;
  SIGNAL and_1166_nl : STD_LOGIC;
  SIGNAL and_1167_nl : STD_LOGIC;
  SIGNAL mux_38_nl : STD_LOGIC;
  SIGNAL nor_497_nl : STD_LOGIC;
  SIGNAL and_1163_nl : STD_LOGIC;
  SIGNAL and_1164_nl : STD_LOGIC;
  SIGNAL and_1165_nl : STD_LOGIC;
  SIGNAL mux_42_nl : STD_LOGIC;
  SIGNAL nor_496_nl : STD_LOGIC;
  SIGNAL and_1159_nl : STD_LOGIC;
  SIGNAL and_1160_nl : STD_LOGIC;
  SIGNAL and_1161_nl : STD_LOGIC;
  SIGNAL and_1162_nl : STD_LOGIC;
  SIGNAL mux_47_nl : STD_LOGIC;
  SIGNAL nor_495_nl : STD_LOGIC;
  SIGNAL nor_493_nl : STD_LOGIC;
  SIGNAL and_1155_nl : STD_LOGIC;
  SIGNAL and_1156_nl : STD_LOGIC;
  SIGNAL and_1157_nl : STD_LOGIC;
  SIGNAL and_1158_nl : STD_LOGIC;
  SIGNAL mux_53_nl : STD_LOGIC;
  SIGNAL nor_494_nl : STD_LOGIC;
  SIGNAL nor_490_nl : STD_LOGIC;
  SIGNAL nor_491_nl : STD_LOGIC;
  SIGNAL and_1151_nl : STD_LOGIC;
  SIGNAL and_1152_nl : STD_LOGIC;
  SIGNAL and_1153_nl : STD_LOGIC;
  SIGNAL and_1154_nl : STD_LOGIC;
  SIGNAL mux_60_nl : STD_LOGIC;
  SIGNAL nor_492_nl : STD_LOGIC;
  SIGNAL nor_486_nl : STD_LOGIC;
  SIGNAL nor_487_nl : STD_LOGIC;
  SIGNAL nor_488_nl : STD_LOGIC;
  SIGNAL and_1147_nl : STD_LOGIC;
  SIGNAL and_1148_nl : STD_LOGIC;
  SIGNAL and_1149_nl : STD_LOGIC;
  SIGNAL and_1150_nl : STD_LOGIC;
  SIGNAL mux_68_nl : STD_LOGIC;
  SIGNAL nor_489_nl : STD_LOGIC;
  SIGNAL nor_481_nl : STD_LOGIC;
  SIGNAL or_165_nl : STD_LOGIC;
  SIGNAL nor_482_nl : STD_LOGIC;
  SIGNAL nor_483_nl : STD_LOGIC;
  SIGNAL nor_484_nl : STD_LOGIC;
  SIGNAL and_1143_nl : STD_LOGIC;
  SIGNAL and_1144_nl : STD_LOGIC;
  SIGNAL and_1145_nl : STD_LOGIC;
  SIGNAL and_1146_nl : STD_LOGIC;
  SIGNAL mux_77_nl : STD_LOGIC;
  SIGNAL nor_485_nl : STD_LOGIC;
  SIGNAL nor_480_nl : STD_LOGIC;
  SIGNAL or_175_nl : STD_LOGIC;
  SIGNAL mux_79_nl : STD_LOGIC;
  SIGNAL nor_479_nl : STD_LOGIC;
  SIGNAL mux_80_nl : STD_LOGIC;
  SIGNAL nor_478_nl : STD_LOGIC;
  SIGNAL mux_81_nl : STD_LOGIC;
  SIGNAL nor_477_nl : STD_LOGIC;
  SIGNAL mux_82_nl : STD_LOGIC;
  SIGNAL nor_476_nl : STD_LOGIC;
  SIGNAL mux_83_nl : STD_LOGIC;
  SIGNAL nor_475_nl : STD_LOGIC;
  SIGNAL mux_84_nl : STD_LOGIC;
  SIGNAL nor_473_nl : STD_LOGIC;
  SIGNAL mux_85_nl : STD_LOGIC;
  SIGNAL nor_474_nl : STD_LOGIC;
  SIGNAL nor_470_nl : STD_LOGIC;
  SIGNAL mux_87_nl : STD_LOGIC;
  SIGNAL nor_471_nl : STD_LOGIC;
  SIGNAL mux_88_nl : STD_LOGIC;
  SIGNAL nor_472_nl : STD_LOGIC;
  SIGNAL nor_466_nl : STD_LOGIC;
  SIGNAL nor_467_nl : STD_LOGIC;
  SIGNAL mux_91_nl : STD_LOGIC;
  SIGNAL nor_468_nl : STD_LOGIC;
  SIGNAL mux_92_nl : STD_LOGIC;
  SIGNAL nor_469_nl : STD_LOGIC;
  SIGNAL nor_461_nl : STD_LOGIC;
  SIGNAL or_250_nl : STD_LOGIC;
  SIGNAL nor_462_nl : STD_LOGIC;
  SIGNAL nor_463_nl : STD_LOGIC;
  SIGNAL mux_96_nl : STD_LOGIC;
  SIGNAL nor_464_nl : STD_LOGIC;
  SIGNAL mux_97_nl : STD_LOGIC;
  SIGNAL nor_465_nl : STD_LOGIC;
  SIGNAL mux_98_nl : STD_LOGIC;
  SIGNAL nor_460_nl : STD_LOGIC;
  SIGNAL and_1142_nl : STD_LOGIC;
  SIGNAL mux_100_nl : STD_LOGIC;
  SIGNAL nor_459_nl : STD_LOGIC;
  SIGNAL and_1140_nl : STD_LOGIC;
  SIGNAL and_1141_nl : STD_LOGIC;
  SIGNAL mux_103_nl : STD_LOGIC;
  SIGNAL nor_458_nl : STD_LOGIC;
  SIGNAL and_1137_nl : STD_LOGIC;
  SIGNAL and_1138_nl : STD_LOGIC;
  SIGNAL and_1139_nl : STD_LOGIC;
  SIGNAL mux_107_nl : STD_LOGIC;
  SIGNAL nor_457_nl : STD_LOGIC;
  SIGNAL and_1133_nl : STD_LOGIC;
  SIGNAL and_1134_nl : STD_LOGIC;
  SIGNAL and_1135_nl : STD_LOGIC;
  SIGNAL and_1136_nl : STD_LOGIC;
  SIGNAL mux_112_nl : STD_LOGIC;
  SIGNAL nor_456_nl : STD_LOGIC;
  SIGNAL nor_454_nl : STD_LOGIC;
  SIGNAL and_1129_nl : STD_LOGIC;
  SIGNAL and_1130_nl : STD_LOGIC;
  SIGNAL and_1131_nl : STD_LOGIC;
  SIGNAL and_1132_nl : STD_LOGIC;
  SIGNAL mux_118_nl : STD_LOGIC;
  SIGNAL nor_455_nl : STD_LOGIC;
  SIGNAL nor_451_nl : STD_LOGIC;
  SIGNAL nor_452_nl : STD_LOGIC;
  SIGNAL and_1125_nl : STD_LOGIC;
  SIGNAL and_1126_nl : STD_LOGIC;
  SIGNAL and_1127_nl : STD_LOGIC;
  SIGNAL and_1128_nl : STD_LOGIC;
  SIGNAL mux_125_nl : STD_LOGIC;
  SIGNAL nor_453_nl : STD_LOGIC;
  SIGNAL nor_447_nl : STD_LOGIC;
  SIGNAL nor_448_nl : STD_LOGIC;
  SIGNAL nor_449_nl : STD_LOGIC;
  SIGNAL and_1121_nl : STD_LOGIC;
  SIGNAL and_1122_nl : STD_LOGIC;
  SIGNAL and_1123_nl : STD_LOGIC;
  SIGNAL and_1124_nl : STD_LOGIC;
  SIGNAL mux_133_nl : STD_LOGIC;
  SIGNAL nor_450_nl : STD_LOGIC;
  SIGNAL nor_442_nl : STD_LOGIC;
  SIGNAL or_352_nl : STD_LOGIC;
  SIGNAL nor_443_nl : STD_LOGIC;
  SIGNAL nor_444_nl : STD_LOGIC;
  SIGNAL nor_445_nl : STD_LOGIC;
  SIGNAL and_1117_nl : STD_LOGIC;
  SIGNAL and_1118_nl : STD_LOGIC;
  SIGNAL and_1119_nl : STD_LOGIC;
  SIGNAL and_1120_nl : STD_LOGIC;
  SIGNAL mux_142_nl : STD_LOGIC;
  SIGNAL nor_446_nl : STD_LOGIC;
  SIGNAL and_1116_nl : STD_LOGIC;
  SIGNAL or_362_nl : STD_LOGIC;
  SIGNAL mux_144_nl : STD_LOGIC;
  SIGNAL and_1172_nl : STD_LOGIC;
  SIGNAL mux_145_nl : STD_LOGIC;
  SIGNAL and_1114_nl : STD_LOGIC;
  SIGNAL mux_146_nl : STD_LOGIC;
  SIGNAL and_1113_nl : STD_LOGIC;
  SIGNAL mux_147_nl : STD_LOGIC;
  SIGNAL and_1112_nl : STD_LOGIC;
  SIGNAL mux_148_nl : STD_LOGIC;
  SIGNAL and_1111_nl : STD_LOGIC;
  SIGNAL mux_149_nl : STD_LOGIC;
  SIGNAL and_1109_nl : STD_LOGIC;
  SIGNAL mux_150_nl : STD_LOGIC;
  SIGNAL and_1110_nl : STD_LOGIC;
  SIGNAL and_1106_nl : STD_LOGIC;
  SIGNAL mux_152_nl : STD_LOGIC;
  SIGNAL and_1107_nl : STD_LOGIC;
  SIGNAL mux_153_nl : STD_LOGIC;
  SIGNAL and_1108_nl : STD_LOGIC;
  SIGNAL and_1102_nl : STD_LOGIC;
  SIGNAL and_1103_nl : STD_LOGIC;
  SIGNAL mux_156_nl : STD_LOGIC;
  SIGNAL and_1104_nl : STD_LOGIC;
  SIGNAL mux_157_nl : STD_LOGIC;
  SIGNAL and_1105_nl : STD_LOGIC;
  SIGNAL and_1097_nl : STD_LOGIC;
  SIGNAL or_437_nl : STD_LOGIC;
  SIGNAL and_1098_nl : STD_LOGIC;
  SIGNAL and_1099_nl : STD_LOGIC;
  SIGNAL mux_161_nl : STD_LOGIC;
  SIGNAL and_1100_nl : STD_LOGIC;
  SIGNAL mux_162_nl : STD_LOGIC;
  SIGNAL and_1101_nl : STD_LOGIC;
  SIGNAL mux_163_nl : STD_LOGIC;
  SIGNAL and_1171_nl : STD_LOGIC;
  SIGNAL and_1094_nl : STD_LOGIC;
  SIGNAL mux_165_nl : STD_LOGIC;
  SIGNAL and_1095_nl : STD_LOGIC;
  SIGNAL and_1091_nl : STD_LOGIC;
  SIGNAL and_1092_nl : STD_LOGIC;
  SIGNAL mux_168_nl : STD_LOGIC;
  SIGNAL and_1093_nl : STD_LOGIC;
  SIGNAL and_1087_nl : STD_LOGIC;
  SIGNAL and_1088_nl : STD_LOGIC;
  SIGNAL and_1089_nl : STD_LOGIC;
  SIGNAL mux_172_nl : STD_LOGIC;
  SIGNAL and_1090_nl : STD_LOGIC;
  SIGNAL and_1082_nl : STD_LOGIC;
  SIGNAL and_1083_nl : STD_LOGIC;
  SIGNAL and_1084_nl : STD_LOGIC;
  SIGNAL and_1085_nl : STD_LOGIC;
  SIGNAL mux_177_nl : STD_LOGIC;
  SIGNAL and_1086_nl : STD_LOGIC;
  SIGNAL and_1076_nl : STD_LOGIC;
  SIGNAL and_1077_nl : STD_LOGIC;
  SIGNAL and_1078_nl : STD_LOGIC;
  SIGNAL and_1079_nl : STD_LOGIC;
  SIGNAL and_1080_nl : STD_LOGIC;
  SIGNAL mux_183_nl : STD_LOGIC;
  SIGNAL and_1081_nl : STD_LOGIC;
  SIGNAL and_1069_nl : STD_LOGIC;
  SIGNAL and_1070_nl : STD_LOGIC;
  SIGNAL and_1071_nl : STD_LOGIC;
  SIGNAL and_1072_nl : STD_LOGIC;
  SIGNAL and_1073_nl : STD_LOGIC;
  SIGNAL and_1074_nl : STD_LOGIC;
  SIGNAL mux_190_nl : STD_LOGIC;
  SIGNAL and_1075_nl : STD_LOGIC;
  SIGNAL and_1061_nl : STD_LOGIC;
  SIGNAL and_1062_nl : STD_LOGIC;
  SIGNAL and_1063_nl : STD_LOGIC;
  SIGNAL and_1064_nl : STD_LOGIC;
  SIGNAL and_1065_nl : STD_LOGIC;
  SIGNAL and_1066_nl : STD_LOGIC;
  SIGNAL and_1067_nl : STD_LOGIC;
  SIGNAL mux_198_nl : STD_LOGIC;
  SIGNAL and_1068_nl : STD_LOGIC;
  SIGNAL and_1052_nl : STD_LOGIC;
  SIGNAL or_540_nl : STD_LOGIC;
  SIGNAL and_1053_nl : STD_LOGIC;
  SIGNAL and_1054_nl : STD_LOGIC;
  SIGNAL and_1055_nl : STD_LOGIC;
  SIGNAL and_1056_nl : STD_LOGIC;
  SIGNAL and_1057_nl : STD_LOGIC;
  SIGNAL and_1058_nl : STD_LOGIC;
  SIGNAL and_1059_nl : STD_LOGIC;
  SIGNAL mux_207_nl : STD_LOGIC;
  SIGNAL and_1060_nl : STD_LOGIC;
  SIGNAL nor_439_nl : STD_LOGIC;
  SIGNAL or_550_nl : STD_LOGIC;
  SIGNAL mux_209_nl : STD_LOGIC;
  SIGNAL and_1170_nl : STD_LOGIC;
  SIGNAL mux_210_nl : STD_LOGIC;
  SIGNAL and_1050_nl : STD_LOGIC;
  SIGNAL mux_211_nl : STD_LOGIC;
  SIGNAL and_1049_nl : STD_LOGIC;
  SIGNAL mux_212_nl : STD_LOGIC;
  SIGNAL and_1048_nl : STD_LOGIC;
  SIGNAL mux_213_nl : STD_LOGIC;
  SIGNAL and_1047_nl : STD_LOGIC;
  SIGNAL mux_214_nl : STD_LOGIC;
  SIGNAL and_1045_nl : STD_LOGIC;
  SIGNAL mux_215_nl : STD_LOGIC;
  SIGNAL and_1046_nl : STD_LOGIC;
  SIGNAL and_1042_nl : STD_LOGIC;
  SIGNAL mux_217_nl : STD_LOGIC;
  SIGNAL and_1043_nl : STD_LOGIC;
  SIGNAL mux_218_nl : STD_LOGIC;
  SIGNAL and_1044_nl : STD_LOGIC;
  SIGNAL and_1038_nl : STD_LOGIC;
  SIGNAL and_1039_nl : STD_LOGIC;
  SIGNAL mux_221_nl : STD_LOGIC;
  SIGNAL and_1040_nl : STD_LOGIC;
  SIGNAL mux_222_nl : STD_LOGIC;
  SIGNAL and_1041_nl : STD_LOGIC;
  SIGNAL and_1033_nl : STD_LOGIC;
  SIGNAL or_624_nl : STD_LOGIC;
  SIGNAL and_1034_nl : STD_LOGIC;
  SIGNAL and_1035_nl : STD_LOGIC;
  SIGNAL mux_226_nl : STD_LOGIC;
  SIGNAL and_1036_nl : STD_LOGIC;
  SIGNAL mux_227_nl : STD_LOGIC;
  SIGNAL and_1037_nl : STD_LOGIC;
  SIGNAL mux_228_nl : STD_LOGIC;
  SIGNAL and_1169_nl : STD_LOGIC;
  SIGNAL and_1030_nl : STD_LOGIC;
  SIGNAL mux_230_nl : STD_LOGIC;
  SIGNAL and_1031_nl : STD_LOGIC;
  SIGNAL and_1027_nl : STD_LOGIC;
  SIGNAL and_1028_nl : STD_LOGIC;
  SIGNAL mux_233_nl : STD_LOGIC;
  SIGNAL and_1029_nl : STD_LOGIC;
  SIGNAL and_1023_nl : STD_LOGIC;
  SIGNAL and_1024_nl : STD_LOGIC;
  SIGNAL and_1025_nl : STD_LOGIC;
  SIGNAL mux_237_nl : STD_LOGIC;
  SIGNAL and_1026_nl : STD_LOGIC;
  SIGNAL and_1018_nl : STD_LOGIC;
  SIGNAL and_1019_nl : STD_LOGIC;
  SIGNAL and_1020_nl : STD_LOGIC;
  SIGNAL and_1021_nl : STD_LOGIC;
  SIGNAL mux_242_nl : STD_LOGIC;
  SIGNAL and_1022_nl : STD_LOGIC;
  SIGNAL and_1012_nl : STD_LOGIC;
  SIGNAL and_1013_nl : STD_LOGIC;
  SIGNAL and_1014_nl : STD_LOGIC;
  SIGNAL and_1015_nl : STD_LOGIC;
  SIGNAL and_1016_nl : STD_LOGIC;
  SIGNAL mux_248_nl : STD_LOGIC;
  SIGNAL and_1017_nl : STD_LOGIC;
  SIGNAL and_1005_nl : STD_LOGIC;
  SIGNAL and_1006_nl : STD_LOGIC;
  SIGNAL and_1007_nl : STD_LOGIC;
  SIGNAL and_1008_nl : STD_LOGIC;
  SIGNAL and_1009_nl : STD_LOGIC;
  SIGNAL and_1010_nl : STD_LOGIC;
  SIGNAL mux_255_nl : STD_LOGIC;
  SIGNAL and_1011_nl : STD_LOGIC;
  SIGNAL and_997_nl : STD_LOGIC;
  SIGNAL and_998_nl : STD_LOGIC;
  SIGNAL and_999_nl : STD_LOGIC;
  SIGNAL and_1000_nl : STD_LOGIC;
  SIGNAL and_1001_nl : STD_LOGIC;
  SIGNAL and_1002_nl : STD_LOGIC;
  SIGNAL and_1003_nl : STD_LOGIC;
  SIGNAL mux_263_nl : STD_LOGIC;
  SIGNAL and_1004_nl : STD_LOGIC;
  SIGNAL and_988_nl : STD_LOGIC;
  SIGNAL or_725_nl : STD_LOGIC;
  SIGNAL and_989_nl : STD_LOGIC;
  SIGNAL and_990_nl : STD_LOGIC;
  SIGNAL and_991_nl : STD_LOGIC;
  SIGNAL and_992_nl : STD_LOGIC;
  SIGNAL and_993_nl : STD_LOGIC;
  SIGNAL and_994_nl : STD_LOGIC;
  SIGNAL and_995_nl : STD_LOGIC;
  SIGNAL mux_272_nl : STD_LOGIC;
  SIGNAL and_996_nl : STD_LOGIC;
  SIGNAL and_987_nl : STD_LOGIC;
  SIGNAL or_735_nl : STD_LOGIC;
  SIGNAL mux_274_nl : STD_LOGIC;
  SIGNAL nor_436_nl : STD_LOGIC;
  SIGNAL mux_275_nl : STD_LOGIC;
  SIGNAL nor_435_nl : STD_LOGIC;
  SIGNAL mux_276_nl : STD_LOGIC;
  SIGNAL nor_434_nl : STD_LOGIC;
  SIGNAL mux_277_nl : STD_LOGIC;
  SIGNAL nor_433_nl : STD_LOGIC;
  SIGNAL mux_278_nl : STD_LOGIC;
  SIGNAL nor_432_nl : STD_LOGIC;
  SIGNAL mux_279_nl : STD_LOGIC;
  SIGNAL nor_430_nl : STD_LOGIC;
  SIGNAL mux_280_nl : STD_LOGIC;
  SIGNAL nor_431_nl : STD_LOGIC;
  SIGNAL nor_427_nl : STD_LOGIC;
  SIGNAL mux_282_nl : STD_LOGIC;
  SIGNAL nor_428_nl : STD_LOGIC;
  SIGNAL mux_283_nl : STD_LOGIC;
  SIGNAL nor_429_nl : STD_LOGIC;
  SIGNAL nor_423_nl : STD_LOGIC;
  SIGNAL nor_424_nl : STD_LOGIC;
  SIGNAL mux_286_nl : STD_LOGIC;
  SIGNAL nor_425_nl : STD_LOGIC;
  SIGNAL mux_287_nl : STD_LOGIC;
  SIGNAL nor_426_nl : STD_LOGIC;
  SIGNAL nor_418_nl : STD_LOGIC;
  SIGNAL or_808_nl : STD_LOGIC;
  SIGNAL nor_419_nl : STD_LOGIC;
  SIGNAL nor_420_nl : STD_LOGIC;
  SIGNAL mux_291_nl : STD_LOGIC;
  SIGNAL nor_421_nl : STD_LOGIC;
  SIGNAL mux_292_nl : STD_LOGIC;
  SIGNAL nor_422_nl : STD_LOGIC;
  SIGNAL nor_409_nl : STD_LOGIC;
  SIGNAL or_823_nl : STD_LOGIC;
  SIGNAL nor_410_nl : STD_LOGIC;
  SIGNAL or_822_nl : STD_LOGIC;
  SIGNAL nor_411_nl : STD_LOGIC;
  SIGNAL or_821_nl : STD_LOGIC;
  SIGNAL nor_412_nl : STD_LOGIC;
  SIGNAL or_820_nl : STD_LOGIC;
  SIGNAL nor_413_nl : STD_LOGIC;
  SIGNAL or_819_nl : STD_LOGIC;
  SIGNAL nor_414_nl : STD_LOGIC;
  SIGNAL or_818_nl : STD_LOGIC;
  SIGNAL nor_415_nl : STD_LOGIC;
  SIGNAL or_817_nl : STD_LOGIC;
  SIGNAL nor_416_nl : STD_LOGIC;
  SIGNAL or_816_nl : STD_LOGIC;
  SIGNAL mux_301_nl : STD_LOGIC;
  SIGNAL nor_417_nl : STD_LOGIC;
  SIGNAL or_815_nl : STD_LOGIC;
  SIGNAL mux_302_nl : STD_LOGIC;
  SIGNAL nor_408_nl : STD_LOGIC;
  SIGNAL and_986_nl : STD_LOGIC;
  SIGNAL mux_304_nl : STD_LOGIC;
  SIGNAL nor_407_nl : STD_LOGIC;
  SIGNAL and_984_nl : STD_LOGIC;
  SIGNAL and_985_nl : STD_LOGIC;
  SIGNAL mux_307_nl : STD_LOGIC;
  SIGNAL nor_406_nl : STD_LOGIC;
  SIGNAL and_981_nl : STD_LOGIC;
  SIGNAL and_982_nl : STD_LOGIC;
  SIGNAL and_983_nl : STD_LOGIC;
  SIGNAL mux_311_nl : STD_LOGIC;
  SIGNAL nor_405_nl : STD_LOGIC;
  SIGNAL and_977_nl : STD_LOGIC;
  SIGNAL and_978_nl : STD_LOGIC;
  SIGNAL and_979_nl : STD_LOGIC;
  SIGNAL and_980_nl : STD_LOGIC;
  SIGNAL mux_316_nl : STD_LOGIC;
  SIGNAL nor_404_nl : STD_LOGIC;
  SIGNAL nor_402_nl : STD_LOGIC;
  SIGNAL and_973_nl : STD_LOGIC;
  SIGNAL and_974_nl : STD_LOGIC;
  SIGNAL and_975_nl : STD_LOGIC;
  SIGNAL and_976_nl : STD_LOGIC;
  SIGNAL mux_322_nl : STD_LOGIC;
  SIGNAL nor_403_nl : STD_LOGIC;
  SIGNAL nor_399_nl : STD_LOGIC;
  SIGNAL nor_400_nl : STD_LOGIC;
  SIGNAL and_969_nl : STD_LOGIC;
  SIGNAL and_970_nl : STD_LOGIC;
  SIGNAL and_971_nl : STD_LOGIC;
  SIGNAL and_972_nl : STD_LOGIC;
  SIGNAL mux_329_nl : STD_LOGIC;
  SIGNAL nor_401_nl : STD_LOGIC;
  SIGNAL nor_395_nl : STD_LOGIC;
  SIGNAL nor_396_nl : STD_LOGIC;
  SIGNAL nor_397_nl : STD_LOGIC;
  SIGNAL and_965_nl : STD_LOGIC;
  SIGNAL and_966_nl : STD_LOGIC;
  SIGNAL and_967_nl : STD_LOGIC;
  SIGNAL and_968_nl : STD_LOGIC;
  SIGNAL mux_337_nl : STD_LOGIC;
  SIGNAL nor_398_nl : STD_LOGIC;
  SIGNAL nor_390_nl : STD_LOGIC;
  SIGNAL or_919_nl : STD_LOGIC;
  SIGNAL nor_391_nl : STD_LOGIC;
  SIGNAL nor_392_nl : STD_LOGIC;
  SIGNAL nor_393_nl : STD_LOGIC;
  SIGNAL and_961_nl : STD_LOGIC;
  SIGNAL and_962_nl : STD_LOGIC;
  SIGNAL and_963_nl : STD_LOGIC;
  SIGNAL and_964_nl : STD_LOGIC;
  SIGNAL mux_346_nl : STD_LOGIC;
  SIGNAL nor_394_nl : STD_LOGIC;
  SIGNAL nor_380_nl : STD_LOGIC;
  SIGNAL or_938_nl : STD_LOGIC;
  SIGNAL nor_381_nl : STD_LOGIC;
  SIGNAL or_937_nl : STD_LOGIC;
  SIGNAL nor_382_nl : STD_LOGIC;
  SIGNAL or_936_nl : STD_LOGIC;
  SIGNAL nor_383_nl : STD_LOGIC;
  SIGNAL or_935_nl : STD_LOGIC;
  SIGNAL nor_384_nl : STD_LOGIC;
  SIGNAL or_934_nl : STD_LOGIC;
  SIGNAL nor_385_nl : STD_LOGIC;
  SIGNAL or_933_nl : STD_LOGIC;
  SIGNAL nor_386_nl : STD_LOGIC;
  SIGNAL or_932_nl : STD_LOGIC;
  SIGNAL nor_387_nl : STD_LOGIC;
  SIGNAL or_931_nl : STD_LOGIC;
  SIGNAL nor_388_nl : STD_LOGIC;
  SIGNAL or_930_nl : STD_LOGIC;
  SIGNAL nor_389_nl : STD_LOGIC;
  SIGNAL or_929_nl : STD_LOGIC;
  SIGNAL mux_357_nl : STD_LOGIC;
  SIGNAL nor_379_nl : STD_LOGIC;
  SIGNAL mux_358_nl : STD_LOGIC;
  SIGNAL nor_378_nl : STD_LOGIC;
  SIGNAL mux_359_nl : STD_LOGIC;
  SIGNAL nor_377_nl : STD_LOGIC;
  SIGNAL mux_360_nl : STD_LOGIC;
  SIGNAL nor_376_nl : STD_LOGIC;
  SIGNAL mux_361_nl : STD_LOGIC;
  SIGNAL nor_375_nl : STD_LOGIC;
  SIGNAL mux_362_nl : STD_LOGIC;
  SIGNAL nor_373_nl : STD_LOGIC;
  SIGNAL mux_363_nl : STD_LOGIC;
  SIGNAL nor_374_nl : STD_LOGIC;
  SIGNAL nor_370_nl : STD_LOGIC;
  SIGNAL mux_365_nl : STD_LOGIC;
  SIGNAL nor_371_nl : STD_LOGIC;
  SIGNAL mux_366_nl : STD_LOGIC;
  SIGNAL nor_372_nl : STD_LOGIC;
  SIGNAL nor_366_nl : STD_LOGIC;
  SIGNAL nor_367_nl : STD_LOGIC;
  SIGNAL mux_369_nl : STD_LOGIC;
  SIGNAL nor_368_nl : STD_LOGIC;
  SIGNAL mux_370_nl : STD_LOGIC;
  SIGNAL nor_369_nl : STD_LOGIC;
  SIGNAL nor_361_nl : STD_LOGIC;
  SIGNAL or_1012_nl : STD_LOGIC;
  SIGNAL nor_362_nl : STD_LOGIC;
  SIGNAL nor_363_nl : STD_LOGIC;
  SIGNAL mux_374_nl : STD_LOGIC;
  SIGNAL nor_364_nl : STD_LOGIC;
  SIGNAL mux_375_nl : STD_LOGIC;
  SIGNAL nor_365_nl : STD_LOGIC;
  SIGNAL nor_352_nl : STD_LOGIC;
  SIGNAL or_1027_nl : STD_LOGIC;
  SIGNAL nor_353_nl : STD_LOGIC;
  SIGNAL or_1026_nl : STD_LOGIC;
  SIGNAL nor_354_nl : STD_LOGIC;
  SIGNAL or_1025_nl : STD_LOGIC;
  SIGNAL nor_355_nl : STD_LOGIC;
  SIGNAL or_1024_nl : STD_LOGIC;
  SIGNAL nor_356_nl : STD_LOGIC;
  SIGNAL or_1023_nl : STD_LOGIC;
  SIGNAL nor_357_nl : STD_LOGIC;
  SIGNAL or_1022_nl : STD_LOGIC;
  SIGNAL nor_358_nl : STD_LOGIC;
  SIGNAL or_1021_nl : STD_LOGIC;
  SIGNAL nor_359_nl : STD_LOGIC;
  SIGNAL or_1020_nl : STD_LOGIC;
  SIGNAL mux_384_nl : STD_LOGIC;
  SIGNAL nor_360_nl : STD_LOGIC;
  SIGNAL or_1019_nl : STD_LOGIC;
  SIGNAL mux_385_nl : STD_LOGIC;
  SIGNAL nor_351_nl : STD_LOGIC;
  SIGNAL and_960_nl : STD_LOGIC;
  SIGNAL mux_387_nl : STD_LOGIC;
  SIGNAL nor_350_nl : STD_LOGIC;
  SIGNAL and_958_nl : STD_LOGIC;
  SIGNAL and_959_nl : STD_LOGIC;
  SIGNAL mux_390_nl : STD_LOGIC;
  SIGNAL nor_349_nl : STD_LOGIC;
  SIGNAL and_955_nl : STD_LOGIC;
  SIGNAL and_956_nl : STD_LOGIC;
  SIGNAL and_957_nl : STD_LOGIC;
  SIGNAL mux_394_nl : STD_LOGIC;
  SIGNAL nor_348_nl : STD_LOGIC;
  SIGNAL and_951_nl : STD_LOGIC;
  SIGNAL and_952_nl : STD_LOGIC;
  SIGNAL and_953_nl : STD_LOGIC;
  SIGNAL and_954_nl : STD_LOGIC;
  SIGNAL mux_399_nl : STD_LOGIC;
  SIGNAL nor_347_nl : STD_LOGIC;
  SIGNAL nor_345_nl : STD_LOGIC;
  SIGNAL and_947_nl : STD_LOGIC;
  SIGNAL and_948_nl : STD_LOGIC;
  SIGNAL and_949_nl : STD_LOGIC;
  SIGNAL and_950_nl : STD_LOGIC;
  SIGNAL mux_405_nl : STD_LOGIC;
  SIGNAL nor_346_nl : STD_LOGIC;
  SIGNAL nor_342_nl : STD_LOGIC;
  SIGNAL nor_343_nl : STD_LOGIC;
  SIGNAL and_943_nl : STD_LOGIC;
  SIGNAL and_944_nl : STD_LOGIC;
  SIGNAL and_945_nl : STD_LOGIC;
  SIGNAL and_946_nl : STD_LOGIC;
  SIGNAL mux_412_nl : STD_LOGIC;
  SIGNAL nor_344_nl : STD_LOGIC;
  SIGNAL nor_338_nl : STD_LOGIC;
  SIGNAL nor_339_nl : STD_LOGIC;
  SIGNAL nor_340_nl : STD_LOGIC;
  SIGNAL and_939_nl : STD_LOGIC;
  SIGNAL and_940_nl : STD_LOGIC;
  SIGNAL and_941_nl : STD_LOGIC;
  SIGNAL and_942_nl : STD_LOGIC;
  SIGNAL mux_420_nl : STD_LOGIC;
  SIGNAL nor_341_nl : STD_LOGIC;
  SIGNAL nor_333_nl : STD_LOGIC;
  SIGNAL nand_12_nl : STD_LOGIC;
  SIGNAL nor_334_nl : STD_LOGIC;
  SIGNAL nor_335_nl : STD_LOGIC;
  SIGNAL nor_336_nl : STD_LOGIC;
  SIGNAL and_935_nl : STD_LOGIC;
  SIGNAL and_936_nl : STD_LOGIC;
  SIGNAL and_937_nl : STD_LOGIC;
  SIGNAL and_938_nl : STD_LOGIC;
  SIGNAL mux_429_nl : STD_LOGIC;
  SIGNAL nor_337_nl : STD_LOGIC;
  SIGNAL nor_324_nl : STD_LOGIC;
  SIGNAL nand_1_nl : STD_LOGIC;
  SIGNAL nor_325_nl : STD_LOGIC;
  SIGNAL nand_2_nl : STD_LOGIC;
  SIGNAL nor_326_nl : STD_LOGIC;
  SIGNAL nand_3_nl : STD_LOGIC;
  SIGNAL nor_327_nl : STD_LOGIC;
  SIGNAL nand_4_nl : STD_LOGIC;
  SIGNAL nor_328_nl : STD_LOGIC;
  SIGNAL nand_5_nl : STD_LOGIC;
  SIGNAL nor_329_nl : STD_LOGIC;
  SIGNAL nand_6_nl : STD_LOGIC;
  SIGNAL nor_330_nl : STD_LOGIC;
  SIGNAL nand_7_nl : STD_LOGIC;
  SIGNAL nor_331_nl : STD_LOGIC;
  SIGNAL nand_8_nl : STD_LOGIC;
  SIGNAL nor_332_nl : STD_LOGIC;
  SIGNAL nand_9_nl : STD_LOGIC;
  SIGNAL and_934_nl : STD_LOGIC;
  SIGNAL nand_11_nl : STD_LOGIC;
  SIGNAL base_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL m_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL return_rsci_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL return_rsci_z : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL ccs_ccore_start_rsci_dat : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL ccs_ccore_start_rsci_idat_1 : STD_LOGIC_VECTOR (0 DOWNTO 0);

  SIGNAL rem_13_cmp_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_1_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_1_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_1_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_2_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_2_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_2_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_3_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_3_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_3_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_4_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_4_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_4_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_5_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_5_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_5_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_6_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_6_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_6_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_7_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_7_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_7_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_8_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_8_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_8_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_9_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_9_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_9_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_10_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_10_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_10_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_11_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_11_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_11_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_v_64_11_2(input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(10 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_13_2(input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(12 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_64_2_2(input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  base_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 1,
      width => 64
      )
    PORT MAP(
      dat => base_rsci_dat,
      idat => base_rsci_idat_1
    );
  base_rsci_dat <= base_rsc_dat;
  base_rsci_idat <= base_rsci_idat_1;

  m_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 2,
      width => 64
      )
    PORT MAP(
      dat => m_rsci_dat,
      idat => m_rsci_idat_1
    );
  m_rsci_dat <= m_rsc_dat;
  m_rsci_idat <= m_rsci_idat_1;

  return_rsci : work.mgc_out_dreg_pkg_v2.mgc_out_dreg_v2
    GENERIC MAP(
      rscid => 3,
      width => 64
      )
    PORT MAP(
      d => return_rsci_d_1,
      z => return_rsci_z
    );
  return_rsci_d_1 <= return_rsci_d;
  return_rsc_z <= return_rsci_z;

  ccs_ccore_start_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 7,
      width => 1
      )
    PORT MAP(
      dat => ccs_ccore_start_rsci_dat,
      idat => ccs_ccore_start_rsci_idat_1
    );
  ccs_ccore_start_rsci_dat(0) <= ccs_ccore_start_rsc_dat;
  ccs_ccore_start_rsci_idat <= ccs_ccore_start_rsci_idat_1(0);

  rem_13_cmp : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_a,
      b => rem_13_cmp_b,
      z => rem_13_cmp_z_1
    );
  rem_13_cmp_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_a_63_0),65));
  rem_13_cmp_b <= '0' & rem_13_cmp_b_63_0;
  rem_13_cmp_z <= rem_13_cmp_z_1;

  rem_13_cmp_1 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_1_a,
      b => rem_13_cmp_1_b,
      z => rem_13_cmp_1_z_1
    );
  rem_13_cmp_1_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_1_a_63_0),65));
  rem_13_cmp_1_b <= '0' & rem_13_cmp_1_b_63_0;
  rem_13_cmp_1_z <= rem_13_cmp_1_z_1;

  rem_13_cmp_2 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_2_a,
      b => rem_13_cmp_2_b,
      z => rem_13_cmp_2_z_1
    );
  rem_13_cmp_2_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_2_a_63_0),65));
  rem_13_cmp_2_b <= '0' & rem_13_cmp_2_b_63_0;
  rem_13_cmp_2_z <= rem_13_cmp_2_z_1;

  rem_13_cmp_3 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_3_a,
      b => rem_13_cmp_3_b,
      z => rem_13_cmp_3_z_1
    );
  rem_13_cmp_3_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_3_a_63_0),65));
  rem_13_cmp_3_b <= '0' & rem_13_cmp_3_b_63_0;
  rem_13_cmp_3_z <= rem_13_cmp_3_z_1;

  rem_13_cmp_4 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_4_a,
      b => rem_13_cmp_4_b,
      z => rem_13_cmp_4_z_1
    );
  rem_13_cmp_4_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_4_a_63_0),65));
  rem_13_cmp_4_b <= '0' & rem_13_cmp_4_b_63_0;
  rem_13_cmp_4_z <= rem_13_cmp_4_z_1;

  rem_13_cmp_5 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_5_a,
      b => rem_13_cmp_5_b,
      z => rem_13_cmp_5_z_1
    );
  rem_13_cmp_5_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_5_a_63_0),65));
  rem_13_cmp_5_b <= '0' & rem_13_cmp_5_b_63_0;
  rem_13_cmp_5_z <= rem_13_cmp_5_z_1;

  rem_13_cmp_6 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_6_a,
      b => rem_13_cmp_6_b,
      z => rem_13_cmp_6_z_1
    );
  rem_13_cmp_6_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_6_a_63_0),65));
  rem_13_cmp_6_b <= '0' & rem_13_cmp_6_b_63_0;
  rem_13_cmp_6_z <= rem_13_cmp_6_z_1;

  rem_13_cmp_7 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_7_a,
      b => rem_13_cmp_7_b,
      z => rem_13_cmp_7_z_1
    );
  rem_13_cmp_7_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_7_a_63_0),65));
  rem_13_cmp_7_b <= '0' & rem_13_cmp_7_b_63_0;
  rem_13_cmp_7_z <= rem_13_cmp_7_z_1;

  rem_13_cmp_8 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_8_a,
      b => rem_13_cmp_8_b,
      z => rem_13_cmp_8_z_1
    );
  rem_13_cmp_8_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_8_a_63_0),65));
  rem_13_cmp_8_b <= '0' & rem_13_cmp_8_b_63_0;
  rem_13_cmp_8_z <= rem_13_cmp_8_z_1;

  rem_13_cmp_9 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_9_a,
      b => rem_13_cmp_9_b,
      z => rem_13_cmp_9_z_1
    );
  rem_13_cmp_9_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_9_a_63_0),65));
  rem_13_cmp_9_b <= '0' & rem_13_cmp_9_b_63_0;
  rem_13_cmp_9_z <= rem_13_cmp_9_z_1;

  rem_13_cmp_10 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_10_a,
      b => rem_13_cmp_10_b,
      z => rem_13_cmp_10_z_1
    );
  rem_13_cmp_10_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_10_a_63_0),65));
  rem_13_cmp_10_b <= '0' & rem_13_cmp_10_b_63_0;
  rem_13_cmp_10_z <= rem_13_cmp_10_z_1;

  rem_13_cmp_11 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_11_a,
      b => rem_13_cmp_11_b,
      z => rem_13_cmp_11_z_1
    );
  rem_13_cmp_11_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_11_a_63_0),65));
  rem_13_cmp_11_b <= '0' & rem_13_cmp_11_b_63_0;
  rem_13_cmp_11_z <= rem_13_cmp_11_z_1;

  and_1203_cse <= ccs_ccore_en AND main_stage_0_12 AND asn_itm_11;
  and_1173_cse <= ccs_ccore_en AND (and_dcpl_294 OR and_dcpl_300 OR and_dcpl_306
      OR and_dcpl_312 OR and_dcpl_318 OR and_dcpl_324 OR and_dcpl_330 OR and_dcpl_336
      OR and_dcpl_342 OR and_dcpl_348 OR and_tmp_35);
  and_1175_cse <= ccs_ccore_en AND (and_dcpl_356 OR and_dcpl_360 OR and_dcpl_364
      OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_376 OR and_dcpl_379 OR and_dcpl_382
      OR and_dcpl_385 OR and_dcpl_388 OR mux_tmp_76);
  and_1177_cse <= ccs_ccore_en AND (and_dcpl_394 OR and_dcpl_397 OR and_dcpl_400
      OR and_dcpl_403 OR and_dcpl_406 OR and_dcpl_409 OR and_dcpl_413 OR and_dcpl_417
      OR and_dcpl_421 OR and_dcpl_425 OR and_tmp_80);
  and_1179_cse <= ccs_ccore_en AND (and_dcpl_431 OR and_dcpl_433 OR and_dcpl_435
      OR and_dcpl_437 OR and_dcpl_439 OR and_dcpl_442 OR and_dcpl_445 OR and_dcpl_448
      OR and_dcpl_451 OR and_dcpl_454 OR mux_tmp_141);
  and_1181_cse <= ccs_ccore_en AND (and_dcpl_461 OR and_dcpl_465 OR and_dcpl_469
      OR and_dcpl_473 OR and_dcpl_477 OR and_dcpl_480 OR and_dcpl_483 OR and_dcpl_486
      OR and_dcpl_489 OR and_dcpl_492 OR and_tmp_125);
  and_1183_cse <= ccs_ccore_en AND (and_dcpl_498 OR and_dcpl_500 OR and_dcpl_502
      OR and_dcpl_504 OR and_dcpl_506 OR and_dcpl_508 OR and_dcpl_510 OR and_dcpl_512
      OR and_dcpl_514 OR and_dcpl_516 OR mux_tmp_206);
  and_1185_cse <= ccs_ccore_en AND (and_dcpl_520 OR and_dcpl_523 OR and_dcpl_526
      OR and_dcpl_529 OR and_dcpl_532 OR and_dcpl_534 OR and_dcpl_536 OR and_dcpl_538
      OR and_dcpl_540 OR and_dcpl_542 OR and_tmp_170);
  and_1187_cse <= ccs_ccore_en AND (and_dcpl_546 OR and_dcpl_548 OR and_dcpl_550
      OR and_dcpl_552 OR and_dcpl_554 OR and_dcpl_556 OR and_dcpl_558 OR and_dcpl_560
      OR and_dcpl_562 OR and_dcpl_564 OR mux_tmp_271);
  and_1189_cse <= ccs_ccore_en AND (and_dcpl_569 OR and_dcpl_573 OR and_dcpl_577
      OR and_dcpl_581 OR and_dcpl_585 OR and_dcpl_589 OR and_dcpl_593 OR and_dcpl_597
      OR and_dcpl_601 OR and_dcpl_605 OR and_tmp_206);
  and_1191_cse <= ccs_ccore_en AND (and_dcpl_610 OR and_dcpl_612 OR and_dcpl_614
      OR and_dcpl_616 OR and_dcpl_618 OR and_dcpl_622 OR and_dcpl_625 OR and_dcpl_628
      OR and_dcpl_631 OR and_dcpl_634 OR mux_tmp_354);
  and_1193_cse <= ccs_ccore_en AND (and_dcpl_638 OR and_dcpl_641 OR and_dcpl_644
      OR and_dcpl_647 OR and_dcpl_650 OR and_dcpl_653 OR and_dcpl_657 OR and_dcpl_661
      OR and_dcpl_665 OR and_dcpl_669 OR and_tmp_233);
  and_1195_cse <= ccs_ccore_en AND (and_dcpl_673 OR and_dcpl_675 OR and_dcpl_677
      OR and_dcpl_679 OR and_dcpl_681 OR and_dcpl_684 OR and_dcpl_687 OR and_dcpl_690
      OR and_dcpl_693 OR and_dcpl_696 OR mux_tmp_437);
  and_1205_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_2;
  and_1207_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_6;
  and_1209_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_9;
  and_1211_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_11;
  and_1213_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_2;
  and_1215_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_6;
  and_1217_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_9;
  and_1219_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_11;
  and_1221_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_18 AND (NOT (rem_12cyc_st_10_1_0(0)));
  and_1223_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_18 AND (rem_12cyc_st_10_1_0(0));
  and_1225_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_23 AND (NOT (rem_12cyc_st_10_1_0(0)));
  and_1227_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_23 AND (rem_12cyc_st_10_1_0(0));
  and_1229_cse <= ccs_ccore_en AND and_dcpl_3;
  and_1231_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_29;
  and_1233_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_33;
  and_1235_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_36;
  and_1237_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_38;
  and_1239_cse <= ccs_ccore_en AND and_dcpl_40 AND and_dcpl_29;
  and_1241_cse <= ccs_ccore_en AND and_dcpl_40 AND and_dcpl_33;
  and_1243_cse <= ccs_ccore_en AND and_dcpl_40 AND and_dcpl_36;
  and_1245_cse <= ccs_ccore_en AND and_dcpl_40 AND and_dcpl_38;
  and_1247_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_45 AND (NOT (rem_12cyc_st_9_1_0(0)));
  and_1249_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_45 AND (rem_12cyc_st_9_1_0(0));
  and_1251_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_50 AND (NOT (rem_12cyc_st_9_1_0(0)));
  and_1253_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_50 AND (rem_12cyc_st_9_1_0(0));
  and_1255_cse <= ccs_ccore_en AND and_dcpl_30;
  and_1257_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_56;
  and_1259_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_60;
  and_1261_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_63;
  and_1263_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_65;
  and_1265_cse <= ccs_ccore_en AND and_dcpl_67 AND and_dcpl_56;
  and_1267_cse <= ccs_ccore_en AND and_dcpl_67 AND and_dcpl_60;
  and_1269_cse <= ccs_ccore_en AND and_dcpl_67 AND and_dcpl_63;
  and_1271_cse <= ccs_ccore_en AND and_dcpl_67 AND and_dcpl_65;
  and_1273_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_72 AND (NOT (rem_12cyc_st_8_1_0(0)));
  and_1275_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_72 AND (rem_12cyc_st_8_1_0(0));
  and_1277_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_77 AND (NOT (rem_12cyc_st_8_1_0(0)));
  and_1279_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_77 AND (rem_12cyc_st_8_1_0(0));
  and_1281_cse <= ccs_ccore_en AND and_dcpl_57;
  and_1283_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_83;
  and_1285_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_87;
  and_1287_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_90;
  and_1289_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_92;
  and_1291_cse <= ccs_ccore_en AND and_dcpl_94 AND and_dcpl_83;
  and_1293_cse <= ccs_ccore_en AND and_dcpl_94 AND and_dcpl_87;
  and_1295_cse <= ccs_ccore_en AND and_dcpl_94 AND and_dcpl_90;
  and_1297_cse <= ccs_ccore_en AND and_dcpl_94 AND and_dcpl_92;
  and_1299_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_99 AND (NOT (rem_12cyc_st_7_1_0(0)));
  and_1301_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_99 AND (rem_12cyc_st_7_1_0(0));
  and_1303_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_104 AND (NOT (rem_12cyc_st_7_1_0(0)));
  and_1305_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_104 AND (rem_12cyc_st_7_1_0(0));
  and_1307_cse <= ccs_ccore_en AND and_dcpl_84;
  and_1309_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_110;
  and_1311_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_115;
  and_1313_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_117;
  and_1315_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_119;
  and_1317_cse <= ccs_ccore_en AND and_dcpl_121 AND and_dcpl_110;
  and_1319_cse <= ccs_ccore_en AND and_dcpl_121 AND and_dcpl_115;
  and_1321_cse <= ccs_ccore_en AND and_dcpl_121 AND and_dcpl_117;
  and_1323_cse <= ccs_ccore_en AND and_dcpl_121 AND and_dcpl_119;
  and_1325_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_126 AND (NOT (rem_12cyc_st_6_1_0(1)));
  and_1327_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_129 AND (NOT (rem_12cyc_st_6_1_0(1)));
  and_1329_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_126 AND (rem_12cyc_st_6_1_0(1));
  and_1331_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_129 AND (rem_12cyc_st_6_1_0(1));
  and_1333_cse <= ccs_ccore_en AND and_dcpl_111;
  and_1335_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_137;
  and_1337_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_141;
  and_1339_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_144;
  and_1341_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_146;
  and_1343_cse <= ccs_ccore_en AND and_dcpl_148 AND and_dcpl_137;
  and_1345_cse <= ccs_ccore_en AND and_dcpl_148 AND and_dcpl_141;
  and_1347_cse <= ccs_ccore_en AND and_dcpl_148 AND and_dcpl_144;
  and_1349_cse <= ccs_ccore_en AND and_dcpl_148 AND and_dcpl_146;
  and_1351_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_153 AND (NOT (rem_12cyc_st_5_1_0(0)));
  and_1353_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_153 AND (rem_12cyc_st_5_1_0(0));
  and_1355_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_158 AND (NOT (rem_12cyc_st_5_1_0(0)));
  and_1357_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_158 AND (rem_12cyc_st_5_1_0(0));
  and_1359_cse <= ccs_ccore_en AND and_dcpl_138;
  and_1361_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_164;
  and_1363_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_168;
  and_1365_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_171;
  and_1367_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_173;
  and_1369_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_175 AND (NOT (rem_12cyc_st_4_1_0(0)));
  and_1371_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_175 AND (rem_12cyc_st_4_1_0(0));
  and_1373_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_180 AND (NOT (rem_12cyc_st_4_1_0(0)));
  and_1375_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_180 AND (rem_12cyc_st_4_1_0(0));
  and_1377_cse <= ccs_ccore_en AND and_dcpl_185 AND and_dcpl_164;
  and_1379_cse <= ccs_ccore_en AND and_dcpl_185 AND and_dcpl_168;
  and_1381_cse <= ccs_ccore_en AND and_dcpl_185 AND and_dcpl_171;
  and_1383_cse <= ccs_ccore_en AND and_dcpl_185 AND and_dcpl_173;
  and_1385_cse <= ccs_ccore_en AND and_dcpl_165;
  and_1387_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_191;
  and_1389_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_195;
  and_1391_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_198;
  and_1393_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_200;
  and_1395_cse <= ccs_ccore_en AND and_dcpl_202 AND and_dcpl_191;
  and_1397_cse <= ccs_ccore_en AND and_dcpl_202 AND and_dcpl_195;
  and_1399_cse <= ccs_ccore_en AND and_dcpl_202 AND and_dcpl_198;
  and_1401_cse <= ccs_ccore_en AND and_dcpl_202 AND and_dcpl_200;
  and_1403_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_207 AND (NOT (rem_12cyc_st_3_1_0(0)));
  and_1405_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_207 AND (rem_12cyc_st_3_1_0(0));
  and_1407_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_212 AND (NOT (rem_12cyc_st_3_1_0(0)));
  and_1409_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_212 AND (rem_12cyc_st_3_1_0(0));
  and_1411_cse <= ccs_ccore_en AND and_dcpl_192;
  and_1413_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_218;
  and_1415_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_222;
  and_1417_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_225;
  and_1419_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_227;
  and_1421_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_229 AND (NOT (rem_12cyc_st_2_1_0(0)));
  and_1423_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_229 AND (rem_12cyc_st_2_1_0(0));
  and_1425_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_234 AND (NOT (rem_12cyc_st_2_1_0(0)));
  and_1427_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_234 AND (rem_12cyc_st_2_1_0(0));
  and_1429_cse <= ccs_ccore_en AND and_dcpl_239 AND and_dcpl_218;
  and_1431_cse <= ccs_ccore_en AND and_dcpl_239 AND and_dcpl_222;
  and_1433_cse <= ccs_ccore_en AND and_dcpl_239 AND and_dcpl_225;
  and_1435_cse <= ccs_ccore_en AND and_dcpl_239 AND and_dcpl_227;
  and_1437_cse <= ccs_ccore_en AND and_dcpl_219;
  and_1439_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_245;
  and_1441_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_249;
  and_1443_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_252;
  and_1445_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_254;
  and_1447_cse <= ccs_ccore_en AND and_dcpl_256 AND and_dcpl_245;
  and_1449_cse <= ccs_ccore_en AND and_dcpl_256 AND and_dcpl_249;
  and_1451_cse <= ccs_ccore_en AND and_dcpl_256 AND and_dcpl_252;
  and_1453_cse <= ccs_ccore_en AND and_dcpl_256 AND and_dcpl_254;
  and_1455_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_261 AND (NOT (rem_12cyc_1_0(0)));
  and_1457_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_261 AND (rem_12cyc_1_0(0));
  and_1459_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_266 AND (NOT (rem_12cyc_1_0(0)));
  and_1461_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_266 AND (rem_12cyc_1_0(0));
  and_1463_cse <= ccs_ccore_en AND and_dcpl_246;
  and_1197_cse <= ccs_ccore_en AND ccs_ccore_start_rsci_idat;
  and_273_nl <= and_dcpl_272 AND and_dcpl_271;
  and_275_nl <= and_dcpl_272 AND and_dcpl_274;
  and_277_nl <= and_dcpl_272 AND and_dcpl_276;
  and_279_nl <= and_dcpl_272 AND and_dcpl_278;
  and_281_nl <= and_dcpl_280 AND and_dcpl_271;
  and_282_nl <= and_dcpl_280 AND and_dcpl_274;
  and_283_nl <= and_dcpl_280 AND and_dcpl_276;
  and_284_nl <= and_dcpl_280 AND and_dcpl_278;
  and_286_nl <= and_dcpl_285 AND and_dcpl_271;
  and_287_nl <= and_dcpl_285 AND and_dcpl_274;
  and_288_nl <= and_dcpl_285 AND and_dcpl_276;
  and_289_nl <= and_dcpl_285 AND and_dcpl_278;
  and_290_nl <= CONV_SL_1_1(rem_12cyc_st_12_3_2=STD_LOGIC_VECTOR'("11"));
  result_sva_duc_mx0 <= MUX1HOT_v_64_13_2((rem_13_cmp_1_z(63 DOWNTO 0)), (rem_13_cmp_2_z(63
      DOWNTO 0)), (rem_13_cmp_3_z(63 DOWNTO 0)), (rem_13_cmp_4_z(63 DOWNTO 0)), (rem_13_cmp_5_z(63
      DOWNTO 0)), (rem_13_cmp_6_z(63 DOWNTO 0)), (rem_13_cmp_7_z(63 DOWNTO 0)), (rem_13_cmp_8_z(63
      DOWNTO 0)), (rem_13_cmp_9_z(63 DOWNTO 0)), (rem_13_cmp_10_z(63 DOWNTO 0)),
      (rem_13_cmp_11_z(63 DOWNTO 0)), (rem_13_cmp_z(63 DOWNTO 0)), result_sva_duc,
      STD_LOGIC_VECTOR'( and_273_nl & and_275_nl & and_277_nl & and_279_nl & and_281_nl
      & and_282_nl & and_283_nl & and_284_nl & and_286_nl & and_287_nl & and_288_nl
      & and_289_nl & and_290_nl));
  acc_1_tmp <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(rem_12cyc_3_2 & rem_12cyc_1_0)
      + UNSIGNED'( "0001"), 4));
  xor_nl <= (acc_1_tmp(2)) XOR (acc_1_tmp(3));
  nor_nl <= NOT(CONV_SL_1_1(acc_1_tmp(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10")));
  acc_tmp <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(xor_nl, 1),
      2) + CONV_UNSIGNED(CONV_UNSIGNED(nor_nl, 1), 2), 2));
  and_dcpl_1 <= NOT((rem_12cyc_st_10_3_2(1)) OR (rem_12cyc_st_10_1_0(1)));
  and_dcpl_2 <= and_dcpl_1 AND (NOT (rem_12cyc_st_10_1_0(0)));
  and_dcpl_3 <= main_stage_0_11 AND asn_itm_10;
  and_dcpl_4 <= and_dcpl_3 AND (NOT (rem_12cyc_st_10_3_2(0)));
  and_dcpl_6 <= and_dcpl_1 AND (rem_12cyc_st_10_1_0(0));
  and_dcpl_8 <= (NOT (rem_12cyc_st_10_3_2(1))) AND (rem_12cyc_st_10_1_0(1));
  and_dcpl_9 <= and_dcpl_8 AND (NOT (rem_12cyc_st_10_1_0(0)));
  and_dcpl_11 <= and_dcpl_8 AND (rem_12cyc_st_10_1_0(0));
  and_dcpl_13 <= and_dcpl_3 AND (rem_12cyc_st_10_3_2(0));
  and_dcpl_18 <= (rem_12cyc_st_10_3_2(1)) AND (NOT (rem_12cyc_st_10_1_0(1)));
  and_dcpl_23 <= (rem_12cyc_st_10_3_2(1)) AND (rem_12cyc_st_10_1_0(1));
  and_dcpl_28 <= NOT((rem_12cyc_st_9_3_2(1)) OR (rem_12cyc_st_9_1_0(1)));
  and_dcpl_29 <= and_dcpl_28 AND (NOT (rem_12cyc_st_9_1_0(0)));
  and_dcpl_30 <= main_stage_0_10 AND asn_itm_9;
  and_dcpl_31 <= and_dcpl_30 AND (NOT (rem_12cyc_st_9_3_2(0)));
  and_dcpl_33 <= and_dcpl_28 AND (rem_12cyc_st_9_1_0(0));
  and_dcpl_35 <= (NOT (rem_12cyc_st_9_3_2(1))) AND (rem_12cyc_st_9_1_0(1));
  and_dcpl_36 <= and_dcpl_35 AND (NOT (rem_12cyc_st_9_1_0(0)));
  and_dcpl_38 <= and_dcpl_35 AND (rem_12cyc_st_9_1_0(0));
  and_dcpl_40 <= and_dcpl_30 AND (rem_12cyc_st_9_3_2(0));
  and_dcpl_45 <= (rem_12cyc_st_9_3_2(1)) AND (NOT (rem_12cyc_st_9_1_0(1)));
  and_dcpl_50 <= (rem_12cyc_st_9_3_2(1)) AND (rem_12cyc_st_9_1_0(1));
  and_dcpl_55 <= NOT((rem_12cyc_st_8_3_2(1)) OR (rem_12cyc_st_8_1_0(1)));
  and_dcpl_56 <= and_dcpl_55 AND (NOT (rem_12cyc_st_8_1_0(0)));
  and_dcpl_57 <= main_stage_0_9 AND asn_itm_8;
  and_dcpl_58 <= and_dcpl_57 AND (NOT (rem_12cyc_st_8_3_2(0)));
  and_dcpl_60 <= and_dcpl_55 AND (rem_12cyc_st_8_1_0(0));
  and_dcpl_62 <= (NOT (rem_12cyc_st_8_3_2(1))) AND (rem_12cyc_st_8_1_0(1));
  and_dcpl_63 <= and_dcpl_62 AND (NOT (rem_12cyc_st_8_1_0(0)));
  and_dcpl_65 <= and_dcpl_62 AND (rem_12cyc_st_8_1_0(0));
  and_dcpl_67 <= and_dcpl_57 AND (rem_12cyc_st_8_3_2(0));
  and_dcpl_72 <= (rem_12cyc_st_8_3_2(1)) AND (NOT (rem_12cyc_st_8_1_0(1)));
  and_dcpl_77 <= (rem_12cyc_st_8_3_2(1)) AND (rem_12cyc_st_8_1_0(1));
  and_dcpl_82 <= NOT((rem_12cyc_st_7_3_2(1)) OR (rem_12cyc_st_7_1_0(1)));
  and_dcpl_83 <= and_dcpl_82 AND (NOT (rem_12cyc_st_7_1_0(0)));
  and_dcpl_84 <= main_stage_0_8 AND asn_itm_7;
  and_dcpl_85 <= and_dcpl_84 AND (NOT (rem_12cyc_st_7_3_2(0)));
  and_dcpl_87 <= and_dcpl_82 AND (rem_12cyc_st_7_1_0(0));
  and_dcpl_89 <= (NOT (rem_12cyc_st_7_3_2(1))) AND (rem_12cyc_st_7_1_0(1));
  and_dcpl_90 <= and_dcpl_89 AND (NOT (rem_12cyc_st_7_1_0(0)));
  and_dcpl_92 <= and_dcpl_89 AND (rem_12cyc_st_7_1_0(0));
  and_dcpl_94 <= and_dcpl_84 AND (rem_12cyc_st_7_3_2(0));
  and_dcpl_99 <= (rem_12cyc_st_7_3_2(1)) AND (NOT (rem_12cyc_st_7_1_0(1)));
  and_dcpl_104 <= (rem_12cyc_st_7_3_2(1)) AND (rem_12cyc_st_7_1_0(1));
  and_dcpl_109 <= NOT((rem_12cyc_st_6_3_2(1)) OR (rem_12cyc_st_6_1_0(0)));
  and_dcpl_110 <= and_dcpl_109 AND (NOT (rem_12cyc_st_6_1_0(1)));
  and_dcpl_111 <= main_stage_0_7 AND asn_itm_6;
  and_dcpl_112 <= and_dcpl_111 AND (NOT (rem_12cyc_st_6_3_2(0)));
  and_dcpl_114 <= (NOT (rem_12cyc_st_6_3_2(1))) AND (rem_12cyc_st_6_1_0(0));
  and_dcpl_115 <= and_dcpl_114 AND (NOT (rem_12cyc_st_6_1_0(1)));
  and_dcpl_117 <= and_dcpl_109 AND (rem_12cyc_st_6_1_0(1));
  and_dcpl_119 <= and_dcpl_114 AND (rem_12cyc_st_6_1_0(1));
  and_dcpl_121 <= and_dcpl_111 AND (rem_12cyc_st_6_3_2(0));
  and_dcpl_126 <= (rem_12cyc_st_6_3_2(1)) AND (NOT (rem_12cyc_st_6_1_0(0)));
  and_dcpl_129 <= (rem_12cyc_st_6_3_2(1)) AND (rem_12cyc_st_6_1_0(0));
  and_dcpl_136 <= NOT((rem_12cyc_st_5_3_2(1)) OR (rem_12cyc_st_5_1_0(1)));
  and_dcpl_137 <= and_dcpl_136 AND (NOT (rem_12cyc_st_5_1_0(0)));
  and_dcpl_138 <= main_stage_0_6 AND asn_itm_5;
  and_dcpl_139 <= and_dcpl_138 AND (NOT (rem_12cyc_st_5_3_2(0)));
  and_dcpl_141 <= and_dcpl_136 AND (rem_12cyc_st_5_1_0(0));
  and_dcpl_143 <= (NOT (rem_12cyc_st_5_3_2(1))) AND (rem_12cyc_st_5_1_0(1));
  and_dcpl_144 <= and_dcpl_143 AND (NOT (rem_12cyc_st_5_1_0(0)));
  and_dcpl_146 <= and_dcpl_143 AND (rem_12cyc_st_5_1_0(0));
  and_dcpl_148 <= and_dcpl_138 AND (rem_12cyc_st_5_3_2(0));
  and_dcpl_153 <= (rem_12cyc_st_5_3_2(1)) AND (NOT (rem_12cyc_st_5_1_0(1)));
  and_dcpl_158 <= (rem_12cyc_st_5_3_2(1)) AND (rem_12cyc_st_5_1_0(1));
  and_dcpl_163 <= NOT((rem_12cyc_st_4_3_2(0)) OR (rem_12cyc_st_4_1_0(1)));
  and_dcpl_164 <= and_dcpl_163 AND (NOT (rem_12cyc_st_4_1_0(0)));
  and_dcpl_165 <= main_stage_0_5 AND asn_itm_4;
  and_dcpl_166 <= and_dcpl_165 AND (NOT (rem_12cyc_st_4_3_2(1)));
  and_dcpl_168 <= and_dcpl_163 AND (rem_12cyc_st_4_1_0(0));
  and_dcpl_170 <= (NOT (rem_12cyc_st_4_3_2(0))) AND (rem_12cyc_st_4_1_0(1));
  and_dcpl_171 <= and_dcpl_170 AND (NOT (rem_12cyc_st_4_1_0(0)));
  and_dcpl_173 <= and_dcpl_170 AND (rem_12cyc_st_4_1_0(0));
  and_dcpl_175 <= (rem_12cyc_st_4_3_2(0)) AND (NOT (rem_12cyc_st_4_1_0(1)));
  and_dcpl_180 <= (rem_12cyc_st_4_3_2(0)) AND (rem_12cyc_st_4_1_0(1));
  and_dcpl_185 <= and_dcpl_165 AND (rem_12cyc_st_4_3_2(1));
  and_dcpl_190 <= NOT((rem_12cyc_st_3_3_2(1)) OR (rem_12cyc_st_3_1_0(1)));
  and_dcpl_191 <= and_dcpl_190 AND (NOT (rem_12cyc_st_3_1_0(0)));
  and_dcpl_192 <= main_stage_0_4 AND asn_itm_3;
  and_dcpl_193 <= and_dcpl_192 AND (NOT (rem_12cyc_st_3_3_2(0)));
  and_dcpl_195 <= and_dcpl_190 AND (rem_12cyc_st_3_1_0(0));
  and_dcpl_197 <= (NOT (rem_12cyc_st_3_3_2(1))) AND (rem_12cyc_st_3_1_0(1));
  and_dcpl_198 <= and_dcpl_197 AND (NOT (rem_12cyc_st_3_1_0(0)));
  and_dcpl_200 <= and_dcpl_197 AND (rem_12cyc_st_3_1_0(0));
  and_dcpl_202 <= and_dcpl_192 AND (rem_12cyc_st_3_3_2(0));
  and_dcpl_207 <= (rem_12cyc_st_3_3_2(1)) AND (NOT (rem_12cyc_st_3_1_0(1)));
  and_dcpl_212 <= (rem_12cyc_st_3_3_2(1)) AND (rem_12cyc_st_3_1_0(1));
  and_dcpl_217 <= NOT((rem_12cyc_st_2_3_2(0)) OR (rem_12cyc_st_2_1_0(1)));
  and_dcpl_218 <= and_dcpl_217 AND (NOT (rem_12cyc_st_2_1_0(0)));
  and_dcpl_219 <= main_stage_0_3 AND asn_itm_2;
  and_dcpl_220 <= and_dcpl_219 AND (NOT (rem_12cyc_st_2_3_2(1)));
  and_dcpl_222 <= and_dcpl_217 AND (rem_12cyc_st_2_1_0(0));
  and_dcpl_224 <= (NOT (rem_12cyc_st_2_3_2(0))) AND (rem_12cyc_st_2_1_0(1));
  and_dcpl_225 <= and_dcpl_224 AND (NOT (rem_12cyc_st_2_1_0(0)));
  and_dcpl_227 <= and_dcpl_224 AND (rem_12cyc_st_2_1_0(0));
  and_dcpl_229 <= (rem_12cyc_st_2_3_2(0)) AND (NOT (rem_12cyc_st_2_1_0(1)));
  and_dcpl_234 <= (rem_12cyc_st_2_3_2(0)) AND (rem_12cyc_st_2_1_0(1));
  and_dcpl_239 <= and_dcpl_219 AND (rem_12cyc_st_2_3_2(1));
  and_dcpl_244 <= NOT((rem_12cyc_3_2(1)) OR (rem_12cyc_1_0(1)));
  and_dcpl_245 <= and_dcpl_244 AND (NOT (rem_12cyc_1_0(0)));
  and_dcpl_246 <= main_stage_0_2 AND asn_itm_1;
  and_dcpl_247 <= and_dcpl_246 AND (NOT (rem_12cyc_3_2(0)));
  and_dcpl_249 <= and_dcpl_244 AND (rem_12cyc_1_0(0));
  and_dcpl_251 <= (NOT (rem_12cyc_3_2(1))) AND (rem_12cyc_1_0(1));
  and_dcpl_252 <= and_dcpl_251 AND (NOT (rem_12cyc_1_0(0)));
  and_dcpl_254 <= and_dcpl_251 AND (rem_12cyc_1_0(0));
  and_dcpl_256 <= and_dcpl_246 AND (rem_12cyc_3_2(0));
  and_dcpl_261 <= (rem_12cyc_3_2(1)) AND (NOT (rem_12cyc_1_0(1)));
  and_dcpl_266 <= (rem_12cyc_3_2(1)) AND (rem_12cyc_1_0(1));
  and_dcpl_271 <= NOT(CONV_SL_1_1(rem_12cyc_st_12_1_0/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_272 <= NOT(CONV_SL_1_1(rem_12cyc_st_12_3_2/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_274 <= CONV_SL_1_1(rem_12cyc_st_12_1_0=STD_LOGIC_VECTOR'("01"));
  and_dcpl_276 <= CONV_SL_1_1(rem_12cyc_st_12_1_0=STD_LOGIC_VECTOR'("10"));
  and_dcpl_278 <= CONV_SL_1_1(rem_12cyc_st_12_1_0=STD_LOGIC_VECTOR'("11"));
  and_dcpl_280 <= CONV_SL_1_1(rem_12cyc_st_12_3_2=STD_LOGIC_VECTOR'("01"));
  and_dcpl_285 <= CONV_SL_1_1(rem_12cyc_st_12_3_2=STD_LOGIC_VECTOR'("10"));
  and_dcpl_291 <= NOT(CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_292 <= ccs_ccore_start_rsci_idat AND (NOT (acc_tmp(0)));
  and_dcpl_293 <= and_dcpl_292 AND (NOT (acc_tmp(1)));
  and_dcpl_294 <= and_dcpl_293 AND and_dcpl_291;
  and_dcpl_295 <= NOT(CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_296 <= and_dcpl_295 AND (NOT (rem_12cyc_st_2_1_0(1)));
  and_dcpl_298 <= (NOT (rem_12cyc_st_2_1_0(0))) AND main_stage_0_3 AND asn_itm_2;
  not_tmp_54 <= NOT(asn_itm_1 AND main_stage_0_2);
  or_tmp_2 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_54;
  or_1_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("00"));
  nor_518_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_2));
  mux_14_nl <= MUX_s_1_2_2(nor_518_nl, or_tmp_2, or_1_cse);
  and_dcpl_300 <= mux_14_nl AND and_dcpl_298 AND and_dcpl_296;
  and_dcpl_301 <= NOT(CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_302 <= and_dcpl_301 AND (NOT (rem_12cyc_st_3_1_0(1)));
  and_dcpl_304 <= (NOT (rem_12cyc_st_3_1_0(0))) AND main_stage_0_4 AND asn_itm_3;
  or_6_cse <= (rem_12cyc_st_2_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp <= or_6_cse AND or_tmp_2;
  nor_517_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp));
  mux_15_nl <= MUX_s_1_2_2(nor_517_nl, and_tmp, or_1_cse);
  and_dcpl_306 <= mux_15_nl AND and_dcpl_304 AND and_dcpl_302;
  and_dcpl_307 <= NOT(CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_308 <= and_dcpl_307 AND (NOT (rem_12cyc_st_4_1_0(1)));
  and_dcpl_310 <= (NOT (rem_12cyc_st_4_1_0(0))) AND main_stage_0_5 AND asn_itm_4;
  or_10_cse <= (rem_12cyc_st_3_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_2 <= or_6_cse AND or_10_cse AND or_tmp_2;
  nor_516_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_2));
  mux_16_nl <= MUX_s_1_2_2(nor_516_nl, and_tmp_2, or_1_cse);
  and_dcpl_312 <= mux_16_nl AND and_dcpl_310 AND and_dcpl_308;
  and_dcpl_313 <= NOT(CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_314 <= and_dcpl_313 AND (NOT (rem_12cyc_st_5_1_0(1)));
  and_dcpl_316 <= (NOT (rem_12cyc_st_5_1_0(0))) AND main_stage_0_6 AND asn_itm_5;
  or_15_cse <= (rem_12cyc_st_4_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_5 <= or_6_cse AND or_10_cse AND or_15_cse AND or_tmp_2;
  nor_515_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_5));
  mux_17_nl <= MUX_s_1_2_2(nor_515_nl, and_tmp_5, or_1_cse);
  and_dcpl_318 <= mux_17_nl AND and_dcpl_316 AND and_dcpl_314;
  or_21_cse <= (rem_12cyc_st_5_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_9 <= or_6_cse AND or_10_cse AND or_15_cse AND or_21_cse AND or_tmp_2;
  nor_514_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_9));
  mux_18_nl <= MUX_s_1_2_2(nor_514_nl, and_tmp_9, or_1_cse);
  and_dcpl_324 <= mux_18_nl AND and_dcpl_112 AND and_dcpl_110;
  or_28_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_512_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_2));
  mux_19_nl <= MUX_s_1_2_2(nor_512_nl, or_tmp_2, or_28_cse);
  and_tmp_13 <= or_6_cse AND or_10_cse AND or_15_cse AND or_21_cse AND mux_19_nl;
  nor_513_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_13));
  mux_20_nl <= MUX_s_1_2_2(nor_513_nl, and_tmp_13, or_1_cse);
  and_dcpl_330 <= mux_20_nl AND and_dcpl_85 AND and_dcpl_83;
  or_37_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_509_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_2));
  mux_tmp_19 <= MUX_s_1_2_2(nor_509_nl, or_tmp_2, or_37_cse);
  nor_510_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_19));
  mux_22_nl <= MUX_s_1_2_2(nor_510_nl, mux_tmp_19, or_28_cse);
  and_tmp_17 <= or_6_cse AND or_10_cse AND or_15_cse AND or_21_cse AND mux_22_nl;
  nor_511_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_17));
  mux_23_nl <= MUX_s_1_2_2(nor_511_nl, and_tmp_17, or_1_cse);
  and_dcpl_336 <= mux_23_nl AND and_dcpl_58 AND and_dcpl_56;
  or_48_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_505_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_2));
  mux_tmp_22 <= MUX_s_1_2_2(nor_505_nl, or_tmp_2, or_48_cse);
  nor_506_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_22));
  mux_tmp_23 <= MUX_s_1_2_2(nor_506_nl, mux_tmp_22, or_37_cse);
  nor_507_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_23));
  mux_26_nl <= MUX_s_1_2_2(nor_507_nl, mux_tmp_23, or_28_cse);
  and_tmp_21 <= or_6_cse AND or_10_cse AND or_15_cse AND or_21_cse AND mux_26_nl;
  nor_508_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_21));
  mux_27_nl <= MUX_s_1_2_2(nor_508_nl, and_tmp_21, or_1_cse);
  and_dcpl_342 <= mux_27_nl AND and_dcpl_31 AND and_dcpl_29;
  nor_500_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_2));
  or_61_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_26 <= MUX_s_1_2_2(nor_500_nl, or_tmp_2, or_61_nl);
  nor_501_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_26));
  mux_tmp_27 <= MUX_s_1_2_2(nor_501_nl, mux_tmp_26, or_48_cse);
  nor_502_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_27));
  mux_tmp_28 <= MUX_s_1_2_2(nor_502_nl, mux_tmp_27, or_37_cse);
  nor_503_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_28));
  mux_31_nl <= MUX_s_1_2_2(nor_503_nl, mux_tmp_28, or_28_cse);
  and_tmp_25 <= or_6_cse AND or_10_cse AND or_15_cse AND or_21_cse AND mux_31_nl;
  nor_504_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_25));
  mux_32_nl <= MUX_s_1_2_2(nor_504_nl, and_tmp_25, or_1_cse);
  and_dcpl_348 <= mux_32_nl AND and_dcpl_4 AND and_dcpl_2;
  and_tmp_35 <= ((NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_8)
      OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_9)
      OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_10)
      OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"))) AND or_6_cse AND
      or_10_cse AND or_15_cse AND or_21_cse AND ((NOT main_stage_0_7) OR (NOT asn_itm_6)
      OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00")))
      AND ((NOT main_stage_0_11) OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("00"))) AND (CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT ccs_ccore_start_rsci_idat));
  and_dcpl_355 <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_356 <= and_dcpl_293 AND and_dcpl_355;
  and_dcpl_358 <= (rem_12cyc_st_2_1_0(0)) AND main_stage_0_3 AND asn_itm_2;
  or_tmp_80 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_54;
  or_83_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("00"));
  nor_499_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_80));
  mux_33_nl <= MUX_s_1_2_2(nor_499_nl, or_tmp_80, or_83_cse);
  and_dcpl_360 <= mux_33_nl AND and_dcpl_358 AND and_dcpl_296;
  and_dcpl_362 <= (rem_12cyc_st_3_1_0(0)) AND main_stage_0_4 AND asn_itm_3;
  nand_276_cse <= NOT(asn_itm_2 AND main_stage_0_3 AND (rem_12cyc_st_2_1_0(0)));
  or_88_cse <= (rem_12cyc_st_2_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1168_nl <= nand_276_cse AND or_tmp_80;
  mux_tmp_32 <= MUX_s_1_2_2(and_1168_nl, or_tmp_80, or_88_cse);
  nor_498_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_32));
  mux_35_nl <= MUX_s_1_2_2(nor_498_nl, mux_tmp_32, or_83_cse);
  and_dcpl_364 <= mux_35_nl AND and_dcpl_362 AND and_dcpl_302;
  and_dcpl_366 <= (rem_12cyc_st_4_1_0(0)) AND main_stage_0_5 AND asn_itm_4;
  nand_274_cse <= NOT(asn_itm_3 AND main_stage_0_4 AND (rem_12cyc_st_3_1_0(0)));
  or_93_cse <= (rem_12cyc_st_3_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1166_nl <= nand_274_cse AND or_tmp_80;
  mux_tmp_34 <= MUX_s_1_2_2(and_1166_nl, or_tmp_80, or_93_cse);
  and_1167_nl <= nand_276_cse AND mux_tmp_34;
  mux_tmp_35 <= MUX_s_1_2_2(and_1167_nl, mux_tmp_34, or_88_cse);
  nor_497_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_35));
  mux_38_nl <= MUX_s_1_2_2(nor_497_nl, mux_tmp_35, or_83_cse);
  and_dcpl_368 <= mux_38_nl AND and_dcpl_366 AND and_dcpl_308;
  and_dcpl_370 <= (rem_12cyc_st_5_1_0(0)) AND main_stage_0_6 AND asn_itm_5;
  nand_271_cse <= NOT(asn_itm_4 AND main_stage_0_5 AND (rem_12cyc_st_4_1_0(0)));
  or_100_cse <= (rem_12cyc_st_4_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1163_nl <= nand_271_cse AND or_tmp_80;
  mux_tmp_37 <= MUX_s_1_2_2(and_1163_nl, or_tmp_80, or_100_cse);
  and_1164_nl <= nand_274_cse AND mux_tmp_37;
  mux_tmp_38 <= MUX_s_1_2_2(and_1164_nl, mux_tmp_37, or_93_cse);
  and_1165_nl <= nand_276_cse AND mux_tmp_38;
  mux_tmp_39 <= MUX_s_1_2_2(and_1165_nl, mux_tmp_38, or_88_cse);
  nor_496_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_39));
  mux_42_nl <= MUX_s_1_2_2(nor_496_nl, mux_tmp_39, or_83_cse);
  and_dcpl_372 <= mux_42_nl AND and_dcpl_370 AND and_dcpl_314;
  nand_267_cse <= NOT(asn_itm_5 AND main_stage_0_6 AND (rem_12cyc_st_5_1_0(0)));
  or_109_cse <= (rem_12cyc_st_5_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1159_nl <= nand_267_cse AND or_tmp_80;
  mux_tmp_41 <= MUX_s_1_2_2(and_1159_nl, or_tmp_80, or_109_cse);
  and_1160_nl <= nand_271_cse AND mux_tmp_41;
  mux_tmp_42 <= MUX_s_1_2_2(and_1160_nl, mux_tmp_41, or_100_cse);
  and_1161_nl <= nand_274_cse AND mux_tmp_42;
  mux_tmp_43 <= MUX_s_1_2_2(and_1161_nl, mux_tmp_42, or_93_cse);
  and_1162_nl <= nand_276_cse AND mux_tmp_43;
  mux_tmp_44 <= MUX_s_1_2_2(and_1162_nl, mux_tmp_43, or_88_cse);
  nor_495_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_44));
  mux_47_nl <= MUX_s_1_2_2(nor_495_nl, mux_tmp_44, or_83_cse);
  and_dcpl_376 <= mux_47_nl AND and_dcpl_112 AND and_dcpl_115;
  or_120_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_493_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_80));
  mux_tmp_46 <= MUX_s_1_2_2(nor_493_nl, or_tmp_80, or_120_cse);
  and_1155_nl <= nand_267_cse AND mux_tmp_46;
  mux_tmp_47 <= MUX_s_1_2_2(and_1155_nl, mux_tmp_46, or_109_cse);
  and_1156_nl <= nand_271_cse AND mux_tmp_47;
  mux_tmp_48 <= MUX_s_1_2_2(and_1156_nl, mux_tmp_47, or_100_cse);
  and_1157_nl <= nand_274_cse AND mux_tmp_48;
  mux_tmp_49 <= MUX_s_1_2_2(and_1157_nl, mux_tmp_48, or_93_cse);
  and_1158_nl <= nand_276_cse AND mux_tmp_49;
  mux_tmp_50 <= MUX_s_1_2_2(and_1158_nl, mux_tmp_49, or_88_cse);
  nor_494_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_50));
  mux_53_nl <= MUX_s_1_2_2(nor_494_nl, mux_tmp_50, or_83_cse);
  and_dcpl_379 <= mux_53_nl AND and_dcpl_85 AND and_dcpl_87;
  or_133_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_490_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_80));
  mux_tmp_52 <= MUX_s_1_2_2(nor_490_nl, or_tmp_80, or_133_cse);
  nor_491_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_52));
  mux_tmp_53 <= MUX_s_1_2_2(nor_491_nl, mux_tmp_52, or_120_cse);
  and_1151_nl <= nand_267_cse AND mux_tmp_53;
  mux_tmp_54 <= MUX_s_1_2_2(and_1151_nl, mux_tmp_53, or_109_cse);
  and_1152_nl <= nand_271_cse AND mux_tmp_54;
  mux_tmp_55 <= MUX_s_1_2_2(and_1152_nl, mux_tmp_54, or_100_cse);
  and_1153_nl <= nand_274_cse AND mux_tmp_55;
  mux_tmp_56 <= MUX_s_1_2_2(and_1153_nl, mux_tmp_55, or_93_cse);
  and_1154_nl <= nand_276_cse AND mux_tmp_56;
  mux_tmp_57 <= MUX_s_1_2_2(and_1154_nl, mux_tmp_56, or_88_cse);
  nor_492_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_57));
  mux_60_nl <= MUX_s_1_2_2(nor_492_nl, mux_tmp_57, or_83_cse);
  and_dcpl_382 <= mux_60_nl AND and_dcpl_58 AND and_dcpl_60;
  or_148_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_486_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_80));
  mux_tmp_59 <= MUX_s_1_2_2(nor_486_nl, or_tmp_80, or_148_cse);
  nor_487_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_59));
  mux_tmp_60 <= MUX_s_1_2_2(nor_487_nl, mux_tmp_59, or_133_cse);
  nor_488_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_60));
  mux_tmp_61 <= MUX_s_1_2_2(nor_488_nl, mux_tmp_60, or_120_cse);
  and_1147_nl <= nand_267_cse AND mux_tmp_61;
  mux_tmp_62 <= MUX_s_1_2_2(and_1147_nl, mux_tmp_61, or_109_cse);
  and_1148_nl <= nand_271_cse AND mux_tmp_62;
  mux_tmp_63 <= MUX_s_1_2_2(and_1148_nl, mux_tmp_62, or_100_cse);
  and_1149_nl <= nand_274_cse AND mux_tmp_63;
  mux_tmp_64 <= MUX_s_1_2_2(and_1149_nl, mux_tmp_63, or_93_cse);
  and_1150_nl <= nand_276_cse AND mux_tmp_64;
  mux_tmp_65 <= MUX_s_1_2_2(and_1150_nl, mux_tmp_64, or_88_cse);
  nor_489_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_65));
  mux_68_nl <= MUX_s_1_2_2(nor_489_nl, mux_tmp_65, or_83_cse);
  and_dcpl_385 <= mux_68_nl AND and_dcpl_31 AND and_dcpl_33;
  nor_481_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_80));
  or_165_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_67 <= MUX_s_1_2_2(nor_481_nl, or_tmp_80, or_165_nl);
  nor_482_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_67));
  mux_tmp_68 <= MUX_s_1_2_2(nor_482_nl, mux_tmp_67, or_148_cse);
  nor_483_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_68));
  mux_tmp_69 <= MUX_s_1_2_2(nor_483_nl, mux_tmp_68, or_133_cse);
  nor_484_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_69));
  mux_tmp_70 <= MUX_s_1_2_2(nor_484_nl, mux_tmp_69, or_120_cse);
  and_1143_nl <= nand_267_cse AND mux_tmp_70;
  mux_tmp_71 <= MUX_s_1_2_2(and_1143_nl, mux_tmp_70, or_109_cse);
  and_1144_nl <= nand_271_cse AND mux_tmp_71;
  mux_tmp_72 <= MUX_s_1_2_2(and_1144_nl, mux_tmp_71, or_100_cse);
  and_1145_nl <= nand_274_cse AND mux_tmp_72;
  mux_tmp_73 <= MUX_s_1_2_2(and_1145_nl, mux_tmp_72, or_93_cse);
  and_1146_nl <= nand_276_cse AND mux_tmp_73;
  mux_tmp_74 <= MUX_s_1_2_2(and_1146_nl, mux_tmp_73, or_88_cse);
  nor_485_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_74));
  mux_77_nl <= MUX_s_1_2_2(nor_485_nl, mux_tmp_74, or_83_cse);
  and_dcpl_388 <= mux_77_nl AND and_dcpl_4 AND and_dcpl_6;
  nand_250_cse <= NOT((acc_1_tmp(0)) AND ccs_ccore_start_rsci_idat);
  and_tmp_44 <= ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_9)
      OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_10)
      OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_3)
      OR (NOT asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_4)
      OR (NOT asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_5)
      OR (NOT asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_6)
      OR (NOT asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_7)
      OR (NOT asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_11)
      OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("00"))) AND (CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("00"))
      OR (acc_1_tmp(1)) OR nand_250_cse);
  nor_480_nl <= NOT((rem_12cyc_1_0(0)) OR (NOT and_tmp_44));
  or_175_nl <= (NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_1_0(1));
  mux_tmp_76 <= MUX_s_1_2_2(nor_480_nl, and_tmp_44, or_175_nl);
  and_dcpl_393 <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_394 <= and_dcpl_293 AND and_dcpl_393;
  and_dcpl_395 <= and_dcpl_295 AND (rem_12cyc_st_2_1_0(1));
  or_tmp_185 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_54;
  or_190_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("00"));
  nor_479_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_185));
  mux_79_nl <= MUX_s_1_2_2(nor_479_nl, or_tmp_185, or_190_cse);
  and_dcpl_397 <= mux_79_nl AND and_dcpl_298 AND and_dcpl_395;
  and_dcpl_398 <= and_dcpl_301 AND (rem_12cyc_st_3_1_0(1));
  or_195_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp_45 <= or_195_cse AND or_tmp_185;
  nor_478_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_45));
  mux_80_nl <= MUX_s_1_2_2(nor_478_nl, and_tmp_45, or_190_cse);
  and_dcpl_400 <= mux_80_nl AND and_dcpl_304 AND and_dcpl_398;
  and_dcpl_401 <= and_dcpl_307 AND (rem_12cyc_st_4_1_0(1));
  or_199_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_47 <= or_195_cse AND or_199_cse AND or_tmp_185;
  nor_477_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_47));
  mux_81_nl <= MUX_s_1_2_2(nor_477_nl, and_tmp_47, or_190_cse);
  and_dcpl_403 <= mux_81_nl AND and_dcpl_310 AND and_dcpl_401;
  and_dcpl_404 <= and_dcpl_313 AND (rem_12cyc_st_5_1_0(1));
  or_204_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_50 <= or_195_cse AND or_199_cse AND or_204_cse AND or_tmp_185;
  nor_476_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_50));
  mux_82_nl <= MUX_s_1_2_2(nor_476_nl, and_tmp_50, or_190_cse);
  and_dcpl_406 <= mux_82_nl AND and_dcpl_316 AND and_dcpl_404;
  or_210_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_54 <= or_195_cse AND or_199_cse AND or_204_cse AND or_210_cse AND or_tmp_185;
  nor_475_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_54));
  mux_83_nl <= MUX_s_1_2_2(nor_475_nl, and_tmp_54, or_190_cse);
  and_dcpl_409 <= mux_83_nl AND and_dcpl_112 AND and_dcpl_117;
  or_217_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_473_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_185));
  mux_84_nl <= MUX_s_1_2_2(nor_473_nl, or_tmp_185, or_217_cse);
  and_tmp_58 <= or_195_cse AND or_199_cse AND or_204_cse AND or_210_cse AND mux_84_nl;
  nor_474_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_58));
  mux_85_nl <= MUX_s_1_2_2(nor_474_nl, and_tmp_58, or_190_cse);
  and_dcpl_413 <= mux_85_nl AND and_dcpl_85 AND and_dcpl_90;
  or_226_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_470_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_185));
  mux_tmp_84 <= MUX_s_1_2_2(nor_470_nl, or_tmp_185, or_226_cse);
  nor_471_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_84));
  mux_87_nl <= MUX_s_1_2_2(nor_471_nl, mux_tmp_84, or_217_cse);
  and_tmp_62 <= or_195_cse AND or_199_cse AND or_204_cse AND or_210_cse AND mux_87_nl;
  nor_472_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_62));
  mux_88_nl <= MUX_s_1_2_2(nor_472_nl, and_tmp_62, or_190_cse);
  and_dcpl_417 <= mux_88_nl AND and_dcpl_58 AND and_dcpl_63;
  or_237_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_466_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_185));
  mux_tmp_87 <= MUX_s_1_2_2(nor_466_nl, or_tmp_185, or_237_cse);
  nor_467_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_87));
  mux_tmp_88 <= MUX_s_1_2_2(nor_467_nl, mux_tmp_87, or_226_cse);
  nor_468_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_88));
  mux_91_nl <= MUX_s_1_2_2(nor_468_nl, mux_tmp_88, or_217_cse);
  and_tmp_66 <= or_195_cse AND or_199_cse AND or_204_cse AND or_210_cse AND mux_91_nl;
  nor_469_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_66));
  mux_92_nl <= MUX_s_1_2_2(nor_469_nl, and_tmp_66, or_190_cse);
  and_dcpl_421 <= mux_92_nl AND and_dcpl_31 AND and_dcpl_36;
  nor_461_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_185));
  or_250_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_91 <= MUX_s_1_2_2(nor_461_nl, or_tmp_185, or_250_nl);
  nor_462_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_91));
  mux_tmp_92 <= MUX_s_1_2_2(nor_462_nl, mux_tmp_91, or_237_cse);
  nor_463_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_92));
  mux_tmp_93 <= MUX_s_1_2_2(nor_463_nl, mux_tmp_92, or_226_cse);
  nor_464_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_93));
  mux_96_nl <= MUX_s_1_2_2(nor_464_nl, mux_tmp_93, or_217_cse);
  and_tmp_70 <= or_195_cse AND or_199_cse AND or_204_cse AND or_210_cse AND mux_96_nl;
  nor_465_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_70));
  mux_97_nl <= MUX_s_1_2_2(nor_465_nl, and_tmp_70, or_190_cse);
  and_dcpl_425 <= mux_97_nl AND and_dcpl_4 AND and_dcpl_9;
  and_tmp_80 <= ((NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10"))) AND ((NOT main_stage_0_8)
      OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_9)
      OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_10)
      OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"))) AND or_195_cse
      AND or_199_cse AND or_204_cse AND or_210_cse AND ((NOT main_stage_0_7) OR (NOT
      asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00")))
      AND ((NOT main_stage_0_11) OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("00"))) AND (CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT ccs_ccore_start_rsci_idat));
  and_dcpl_430 <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_431 <= and_dcpl_293 AND and_dcpl_430;
  or_tmp_263 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_54;
  or_270_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("00"));
  nor_460_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_263));
  mux_98_nl <= MUX_s_1_2_2(nor_460_nl, or_tmp_263, or_270_cse);
  and_dcpl_433 <= mux_98_nl AND and_dcpl_358 AND and_dcpl_395;
  or_275_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1142_nl <= nand_276_cse AND or_tmp_263;
  mux_tmp_97 <= MUX_s_1_2_2(and_1142_nl, or_tmp_263, or_275_cse);
  nor_459_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_97));
  mux_100_nl <= MUX_s_1_2_2(nor_459_nl, mux_tmp_97, or_270_cse);
  and_dcpl_435 <= mux_100_nl AND and_dcpl_362 AND and_dcpl_398;
  or_280_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1140_nl <= nand_274_cse AND or_tmp_263;
  mux_tmp_99 <= MUX_s_1_2_2(and_1140_nl, or_tmp_263, or_280_cse);
  and_1141_nl <= nand_276_cse AND mux_tmp_99;
  mux_tmp_100 <= MUX_s_1_2_2(and_1141_nl, mux_tmp_99, or_275_cse);
  nor_458_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_100));
  mux_103_nl <= MUX_s_1_2_2(nor_458_nl, mux_tmp_100, or_270_cse);
  and_dcpl_437 <= mux_103_nl AND and_dcpl_366 AND and_dcpl_401;
  or_287_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1137_nl <= nand_271_cse AND or_tmp_263;
  mux_tmp_102 <= MUX_s_1_2_2(and_1137_nl, or_tmp_263, or_287_cse);
  and_1138_nl <= nand_274_cse AND mux_tmp_102;
  mux_tmp_103 <= MUX_s_1_2_2(and_1138_nl, mux_tmp_102, or_280_cse);
  and_1139_nl <= nand_276_cse AND mux_tmp_103;
  mux_tmp_104 <= MUX_s_1_2_2(and_1139_nl, mux_tmp_103, or_275_cse);
  nor_457_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_104));
  mux_107_nl <= MUX_s_1_2_2(nor_457_nl, mux_tmp_104, or_270_cse);
  and_dcpl_439 <= mux_107_nl AND and_dcpl_370 AND and_dcpl_404;
  or_296_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1133_nl <= nand_267_cse AND or_tmp_263;
  mux_tmp_106 <= MUX_s_1_2_2(and_1133_nl, or_tmp_263, or_296_cse);
  and_1134_nl <= nand_271_cse AND mux_tmp_106;
  mux_tmp_107 <= MUX_s_1_2_2(and_1134_nl, mux_tmp_106, or_287_cse);
  and_1135_nl <= nand_274_cse AND mux_tmp_107;
  mux_tmp_108 <= MUX_s_1_2_2(and_1135_nl, mux_tmp_107, or_280_cse);
  and_1136_nl <= nand_276_cse AND mux_tmp_108;
  mux_tmp_109 <= MUX_s_1_2_2(and_1136_nl, mux_tmp_108, or_275_cse);
  nor_456_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_109));
  mux_112_nl <= MUX_s_1_2_2(nor_456_nl, mux_tmp_109, or_270_cse);
  and_dcpl_442 <= mux_112_nl AND and_dcpl_112 AND and_dcpl_119;
  or_307_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_454_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_263));
  mux_tmp_111 <= MUX_s_1_2_2(nor_454_nl, or_tmp_263, or_307_cse);
  and_1129_nl <= nand_267_cse AND mux_tmp_111;
  mux_tmp_112 <= MUX_s_1_2_2(and_1129_nl, mux_tmp_111, or_296_cse);
  and_1130_nl <= nand_271_cse AND mux_tmp_112;
  mux_tmp_113 <= MUX_s_1_2_2(and_1130_nl, mux_tmp_112, or_287_cse);
  and_1131_nl <= nand_274_cse AND mux_tmp_113;
  mux_tmp_114 <= MUX_s_1_2_2(and_1131_nl, mux_tmp_113, or_280_cse);
  and_1132_nl <= nand_276_cse AND mux_tmp_114;
  mux_tmp_115 <= MUX_s_1_2_2(and_1132_nl, mux_tmp_114, or_275_cse);
  nor_455_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_115));
  mux_118_nl <= MUX_s_1_2_2(nor_455_nl, mux_tmp_115, or_270_cse);
  and_dcpl_445 <= mux_118_nl AND and_dcpl_85 AND and_dcpl_92;
  or_320_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_451_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_263));
  mux_tmp_117 <= MUX_s_1_2_2(nor_451_nl, or_tmp_263, or_320_cse);
  nor_452_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_117));
  mux_tmp_118 <= MUX_s_1_2_2(nor_452_nl, mux_tmp_117, or_307_cse);
  and_1125_nl <= nand_267_cse AND mux_tmp_118;
  mux_tmp_119 <= MUX_s_1_2_2(and_1125_nl, mux_tmp_118, or_296_cse);
  and_1126_nl <= nand_271_cse AND mux_tmp_119;
  mux_tmp_120 <= MUX_s_1_2_2(and_1126_nl, mux_tmp_119, or_287_cse);
  and_1127_nl <= nand_274_cse AND mux_tmp_120;
  mux_tmp_121 <= MUX_s_1_2_2(and_1127_nl, mux_tmp_120, or_280_cse);
  and_1128_nl <= nand_276_cse AND mux_tmp_121;
  mux_tmp_122 <= MUX_s_1_2_2(and_1128_nl, mux_tmp_121, or_275_cse);
  nor_453_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_122));
  mux_125_nl <= MUX_s_1_2_2(nor_453_nl, mux_tmp_122, or_270_cse);
  and_dcpl_448 <= mux_125_nl AND and_dcpl_58 AND and_dcpl_65;
  or_335_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_447_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_263));
  mux_tmp_124 <= MUX_s_1_2_2(nor_447_nl, or_tmp_263, or_335_cse);
  nor_448_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_124));
  mux_tmp_125 <= MUX_s_1_2_2(nor_448_nl, mux_tmp_124, or_320_cse);
  nor_449_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_125));
  mux_tmp_126 <= MUX_s_1_2_2(nor_449_nl, mux_tmp_125, or_307_cse);
  and_1121_nl <= nand_267_cse AND mux_tmp_126;
  mux_tmp_127 <= MUX_s_1_2_2(and_1121_nl, mux_tmp_126, or_296_cse);
  and_1122_nl <= nand_271_cse AND mux_tmp_127;
  mux_tmp_128 <= MUX_s_1_2_2(and_1122_nl, mux_tmp_127, or_287_cse);
  and_1123_nl <= nand_274_cse AND mux_tmp_128;
  mux_tmp_129 <= MUX_s_1_2_2(and_1123_nl, mux_tmp_128, or_280_cse);
  and_1124_nl <= nand_276_cse AND mux_tmp_129;
  mux_tmp_130 <= MUX_s_1_2_2(and_1124_nl, mux_tmp_129, or_275_cse);
  nor_450_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_130));
  mux_133_nl <= MUX_s_1_2_2(nor_450_nl, mux_tmp_130, or_270_cse);
  and_dcpl_451 <= mux_133_nl AND and_dcpl_31 AND and_dcpl_38;
  nor_442_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_263));
  or_352_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_132 <= MUX_s_1_2_2(nor_442_nl, or_tmp_263, or_352_nl);
  nor_443_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_132));
  mux_tmp_133 <= MUX_s_1_2_2(nor_443_nl, mux_tmp_132, or_335_cse);
  nor_444_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_133));
  mux_tmp_134 <= MUX_s_1_2_2(nor_444_nl, mux_tmp_133, or_320_cse);
  nor_445_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_134));
  mux_tmp_135 <= MUX_s_1_2_2(nor_445_nl, mux_tmp_134, or_307_cse);
  and_1117_nl <= nand_267_cse AND mux_tmp_135;
  mux_tmp_136 <= MUX_s_1_2_2(and_1117_nl, mux_tmp_135, or_296_cse);
  and_1118_nl <= nand_271_cse AND mux_tmp_136;
  mux_tmp_137 <= MUX_s_1_2_2(and_1118_nl, mux_tmp_136, or_287_cse);
  and_1119_nl <= nand_274_cse AND mux_tmp_137;
  mux_tmp_138 <= MUX_s_1_2_2(and_1119_nl, mux_tmp_137, or_280_cse);
  and_1120_nl <= nand_276_cse AND mux_tmp_138;
  mux_tmp_139 <= MUX_s_1_2_2(and_1120_nl, mux_tmp_138, or_275_cse);
  nor_446_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_139));
  mux_142_nl <= MUX_s_1_2_2(nor_446_nl, mux_tmp_139, or_270_cse);
  and_dcpl_454 <= mux_142_nl AND and_dcpl_4 AND and_dcpl_11;
  nand_222_cse <= NOT(CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND ccs_ccore_start_rsci_idat);
  and_tmp_89 <= ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_9)
      OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_10)
      OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_3)
      OR (NOT asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_4)
      OR (NOT asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_5)
      OR (NOT asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_6)
      OR (NOT asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_7)
      OR (NOT asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_11)
      OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("00"))) AND (CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("00"))
      OR nand_222_cse);
  nand_223_cse <= NOT(CONV_SL_1_1(rem_12cyc_1_0=STD_LOGIC_VECTOR'("11")));
  and_1116_nl <= nand_223_cse AND and_tmp_89;
  or_362_nl <= (NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_141 <= MUX_s_1_2_2(and_1116_nl, and_tmp_89, or_362_nl);
  and_dcpl_460 <= ccs_ccore_start_rsci_idat AND CONV_SL_1_1(acc_tmp=STD_LOGIC_VECTOR'("01"));
  and_dcpl_461 <= and_dcpl_460 AND and_dcpl_291;
  and_dcpl_462 <= CONV_SL_1_1(rem_12cyc_st_2_3_2=STD_LOGIC_VECTOR'("01"));
  and_dcpl_463 <= and_dcpl_462 AND (NOT (rem_12cyc_st_2_1_0(1)));
  not_tmp_332 <= NOT((rem_12cyc_3_2(0)) AND asn_itm_1 AND main_stage_0_2);
  or_tmp_368 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00")) OR (rem_12cyc_3_2(1))
      OR not_tmp_332;
  nand_281_cse <= NOT((acc_tmp(0)) AND ccs_ccore_start_rsci_idat);
  or_377_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (acc_tmp(1));
  and_1172_nl <= nand_281_cse AND or_tmp_368;
  mux_144_nl <= MUX_s_1_2_2(and_1172_nl, or_tmp_368, or_377_cse);
  and_dcpl_465 <= mux_144_nl AND and_dcpl_298 AND and_dcpl_463;
  and_dcpl_466 <= CONV_SL_1_1(rem_12cyc_st_3_3_2=STD_LOGIC_VECTOR'("01"));
  and_dcpl_467 <= and_dcpl_466 AND (NOT (rem_12cyc_st_3_1_0(1)));
  or_382_cse <= (rem_12cyc_st_2_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp_90 <= or_382_cse AND or_tmp_368;
  and_1114_nl <= nand_281_cse AND and_tmp_90;
  mux_145_nl <= MUX_s_1_2_2(and_1114_nl, and_tmp_90, or_377_cse);
  and_dcpl_469 <= mux_145_nl AND and_dcpl_304 AND and_dcpl_467;
  and_dcpl_470 <= CONV_SL_1_1(rem_12cyc_st_4_3_2=STD_LOGIC_VECTOR'("01"));
  and_dcpl_471 <= and_dcpl_470 AND (NOT (rem_12cyc_st_4_1_0(1)));
  or_386_cse <= (rem_12cyc_st_3_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_92 <= or_382_cse AND or_386_cse AND or_tmp_368;
  and_1113_nl <= nand_281_cse AND and_tmp_92;
  mux_146_nl <= MUX_s_1_2_2(and_1113_nl, and_tmp_92, or_377_cse);
  and_dcpl_473 <= mux_146_nl AND and_dcpl_310 AND and_dcpl_471;
  and_dcpl_474 <= CONV_SL_1_1(rem_12cyc_st_5_3_2=STD_LOGIC_VECTOR'("01"));
  and_dcpl_475 <= and_dcpl_474 AND (NOT (rem_12cyc_st_5_1_0(1)));
  or_391_cse <= (rem_12cyc_st_4_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_95 <= or_382_cse AND or_386_cse AND or_391_cse AND or_tmp_368;
  and_1112_nl <= nand_281_cse AND and_tmp_95;
  mux_147_nl <= MUX_s_1_2_2(and_1112_nl, and_tmp_95, or_377_cse);
  and_dcpl_477 <= mux_147_nl AND and_dcpl_316 AND and_dcpl_475;
  or_397_cse <= (rem_12cyc_st_5_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_99 <= or_382_cse AND or_386_cse AND or_391_cse AND or_397_cse AND or_tmp_368;
  and_1111_nl <= nand_281_cse AND and_tmp_99;
  mux_148_nl <= MUX_s_1_2_2(and_1111_nl, and_tmp_99, or_377_cse);
  and_dcpl_480 <= mux_148_nl AND and_dcpl_121 AND and_dcpl_110;
  nand_215_cse <= NOT((rem_12cyc_st_6_3_2(0)) AND asn_itm_6 AND main_stage_0_7);
  or_404_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00")) OR (rem_12cyc_st_6_3_2(1));
  and_1109_nl <= nand_215_cse AND or_tmp_368;
  mux_149_nl <= MUX_s_1_2_2(and_1109_nl, or_tmp_368, or_404_cse);
  and_tmp_103 <= or_382_cse AND or_386_cse AND or_391_cse AND or_397_cse AND mux_149_nl;
  and_1110_nl <= nand_281_cse AND and_tmp_103;
  mux_150_nl <= MUX_s_1_2_2(and_1110_nl, and_tmp_103, or_377_cse);
  and_dcpl_483 <= mux_150_nl AND and_dcpl_94 AND and_dcpl_83;
  nand_212_cse <= NOT((rem_12cyc_st_7_3_2(0)) AND asn_itm_7 AND main_stage_0_8);
  or_413_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00")) OR (rem_12cyc_st_7_3_2(1));
  and_1106_nl <= nand_212_cse AND or_tmp_368;
  mux_tmp_149 <= MUX_s_1_2_2(and_1106_nl, or_tmp_368, or_413_cse);
  and_1107_nl <= nand_215_cse AND mux_tmp_149;
  mux_152_nl <= MUX_s_1_2_2(and_1107_nl, mux_tmp_149, or_404_cse);
  and_tmp_107 <= or_382_cse AND or_386_cse AND or_391_cse AND or_397_cse AND mux_152_nl;
  and_1108_nl <= nand_281_cse AND and_tmp_107;
  mux_153_nl <= MUX_s_1_2_2(and_1108_nl, and_tmp_107, or_377_cse);
  and_dcpl_486 <= mux_153_nl AND and_dcpl_67 AND and_dcpl_56;
  nand_208_cse <= NOT((rem_12cyc_st_8_3_2(0)) AND asn_itm_8 AND main_stage_0_9);
  or_424_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00")) OR (rem_12cyc_st_8_3_2(1));
  and_1102_nl <= nand_208_cse AND or_tmp_368;
  mux_tmp_152 <= MUX_s_1_2_2(and_1102_nl, or_tmp_368, or_424_cse);
  and_1103_nl <= nand_212_cse AND mux_tmp_152;
  mux_tmp_153 <= MUX_s_1_2_2(and_1103_nl, mux_tmp_152, or_413_cse);
  and_1104_nl <= nand_215_cse AND mux_tmp_153;
  mux_156_nl <= MUX_s_1_2_2(and_1104_nl, mux_tmp_153, or_404_cse);
  and_tmp_111 <= or_382_cse AND or_386_cse AND or_391_cse AND or_397_cse AND mux_156_nl;
  and_1105_nl <= nand_281_cse AND and_tmp_111;
  mux_157_nl <= MUX_s_1_2_2(and_1105_nl, and_tmp_111, or_377_cse);
  and_dcpl_489 <= mux_157_nl AND and_dcpl_40 AND and_dcpl_29;
  nand_203_cse <= NOT((rem_12cyc_st_9_3_2(0)) AND asn_itm_9 AND main_stage_0_10);
  and_1097_nl <= nand_203_cse AND or_tmp_368;
  or_437_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00")) OR (rem_12cyc_st_9_3_2(1));
  mux_tmp_156 <= MUX_s_1_2_2(and_1097_nl, or_tmp_368, or_437_nl);
  and_1098_nl <= nand_208_cse AND mux_tmp_156;
  mux_tmp_157 <= MUX_s_1_2_2(and_1098_nl, mux_tmp_156, or_424_cse);
  and_1099_nl <= nand_212_cse AND mux_tmp_157;
  mux_tmp_158 <= MUX_s_1_2_2(and_1099_nl, mux_tmp_157, or_413_cse);
  and_1100_nl <= nand_215_cse AND mux_tmp_158;
  mux_161_nl <= MUX_s_1_2_2(and_1100_nl, mux_tmp_158, or_404_cse);
  and_tmp_115 <= or_382_cse AND or_386_cse AND or_391_cse AND or_397_cse AND mux_161_nl;
  and_1101_nl <= nand_281_cse AND and_tmp_115;
  mux_162_nl <= MUX_s_1_2_2(and_1101_nl, and_tmp_115, or_377_cse);
  and_dcpl_492 <= mux_162_nl AND and_dcpl_13 AND and_dcpl_2;
  and_tmp_125 <= ((NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_8)
      OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_9)
      OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_10)
      OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("01"))) AND or_382_cse
      AND or_386_cse AND or_391_cse AND or_397_cse AND ((NOT main_stage_0_7) OR (NOT
      asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("01")))
      AND ((NOT main_stage_0_11) OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("01"))) AND (CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT ccs_ccore_start_rsci_idat));
  and_dcpl_498 <= and_dcpl_460 AND and_dcpl_355;
  or_tmp_446 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("01")) OR (rem_12cyc_3_2(1))
      OR not_tmp_332;
  or_458_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (acc_tmp(1));
  and_1171_nl <= nand_281_cse AND or_tmp_446;
  mux_163_nl <= MUX_s_1_2_2(and_1171_nl, or_tmp_446, or_458_cse);
  and_dcpl_500 <= mux_163_nl AND and_dcpl_358 AND and_dcpl_463;
  or_463_cse <= (rem_12cyc_st_2_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("01"));
  and_1094_nl <= nand_276_cse AND or_tmp_446;
  mux_tmp_162 <= MUX_s_1_2_2(and_1094_nl, or_tmp_446, or_463_cse);
  and_1095_nl <= nand_281_cse AND mux_tmp_162;
  mux_165_nl <= MUX_s_1_2_2(and_1095_nl, mux_tmp_162, or_458_cse);
  and_dcpl_502 <= mux_165_nl AND and_dcpl_362 AND and_dcpl_467;
  nand_198_cse <= NOT((rem_12cyc_st_3_3_2(0)) AND asn_itm_3 AND main_stage_0_4 AND
      (rem_12cyc_st_3_1_0(0)));
  or_468_cse <= (rem_12cyc_st_3_1_0(1)) OR (rem_12cyc_st_3_3_2(1));
  and_1091_nl <= nand_198_cse AND or_tmp_446;
  mux_tmp_164 <= MUX_s_1_2_2(and_1091_nl, or_tmp_446, or_468_cse);
  and_1092_nl <= nand_276_cse AND mux_tmp_164;
  mux_tmp_165 <= MUX_s_1_2_2(and_1092_nl, mux_tmp_164, or_463_cse);
  and_1093_nl <= nand_281_cse AND mux_tmp_165;
  mux_168_nl <= MUX_s_1_2_2(and_1093_nl, mux_tmp_165, or_458_cse);
  and_dcpl_504 <= mux_168_nl AND and_dcpl_366 AND and_dcpl_471;
  or_475_cse <= (rem_12cyc_st_4_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("01"));
  and_1087_nl <= nand_271_cse AND or_tmp_446;
  mux_tmp_167 <= MUX_s_1_2_2(and_1087_nl, or_tmp_446, or_475_cse);
  and_1088_nl <= nand_198_cse AND mux_tmp_167;
  mux_tmp_168 <= MUX_s_1_2_2(and_1088_nl, mux_tmp_167, or_468_cse);
  and_1089_nl <= nand_276_cse AND mux_tmp_168;
  mux_tmp_169 <= MUX_s_1_2_2(and_1089_nl, mux_tmp_168, or_463_cse);
  and_1090_nl <= nand_281_cse AND mux_tmp_169;
  mux_172_nl <= MUX_s_1_2_2(and_1090_nl, mux_tmp_169, or_458_cse);
  and_dcpl_506 <= mux_172_nl AND and_dcpl_370 AND and_dcpl_475;
  nand_189_cse <= NOT((rem_12cyc_st_5_3_2(0)) AND asn_itm_5 AND main_stage_0_6 AND
      (rem_12cyc_st_5_1_0(0)));
  or_484_cse <= (rem_12cyc_st_5_1_0(1)) OR (rem_12cyc_st_5_3_2(1));
  and_1082_nl <= nand_189_cse AND or_tmp_446;
  mux_tmp_171 <= MUX_s_1_2_2(and_1082_nl, or_tmp_446, or_484_cse);
  and_1083_nl <= nand_271_cse AND mux_tmp_171;
  mux_tmp_172 <= MUX_s_1_2_2(and_1083_nl, mux_tmp_171, or_475_cse);
  and_1084_nl <= nand_198_cse AND mux_tmp_172;
  mux_tmp_173 <= MUX_s_1_2_2(and_1084_nl, mux_tmp_172, or_468_cse);
  and_1085_nl <= nand_276_cse AND mux_tmp_173;
  mux_tmp_174 <= MUX_s_1_2_2(and_1085_nl, mux_tmp_173, or_463_cse);
  and_1086_nl <= nand_281_cse AND mux_tmp_174;
  mux_177_nl <= MUX_s_1_2_2(and_1086_nl, mux_tmp_174, or_458_cse);
  and_dcpl_508 <= mux_177_nl AND and_dcpl_121 AND and_dcpl_115;
  or_495_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01")) OR (rem_12cyc_st_6_3_2(1));
  and_1076_nl <= nand_215_cse AND or_tmp_446;
  mux_tmp_176 <= MUX_s_1_2_2(and_1076_nl, or_tmp_446, or_495_cse);
  and_1077_nl <= nand_189_cse AND mux_tmp_176;
  mux_tmp_177 <= MUX_s_1_2_2(and_1077_nl, mux_tmp_176, or_484_cse);
  and_1078_nl <= nand_271_cse AND mux_tmp_177;
  mux_tmp_178 <= MUX_s_1_2_2(and_1078_nl, mux_tmp_177, or_475_cse);
  and_1079_nl <= nand_198_cse AND mux_tmp_178;
  mux_tmp_179 <= MUX_s_1_2_2(and_1079_nl, mux_tmp_178, or_468_cse);
  and_1080_nl <= nand_276_cse AND mux_tmp_179;
  mux_tmp_180 <= MUX_s_1_2_2(and_1080_nl, mux_tmp_179, or_463_cse);
  and_1081_nl <= nand_281_cse AND mux_tmp_180;
  mux_183_nl <= MUX_s_1_2_2(and_1081_nl, mux_tmp_180, or_458_cse);
  and_dcpl_510 <= mux_183_nl AND and_dcpl_94 AND and_dcpl_87;
  or_508_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01")) OR (rem_12cyc_st_7_3_2(1));
  and_1069_nl <= nand_212_cse AND or_tmp_446;
  mux_tmp_182 <= MUX_s_1_2_2(and_1069_nl, or_tmp_446, or_508_cse);
  and_1070_nl <= nand_215_cse AND mux_tmp_182;
  mux_tmp_183 <= MUX_s_1_2_2(and_1070_nl, mux_tmp_182, or_495_cse);
  and_1071_nl <= nand_189_cse AND mux_tmp_183;
  mux_tmp_184 <= MUX_s_1_2_2(and_1071_nl, mux_tmp_183, or_484_cse);
  and_1072_nl <= nand_271_cse AND mux_tmp_184;
  mux_tmp_185 <= MUX_s_1_2_2(and_1072_nl, mux_tmp_184, or_475_cse);
  and_1073_nl <= nand_198_cse AND mux_tmp_185;
  mux_tmp_186 <= MUX_s_1_2_2(and_1073_nl, mux_tmp_185, or_468_cse);
  and_1074_nl <= nand_276_cse AND mux_tmp_186;
  mux_tmp_187 <= MUX_s_1_2_2(and_1074_nl, mux_tmp_186, or_463_cse);
  and_1075_nl <= nand_281_cse AND mux_tmp_187;
  mux_190_nl <= MUX_s_1_2_2(and_1075_nl, mux_tmp_187, or_458_cse);
  and_dcpl_512 <= mux_190_nl AND and_dcpl_67 AND and_dcpl_60;
  or_523_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01")) OR (rem_12cyc_st_8_3_2(1));
  and_1061_nl <= nand_208_cse AND or_tmp_446;
  mux_tmp_189 <= MUX_s_1_2_2(and_1061_nl, or_tmp_446, or_523_cse);
  and_1062_nl <= nand_212_cse AND mux_tmp_189;
  mux_tmp_190 <= MUX_s_1_2_2(and_1062_nl, mux_tmp_189, or_508_cse);
  and_1063_nl <= nand_215_cse AND mux_tmp_190;
  mux_tmp_191 <= MUX_s_1_2_2(and_1063_nl, mux_tmp_190, or_495_cse);
  and_1064_nl <= nand_189_cse AND mux_tmp_191;
  mux_tmp_192 <= MUX_s_1_2_2(and_1064_nl, mux_tmp_191, or_484_cse);
  and_1065_nl <= nand_271_cse AND mux_tmp_192;
  mux_tmp_193 <= MUX_s_1_2_2(and_1065_nl, mux_tmp_192, or_475_cse);
  and_1066_nl <= nand_198_cse AND mux_tmp_193;
  mux_tmp_194 <= MUX_s_1_2_2(and_1066_nl, mux_tmp_193, or_468_cse);
  and_1067_nl <= nand_276_cse AND mux_tmp_194;
  mux_tmp_195 <= MUX_s_1_2_2(and_1067_nl, mux_tmp_194, or_463_cse);
  and_1068_nl <= nand_281_cse AND mux_tmp_195;
  mux_198_nl <= MUX_s_1_2_2(and_1068_nl, mux_tmp_195, or_458_cse);
  and_dcpl_514 <= mux_198_nl AND and_dcpl_40 AND and_dcpl_33;
  and_1052_nl <= nand_203_cse AND or_tmp_446;
  or_540_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01")) OR (rem_12cyc_st_9_3_2(1));
  mux_tmp_197 <= MUX_s_1_2_2(and_1052_nl, or_tmp_446, or_540_nl);
  and_1053_nl <= nand_208_cse AND mux_tmp_197;
  mux_tmp_198 <= MUX_s_1_2_2(and_1053_nl, mux_tmp_197, or_523_cse);
  and_1054_nl <= nand_212_cse AND mux_tmp_198;
  mux_tmp_199 <= MUX_s_1_2_2(and_1054_nl, mux_tmp_198, or_508_cse);
  and_1055_nl <= nand_215_cse AND mux_tmp_199;
  mux_tmp_200 <= MUX_s_1_2_2(and_1055_nl, mux_tmp_199, or_495_cse);
  and_1056_nl <= nand_189_cse AND mux_tmp_200;
  mux_tmp_201 <= MUX_s_1_2_2(and_1056_nl, mux_tmp_200, or_484_cse);
  and_1057_nl <= nand_271_cse AND mux_tmp_201;
  mux_tmp_202 <= MUX_s_1_2_2(and_1057_nl, mux_tmp_201, or_475_cse);
  and_1058_nl <= nand_198_cse AND mux_tmp_202;
  mux_tmp_203 <= MUX_s_1_2_2(and_1058_nl, mux_tmp_202, or_468_cse);
  and_1059_nl <= nand_276_cse AND mux_tmp_203;
  mux_tmp_204 <= MUX_s_1_2_2(and_1059_nl, mux_tmp_203, or_463_cse);
  and_1060_nl <= nand_281_cse AND mux_tmp_204;
  mux_207_nl <= MUX_s_1_2_2(and_1060_nl, mux_tmp_204, or_458_cse);
  and_dcpl_516 <= mux_207_nl AND and_dcpl_13 AND and_dcpl_6;
  and_tmp_134 <= ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_9)
      OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_10)
      OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_3)
      OR (NOT asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_4)
      OR (NOT asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_5)
      OR (NOT asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_6)
      OR (NOT asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_7)
      OR (NOT asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_11)
      OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("01"))) AND (CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("01"))
      OR (acc_1_tmp(1)) OR nand_250_cse);
  nor_439_nl <= NOT((rem_12cyc_1_0(0)) OR (NOT and_tmp_134));
  or_550_nl <= (NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_1_0(1));
  mux_tmp_206 <= MUX_s_1_2_2(nor_439_nl, and_tmp_134, or_550_nl);
  and_dcpl_520 <= and_dcpl_460 AND and_dcpl_393;
  and_dcpl_521 <= and_dcpl_462 AND (rem_12cyc_st_2_1_0(1));
  or_tmp_551 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10")) OR (rem_12cyc_3_2(1))
      OR not_tmp_332;
  or_564_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (acc_tmp(1));
  and_1170_nl <= nand_281_cse AND or_tmp_551;
  mux_209_nl <= MUX_s_1_2_2(and_1170_nl, or_tmp_551, or_564_cse);
  and_dcpl_523 <= mux_209_nl AND and_dcpl_298 AND and_dcpl_521;
  and_dcpl_524 <= and_dcpl_466 AND (rem_12cyc_st_3_1_0(1));
  or_569_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp_135 <= or_569_cse AND or_tmp_551;
  and_1050_nl <= nand_281_cse AND and_tmp_135;
  mux_210_nl <= MUX_s_1_2_2(and_1050_nl, and_tmp_135, or_564_cse);
  and_dcpl_526 <= mux_210_nl AND and_dcpl_304 AND and_dcpl_524;
  and_dcpl_527 <= and_dcpl_470 AND (rem_12cyc_st_4_1_0(1));
  or_573_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_137 <= or_569_cse AND or_573_cse AND or_tmp_551;
  and_1049_nl <= nand_281_cse AND and_tmp_137;
  mux_211_nl <= MUX_s_1_2_2(and_1049_nl, and_tmp_137, or_564_cse);
  and_dcpl_529 <= mux_211_nl AND and_dcpl_310 AND and_dcpl_527;
  and_dcpl_530 <= and_dcpl_474 AND (rem_12cyc_st_5_1_0(1));
  or_578_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_140 <= or_569_cse AND or_573_cse AND or_578_cse AND or_tmp_551;
  and_1048_nl <= nand_281_cse AND and_tmp_140;
  mux_212_nl <= MUX_s_1_2_2(and_1048_nl, and_tmp_140, or_564_cse);
  and_dcpl_532 <= mux_212_nl AND and_dcpl_316 AND and_dcpl_530;
  or_584_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_144 <= or_569_cse AND or_573_cse AND or_578_cse AND or_584_cse AND or_tmp_551;
  and_1047_nl <= nand_281_cse AND and_tmp_144;
  mux_213_nl <= MUX_s_1_2_2(and_1047_nl, and_tmp_144, or_564_cse);
  and_dcpl_534 <= mux_213_nl AND and_dcpl_121 AND and_dcpl_117;
  or_591_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10")) OR (rem_12cyc_st_6_3_2(1));
  and_1045_nl <= nand_215_cse AND or_tmp_551;
  mux_214_nl <= MUX_s_1_2_2(and_1045_nl, or_tmp_551, or_591_cse);
  and_tmp_148 <= or_569_cse AND or_573_cse AND or_578_cse AND or_584_cse AND mux_214_nl;
  and_1046_nl <= nand_281_cse AND and_tmp_148;
  mux_215_nl <= MUX_s_1_2_2(and_1046_nl, and_tmp_148, or_564_cse);
  and_dcpl_536 <= mux_215_nl AND and_dcpl_94 AND and_dcpl_90;
  or_600_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10")) OR (rem_12cyc_st_7_3_2(1));
  and_1042_nl <= nand_212_cse AND or_tmp_551;
  mux_tmp_214 <= MUX_s_1_2_2(and_1042_nl, or_tmp_551, or_600_cse);
  and_1043_nl <= nand_215_cse AND mux_tmp_214;
  mux_217_nl <= MUX_s_1_2_2(and_1043_nl, mux_tmp_214, or_591_cse);
  and_tmp_152 <= or_569_cse AND or_573_cse AND or_578_cse AND or_584_cse AND mux_217_nl;
  and_1044_nl <= nand_281_cse AND and_tmp_152;
  mux_218_nl <= MUX_s_1_2_2(and_1044_nl, and_tmp_152, or_564_cse);
  and_dcpl_538 <= mux_218_nl AND and_dcpl_67 AND and_dcpl_63;
  or_611_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10")) OR (rem_12cyc_st_8_3_2(1));
  and_1038_nl <= nand_208_cse AND or_tmp_551;
  mux_tmp_217 <= MUX_s_1_2_2(and_1038_nl, or_tmp_551, or_611_cse);
  and_1039_nl <= nand_212_cse AND mux_tmp_217;
  mux_tmp_218 <= MUX_s_1_2_2(and_1039_nl, mux_tmp_217, or_600_cse);
  and_1040_nl <= nand_215_cse AND mux_tmp_218;
  mux_221_nl <= MUX_s_1_2_2(and_1040_nl, mux_tmp_218, or_591_cse);
  and_tmp_156 <= or_569_cse AND or_573_cse AND or_578_cse AND or_584_cse AND mux_221_nl;
  and_1041_nl <= nand_281_cse AND and_tmp_156;
  mux_222_nl <= MUX_s_1_2_2(and_1041_nl, and_tmp_156, or_564_cse);
  and_dcpl_540 <= mux_222_nl AND and_dcpl_40 AND and_dcpl_36;
  and_1033_nl <= nand_203_cse AND or_tmp_551;
  or_624_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10")) OR (rem_12cyc_st_9_3_2(1));
  mux_tmp_221 <= MUX_s_1_2_2(and_1033_nl, or_tmp_551, or_624_nl);
  and_1034_nl <= nand_208_cse AND mux_tmp_221;
  mux_tmp_222 <= MUX_s_1_2_2(and_1034_nl, mux_tmp_221, or_611_cse);
  and_1035_nl <= nand_212_cse AND mux_tmp_222;
  mux_tmp_223 <= MUX_s_1_2_2(and_1035_nl, mux_tmp_222, or_600_cse);
  and_1036_nl <= nand_215_cse AND mux_tmp_223;
  mux_226_nl <= MUX_s_1_2_2(and_1036_nl, mux_tmp_223, or_591_cse);
  and_tmp_160 <= or_569_cse AND or_573_cse AND or_578_cse AND or_584_cse AND mux_226_nl;
  and_1037_nl <= nand_281_cse AND and_tmp_160;
  mux_227_nl <= MUX_s_1_2_2(and_1037_nl, and_tmp_160, or_564_cse);
  and_dcpl_542 <= mux_227_nl AND and_dcpl_13 AND and_dcpl_9;
  and_tmp_170 <= ((NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10"))) AND ((NOT main_stage_0_8)
      OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_9)
      OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_10)
      OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("01"))) AND or_569_cse
      AND or_573_cse AND or_578_cse AND or_584_cse AND ((NOT main_stage_0_7) OR (NOT
      asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("01")))
      AND ((NOT main_stage_0_11) OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("01"))) AND (CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT ccs_ccore_start_rsci_idat));
  and_dcpl_546 <= and_dcpl_460 AND and_dcpl_430;
  or_tmp_629 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("11")) OR (rem_12cyc_3_2(1))
      OR not_tmp_332;
  or_643_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (acc_tmp(1));
  and_1169_nl <= nand_281_cse AND or_tmp_629;
  mux_228_nl <= MUX_s_1_2_2(and_1169_nl, or_tmp_629, or_643_cse);
  and_dcpl_548 <= mux_228_nl AND and_dcpl_358 AND and_dcpl_521;
  or_648_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("01"));
  and_1030_nl <= nand_276_cse AND or_tmp_629;
  mux_tmp_227 <= MUX_s_1_2_2(and_1030_nl, or_tmp_629, or_648_cse);
  and_1031_nl <= nand_281_cse AND mux_tmp_227;
  mux_230_nl <= MUX_s_1_2_2(and_1031_nl, mux_tmp_227, or_643_cse);
  and_dcpl_550 <= mux_230_nl AND and_dcpl_362 AND and_dcpl_524;
  or_653_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR (rem_12cyc_st_3_3_2(1));
  and_1027_nl <= nand_198_cse AND or_tmp_629;
  mux_tmp_229 <= MUX_s_1_2_2(and_1027_nl, or_tmp_629, or_653_cse);
  and_1028_nl <= nand_276_cse AND mux_tmp_229;
  mux_tmp_230 <= MUX_s_1_2_2(and_1028_nl, mux_tmp_229, or_648_cse);
  and_1029_nl <= nand_281_cse AND mux_tmp_230;
  mux_233_nl <= MUX_s_1_2_2(and_1029_nl, mux_tmp_230, or_643_cse);
  and_dcpl_552 <= mux_233_nl AND and_dcpl_366 AND and_dcpl_527;
  or_660_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("01"));
  and_1023_nl <= nand_271_cse AND or_tmp_629;
  mux_tmp_232 <= MUX_s_1_2_2(and_1023_nl, or_tmp_629, or_660_cse);
  and_1024_nl <= nand_198_cse AND mux_tmp_232;
  mux_tmp_233 <= MUX_s_1_2_2(and_1024_nl, mux_tmp_232, or_653_cse);
  and_1025_nl <= nand_276_cse AND mux_tmp_233;
  mux_tmp_234 <= MUX_s_1_2_2(and_1025_nl, mux_tmp_233, or_648_cse);
  and_1026_nl <= nand_281_cse AND mux_tmp_234;
  mux_237_nl <= MUX_s_1_2_2(and_1026_nl, mux_tmp_234, or_643_cse);
  and_dcpl_554 <= mux_237_nl AND and_dcpl_370 AND and_dcpl_530;
  or_669_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR (rem_12cyc_st_5_3_2(1));
  and_1018_nl <= nand_189_cse AND or_tmp_629;
  mux_tmp_236 <= MUX_s_1_2_2(and_1018_nl, or_tmp_629, or_669_cse);
  and_1019_nl <= nand_271_cse AND mux_tmp_236;
  mux_tmp_237 <= MUX_s_1_2_2(and_1019_nl, mux_tmp_236, or_660_cse);
  and_1020_nl <= nand_198_cse AND mux_tmp_237;
  mux_tmp_238 <= MUX_s_1_2_2(and_1020_nl, mux_tmp_237, or_653_cse);
  and_1021_nl <= nand_276_cse AND mux_tmp_238;
  mux_tmp_239 <= MUX_s_1_2_2(and_1021_nl, mux_tmp_238, or_648_cse);
  and_1022_nl <= nand_281_cse AND mux_tmp_239;
  mux_242_nl <= MUX_s_1_2_2(and_1022_nl, mux_tmp_239, or_643_cse);
  and_dcpl_556 <= mux_242_nl AND and_dcpl_121 AND and_dcpl_119;
  or_680_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("11")) OR (rem_12cyc_st_6_3_2(1));
  and_1012_nl <= nand_215_cse AND or_tmp_629;
  mux_tmp_241 <= MUX_s_1_2_2(and_1012_nl, or_tmp_629, or_680_cse);
  and_1013_nl <= nand_189_cse AND mux_tmp_241;
  mux_tmp_242 <= MUX_s_1_2_2(and_1013_nl, mux_tmp_241, or_669_cse);
  and_1014_nl <= nand_271_cse AND mux_tmp_242;
  mux_tmp_243 <= MUX_s_1_2_2(and_1014_nl, mux_tmp_242, or_660_cse);
  and_1015_nl <= nand_198_cse AND mux_tmp_243;
  mux_tmp_244 <= MUX_s_1_2_2(and_1015_nl, mux_tmp_243, or_653_cse);
  and_1016_nl <= nand_276_cse AND mux_tmp_244;
  mux_tmp_245 <= MUX_s_1_2_2(and_1016_nl, mux_tmp_244, or_648_cse);
  and_1017_nl <= nand_281_cse AND mux_tmp_245;
  mux_248_nl <= MUX_s_1_2_2(and_1017_nl, mux_tmp_245, or_643_cse);
  and_dcpl_558 <= mux_248_nl AND and_dcpl_94 AND and_dcpl_92;
  or_693_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("11")) OR (rem_12cyc_st_7_3_2(1));
  and_1005_nl <= nand_212_cse AND or_tmp_629;
  mux_tmp_247 <= MUX_s_1_2_2(and_1005_nl, or_tmp_629, or_693_cse);
  and_1006_nl <= nand_215_cse AND mux_tmp_247;
  mux_tmp_248 <= MUX_s_1_2_2(and_1006_nl, mux_tmp_247, or_680_cse);
  and_1007_nl <= nand_189_cse AND mux_tmp_248;
  mux_tmp_249 <= MUX_s_1_2_2(and_1007_nl, mux_tmp_248, or_669_cse);
  and_1008_nl <= nand_271_cse AND mux_tmp_249;
  mux_tmp_250 <= MUX_s_1_2_2(and_1008_nl, mux_tmp_249, or_660_cse);
  and_1009_nl <= nand_198_cse AND mux_tmp_250;
  mux_tmp_251 <= MUX_s_1_2_2(and_1009_nl, mux_tmp_250, or_653_cse);
  and_1010_nl <= nand_276_cse AND mux_tmp_251;
  mux_tmp_252 <= MUX_s_1_2_2(and_1010_nl, mux_tmp_251, or_648_cse);
  and_1011_nl <= nand_281_cse AND mux_tmp_252;
  mux_255_nl <= MUX_s_1_2_2(and_1011_nl, mux_tmp_252, or_643_cse);
  and_dcpl_560 <= mux_255_nl AND and_dcpl_67 AND and_dcpl_65;
  or_708_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("11")) OR (rem_12cyc_st_8_3_2(1));
  and_997_nl <= nand_208_cse AND or_tmp_629;
  mux_tmp_254 <= MUX_s_1_2_2(and_997_nl, or_tmp_629, or_708_cse);
  and_998_nl <= nand_212_cse AND mux_tmp_254;
  mux_tmp_255 <= MUX_s_1_2_2(and_998_nl, mux_tmp_254, or_693_cse);
  and_999_nl <= nand_215_cse AND mux_tmp_255;
  mux_tmp_256 <= MUX_s_1_2_2(and_999_nl, mux_tmp_255, or_680_cse);
  and_1000_nl <= nand_189_cse AND mux_tmp_256;
  mux_tmp_257 <= MUX_s_1_2_2(and_1000_nl, mux_tmp_256, or_669_cse);
  and_1001_nl <= nand_271_cse AND mux_tmp_257;
  mux_tmp_258 <= MUX_s_1_2_2(and_1001_nl, mux_tmp_257, or_660_cse);
  and_1002_nl <= nand_198_cse AND mux_tmp_258;
  mux_tmp_259 <= MUX_s_1_2_2(and_1002_nl, mux_tmp_258, or_653_cse);
  and_1003_nl <= nand_276_cse AND mux_tmp_259;
  mux_tmp_260 <= MUX_s_1_2_2(and_1003_nl, mux_tmp_259, or_648_cse);
  and_1004_nl <= nand_281_cse AND mux_tmp_260;
  mux_263_nl <= MUX_s_1_2_2(and_1004_nl, mux_tmp_260, or_643_cse);
  and_dcpl_562 <= mux_263_nl AND and_dcpl_40 AND and_dcpl_38;
  and_988_nl <= nand_203_cse AND or_tmp_629;
  or_725_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("11")) OR (rem_12cyc_st_9_3_2(1));
  mux_tmp_262 <= MUX_s_1_2_2(and_988_nl, or_tmp_629, or_725_nl);
  and_989_nl <= nand_208_cse AND mux_tmp_262;
  mux_tmp_263 <= MUX_s_1_2_2(and_989_nl, mux_tmp_262, or_708_cse);
  and_990_nl <= nand_212_cse AND mux_tmp_263;
  mux_tmp_264 <= MUX_s_1_2_2(and_990_nl, mux_tmp_263, or_693_cse);
  and_991_nl <= nand_215_cse AND mux_tmp_264;
  mux_tmp_265 <= MUX_s_1_2_2(and_991_nl, mux_tmp_264, or_680_cse);
  and_992_nl <= nand_189_cse AND mux_tmp_265;
  mux_tmp_266 <= MUX_s_1_2_2(and_992_nl, mux_tmp_265, or_669_cse);
  and_993_nl <= nand_271_cse AND mux_tmp_266;
  mux_tmp_267 <= MUX_s_1_2_2(and_993_nl, mux_tmp_266, or_660_cse);
  and_994_nl <= nand_198_cse AND mux_tmp_267;
  mux_tmp_268 <= MUX_s_1_2_2(and_994_nl, mux_tmp_267, or_653_cse);
  and_995_nl <= nand_276_cse AND mux_tmp_268;
  mux_tmp_269 <= MUX_s_1_2_2(and_995_nl, mux_tmp_268, or_648_cse);
  and_996_nl <= nand_281_cse AND mux_tmp_269;
  mux_272_nl <= MUX_s_1_2_2(and_996_nl, mux_tmp_269, or_643_cse);
  and_dcpl_564 <= mux_272_nl AND and_dcpl_13 AND and_dcpl_11;
  and_tmp_179 <= (NOT(main_stage_0_8 AND asn_itm_7 AND CONV_SL_1_1(rem_12cyc_st_7_1_0=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(rem_12cyc_st_7_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_9
      AND asn_itm_8 AND CONV_SL_1_1(rem_12cyc_st_8_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_8_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_10
      AND asn_itm_9 AND CONV_SL_1_1(rem_12cyc_st_9_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_9_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_3
      AND asn_itm_2 AND CONV_SL_1_1(rem_12cyc_st_2_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_2_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_4
      AND asn_itm_3 AND CONV_SL_1_1(rem_12cyc_st_3_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_3_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_5
      AND asn_itm_4 AND CONV_SL_1_1(rem_12cyc_st_4_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_4_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_6
      AND asn_itm_5 AND CONV_SL_1_1(rem_12cyc_st_5_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_5_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_7
      AND asn_itm_6 AND CONV_SL_1_1(rem_12cyc_st_6_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_6_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_11
      AND asn_itm_10 AND CONV_SL_1_1(rem_12cyc_st_10_1_0=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(rem_12cyc_st_10_3_2=STD_LOGIC_VECTOR'("01")))) AND ((acc_tmp(1))
      OR (NOT((acc_tmp(0)) AND CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND ccs_ccore_start_rsci_idat)));
  and_987_nl <= (NOT((rem_12cyc_3_2(0)) AND CONV_SL_1_1(rem_12cyc_1_0=STD_LOGIC_VECTOR'("11"))))
      AND and_tmp_179;
  or_735_nl <= (NOT main_stage_0_2) OR (NOT asn_itm_1) OR (rem_12cyc_3_2(1));
  mux_tmp_271 <= MUX_s_1_2_2(and_987_nl, and_tmp_179, or_735_nl);
  and_dcpl_568 <= and_dcpl_292 AND (acc_tmp(1));
  and_dcpl_569 <= and_dcpl_568 AND and_dcpl_291;
  and_dcpl_570 <= CONV_SL_1_1(rem_12cyc_st_2_3_2=STD_LOGIC_VECTOR'("10"));
  and_dcpl_571 <= and_dcpl_570 AND (NOT (rem_12cyc_st_2_1_0(1)));
  or_tmp_733 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR not_tmp_54;
  or_748_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("10"));
  nor_436_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_733));
  mux_274_nl <= MUX_s_1_2_2(nor_436_nl, or_tmp_733, or_748_cse);
  and_dcpl_573 <= mux_274_nl AND and_dcpl_298 AND and_dcpl_571;
  and_dcpl_574 <= CONV_SL_1_1(rem_12cyc_st_3_3_2=STD_LOGIC_VECTOR'("10"));
  and_dcpl_575 <= and_dcpl_574 AND (NOT (rem_12cyc_st_3_1_0(1)));
  or_753_cse <= (rem_12cyc_st_2_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp_180 <= or_753_cse AND or_tmp_733;
  nor_435_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_180));
  mux_275_nl <= MUX_s_1_2_2(nor_435_nl, and_tmp_180, or_748_cse);
  and_dcpl_577 <= mux_275_nl AND and_dcpl_304 AND and_dcpl_575;
  and_dcpl_578 <= CONV_SL_1_1(rem_12cyc_st_4_3_2=STD_LOGIC_VECTOR'("10"));
  and_dcpl_579 <= and_dcpl_578 AND (NOT (rem_12cyc_st_4_1_0(1)));
  or_757_cse <= (rem_12cyc_st_3_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_182 <= or_753_cse AND or_757_cse AND or_tmp_733;
  nor_434_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_182));
  mux_276_nl <= MUX_s_1_2_2(nor_434_nl, and_tmp_182, or_748_cse);
  and_dcpl_581 <= mux_276_nl AND and_dcpl_310 AND and_dcpl_579;
  and_dcpl_582 <= CONV_SL_1_1(rem_12cyc_st_5_3_2=STD_LOGIC_VECTOR'("10"));
  and_dcpl_583 <= and_dcpl_582 AND (NOT (rem_12cyc_st_5_1_0(1)));
  or_762_cse <= (rem_12cyc_st_4_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_185 <= or_753_cse AND or_757_cse AND or_762_cse AND or_tmp_733;
  nor_433_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_185));
  mux_277_nl <= MUX_s_1_2_2(nor_433_nl, and_tmp_185, or_748_cse);
  and_dcpl_585 <= mux_277_nl AND and_dcpl_316 AND and_dcpl_583;
  or_768_cse <= (rem_12cyc_st_5_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_189 <= or_753_cse AND or_757_cse AND or_762_cse AND or_768_cse AND or_tmp_733;
  nor_432_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_189));
  mux_278_nl <= MUX_s_1_2_2(nor_432_nl, and_tmp_189, or_748_cse);
  and_dcpl_589 <= mux_278_nl AND and_dcpl_112 AND and_dcpl_126 AND (NOT (rem_12cyc_st_6_1_0(1)));
  or_775_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_430_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_733));
  mux_279_nl <= MUX_s_1_2_2(nor_430_nl, or_tmp_733, or_775_cse);
  and_tmp_193 <= or_753_cse AND or_757_cse AND or_762_cse AND or_768_cse AND mux_279_nl;
  nor_431_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_193));
  mux_280_nl <= MUX_s_1_2_2(nor_431_nl, and_tmp_193, or_748_cse);
  and_dcpl_593 <= mux_280_nl AND and_dcpl_85 AND and_dcpl_99 AND (NOT (rem_12cyc_st_7_1_0(0)));
  or_784_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_427_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_733));
  mux_tmp_279 <= MUX_s_1_2_2(nor_427_nl, or_tmp_733, or_784_cse);
  nor_428_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_279));
  mux_282_nl <= MUX_s_1_2_2(nor_428_nl, mux_tmp_279, or_775_cse);
  and_tmp_197 <= or_753_cse AND or_757_cse AND or_762_cse AND or_768_cse AND mux_282_nl;
  nor_429_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_197));
  mux_283_nl <= MUX_s_1_2_2(nor_429_nl, and_tmp_197, or_748_cse);
  and_dcpl_597 <= mux_283_nl AND and_dcpl_58 AND and_dcpl_72 AND (NOT (rem_12cyc_st_8_1_0(0)));
  or_795_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_423_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_733));
  mux_tmp_282 <= MUX_s_1_2_2(nor_423_nl, or_tmp_733, or_795_cse);
  nor_424_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_282));
  mux_tmp_283 <= MUX_s_1_2_2(nor_424_nl, mux_tmp_282, or_784_cse);
  nor_425_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_283));
  mux_286_nl <= MUX_s_1_2_2(nor_425_nl, mux_tmp_283, or_775_cse);
  and_tmp_201 <= or_753_cse AND or_757_cse AND or_762_cse AND or_768_cse AND mux_286_nl;
  nor_426_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_201));
  mux_287_nl <= MUX_s_1_2_2(nor_426_nl, and_tmp_201, or_748_cse);
  and_dcpl_601 <= mux_287_nl AND and_dcpl_31 AND and_dcpl_45 AND (NOT (rem_12cyc_st_9_1_0(0)));
  nor_418_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_733));
  or_808_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("10"));
  mux_tmp_286 <= MUX_s_1_2_2(nor_418_nl, or_tmp_733, or_808_nl);
  nor_419_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_286));
  mux_tmp_287 <= MUX_s_1_2_2(nor_419_nl, mux_tmp_286, or_795_cse);
  nor_420_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_287));
  mux_tmp_288 <= MUX_s_1_2_2(nor_420_nl, mux_tmp_287, or_784_cse);
  nor_421_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_288));
  mux_291_nl <= MUX_s_1_2_2(nor_421_nl, mux_tmp_288, or_775_cse);
  and_tmp_205 <= or_753_cse AND or_757_cse AND or_762_cse AND or_768_cse AND mux_291_nl;
  nor_422_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_205));
  mux_292_nl <= MUX_s_1_2_2(nor_422_nl, and_tmp_205, or_748_cse);
  and_dcpl_605 <= mux_292_nl AND and_dcpl_4 AND and_dcpl_18 AND (NOT (rem_12cyc_st_10_1_0(0)));
  or_tmp_808 <= CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(acc_1_tmp(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT ccs_ccore_start_rsci_idat);
  nor_409_nl <= NOT((rem_12cyc_st_10_3_2(1)) OR (NOT or_tmp_808));
  or_823_nl <= (NOT main_stage_0_11) OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_10_3_2(0));
  mux_tmp_291 <= MUX_s_1_2_2(nor_409_nl, or_tmp_808, or_823_nl);
  nor_410_nl <= NOT((rem_12cyc_st_6_3_2(1)) OR (NOT mux_tmp_291));
  or_822_nl <= (NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_6_3_2(0));
  mux_tmp_292 <= MUX_s_1_2_2(nor_410_nl, mux_tmp_291, or_822_nl);
  nor_411_nl <= NOT((rem_12cyc_st_5_3_2(1)) OR (NOT mux_tmp_292));
  or_821_nl <= (NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_5_3_2(0));
  mux_tmp_293 <= MUX_s_1_2_2(nor_411_nl, mux_tmp_292, or_821_nl);
  nor_412_nl <= NOT((rem_12cyc_st_4_3_2(1)) OR (NOT mux_tmp_293));
  or_820_nl <= (NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_4_3_2(0));
  mux_tmp_294 <= MUX_s_1_2_2(nor_412_nl, mux_tmp_293, or_820_nl);
  nor_413_nl <= NOT((rem_12cyc_st_3_3_2(1)) OR (NOT mux_tmp_294));
  or_819_nl <= (NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_3_3_2(0));
  mux_tmp_295 <= MUX_s_1_2_2(nor_413_nl, mux_tmp_294, or_819_nl);
  nor_414_nl <= NOT((rem_12cyc_st_2_3_2(1)) OR (NOT mux_tmp_295));
  or_818_nl <= (NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_2_3_2(0));
  mux_tmp_296 <= MUX_s_1_2_2(nor_414_nl, mux_tmp_295, or_818_nl);
  nor_415_nl <= NOT((rem_12cyc_st_9_3_2(1)) OR (NOT mux_tmp_296));
  or_817_nl <= (NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_9_3_2(0));
  mux_tmp_297 <= MUX_s_1_2_2(nor_415_nl, mux_tmp_296, or_817_nl);
  nor_416_nl <= NOT((rem_12cyc_st_8_3_2(1)) OR (NOT mux_tmp_297));
  or_816_nl <= (NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_8_3_2(0));
  mux_tmp_298 <= MUX_s_1_2_2(nor_416_nl, mux_tmp_297, or_816_nl);
  nor_417_nl <= NOT((rem_12cyc_st_7_3_2(1)) OR (NOT mux_tmp_298));
  or_815_nl <= (NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_7_3_2(0));
  mux_301_nl <= MUX_s_1_2_2(nor_417_nl, mux_tmp_298, or_815_nl);
  and_tmp_206 <= ((NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00"))) AND mux_301_nl;
  and_dcpl_610 <= and_dcpl_568 AND and_dcpl_355;
  or_tmp_820 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR not_tmp_54;
  or_837_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("10"));
  nor_408_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_820));
  mux_302_nl <= MUX_s_1_2_2(nor_408_nl, or_tmp_820, or_837_cse);
  and_dcpl_612 <= mux_302_nl AND and_dcpl_358 AND and_dcpl_571;
  nand_84_cse <= NOT((rem_12cyc_st_2_3_2(1)) AND asn_itm_2 AND main_stage_0_3 AND
      (rem_12cyc_st_2_1_0(0)));
  or_842_cse <= (rem_12cyc_st_2_1_0(1)) OR (rem_12cyc_st_2_3_2(0));
  and_986_nl <= nand_84_cse AND or_tmp_820;
  mux_tmp_301 <= MUX_s_1_2_2(and_986_nl, or_tmp_820, or_842_cse);
  nor_407_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_301));
  mux_304_nl <= MUX_s_1_2_2(nor_407_nl, mux_tmp_301, or_837_cse);
  and_dcpl_614 <= mux_304_nl AND and_dcpl_362 AND and_dcpl_575;
  or_847_cse <= (rem_12cyc_st_3_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("10"));
  and_984_nl <= nand_274_cse AND or_tmp_820;
  mux_tmp_303 <= MUX_s_1_2_2(and_984_nl, or_tmp_820, or_847_cse);
  and_985_nl <= nand_84_cse AND mux_tmp_303;
  mux_tmp_304 <= MUX_s_1_2_2(and_985_nl, mux_tmp_303, or_842_cse);
  nor_406_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_304));
  mux_307_nl <= MUX_s_1_2_2(nor_406_nl, mux_tmp_304, or_837_cse);
  and_dcpl_616 <= mux_307_nl AND and_dcpl_366 AND and_dcpl_579;
  nand_79_cse <= NOT((rem_12cyc_st_4_3_2(1)) AND asn_itm_4 AND main_stage_0_5 AND
      (rem_12cyc_st_4_1_0(0)));
  or_854_cse <= (rem_12cyc_st_4_1_0(1)) OR (rem_12cyc_st_4_3_2(0));
  and_981_nl <= nand_79_cse AND or_tmp_820;
  mux_tmp_306 <= MUX_s_1_2_2(and_981_nl, or_tmp_820, or_854_cse);
  and_982_nl <= nand_274_cse AND mux_tmp_306;
  mux_tmp_307 <= MUX_s_1_2_2(and_982_nl, mux_tmp_306, or_847_cse);
  and_983_nl <= nand_84_cse AND mux_tmp_307;
  mux_tmp_308 <= MUX_s_1_2_2(and_983_nl, mux_tmp_307, or_842_cse);
  nor_405_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_308));
  mux_311_nl <= MUX_s_1_2_2(nor_405_nl, mux_tmp_308, or_837_cse);
  and_dcpl_618 <= mux_311_nl AND and_dcpl_370 AND and_dcpl_583;
  or_863_cse <= (rem_12cyc_st_5_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("10"));
  and_977_nl <= nand_267_cse AND or_tmp_820;
  mux_tmp_310 <= MUX_s_1_2_2(and_977_nl, or_tmp_820, or_863_cse);
  and_978_nl <= nand_79_cse AND mux_tmp_310;
  mux_tmp_311 <= MUX_s_1_2_2(and_978_nl, mux_tmp_310, or_854_cse);
  and_979_nl <= nand_274_cse AND mux_tmp_311;
  mux_tmp_312 <= MUX_s_1_2_2(and_979_nl, mux_tmp_311, or_847_cse);
  and_980_nl <= nand_84_cse AND mux_tmp_312;
  mux_tmp_313 <= MUX_s_1_2_2(and_980_nl, mux_tmp_312, or_842_cse);
  nor_404_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_313));
  mux_316_nl <= MUX_s_1_2_2(nor_404_nl, mux_tmp_313, or_837_cse);
  and_dcpl_622 <= mux_316_nl AND and_dcpl_112 AND and_dcpl_129 AND (NOT (rem_12cyc_st_6_1_0(1)));
  or_874_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_402_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_820));
  mux_tmp_315 <= MUX_s_1_2_2(nor_402_nl, or_tmp_820, or_874_cse);
  and_973_nl <= nand_267_cse AND mux_tmp_315;
  mux_tmp_316 <= MUX_s_1_2_2(and_973_nl, mux_tmp_315, or_863_cse);
  and_974_nl <= nand_79_cse AND mux_tmp_316;
  mux_tmp_317 <= MUX_s_1_2_2(and_974_nl, mux_tmp_316, or_854_cse);
  and_975_nl <= nand_274_cse AND mux_tmp_317;
  mux_tmp_318 <= MUX_s_1_2_2(and_975_nl, mux_tmp_317, or_847_cse);
  and_976_nl <= nand_84_cse AND mux_tmp_318;
  mux_tmp_319 <= MUX_s_1_2_2(and_976_nl, mux_tmp_318, or_842_cse);
  nor_403_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_319));
  mux_322_nl <= MUX_s_1_2_2(nor_403_nl, mux_tmp_319, or_837_cse);
  and_dcpl_625 <= mux_322_nl AND and_dcpl_85 AND and_dcpl_99 AND (rem_12cyc_st_7_1_0(0));
  or_887_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_399_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_820));
  mux_tmp_321 <= MUX_s_1_2_2(nor_399_nl, or_tmp_820, or_887_cse);
  nor_400_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_321));
  mux_tmp_322 <= MUX_s_1_2_2(nor_400_nl, mux_tmp_321, or_874_cse);
  and_969_nl <= nand_267_cse AND mux_tmp_322;
  mux_tmp_323 <= MUX_s_1_2_2(and_969_nl, mux_tmp_322, or_863_cse);
  and_970_nl <= nand_79_cse AND mux_tmp_323;
  mux_tmp_324 <= MUX_s_1_2_2(and_970_nl, mux_tmp_323, or_854_cse);
  and_971_nl <= nand_274_cse AND mux_tmp_324;
  mux_tmp_325 <= MUX_s_1_2_2(and_971_nl, mux_tmp_324, or_847_cse);
  and_972_nl <= nand_84_cse AND mux_tmp_325;
  mux_tmp_326 <= MUX_s_1_2_2(and_972_nl, mux_tmp_325, or_842_cse);
  nor_401_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_326));
  mux_329_nl <= MUX_s_1_2_2(nor_401_nl, mux_tmp_326, or_837_cse);
  and_dcpl_628 <= mux_329_nl AND and_dcpl_58 AND and_dcpl_72 AND (rem_12cyc_st_8_1_0(0));
  or_902_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_395_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_820));
  mux_tmp_328 <= MUX_s_1_2_2(nor_395_nl, or_tmp_820, or_902_cse);
  nor_396_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_328));
  mux_tmp_329 <= MUX_s_1_2_2(nor_396_nl, mux_tmp_328, or_887_cse);
  nor_397_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_329));
  mux_tmp_330 <= MUX_s_1_2_2(nor_397_nl, mux_tmp_329, or_874_cse);
  and_965_nl <= nand_267_cse AND mux_tmp_330;
  mux_tmp_331 <= MUX_s_1_2_2(and_965_nl, mux_tmp_330, or_863_cse);
  and_966_nl <= nand_79_cse AND mux_tmp_331;
  mux_tmp_332 <= MUX_s_1_2_2(and_966_nl, mux_tmp_331, or_854_cse);
  and_967_nl <= nand_274_cse AND mux_tmp_332;
  mux_tmp_333 <= MUX_s_1_2_2(and_967_nl, mux_tmp_332, or_847_cse);
  and_968_nl <= nand_84_cse AND mux_tmp_333;
  mux_tmp_334 <= MUX_s_1_2_2(and_968_nl, mux_tmp_333, or_842_cse);
  nor_398_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_334));
  mux_337_nl <= MUX_s_1_2_2(nor_398_nl, mux_tmp_334, or_837_cse);
  and_dcpl_631 <= mux_337_nl AND and_dcpl_31 AND and_dcpl_45 AND (rem_12cyc_st_9_1_0(0));
  nor_390_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_820));
  or_919_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("10"));
  mux_tmp_336 <= MUX_s_1_2_2(nor_390_nl, or_tmp_820, or_919_nl);
  nor_391_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_336));
  mux_tmp_337 <= MUX_s_1_2_2(nor_391_nl, mux_tmp_336, or_902_cse);
  nor_392_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_337));
  mux_tmp_338 <= MUX_s_1_2_2(nor_392_nl, mux_tmp_337, or_887_cse);
  nor_393_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_338));
  mux_tmp_339 <= MUX_s_1_2_2(nor_393_nl, mux_tmp_338, or_874_cse);
  and_961_nl <= nand_267_cse AND mux_tmp_339;
  mux_tmp_340 <= MUX_s_1_2_2(and_961_nl, mux_tmp_339, or_863_cse);
  and_962_nl <= nand_79_cse AND mux_tmp_340;
  mux_tmp_341 <= MUX_s_1_2_2(and_962_nl, mux_tmp_340, or_854_cse);
  and_963_nl <= nand_274_cse AND mux_tmp_341;
  mux_tmp_342 <= MUX_s_1_2_2(and_963_nl, mux_tmp_341, or_847_cse);
  and_964_nl <= nand_84_cse AND mux_tmp_342;
  mux_tmp_343 <= MUX_s_1_2_2(and_964_nl, mux_tmp_342, or_842_cse);
  nor_394_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_343));
  mux_346_nl <= MUX_s_1_2_2(nor_394_nl, mux_tmp_343, or_837_cse);
  and_dcpl_634 <= mux_346_nl AND and_dcpl_4 AND and_dcpl_18 AND (rem_12cyc_st_10_1_0(0));
  or_tmp_921 <= CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("10")) OR (acc_1_tmp(1)) OR
      nand_250_cse;
  nor_380_nl <= NOT((rem_12cyc_st_10_3_2(1)) OR (NOT or_tmp_921));
  or_938_nl <= (NOT main_stage_0_11) OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_10_3_2(0));
  mux_tmp_345 <= MUX_s_1_2_2(nor_380_nl, or_tmp_921, or_938_nl);
  nor_381_nl <= NOT((rem_12cyc_st_6_3_2(1)) OR (NOT mux_tmp_345));
  or_937_nl <= (NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_6_3_2(0));
  mux_tmp_346 <= MUX_s_1_2_2(nor_381_nl, mux_tmp_345, or_937_nl);
  nor_382_nl <= NOT((rem_12cyc_st_5_3_2(1)) OR (NOT mux_tmp_346));
  or_936_nl <= (NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_5_3_2(0));
  mux_tmp_347 <= MUX_s_1_2_2(nor_382_nl, mux_tmp_346, or_936_nl);
  nor_383_nl <= NOT((rem_12cyc_st_4_3_2(1)) OR (NOT mux_tmp_347));
  or_935_nl <= (NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_4_3_2(0));
  mux_tmp_348 <= MUX_s_1_2_2(nor_383_nl, mux_tmp_347, or_935_nl);
  nor_384_nl <= NOT((rem_12cyc_st_3_3_2(1)) OR (NOT mux_tmp_348));
  or_934_nl <= (NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_3_3_2(0));
  mux_tmp_349 <= MUX_s_1_2_2(nor_384_nl, mux_tmp_348, or_934_nl);
  nor_385_nl <= NOT((rem_12cyc_st_2_3_2(1)) OR (NOT mux_tmp_349));
  or_933_nl <= (NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_2_3_2(0));
  mux_tmp_350 <= MUX_s_1_2_2(nor_385_nl, mux_tmp_349, or_933_nl);
  nor_386_nl <= NOT((rem_12cyc_st_9_3_2(1)) OR (NOT mux_tmp_350));
  or_932_nl <= (NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_9_3_2(0));
  mux_tmp_351 <= MUX_s_1_2_2(nor_386_nl, mux_tmp_350, or_932_nl);
  nor_387_nl <= NOT((rem_12cyc_st_8_3_2(1)) OR (NOT mux_tmp_351));
  or_931_nl <= (NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_8_3_2(0));
  mux_tmp_352 <= MUX_s_1_2_2(nor_387_nl, mux_tmp_351, or_931_nl);
  nor_388_nl <= NOT((rem_12cyc_st_7_3_2(1)) OR (NOT mux_tmp_352));
  or_930_nl <= (NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_7_3_2(0));
  mux_tmp_353 <= MUX_s_1_2_2(nor_388_nl, mux_tmp_352, or_930_nl);
  nor_389_nl <= NOT((rem_12cyc_1_0(0)) OR (NOT mux_tmp_353));
  or_929_nl <= (NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_1_0(1));
  mux_tmp_354 <= MUX_s_1_2_2(nor_389_nl, mux_tmp_353, or_929_nl);
  and_dcpl_638 <= and_dcpl_568 AND and_dcpl_393;
  and_dcpl_639 <= and_dcpl_570 AND (rem_12cyc_st_2_1_0(1));
  or_tmp_934 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR not_tmp_54;
  or_952_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("10"));
  nor_379_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_934));
  mux_357_nl <= MUX_s_1_2_2(nor_379_nl, or_tmp_934, or_952_cse);
  and_dcpl_641 <= mux_357_nl AND and_dcpl_298 AND and_dcpl_639;
  and_dcpl_642 <= and_dcpl_574 AND (rem_12cyc_st_3_1_0(1));
  or_957_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp_207 <= or_957_cse AND or_tmp_934;
  nor_378_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_207));
  mux_358_nl <= MUX_s_1_2_2(nor_378_nl, and_tmp_207, or_952_cse);
  and_dcpl_644 <= mux_358_nl AND and_dcpl_304 AND and_dcpl_642;
  and_dcpl_645 <= and_dcpl_578 AND (rem_12cyc_st_4_1_0(1));
  or_961_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_209 <= or_957_cse AND or_961_cse AND or_tmp_934;
  nor_377_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_209));
  mux_359_nl <= MUX_s_1_2_2(nor_377_nl, and_tmp_209, or_952_cse);
  and_dcpl_647 <= mux_359_nl AND and_dcpl_310 AND and_dcpl_645;
  and_dcpl_648 <= and_dcpl_582 AND (rem_12cyc_st_5_1_0(1));
  or_966_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_212 <= or_957_cse AND or_961_cse AND or_966_cse AND or_tmp_934;
  nor_376_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_212));
  mux_360_nl <= MUX_s_1_2_2(nor_376_nl, and_tmp_212, or_952_cse);
  and_dcpl_650 <= mux_360_nl AND and_dcpl_316 AND and_dcpl_648;
  or_972_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_216 <= or_957_cse AND or_961_cse AND or_966_cse AND or_972_cse AND or_tmp_934;
  nor_375_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_216));
  mux_361_nl <= MUX_s_1_2_2(nor_375_nl, and_tmp_216, or_952_cse);
  and_dcpl_653 <= mux_361_nl AND and_dcpl_112 AND and_dcpl_126 AND (rem_12cyc_st_6_1_0(1));
  or_979_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_373_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_934));
  mux_362_nl <= MUX_s_1_2_2(nor_373_nl, or_tmp_934, or_979_cse);
  and_tmp_220 <= or_957_cse AND or_961_cse AND or_966_cse AND or_972_cse AND mux_362_nl;
  nor_374_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_220));
  mux_363_nl <= MUX_s_1_2_2(nor_374_nl, and_tmp_220, or_952_cse);
  and_dcpl_657 <= mux_363_nl AND and_dcpl_85 AND and_dcpl_104 AND (NOT (rem_12cyc_st_7_1_0(0)));
  or_988_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_370_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_934));
  mux_tmp_362 <= MUX_s_1_2_2(nor_370_nl, or_tmp_934, or_988_cse);
  nor_371_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_362));
  mux_365_nl <= MUX_s_1_2_2(nor_371_nl, mux_tmp_362, or_979_cse);
  and_tmp_224 <= or_957_cse AND or_961_cse AND or_966_cse AND or_972_cse AND mux_365_nl;
  nor_372_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_224));
  mux_366_nl <= MUX_s_1_2_2(nor_372_nl, and_tmp_224, or_952_cse);
  and_dcpl_661 <= mux_366_nl AND and_dcpl_58 AND and_dcpl_77 AND (NOT (rem_12cyc_st_8_1_0(0)));
  or_999_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_366_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_934));
  mux_tmp_365 <= MUX_s_1_2_2(nor_366_nl, or_tmp_934, or_999_cse);
  nor_367_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_365));
  mux_tmp_366 <= MUX_s_1_2_2(nor_367_nl, mux_tmp_365, or_988_cse);
  nor_368_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_366));
  mux_369_nl <= MUX_s_1_2_2(nor_368_nl, mux_tmp_366, or_979_cse);
  and_tmp_228 <= or_957_cse AND or_961_cse AND or_966_cse AND or_972_cse AND mux_369_nl;
  nor_369_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_228));
  mux_370_nl <= MUX_s_1_2_2(nor_369_nl, and_tmp_228, or_952_cse);
  and_dcpl_665 <= mux_370_nl AND and_dcpl_31 AND and_dcpl_50 AND (NOT (rem_12cyc_st_9_1_0(0)));
  nor_361_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_934));
  or_1012_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("10"));
  mux_tmp_369 <= MUX_s_1_2_2(nor_361_nl, or_tmp_934, or_1012_nl);
  nor_362_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_369));
  mux_tmp_370 <= MUX_s_1_2_2(nor_362_nl, mux_tmp_369, or_999_cse);
  nor_363_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_370));
  mux_tmp_371 <= MUX_s_1_2_2(nor_363_nl, mux_tmp_370, or_988_cse);
  nor_364_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_371));
  mux_374_nl <= MUX_s_1_2_2(nor_364_nl, mux_tmp_371, or_979_cse);
  and_tmp_232 <= or_957_cse AND or_961_cse AND or_966_cse AND or_972_cse AND mux_374_nl;
  nor_365_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_232));
  mux_375_nl <= MUX_s_1_2_2(nor_365_nl, and_tmp_232, or_952_cse);
  and_dcpl_669 <= mux_375_nl AND and_dcpl_4 AND and_dcpl_23 AND (NOT (rem_12cyc_st_10_1_0(0)));
  or_tmp_1009 <= CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(acc_1_tmp(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT ccs_ccore_start_rsci_idat);
  nor_352_nl <= NOT((rem_12cyc_st_10_3_2(1)) OR (NOT or_tmp_1009));
  or_1027_nl <= (NOT main_stage_0_11) OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_10_3_2(0));
  mux_tmp_374 <= MUX_s_1_2_2(nor_352_nl, or_tmp_1009, or_1027_nl);
  nor_353_nl <= NOT((rem_12cyc_st_6_3_2(1)) OR (NOT mux_tmp_374));
  or_1026_nl <= (NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_6_3_2(0));
  mux_tmp_375 <= MUX_s_1_2_2(nor_353_nl, mux_tmp_374, or_1026_nl);
  nor_354_nl <= NOT((rem_12cyc_st_5_3_2(1)) OR (NOT mux_tmp_375));
  or_1025_nl <= (NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_5_3_2(0));
  mux_tmp_376 <= MUX_s_1_2_2(nor_354_nl, mux_tmp_375, or_1025_nl);
  nor_355_nl <= NOT((rem_12cyc_st_4_3_2(1)) OR (NOT mux_tmp_376));
  or_1024_nl <= (NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_4_3_2(0));
  mux_tmp_377 <= MUX_s_1_2_2(nor_355_nl, mux_tmp_376, or_1024_nl);
  nor_356_nl <= NOT((rem_12cyc_st_3_3_2(1)) OR (NOT mux_tmp_377));
  or_1023_nl <= (NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_3_3_2(0));
  mux_tmp_378 <= MUX_s_1_2_2(nor_356_nl, mux_tmp_377, or_1023_nl);
  nor_357_nl <= NOT((rem_12cyc_st_2_3_2(1)) OR (NOT mux_tmp_378));
  or_1022_nl <= (NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_2_3_2(0));
  mux_tmp_379 <= MUX_s_1_2_2(nor_357_nl, mux_tmp_378, or_1022_nl);
  nor_358_nl <= NOT((rem_12cyc_st_9_3_2(1)) OR (NOT mux_tmp_379));
  or_1021_nl <= (NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_9_3_2(0));
  mux_tmp_380 <= MUX_s_1_2_2(nor_358_nl, mux_tmp_379, or_1021_nl);
  nor_359_nl <= NOT((rem_12cyc_st_8_3_2(1)) OR (NOT mux_tmp_380));
  or_1020_nl <= (NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_8_3_2(0));
  mux_tmp_381 <= MUX_s_1_2_2(nor_359_nl, mux_tmp_380, or_1020_nl);
  nor_360_nl <= NOT((rem_12cyc_st_7_3_2(1)) OR (NOT mux_tmp_381));
  or_1019_nl <= (NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_7_3_2(0));
  mux_384_nl <= MUX_s_1_2_2(nor_360_nl, mux_tmp_381, or_1019_nl);
  and_tmp_233 <= ((NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10"))) AND mux_384_nl;
  and_dcpl_673 <= and_dcpl_568 AND and_dcpl_430;
  or_tmp_1021 <= (NOT(CONV_SL_1_1(rem_12cyc_1_0=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(rem_12cyc_3_2=STD_LOGIC_VECTOR'("10"))))
      OR not_tmp_54;
  nand_57_cse <= NOT(CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(acc_tmp=STD_LOGIC_VECTOR'("10")));
  nor_351_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_1021));
  mux_385_nl <= MUX_s_1_2_2(nor_351_nl, or_tmp_1021, nand_57_cse);
  and_dcpl_675 <= mux_385_nl AND and_dcpl_358 AND and_dcpl_639;
  or_1045_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR (rem_12cyc_st_2_3_2(0));
  and_960_nl <= nand_84_cse AND or_tmp_1021;
  mux_tmp_384 <= MUX_s_1_2_2(and_960_nl, or_tmp_1021, or_1045_cse);
  nor_350_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_384));
  mux_387_nl <= MUX_s_1_2_2(nor_350_nl, mux_tmp_384, nand_57_cse);
  and_dcpl_677 <= mux_387_nl AND and_dcpl_362 AND and_dcpl_642;
  or_1050_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("10"));
  and_958_nl <= nand_274_cse AND or_tmp_1021;
  mux_tmp_386 <= MUX_s_1_2_2(and_958_nl, or_tmp_1021, or_1050_cse);
  and_959_nl <= nand_84_cse AND mux_tmp_386;
  mux_tmp_387 <= MUX_s_1_2_2(and_959_nl, mux_tmp_386, or_1045_cse);
  nor_349_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_387));
  mux_390_nl <= MUX_s_1_2_2(nor_349_nl, mux_tmp_387, nand_57_cse);
  and_dcpl_679 <= mux_390_nl AND and_dcpl_366 AND and_dcpl_645;
  or_1057_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR (rem_12cyc_st_4_3_2(0));
  and_955_nl <= nand_79_cse AND or_tmp_1021;
  mux_tmp_389 <= MUX_s_1_2_2(and_955_nl, or_tmp_1021, or_1057_cse);
  and_956_nl <= nand_274_cse AND mux_tmp_389;
  mux_tmp_390 <= MUX_s_1_2_2(and_956_nl, mux_tmp_389, or_1050_cse);
  and_957_nl <= nand_84_cse AND mux_tmp_390;
  mux_tmp_391 <= MUX_s_1_2_2(and_957_nl, mux_tmp_390, or_1045_cse);
  nor_348_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_391));
  mux_394_nl <= MUX_s_1_2_2(nor_348_nl, mux_tmp_391, nand_57_cse);
  and_dcpl_681 <= mux_394_nl AND and_dcpl_370 AND and_dcpl_648;
  or_1066_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("10"));
  and_951_nl <= nand_267_cse AND or_tmp_1021;
  mux_tmp_393 <= MUX_s_1_2_2(and_951_nl, or_tmp_1021, or_1066_cse);
  and_952_nl <= nand_79_cse AND mux_tmp_393;
  mux_tmp_394 <= MUX_s_1_2_2(and_952_nl, mux_tmp_393, or_1057_cse);
  and_953_nl <= nand_274_cse AND mux_tmp_394;
  mux_tmp_395 <= MUX_s_1_2_2(and_953_nl, mux_tmp_394, or_1050_cse);
  and_954_nl <= nand_84_cse AND mux_tmp_395;
  mux_tmp_396 <= MUX_s_1_2_2(and_954_nl, mux_tmp_395, or_1045_cse);
  nor_347_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_396));
  mux_399_nl <= MUX_s_1_2_2(nor_347_nl, mux_tmp_396, nand_57_cse);
  and_dcpl_684 <= mux_399_nl AND and_dcpl_112 AND and_dcpl_129 AND (rem_12cyc_st_6_1_0(1));
  nand_36_cse <= NOT(CONV_SL_1_1(rem_12cyc_st_6_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_6_3_2=STD_LOGIC_VECTOR'("10")));
  nor_345_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_1021));
  mux_tmp_398 <= MUX_s_1_2_2(nor_345_nl, or_tmp_1021, nand_36_cse);
  and_947_nl <= nand_267_cse AND mux_tmp_398;
  mux_tmp_399 <= MUX_s_1_2_2(and_947_nl, mux_tmp_398, or_1066_cse);
  and_948_nl <= nand_79_cse AND mux_tmp_399;
  mux_tmp_400 <= MUX_s_1_2_2(and_948_nl, mux_tmp_399, or_1057_cse);
  and_949_nl <= nand_274_cse AND mux_tmp_400;
  mux_tmp_401 <= MUX_s_1_2_2(and_949_nl, mux_tmp_400, or_1050_cse);
  and_950_nl <= nand_84_cse AND mux_tmp_401;
  mux_tmp_402 <= MUX_s_1_2_2(and_950_nl, mux_tmp_401, or_1045_cse);
  nor_346_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_402));
  mux_405_nl <= MUX_s_1_2_2(nor_346_nl, mux_tmp_402, nand_57_cse);
  and_dcpl_687 <= mux_405_nl AND and_dcpl_85 AND and_dcpl_104 AND (rem_12cyc_st_7_1_0(0));
  nand_29_cse <= NOT(CONV_SL_1_1(rem_12cyc_st_7_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_7_3_2=STD_LOGIC_VECTOR'("10")));
  nor_342_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_1021));
  mux_tmp_404 <= MUX_s_1_2_2(nor_342_nl, or_tmp_1021, nand_29_cse);
  nor_343_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_404));
  mux_tmp_405 <= MUX_s_1_2_2(nor_343_nl, mux_tmp_404, nand_36_cse);
  and_943_nl <= nand_267_cse AND mux_tmp_405;
  mux_tmp_406 <= MUX_s_1_2_2(and_943_nl, mux_tmp_405, or_1066_cse);
  and_944_nl <= nand_79_cse AND mux_tmp_406;
  mux_tmp_407 <= MUX_s_1_2_2(and_944_nl, mux_tmp_406, or_1057_cse);
  and_945_nl <= nand_274_cse AND mux_tmp_407;
  mux_tmp_408 <= MUX_s_1_2_2(and_945_nl, mux_tmp_407, or_1050_cse);
  and_946_nl <= nand_84_cse AND mux_tmp_408;
  mux_tmp_409 <= MUX_s_1_2_2(and_946_nl, mux_tmp_408, or_1045_cse);
  nor_344_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_409));
  mux_412_nl <= MUX_s_1_2_2(nor_344_nl, mux_tmp_409, nand_57_cse);
  and_dcpl_690 <= mux_412_nl AND and_dcpl_58 AND and_dcpl_77 AND (rem_12cyc_st_8_1_0(0));
  nand_21_cse <= NOT(CONV_SL_1_1(rem_12cyc_st_8_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_8_3_2=STD_LOGIC_VECTOR'("10")));
  nor_338_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_1021));
  mux_tmp_411 <= MUX_s_1_2_2(nor_338_nl, or_tmp_1021, nand_21_cse);
  nor_339_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_411));
  mux_tmp_412 <= MUX_s_1_2_2(nor_339_nl, mux_tmp_411, nand_29_cse);
  nor_340_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_412));
  mux_tmp_413 <= MUX_s_1_2_2(nor_340_nl, mux_tmp_412, nand_36_cse);
  and_939_nl <= nand_267_cse AND mux_tmp_413;
  mux_tmp_414 <= MUX_s_1_2_2(and_939_nl, mux_tmp_413, or_1066_cse);
  and_940_nl <= nand_79_cse AND mux_tmp_414;
  mux_tmp_415 <= MUX_s_1_2_2(and_940_nl, mux_tmp_414, or_1057_cse);
  and_941_nl <= nand_274_cse AND mux_tmp_415;
  mux_tmp_416 <= MUX_s_1_2_2(and_941_nl, mux_tmp_415, or_1050_cse);
  and_942_nl <= nand_84_cse AND mux_tmp_416;
  mux_tmp_417 <= MUX_s_1_2_2(and_942_nl, mux_tmp_416, or_1045_cse);
  nor_341_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_417));
  mux_420_nl <= MUX_s_1_2_2(nor_341_nl, mux_tmp_417, nand_57_cse);
  and_dcpl_693 <= mux_420_nl AND and_dcpl_31 AND and_dcpl_50 AND (rem_12cyc_st_9_1_0(0));
  nor_333_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_1021));
  nand_12_nl <= NOT(CONV_SL_1_1(rem_12cyc_st_9_1_0=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(rem_12cyc_st_9_3_2=STD_LOGIC_VECTOR'("10")));
  mux_tmp_419 <= MUX_s_1_2_2(nor_333_nl, or_tmp_1021, nand_12_nl);
  nor_334_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_419));
  mux_tmp_420 <= MUX_s_1_2_2(nor_334_nl, mux_tmp_419, nand_21_cse);
  nor_335_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_420));
  mux_tmp_421 <= MUX_s_1_2_2(nor_335_nl, mux_tmp_420, nand_29_cse);
  nor_336_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_421));
  mux_tmp_422 <= MUX_s_1_2_2(nor_336_nl, mux_tmp_421, nand_36_cse);
  and_935_nl <= nand_267_cse AND mux_tmp_422;
  mux_tmp_423 <= MUX_s_1_2_2(and_935_nl, mux_tmp_422, or_1066_cse);
  and_936_nl <= nand_79_cse AND mux_tmp_423;
  mux_tmp_424 <= MUX_s_1_2_2(and_936_nl, mux_tmp_423, or_1057_cse);
  and_937_nl <= nand_274_cse AND mux_tmp_424;
  mux_tmp_425 <= MUX_s_1_2_2(and_937_nl, mux_tmp_424, or_1050_cse);
  and_938_nl <= nand_84_cse AND mux_tmp_425;
  mux_tmp_426 <= MUX_s_1_2_2(and_938_nl, mux_tmp_425, or_1045_cse);
  nor_337_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_426));
  mux_429_nl <= MUX_s_1_2_2(nor_337_nl, mux_tmp_426, nand_57_cse);
  and_dcpl_696 <= mux_429_nl AND and_dcpl_4 AND and_dcpl_23 AND (rem_12cyc_st_10_1_0(0));
  or_tmp_1122 <= CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("10")) OR nand_222_cse;
  nor_324_nl <= NOT((rem_12cyc_st_10_3_2(1)) OR (NOT or_tmp_1122));
  nand_1_nl <= NOT(main_stage_0_11 AND asn_itm_10 AND CONV_SL_1_1(rem_12cyc_st_10_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_10_3_2(0))));
  mux_tmp_428 <= MUX_s_1_2_2(nor_324_nl, or_tmp_1122, nand_1_nl);
  nor_325_nl <= NOT((rem_12cyc_st_6_3_2(1)) OR (NOT mux_tmp_428));
  nand_2_nl <= NOT(main_stage_0_7 AND asn_itm_6 AND CONV_SL_1_1(rem_12cyc_st_6_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_6_3_2(0))));
  mux_tmp_429 <= MUX_s_1_2_2(nor_325_nl, mux_tmp_428, nand_2_nl);
  nor_326_nl <= NOT((rem_12cyc_st_5_3_2(1)) OR (NOT mux_tmp_429));
  nand_3_nl <= NOT(main_stage_0_6 AND asn_itm_5 AND CONV_SL_1_1(rem_12cyc_st_5_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_5_3_2(0))));
  mux_tmp_430 <= MUX_s_1_2_2(nor_326_nl, mux_tmp_429, nand_3_nl);
  nor_327_nl <= NOT((rem_12cyc_st_4_3_2(1)) OR (NOT mux_tmp_430));
  nand_4_nl <= NOT(main_stage_0_5 AND asn_itm_4 AND CONV_SL_1_1(rem_12cyc_st_4_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_4_3_2(0))));
  mux_tmp_431 <= MUX_s_1_2_2(nor_327_nl, mux_tmp_430, nand_4_nl);
  nor_328_nl <= NOT((rem_12cyc_st_3_3_2(1)) OR (NOT mux_tmp_431));
  nand_5_nl <= NOT(main_stage_0_4 AND asn_itm_3 AND CONV_SL_1_1(rem_12cyc_st_3_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_3_3_2(0))));
  mux_tmp_432 <= MUX_s_1_2_2(nor_328_nl, mux_tmp_431, nand_5_nl);
  nor_329_nl <= NOT((rem_12cyc_st_2_3_2(1)) OR (NOT mux_tmp_432));
  nand_6_nl <= NOT(main_stage_0_3 AND asn_itm_2 AND CONV_SL_1_1(rem_12cyc_st_2_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_2_3_2(0))));
  mux_tmp_433 <= MUX_s_1_2_2(nor_329_nl, mux_tmp_432, nand_6_nl);
  nor_330_nl <= NOT((rem_12cyc_st_9_3_2(1)) OR (NOT mux_tmp_433));
  nand_7_nl <= NOT(main_stage_0_10 AND asn_itm_9 AND CONV_SL_1_1(rem_12cyc_st_9_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_9_3_2(0))));
  mux_tmp_434 <= MUX_s_1_2_2(nor_330_nl, mux_tmp_433, nand_7_nl);
  nor_331_nl <= NOT((rem_12cyc_st_8_3_2(1)) OR (NOT mux_tmp_434));
  nand_8_nl <= NOT(main_stage_0_9 AND asn_itm_8 AND CONV_SL_1_1(rem_12cyc_st_8_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_8_3_2(0))));
  mux_tmp_435 <= MUX_s_1_2_2(nor_331_nl, mux_tmp_434, nand_8_nl);
  nor_332_nl <= NOT((rem_12cyc_st_7_3_2(1)) OR (NOT mux_tmp_435));
  nand_9_nl <= NOT(main_stage_0_8 AND asn_itm_7 AND CONV_SL_1_1(rem_12cyc_st_7_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_7_3_2(0))));
  mux_tmp_436 <= MUX_s_1_2_2(nor_332_nl, mux_tmp_435, nand_9_nl);
  and_934_nl <= nand_223_cse AND mux_tmp_436;
  nand_11_nl <= NOT(main_stage_0_2 AND asn_itm_1 AND CONV_SL_1_1(rem_12cyc_3_2=STD_LOGIC_VECTOR'("10")));
  mux_tmp_437 <= MUX_s_1_2_2(and_934_nl, mux_tmp_436, nand_11_nl);
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( ccs_ccore_en = '1' ) THEN
        return_rsci_d <= MUX_v_64_2_2(result_sva_duc_mx0, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(qelse_acc_nl),
            64)), mux_13_nl);
        m_buf_sva_12 <= m_buf_sva_11;
        m_buf_sva_11 <= m_buf_sva_10;
        m_buf_sva_10 <= m_buf_sva_9;
        m_buf_sva_9 <= m_buf_sva_8;
        m_buf_sva_8 <= m_buf_sva_7;
        m_buf_sva_7 <= m_buf_sva_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        asn_itm_12 <= '0';
        asn_itm_11 <= '0';
        asn_itm_10 <= '0';
        asn_itm_9 <= '0';
        asn_itm_8 <= '0';
        asn_itm_7 <= '0';
        asn_itm_6 <= '0';
        asn_itm_5 <= '0';
        asn_itm_4 <= '0';
        asn_itm_3 <= '0';
        asn_itm_2 <= '0';
        asn_itm_1 <= '0';
        main_stage_0_2 <= '0';
        main_stage_0_3 <= '0';
        main_stage_0_4 <= '0';
        main_stage_0_5 <= '0';
        main_stage_0_6 <= '0';
        main_stage_0_7 <= '0';
        main_stage_0_8 <= '0';
        main_stage_0_9 <= '0';
        main_stage_0_10 <= '0';
        main_stage_0_11 <= '0';
        main_stage_0_12 <= '0';
        main_stage_0_13 <= '0';
      ELSIF ( ccs_ccore_en = '1' ) THEN
        asn_itm_12 <= asn_itm_11;
        asn_itm_11 <= asn_itm_10;
        asn_itm_10 <= asn_itm_9;
        asn_itm_9 <= asn_itm_8;
        asn_itm_8 <= asn_itm_7;
        asn_itm_7 <= asn_itm_6;
        asn_itm_6 <= asn_itm_5;
        asn_itm_5 <= asn_itm_4;
        asn_itm_4 <= asn_itm_3;
        asn_itm_3 <= asn_itm_2;
        asn_itm_2 <= asn_itm_1;
        asn_itm_1 <= ccs_ccore_start_rsci_idat;
        main_stage_0_2 <= '1';
        main_stage_0_3 <= main_stage_0_2;
        main_stage_0_4 <= main_stage_0_3;
        main_stage_0_5 <= main_stage_0_4;
        main_stage_0_6 <= main_stage_0_5;
        main_stage_0_7 <= main_stage_0_6;
        main_stage_0_8 <= main_stage_0_7;
        main_stage_0_9 <= main_stage_0_8;
        main_stage_0_10 <= main_stage_0_9;
        main_stage_0_11 <= main_stage_0_10;
        main_stage_0_12 <= main_stage_0_11;
        main_stage_0_13 <= main_stage_0_12;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_sva_duc <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
      ELSIF ( (asn_itm_12 AND main_stage_0_13 AND ccs_ccore_en AND (NOT(CONV_SL_1_1(rem_12cyc_st_12_3_2=STD_LOGIC_VECTOR'("11")))))
          = '1' ) THEN
        result_sva_duc <= result_sva_duc_mx0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_12_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_12_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1203_cse = '1' ) THEN
        rem_12cyc_st_12_3_2 <= rem_12cyc_st_11_3_2;
        rem_12cyc_st_12_1_0 <= rem_12cyc_st_11_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1173_cse = '1' ) THEN
        rem_13_cmp_1_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_3_2_63_0, mut_3_3_63_0,
            mut_3_4_63_0, mut_3_5_63_0, mut_3_6_63_0, mut_3_7_63_0, mut_3_8_63_0,
            mut_3_9_63_0, mut_3_10_63_0, mut_3_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_294
            & and_dcpl_300 & and_dcpl_306 & and_dcpl_312 & and_dcpl_318 & and_dcpl_324
            & and_dcpl_330 & and_dcpl_336 & and_dcpl_342 & and_dcpl_348 & and_tmp_35));
        rem_13_cmp_1_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_2_2_63_0, mut_2_3_63_0,
            mut_2_4_63_0, mut_2_5_63_0, mut_2_6_63_0, mut_2_7_63_0, mut_2_8_63_0,
            mut_2_9_63_0, mut_2_10_63_0, mut_2_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_294
            & and_dcpl_300 & and_dcpl_306 & and_dcpl_312 & and_dcpl_318 & and_dcpl_324
            & and_dcpl_330 & and_dcpl_336 & and_dcpl_342 & and_dcpl_348 & and_tmp_35));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1175_cse = '1' ) THEN
        rem_13_cmp_2_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_5_2_63_0, mut_5_3_63_0,
            mut_5_4_63_0, mut_5_5_63_0, mut_5_6_63_0, mut_5_7_63_0, mut_5_8_63_0,
            mut_5_9_63_0, mut_5_10_63_0, mut_5_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_356
            & and_dcpl_360 & and_dcpl_364 & and_dcpl_368 & and_dcpl_372 & and_dcpl_376
            & and_dcpl_379 & and_dcpl_382 & and_dcpl_385 & and_dcpl_388 & mux_tmp_76));
        rem_13_cmp_2_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_4_2_63_0, mut_4_3_63_0,
            mut_4_4_63_0, mut_4_5_63_0, mut_4_6_63_0, mut_4_7_63_0, mut_4_8_63_0,
            mut_4_9_63_0, mut_4_10_63_0, mut_4_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_356
            & and_dcpl_360 & and_dcpl_364 & and_dcpl_368 & and_dcpl_372 & and_dcpl_376
            & and_dcpl_379 & and_dcpl_382 & and_dcpl_385 & and_dcpl_388 & mux_tmp_76));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1177_cse = '1' ) THEN
        rem_13_cmp_3_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_7_2_63_0, mut_7_3_63_0,
            mut_7_4_63_0, mut_7_5_63_0, mut_7_6_63_0, mut_7_7_63_0, mut_7_8_63_0,
            mut_7_9_63_0, mut_7_10_63_0, mut_7_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_394
            & and_dcpl_397 & and_dcpl_400 & and_dcpl_403 & and_dcpl_406 & and_dcpl_409
            & and_dcpl_413 & and_dcpl_417 & and_dcpl_421 & and_dcpl_425 & and_tmp_80));
        rem_13_cmp_3_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_6_2_63_0, mut_6_3_63_0,
            mut_6_4_63_0, mut_6_5_63_0, mut_6_6_63_0, mut_6_7_63_0, mut_6_8_63_0,
            mut_6_9_63_0, mut_6_10_63_0, mut_6_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_394
            & and_dcpl_397 & and_dcpl_400 & and_dcpl_403 & and_dcpl_406 & and_dcpl_409
            & and_dcpl_413 & and_dcpl_417 & and_dcpl_421 & and_dcpl_425 & and_tmp_80));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1179_cse = '1' ) THEN
        rem_13_cmp_4_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_9_2_63_0, mut_9_3_63_0,
            mut_9_4_63_0, mut_9_5_63_0, mut_9_6_63_0, mut_9_7_63_0, mut_9_8_63_0,
            mut_9_9_63_0, mut_9_10_63_0, mut_9_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_431
            & and_dcpl_433 & and_dcpl_435 & and_dcpl_437 & and_dcpl_439 & and_dcpl_442
            & and_dcpl_445 & and_dcpl_448 & and_dcpl_451 & and_dcpl_454 & mux_tmp_141));
        rem_13_cmp_4_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_8_2_63_0, mut_8_3_63_0,
            mut_8_4_63_0, mut_8_5_63_0, mut_8_6_63_0, mut_8_7_63_0, mut_8_8_63_0,
            mut_8_9_63_0, mut_8_10_63_0, mut_8_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_431
            & and_dcpl_433 & and_dcpl_435 & and_dcpl_437 & and_dcpl_439 & and_dcpl_442
            & and_dcpl_445 & and_dcpl_448 & and_dcpl_451 & and_dcpl_454 & mux_tmp_141));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1181_cse = '1' ) THEN
        rem_13_cmp_5_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_11_2_63_0, mut_11_3_63_0,
            mut_11_4_63_0, mut_11_5_63_0, mut_11_6_63_0, mut_11_7_63_0, mut_11_8_63_0,
            mut_11_9_63_0, mut_11_10_63_0, mut_11_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_461
            & and_dcpl_465 & and_dcpl_469 & and_dcpl_473 & and_dcpl_477 & and_dcpl_480
            & and_dcpl_483 & and_dcpl_486 & and_dcpl_489 & and_dcpl_492 & and_tmp_125));
        rem_13_cmp_5_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_10_2_63_0, mut_10_3_63_0,
            mut_10_4_63_0, mut_10_5_63_0, mut_10_6_63_0, mut_10_7_63_0, mut_10_8_63_0,
            mut_10_9_63_0, mut_10_10_63_0, mut_10_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_461
            & and_dcpl_465 & and_dcpl_469 & and_dcpl_473 & and_dcpl_477 & and_dcpl_480
            & and_dcpl_483 & and_dcpl_486 & and_dcpl_489 & and_dcpl_492 & and_tmp_125));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1183_cse = '1' ) THEN
        rem_13_cmp_6_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_13_2_63_0, mut_13_3_63_0,
            mut_13_4_63_0, mut_13_5_63_0, mut_13_6_63_0, mut_13_7_63_0, mut_13_8_63_0,
            mut_13_9_63_0, mut_13_10_63_0, mut_13_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_498
            & and_dcpl_500 & and_dcpl_502 & and_dcpl_504 & and_dcpl_506 & and_dcpl_508
            & and_dcpl_510 & and_dcpl_512 & and_dcpl_514 & and_dcpl_516 & mux_tmp_206));
        rem_13_cmp_6_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_12_2_63_0, mut_12_3_63_0,
            mut_12_4_63_0, mut_12_5_63_0, mut_12_6_63_0, mut_12_7_63_0, mut_12_8_63_0,
            mut_12_9_63_0, mut_12_10_63_0, mut_12_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_498
            & and_dcpl_500 & and_dcpl_502 & and_dcpl_504 & and_dcpl_506 & and_dcpl_508
            & and_dcpl_510 & and_dcpl_512 & and_dcpl_514 & and_dcpl_516 & mux_tmp_206));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1185_cse = '1' ) THEN
        rem_13_cmp_7_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_15_2_63_0, mut_15_3_63_0,
            mut_15_4_63_0, mut_15_5_63_0, mut_15_6_63_0, mut_15_7_63_0, mut_15_8_63_0,
            mut_15_9_63_0, mut_15_10_63_0, mut_15_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_520
            & and_dcpl_523 & and_dcpl_526 & and_dcpl_529 & and_dcpl_532 & and_dcpl_534
            & and_dcpl_536 & and_dcpl_538 & and_dcpl_540 & and_dcpl_542 & and_tmp_170));
        rem_13_cmp_7_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_14_2_63_0, mut_14_3_63_0,
            mut_14_4_63_0, mut_14_5_63_0, mut_14_6_63_0, mut_14_7_63_0, mut_14_8_63_0,
            mut_14_9_63_0, mut_14_10_63_0, mut_14_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_520
            & and_dcpl_523 & and_dcpl_526 & and_dcpl_529 & and_dcpl_532 & and_dcpl_534
            & and_dcpl_536 & and_dcpl_538 & and_dcpl_540 & and_dcpl_542 & and_tmp_170));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1187_cse = '1' ) THEN
        rem_13_cmp_8_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_17_2_63_0, mut_17_3_63_0,
            mut_17_4_63_0, mut_17_5_63_0, mut_17_6_63_0, mut_17_7_63_0, mut_17_8_63_0,
            mut_17_9_63_0, mut_17_10_63_0, mut_17_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_546
            & and_dcpl_548 & and_dcpl_550 & and_dcpl_552 & and_dcpl_554 & and_dcpl_556
            & and_dcpl_558 & and_dcpl_560 & and_dcpl_562 & and_dcpl_564 & mux_tmp_271));
        rem_13_cmp_8_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_16_2_63_0, mut_16_3_63_0,
            mut_16_4_63_0, mut_16_5_63_0, mut_16_6_63_0, mut_16_7_63_0, mut_16_8_63_0,
            mut_16_9_63_0, mut_16_10_63_0, mut_16_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_546
            & and_dcpl_548 & and_dcpl_550 & and_dcpl_552 & and_dcpl_554 & and_dcpl_556
            & and_dcpl_558 & and_dcpl_560 & and_dcpl_562 & and_dcpl_564 & mux_tmp_271));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1189_cse = '1' ) THEN
        rem_13_cmp_9_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_19_2_63_0, mut_19_3_63_0,
            mut_19_4_63_0, mut_19_5_63_0, mut_19_6_63_0, mut_19_7_63_0, mut_19_8_63_0,
            mut_19_9_63_0, mut_19_10_63_0, mut_19_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_569
            & and_dcpl_573 & and_dcpl_577 & and_dcpl_581 & and_dcpl_585 & and_dcpl_589
            & and_dcpl_593 & and_dcpl_597 & and_dcpl_601 & and_dcpl_605 & and_tmp_206));
        rem_13_cmp_9_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_18_2_63_0, mut_18_3_63_0,
            mut_18_4_63_0, mut_18_5_63_0, mut_18_6_63_0, mut_18_7_63_0, mut_18_8_63_0,
            mut_18_9_63_0, mut_18_10_63_0, mut_18_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_569
            & and_dcpl_573 & and_dcpl_577 & and_dcpl_581 & and_dcpl_585 & and_dcpl_589
            & and_dcpl_593 & and_dcpl_597 & and_dcpl_601 & and_dcpl_605 & and_tmp_206));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1191_cse = '1' ) THEN
        rem_13_cmp_10_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_21_2_63_0, mut_21_3_63_0,
            mut_21_4_63_0, mut_21_5_63_0, mut_21_6_63_0, mut_21_7_63_0, mut_21_8_63_0,
            mut_21_9_63_0, mut_21_10_63_0, mut_21_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_610
            & and_dcpl_612 & and_dcpl_614 & and_dcpl_616 & and_dcpl_618 & and_dcpl_622
            & and_dcpl_625 & and_dcpl_628 & and_dcpl_631 & and_dcpl_634 & mux_tmp_354));
        rem_13_cmp_10_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_20_2_63_0,
            mut_20_3_63_0, mut_20_4_63_0, mut_20_5_63_0, mut_20_6_63_0, mut_20_7_63_0,
            mut_20_8_63_0, mut_20_9_63_0, mut_20_10_63_0, mut_20_11_63_0, STD_LOGIC_VECTOR'(
            and_dcpl_610 & and_dcpl_612 & and_dcpl_614 & and_dcpl_616 & and_dcpl_618
            & and_dcpl_622 & and_dcpl_625 & and_dcpl_628 & and_dcpl_631 & and_dcpl_634
            & mux_tmp_354));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1193_cse = '1' ) THEN
        rem_13_cmp_11_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_23_2_63_0, mut_23_3_63_0,
            mut_23_4_63_0, mut_23_5_63_0, mut_23_6_63_0, mut_23_7_63_0, mut_23_8_63_0,
            mut_23_9_63_0, mut_23_10_63_0, mut_23_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_638
            & and_dcpl_641 & and_dcpl_644 & and_dcpl_647 & and_dcpl_650 & and_dcpl_653
            & and_dcpl_657 & and_dcpl_661 & and_dcpl_665 & and_dcpl_669 & and_tmp_233));
        rem_13_cmp_11_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_22_2_63_0,
            mut_22_3_63_0, mut_22_4_63_0, mut_22_5_63_0, mut_22_6_63_0, mut_22_7_63_0,
            mut_22_8_63_0, mut_22_9_63_0, mut_22_10_63_0, mut_22_11_63_0, STD_LOGIC_VECTOR'(
            and_dcpl_638 & and_dcpl_641 & and_dcpl_644 & and_dcpl_647 & and_dcpl_650
            & and_dcpl_653 & and_dcpl_657 & and_dcpl_661 & and_dcpl_665 & and_dcpl_669
            & and_tmp_233));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1195_cse = '1' ) THEN
        rem_13_cmp_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_1_2_63_0, mut_1_3_63_0,
            mut_1_4_63_0, mut_1_5_63_0, mut_1_6_63_0, mut_1_7_63_0, mut_1_8_63_0,
            mut_1_9_63_0, mut_1_10_63_0, mut_1_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_673
            & and_dcpl_675 & and_dcpl_677 & and_dcpl_679 & and_dcpl_681 & and_dcpl_684
            & and_dcpl_687 & and_dcpl_690 & and_dcpl_693 & and_dcpl_696 & mux_tmp_437));
        rem_13_cmp_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_2_63_0, mut_3_63_0,
            mut_4_63_0, mut_5_63_0, mut_6_63_0, mut_7_63_0, mut_8_63_0, mut_9_63_0,
            mut_10_63_0, mut_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_673 & and_dcpl_675
            & and_dcpl_677 & and_dcpl_679 & and_dcpl_681 & and_dcpl_684 & and_dcpl_687
            & and_dcpl_690 & and_dcpl_693 & and_dcpl_696 & mux_tmp_437));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1205_cse = '1' ) THEN
        mut_3_11_63_0 <= mut_3_10_63_0;
        mut_2_11_63_0 <= mut_2_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1207_cse = '1' ) THEN
        mut_5_11_63_0 <= mut_5_10_63_0;
        mut_4_11_63_0 <= mut_4_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1209_cse = '1' ) THEN
        mut_7_11_63_0 <= mut_7_10_63_0;
        mut_6_11_63_0 <= mut_6_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1211_cse = '1' ) THEN
        mut_9_11_63_0 <= mut_9_10_63_0;
        mut_8_11_63_0 <= mut_8_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1213_cse = '1' ) THEN
        mut_11_11_63_0 <= mut_11_10_63_0;
        mut_10_11_63_0 <= mut_10_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1215_cse = '1' ) THEN
        mut_13_11_63_0 <= mut_13_10_63_0;
        mut_12_11_63_0 <= mut_12_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1217_cse = '1' ) THEN
        mut_15_11_63_0 <= mut_15_10_63_0;
        mut_14_11_63_0 <= mut_14_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1219_cse = '1' ) THEN
        mut_17_11_63_0 <= mut_17_10_63_0;
        mut_16_11_63_0 <= mut_16_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1221_cse = '1' ) THEN
        mut_19_11_63_0 <= mut_19_10_63_0;
        mut_18_11_63_0 <= mut_18_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1223_cse = '1' ) THEN
        mut_21_11_63_0 <= mut_21_10_63_0;
        mut_20_11_63_0 <= mut_20_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1225_cse = '1' ) THEN
        mut_23_11_63_0 <= mut_23_10_63_0;
        mut_22_11_63_0 <= mut_22_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1227_cse = '1' ) THEN
        mut_1_11_63_0 <= mut_1_10_63_0;
        mut_11_63_0 <= mut_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_11_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_11_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1229_cse = '1' ) THEN
        rem_12cyc_st_11_3_2 <= rem_12cyc_st_10_3_2;
        rem_12cyc_st_11_1_0 <= rem_12cyc_st_10_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1231_cse = '1' ) THEN
        mut_3_10_63_0 <= mut_3_9_63_0;
        mut_2_10_63_0 <= mut_2_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1233_cse = '1' ) THEN
        mut_5_10_63_0 <= mut_5_9_63_0;
        mut_4_10_63_0 <= mut_4_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1235_cse = '1' ) THEN
        mut_7_10_63_0 <= mut_7_9_63_0;
        mut_6_10_63_0 <= mut_6_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1237_cse = '1' ) THEN
        mut_9_10_63_0 <= mut_9_9_63_0;
        mut_8_10_63_0 <= mut_8_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1239_cse = '1' ) THEN
        mut_11_10_63_0 <= mut_11_9_63_0;
        mut_10_10_63_0 <= mut_10_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1241_cse = '1' ) THEN
        mut_13_10_63_0 <= mut_13_9_63_0;
        mut_12_10_63_0 <= mut_12_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1243_cse = '1' ) THEN
        mut_15_10_63_0 <= mut_15_9_63_0;
        mut_14_10_63_0 <= mut_14_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1245_cse = '1' ) THEN
        mut_17_10_63_0 <= mut_17_9_63_0;
        mut_16_10_63_0 <= mut_16_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1247_cse = '1' ) THEN
        mut_19_10_63_0 <= mut_19_9_63_0;
        mut_18_10_63_0 <= mut_18_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1249_cse = '1' ) THEN
        mut_21_10_63_0 <= mut_21_9_63_0;
        mut_20_10_63_0 <= mut_20_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1251_cse = '1' ) THEN
        mut_23_10_63_0 <= mut_23_9_63_0;
        mut_22_10_63_0 <= mut_22_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1253_cse = '1' ) THEN
        mut_1_10_63_0 <= mut_1_9_63_0;
        mut_10_63_0 <= mut_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_10_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_10_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1255_cse = '1' ) THEN
        rem_12cyc_st_10_3_2 <= rem_12cyc_st_9_3_2;
        rem_12cyc_st_10_1_0 <= rem_12cyc_st_9_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1257_cse = '1' ) THEN
        mut_3_9_63_0 <= mut_3_8_63_0;
        mut_2_9_63_0 <= mut_2_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1259_cse = '1' ) THEN
        mut_5_9_63_0 <= mut_5_8_63_0;
        mut_4_9_63_0 <= mut_4_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1261_cse = '1' ) THEN
        mut_7_9_63_0 <= mut_7_8_63_0;
        mut_6_9_63_0 <= mut_6_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1263_cse = '1' ) THEN
        mut_9_9_63_0 <= mut_9_8_63_0;
        mut_8_9_63_0 <= mut_8_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1265_cse = '1' ) THEN
        mut_11_9_63_0 <= mut_11_8_63_0;
        mut_10_9_63_0 <= mut_10_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1267_cse = '1' ) THEN
        mut_13_9_63_0 <= mut_13_8_63_0;
        mut_12_9_63_0 <= mut_12_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1269_cse = '1' ) THEN
        mut_15_9_63_0 <= mut_15_8_63_0;
        mut_14_9_63_0 <= mut_14_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1271_cse = '1' ) THEN
        mut_17_9_63_0 <= mut_17_8_63_0;
        mut_16_9_63_0 <= mut_16_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1273_cse = '1' ) THEN
        mut_19_9_63_0 <= mut_19_8_63_0;
        mut_18_9_63_0 <= mut_18_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1275_cse = '1' ) THEN
        mut_21_9_63_0 <= mut_21_8_63_0;
        mut_20_9_63_0 <= mut_20_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1277_cse = '1' ) THEN
        mut_23_9_63_0 <= mut_23_8_63_0;
        mut_22_9_63_0 <= mut_22_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1279_cse = '1' ) THEN
        mut_1_9_63_0 <= mut_1_8_63_0;
        mut_9_63_0 <= mut_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_9_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_9_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1281_cse = '1' ) THEN
        rem_12cyc_st_9_3_2 <= rem_12cyc_st_8_3_2;
        rem_12cyc_st_9_1_0 <= rem_12cyc_st_8_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1283_cse = '1' ) THEN
        mut_3_8_63_0 <= mut_3_7_63_0;
        mut_2_8_63_0 <= mut_2_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1285_cse = '1' ) THEN
        mut_5_8_63_0 <= mut_5_7_63_0;
        mut_4_8_63_0 <= mut_4_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1287_cse = '1' ) THEN
        mut_7_8_63_0 <= mut_7_7_63_0;
        mut_6_8_63_0 <= mut_6_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1289_cse = '1' ) THEN
        mut_9_8_63_0 <= mut_9_7_63_0;
        mut_8_8_63_0 <= mut_8_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1291_cse = '1' ) THEN
        mut_11_8_63_0 <= mut_11_7_63_0;
        mut_10_8_63_0 <= mut_10_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1293_cse = '1' ) THEN
        mut_13_8_63_0 <= mut_13_7_63_0;
        mut_12_8_63_0 <= mut_12_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1295_cse = '1' ) THEN
        mut_15_8_63_0 <= mut_15_7_63_0;
        mut_14_8_63_0 <= mut_14_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1297_cse = '1' ) THEN
        mut_17_8_63_0 <= mut_17_7_63_0;
        mut_16_8_63_0 <= mut_16_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1299_cse = '1' ) THEN
        mut_19_8_63_0 <= mut_19_7_63_0;
        mut_18_8_63_0 <= mut_18_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1301_cse = '1' ) THEN
        mut_21_8_63_0 <= mut_21_7_63_0;
        mut_20_8_63_0 <= mut_20_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1303_cse = '1' ) THEN
        mut_23_8_63_0 <= mut_23_7_63_0;
        mut_22_8_63_0 <= mut_22_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1305_cse = '1' ) THEN
        mut_1_8_63_0 <= mut_1_7_63_0;
        mut_8_63_0 <= mut_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_8_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_8_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1307_cse = '1' ) THEN
        rem_12cyc_st_8_3_2 <= rem_12cyc_st_7_3_2;
        rem_12cyc_st_8_1_0 <= rem_12cyc_st_7_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1309_cse = '1' ) THEN
        mut_3_7_63_0 <= mut_3_6_63_0;
        mut_2_7_63_0 <= mut_2_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1311_cse = '1' ) THEN
        mut_5_7_63_0 <= mut_5_6_63_0;
        mut_4_7_63_0 <= mut_4_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1313_cse = '1' ) THEN
        mut_7_7_63_0 <= mut_7_6_63_0;
        mut_6_7_63_0 <= mut_6_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1315_cse = '1' ) THEN
        mut_9_7_63_0 <= mut_9_6_63_0;
        mut_8_7_63_0 <= mut_8_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1317_cse = '1' ) THEN
        mut_11_7_63_0 <= mut_11_6_63_0;
        mut_10_7_63_0 <= mut_10_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1319_cse = '1' ) THEN
        mut_13_7_63_0 <= mut_13_6_63_0;
        mut_12_7_63_0 <= mut_12_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1321_cse = '1' ) THEN
        mut_15_7_63_0 <= mut_15_6_63_0;
        mut_14_7_63_0 <= mut_14_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1323_cse = '1' ) THEN
        mut_17_7_63_0 <= mut_17_6_63_0;
        mut_16_7_63_0 <= mut_16_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1325_cse = '1' ) THEN
        mut_19_7_63_0 <= mut_19_6_63_0;
        mut_18_7_63_0 <= mut_18_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1327_cse = '1' ) THEN
        mut_21_7_63_0 <= mut_21_6_63_0;
        mut_20_7_63_0 <= mut_20_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1329_cse = '1' ) THEN
        mut_23_7_63_0 <= mut_23_6_63_0;
        mut_22_7_63_0 <= mut_22_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1331_cse = '1' ) THEN
        mut_1_7_63_0 <= mut_1_6_63_0;
        mut_7_63_0 <= mut_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_7_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_7_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1333_cse = '1' ) THEN
        rem_12cyc_st_7_3_2 <= rem_12cyc_st_6_3_2;
        rem_12cyc_st_7_1_0 <= rem_12cyc_st_6_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1335_cse = '1' ) THEN
        mut_3_6_63_0 <= mut_3_5_63_0;
        mut_2_6_63_0 <= mut_2_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1337_cse = '1' ) THEN
        mut_5_6_63_0 <= mut_5_5_63_0;
        mut_4_6_63_0 <= mut_4_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1339_cse = '1' ) THEN
        mut_7_6_63_0 <= mut_7_5_63_0;
        mut_6_6_63_0 <= mut_6_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1341_cse = '1' ) THEN
        mut_9_6_63_0 <= mut_9_5_63_0;
        mut_8_6_63_0 <= mut_8_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1343_cse = '1' ) THEN
        mut_11_6_63_0 <= mut_11_5_63_0;
        mut_10_6_63_0 <= mut_10_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1345_cse = '1' ) THEN
        mut_13_6_63_0 <= mut_13_5_63_0;
        mut_12_6_63_0 <= mut_12_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1347_cse = '1' ) THEN
        mut_15_6_63_0 <= mut_15_5_63_0;
        mut_14_6_63_0 <= mut_14_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1349_cse = '1' ) THEN
        mut_17_6_63_0 <= mut_17_5_63_0;
        mut_16_6_63_0 <= mut_16_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1351_cse = '1' ) THEN
        mut_19_6_63_0 <= mut_19_5_63_0;
        mut_18_6_63_0 <= mut_18_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1353_cse = '1' ) THEN
        mut_21_6_63_0 <= mut_21_5_63_0;
        mut_20_6_63_0 <= mut_20_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1355_cse = '1' ) THEN
        mut_23_6_63_0 <= mut_23_5_63_0;
        mut_22_6_63_0 <= mut_22_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1357_cse = '1' ) THEN
        mut_1_6_63_0 <= mut_1_5_63_0;
        mut_6_63_0 <= mut_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1359_cse = '1' ) THEN
        m_buf_sva_6 <= m_buf_sva_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_6_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_6_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1359_cse = '1' ) THEN
        rem_12cyc_st_6_3_2 <= rem_12cyc_st_5_3_2;
        rem_12cyc_st_6_1_0 <= rem_12cyc_st_5_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1361_cse = '1' ) THEN
        mut_3_5_63_0 <= mut_3_4_63_0;
        mut_2_5_63_0 <= mut_2_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1363_cse = '1' ) THEN
        mut_5_5_63_0 <= mut_5_4_63_0;
        mut_4_5_63_0 <= mut_4_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1365_cse = '1' ) THEN
        mut_7_5_63_0 <= mut_7_4_63_0;
        mut_6_5_63_0 <= mut_6_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1367_cse = '1' ) THEN
        mut_9_5_63_0 <= mut_9_4_63_0;
        mut_8_5_63_0 <= mut_8_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1369_cse = '1' ) THEN
        mut_11_5_63_0 <= mut_11_4_63_0;
        mut_10_5_63_0 <= mut_10_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1371_cse = '1' ) THEN
        mut_13_5_63_0 <= mut_13_4_63_0;
        mut_12_5_63_0 <= mut_12_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1373_cse = '1' ) THEN
        mut_15_5_63_0 <= mut_15_4_63_0;
        mut_14_5_63_0 <= mut_14_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1375_cse = '1' ) THEN
        mut_17_5_63_0 <= mut_17_4_63_0;
        mut_16_5_63_0 <= mut_16_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1377_cse = '1' ) THEN
        mut_19_5_63_0 <= mut_19_4_63_0;
        mut_18_5_63_0 <= mut_18_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1379_cse = '1' ) THEN
        mut_21_5_63_0 <= mut_21_4_63_0;
        mut_20_5_63_0 <= mut_20_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1381_cse = '1' ) THEN
        mut_23_5_63_0 <= mut_23_4_63_0;
        mut_22_5_63_0 <= mut_22_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1383_cse = '1' ) THEN
        mut_1_5_63_0 <= mut_1_4_63_0;
        mut_5_63_0 <= mut_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1385_cse = '1' ) THEN
        m_buf_sva_5 <= m_buf_sva_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_5_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_5_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1385_cse = '1' ) THEN
        rem_12cyc_st_5_3_2 <= rem_12cyc_st_4_3_2;
        rem_12cyc_st_5_1_0 <= rem_12cyc_st_4_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1387_cse = '1' ) THEN
        mut_3_4_63_0 <= mut_3_3_63_0;
        mut_2_4_63_0 <= mut_2_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1389_cse = '1' ) THEN
        mut_5_4_63_0 <= mut_5_3_63_0;
        mut_4_4_63_0 <= mut_4_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1391_cse = '1' ) THEN
        mut_7_4_63_0 <= mut_7_3_63_0;
        mut_6_4_63_0 <= mut_6_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1393_cse = '1' ) THEN
        mut_9_4_63_0 <= mut_9_3_63_0;
        mut_8_4_63_0 <= mut_8_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1395_cse = '1' ) THEN
        mut_11_4_63_0 <= mut_11_3_63_0;
        mut_10_4_63_0 <= mut_10_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1397_cse = '1' ) THEN
        mut_13_4_63_0 <= mut_13_3_63_0;
        mut_12_4_63_0 <= mut_12_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1399_cse = '1' ) THEN
        mut_15_4_63_0 <= mut_15_3_63_0;
        mut_14_4_63_0 <= mut_14_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1401_cse = '1' ) THEN
        mut_17_4_63_0 <= mut_17_3_63_0;
        mut_16_4_63_0 <= mut_16_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1403_cse = '1' ) THEN
        mut_19_4_63_0 <= mut_19_3_63_0;
        mut_18_4_63_0 <= mut_18_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1405_cse = '1' ) THEN
        mut_21_4_63_0 <= mut_21_3_63_0;
        mut_20_4_63_0 <= mut_20_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1407_cse = '1' ) THEN
        mut_23_4_63_0 <= mut_23_3_63_0;
        mut_22_4_63_0 <= mut_22_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1409_cse = '1' ) THEN
        mut_1_4_63_0 <= mut_1_3_63_0;
        mut_4_63_0 <= mut_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1411_cse = '1' ) THEN
        m_buf_sva_4 <= m_buf_sva_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_4_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_4_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1411_cse = '1' ) THEN
        rem_12cyc_st_4_3_2 <= rem_12cyc_st_3_3_2;
        rem_12cyc_st_4_1_0 <= rem_12cyc_st_3_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1413_cse = '1' ) THEN
        mut_3_3_63_0 <= mut_3_2_63_0;
        mut_2_3_63_0 <= mut_2_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1415_cse = '1' ) THEN
        mut_5_3_63_0 <= mut_5_2_63_0;
        mut_4_3_63_0 <= mut_4_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1417_cse = '1' ) THEN
        mut_7_3_63_0 <= mut_7_2_63_0;
        mut_6_3_63_0 <= mut_6_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1419_cse = '1' ) THEN
        mut_9_3_63_0 <= mut_9_2_63_0;
        mut_8_3_63_0 <= mut_8_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1421_cse = '1' ) THEN
        mut_11_3_63_0 <= mut_11_2_63_0;
        mut_10_3_63_0 <= mut_10_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1423_cse = '1' ) THEN
        mut_13_3_63_0 <= mut_13_2_63_0;
        mut_12_3_63_0 <= mut_12_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1425_cse = '1' ) THEN
        mut_15_3_63_0 <= mut_15_2_63_0;
        mut_14_3_63_0 <= mut_14_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1427_cse = '1' ) THEN
        mut_17_3_63_0 <= mut_17_2_63_0;
        mut_16_3_63_0 <= mut_16_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1429_cse = '1' ) THEN
        mut_19_3_63_0 <= mut_19_2_63_0;
        mut_18_3_63_0 <= mut_18_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1431_cse = '1' ) THEN
        mut_21_3_63_0 <= mut_21_2_63_0;
        mut_20_3_63_0 <= mut_20_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1433_cse = '1' ) THEN
        mut_23_3_63_0 <= mut_23_2_63_0;
        mut_22_3_63_0 <= mut_22_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1435_cse = '1' ) THEN
        mut_1_3_63_0 <= mut_1_2_63_0;
        mut_3_63_0 <= mut_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1437_cse = '1' ) THEN
        m_buf_sva_3 <= m_buf_sva_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_3_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_3_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1437_cse = '1' ) THEN
        rem_12cyc_st_3_3_2 <= rem_12cyc_st_2_3_2;
        rem_12cyc_st_3_1_0 <= rem_12cyc_st_2_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1439_cse = '1' ) THEN
        mut_3_2_63_0 <= rem_13_cmp_1_b_63_0;
        mut_2_2_63_0 <= rem_13_cmp_1_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1441_cse = '1' ) THEN
        mut_5_2_63_0 <= rem_13_cmp_2_b_63_0;
        mut_4_2_63_0 <= rem_13_cmp_2_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1443_cse = '1' ) THEN
        mut_7_2_63_0 <= rem_13_cmp_3_b_63_0;
        mut_6_2_63_0 <= rem_13_cmp_3_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1445_cse = '1' ) THEN
        mut_9_2_63_0 <= rem_13_cmp_4_b_63_0;
        mut_8_2_63_0 <= rem_13_cmp_4_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1447_cse = '1' ) THEN
        mut_11_2_63_0 <= rem_13_cmp_5_b_63_0;
        mut_10_2_63_0 <= rem_13_cmp_5_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1449_cse = '1' ) THEN
        mut_13_2_63_0 <= rem_13_cmp_6_b_63_0;
        mut_12_2_63_0 <= rem_13_cmp_6_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1451_cse = '1' ) THEN
        mut_15_2_63_0 <= rem_13_cmp_7_b_63_0;
        mut_14_2_63_0 <= rem_13_cmp_7_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1453_cse = '1' ) THEN
        mut_17_2_63_0 <= rem_13_cmp_8_b_63_0;
        mut_16_2_63_0 <= rem_13_cmp_8_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1455_cse = '1' ) THEN
        mut_19_2_63_0 <= rem_13_cmp_9_b_63_0;
        mut_18_2_63_0 <= rem_13_cmp_9_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1457_cse = '1' ) THEN
        mut_21_2_63_0 <= rem_13_cmp_10_b_63_0;
        mut_20_2_63_0 <= rem_13_cmp_10_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1459_cse = '1' ) THEN
        mut_23_2_63_0 <= rem_13_cmp_11_b_63_0;
        mut_22_2_63_0 <= rem_13_cmp_11_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1461_cse = '1' ) THEN
        mut_1_2_63_0 <= rem_13_cmp_b_63_0;
        mut_2_63_0 <= rem_13_cmp_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1463_cse = '1' ) THEN
        m_buf_sva_2 <= m_buf_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_2_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_2_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1463_cse = '1' ) THEN
        rem_12cyc_st_2_3_2 <= rem_12cyc_3_2;
        rem_12cyc_st_2_1_0 <= rem_12cyc_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1197_cse = '1' ) THEN
        m_buf_sva_1 <= m_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1197_cse = '1' ) THEN
        rem_12cyc_3_2 <= acc_tmp;
        rem_12cyc_1_0 <= acc_1_tmp(1 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  qelse_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(result_sva_duc_mx0) + UNSIGNED(m_buf_sva_12),
      64));
  mux_10_nl <= MUX_s_1_2_2((rem_13_cmp_1_z(63)), (rem_13_cmp_3_z(63)), rem_12cyc_st_12_1_0(1));
  mux_9_nl <= MUX_s_1_2_2((rem_13_cmp_2_z(63)), (rem_13_cmp_4_z(63)), rem_12cyc_st_12_1_0(1));
  mux_11_nl <= MUX_s_1_2_2(mux_10_nl, mux_9_nl, rem_12cyc_st_12_1_0(0));
  mux_7_nl <= MUX_s_1_2_2((rem_13_cmp_9_z(63)), (rem_13_cmp_11_z(63)), rem_12cyc_st_12_1_0(1));
  mux_6_nl <= MUX_s_1_2_2((rem_13_cmp_10_z(63)), (rem_13_cmp_z(63)), rem_12cyc_st_12_1_0(1));
  mux_8_nl <= MUX_s_1_2_2(mux_7_nl, mux_6_nl, rem_12cyc_st_12_1_0(0));
  mux_12_nl <= MUX_s_1_2_2(mux_11_nl, mux_8_nl, rem_12cyc_st_12_3_2(1));
  mux_3_nl <= MUX_s_1_2_2((rem_13_cmp_5_z(63)), (rem_13_cmp_7_z(63)), rem_12cyc_st_12_1_0(1));
  mux_2_nl <= MUX_s_1_2_2((rem_13_cmp_6_z(63)), (rem_13_cmp_8_z(63)), rem_12cyc_st_12_1_0(1));
  mux_4_nl <= MUX_s_1_2_2(mux_3_nl, mux_2_nl, rem_12cyc_st_12_1_0(0));
  mux_5_nl <= MUX_s_1_2_2(mux_4_nl, (result_sva_duc(63)), rem_12cyc_st_12_3_2(1));
  mux_13_nl <= MUX_s_1_2_2(mux_12_nl, mux_5_nl, rem_12cyc_st_12_3_2(0));
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    modulo_dev
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;
USE work.mgc_comps.ALL;


ENTITY modulo_dev IS
  PORT(
    base_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    m_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    return_rsc_z : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    ccs_ccore_start_rsc_dat : IN STD_LOGIC;
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_srst : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC
  );
END modulo_dev;

ARCHITECTURE v1 OF modulo_dev IS
  -- Default Constants

  COMPONENT modulo_dev_core
    PORT(
      base_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      m_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      return_rsc_z : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      ccs_ccore_start_rsc_dat : IN STD_LOGIC;
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_srst : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL modulo_dev_core_inst_base_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_dev_core_inst_m_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_dev_core_inst_return_rsc_z : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  modulo_dev_core_inst : modulo_dev_core
    PORT MAP(
      base_rsc_dat => modulo_dev_core_inst_base_rsc_dat,
      m_rsc_dat => modulo_dev_core_inst_m_rsc_dat,
      return_rsc_z => modulo_dev_core_inst_return_rsc_z,
      ccs_ccore_start_rsc_dat => ccs_ccore_start_rsc_dat,
      ccs_ccore_clk => ccs_ccore_clk,
      ccs_ccore_srst => ccs_ccore_srst,
      ccs_ccore_en => ccs_ccore_en
    );
  modulo_dev_core_inst_base_rsc_dat <= base_rsc_dat;
  modulo_dev_core_inst_m_rsc_dat <= m_rsc_dat;
  return_rsc_z <= modulo_dev_core_inst_return_rsc_z;

END v1;




--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_div IS
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END mgc_div;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

USE work.funcs.all;

ARCHITECTURE beh OF mgc_div IS
BEGIN
  z <= std_logic_vector(unsigned(a) / unsigned(b)) WHEN signd = 0 ELSE
       std_logic_vector(  signed(a) /   signed(b));
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_comps_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_shift_comps_v5 IS

COMPONENT mgc_shift_l_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_shift_comps_v5;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_shift_l_v5 IS
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_shift_l_v5;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_shift_l_v5 IS

  FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1 > arg2) THEN
      RETURN(arg1) ;
    ELSE
      RETURN(arg2) ;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(SIGNED(result), arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE)
  RETURN UNSIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, '0', olen);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE)
  RETURN SIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen);
  END;

BEGIN
UNSGNED:  IF signd_a = 0 GENERATE
    z <= std_logic_vector(fshl_stdar(unsigned(a), unsigned(s), width_z));
  END GENERATE;
SGNED:  IF signd_a /= 0 GENERATE
    z <= std_logic_vector(fshl_stdar(  signed(a), unsigned(s), width_z));
  END GENERATE;
END beh;

--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Wed Jul 21 01:48:05 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_23_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_23_6_64_64_64_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_23_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_23_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_22_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_22_6_64_64_64_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_22_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_22_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_21_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_21_6_64_64_64_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_21_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_21_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_20_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_20_6_64_64_64_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_20_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_20_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_6_64_64_64_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_6_64_64_64_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_6_64_64_64_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_6_64_64_64_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_6_64_64_64_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_6_64_64_64_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_6_64_64_64_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_6_64_64_64_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_6_64_64_64_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_6_64_64_64_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_6_64_64_64_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_6_64_64_64_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    STAGE_MAIN_LOOP_C_3_tr0 : IN STD_LOGIC;
    modExp_dev_while_C_11_tr0 : IN STD_LOGIC;
    STAGE_VEC_LOOP_C_0_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_16_tr0 : IN STD_LOGIC;
    COMP_LOOP_1_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_45_tr0 : IN STD_LOGIC;
    COMP_LOOP_2_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_90_tr0 : IN STD_LOGIC;
    COMP_LOOP_3_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_135_tr0 : IN STD_LOGIC;
    COMP_LOOP_4_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_180_tr0 : IN STD_LOGIC;
    COMP_LOOP_5_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_225_tr0 : IN STD_LOGIC;
    COMP_LOOP_6_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_270_tr0 : IN STD_LOGIC;
    COMP_LOOP_7_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_315_tr0 : IN STD_LOGIC;
    COMP_LOOP_8_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_360_tr0 : IN STD_LOGIC;
    COMP_LOOP_9_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_405_tr0 : IN STD_LOGIC;
    COMP_LOOP_10_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_450_tr0 : IN STD_LOGIC;
    COMP_LOOP_11_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_495_tr0 : IN STD_LOGIC;
    COMP_LOOP_12_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_540_tr0 : IN STD_LOGIC;
    COMP_LOOP_13_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_585_tr0 : IN STD_LOGIC;
    COMP_LOOP_14_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_630_tr0 : IN STD_LOGIC;
    COMP_LOOP_15_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_675_tr0 : IN STD_LOGIC;
    COMP_LOOP_16_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_720_tr0 : IN STD_LOGIC;
    STAGE_VEC_LOOP_C_1_tr0 : IN STD_LOGIC;
    STAGE_MAIN_LOOP_C_4_tr0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_core_core_fsm;

ARCHITECTURE v7 OF inPlaceNTT_DIF_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for inPlaceNTT_DIF_core_core_fsm_1
  TYPE inPlaceNTT_DIF_core_core_fsm_1_ST IS (main_C_0, STAGE_MAIN_LOOP_C_0, STAGE_MAIN_LOOP_C_1,
      STAGE_MAIN_LOOP_C_2, STAGE_MAIN_LOOP_C_3, modExp_dev_while_C_0, modExp_dev_while_C_1,
      modExp_dev_while_C_2, modExp_dev_while_C_3, modExp_dev_while_C_4, modExp_dev_while_C_5,
      modExp_dev_while_C_6, modExp_dev_while_C_7, modExp_dev_while_C_8, modExp_dev_while_C_9,
      modExp_dev_while_C_10, modExp_dev_while_C_11, STAGE_VEC_LOOP_C_0, COMP_LOOP_C_0,
      COMP_LOOP_C_1, COMP_LOOP_C_2, COMP_LOOP_C_3, COMP_LOOP_C_4, COMP_LOOP_C_5,
      COMP_LOOP_C_6, COMP_LOOP_C_7, COMP_LOOP_C_8, COMP_LOOP_C_9, COMP_LOOP_C_10,
      COMP_LOOP_C_11, COMP_LOOP_C_12, COMP_LOOP_C_13, COMP_LOOP_C_14, COMP_LOOP_C_15,
      COMP_LOOP_C_16, COMP_LOOP_1_modExp_dev_1_while_C_0, COMP_LOOP_1_modExp_dev_1_while_C_1,
      COMP_LOOP_1_modExp_dev_1_while_C_2, COMP_LOOP_1_modExp_dev_1_while_C_3, COMP_LOOP_1_modExp_dev_1_while_C_4,
      COMP_LOOP_1_modExp_dev_1_while_C_5, COMP_LOOP_1_modExp_dev_1_while_C_6, COMP_LOOP_1_modExp_dev_1_while_C_7,
      COMP_LOOP_1_modExp_dev_1_while_C_8, COMP_LOOP_1_modExp_dev_1_while_C_9, COMP_LOOP_1_modExp_dev_1_while_C_10,
      COMP_LOOP_1_modExp_dev_1_while_C_11, COMP_LOOP_C_17, COMP_LOOP_C_18, COMP_LOOP_C_19,
      COMP_LOOP_C_20, COMP_LOOP_C_21, COMP_LOOP_C_22, COMP_LOOP_C_23, COMP_LOOP_C_24,
      COMP_LOOP_C_25, COMP_LOOP_C_26, COMP_LOOP_C_27, COMP_LOOP_C_28, COMP_LOOP_C_29,
      COMP_LOOP_C_30, COMP_LOOP_C_31, COMP_LOOP_C_32, COMP_LOOP_C_33, COMP_LOOP_C_34,
      COMP_LOOP_C_35, COMP_LOOP_C_36, COMP_LOOP_C_37, COMP_LOOP_C_38, COMP_LOOP_C_39,
      COMP_LOOP_C_40, COMP_LOOP_C_41, COMP_LOOP_C_42, COMP_LOOP_C_43, COMP_LOOP_C_44,
      COMP_LOOP_C_45, COMP_LOOP_C_46, COMP_LOOP_C_47, COMP_LOOP_C_48, COMP_LOOP_C_49,
      COMP_LOOP_C_50, COMP_LOOP_C_51, COMP_LOOP_C_52, COMP_LOOP_C_53, COMP_LOOP_C_54,
      COMP_LOOP_C_55, COMP_LOOP_C_56, COMP_LOOP_C_57, COMP_LOOP_C_58, COMP_LOOP_C_59,
      COMP_LOOP_C_60, COMP_LOOP_C_61, COMP_LOOP_2_modExp_dev_1_while_C_0, COMP_LOOP_2_modExp_dev_1_while_C_1,
      COMP_LOOP_2_modExp_dev_1_while_C_2, COMP_LOOP_2_modExp_dev_1_while_C_3, COMP_LOOP_2_modExp_dev_1_while_C_4,
      COMP_LOOP_2_modExp_dev_1_while_C_5, COMP_LOOP_2_modExp_dev_1_while_C_6, COMP_LOOP_2_modExp_dev_1_while_C_7,
      COMP_LOOP_2_modExp_dev_1_while_C_8, COMP_LOOP_2_modExp_dev_1_while_C_9, COMP_LOOP_2_modExp_dev_1_while_C_10,
      COMP_LOOP_2_modExp_dev_1_while_C_11, COMP_LOOP_C_62, COMP_LOOP_C_63, COMP_LOOP_C_64,
      COMP_LOOP_C_65, COMP_LOOP_C_66, COMP_LOOP_C_67, COMP_LOOP_C_68, COMP_LOOP_C_69,
      COMP_LOOP_C_70, COMP_LOOP_C_71, COMP_LOOP_C_72, COMP_LOOP_C_73, COMP_LOOP_C_74,
      COMP_LOOP_C_75, COMP_LOOP_C_76, COMP_LOOP_C_77, COMP_LOOP_C_78, COMP_LOOP_C_79,
      COMP_LOOP_C_80, COMP_LOOP_C_81, COMP_LOOP_C_82, COMP_LOOP_C_83, COMP_LOOP_C_84,
      COMP_LOOP_C_85, COMP_LOOP_C_86, COMP_LOOP_C_87, COMP_LOOP_C_88, COMP_LOOP_C_89,
      COMP_LOOP_C_90, COMP_LOOP_C_91, COMP_LOOP_C_92, COMP_LOOP_C_93, COMP_LOOP_C_94,
      COMP_LOOP_C_95, COMP_LOOP_C_96, COMP_LOOP_C_97, COMP_LOOP_C_98, COMP_LOOP_C_99,
      COMP_LOOP_C_100, COMP_LOOP_C_101, COMP_LOOP_C_102, COMP_LOOP_C_103, COMP_LOOP_C_104,
      COMP_LOOP_C_105, COMP_LOOP_C_106, COMP_LOOP_3_modExp_dev_1_while_C_0, COMP_LOOP_3_modExp_dev_1_while_C_1,
      COMP_LOOP_3_modExp_dev_1_while_C_2, COMP_LOOP_3_modExp_dev_1_while_C_3, COMP_LOOP_3_modExp_dev_1_while_C_4,
      COMP_LOOP_3_modExp_dev_1_while_C_5, COMP_LOOP_3_modExp_dev_1_while_C_6, COMP_LOOP_3_modExp_dev_1_while_C_7,
      COMP_LOOP_3_modExp_dev_1_while_C_8, COMP_LOOP_3_modExp_dev_1_while_C_9, COMP_LOOP_3_modExp_dev_1_while_C_10,
      COMP_LOOP_3_modExp_dev_1_while_C_11, COMP_LOOP_C_107, COMP_LOOP_C_108, COMP_LOOP_C_109,
      COMP_LOOP_C_110, COMP_LOOP_C_111, COMP_LOOP_C_112, COMP_LOOP_C_113, COMP_LOOP_C_114,
      COMP_LOOP_C_115, COMP_LOOP_C_116, COMP_LOOP_C_117, COMP_LOOP_C_118, COMP_LOOP_C_119,
      COMP_LOOP_C_120, COMP_LOOP_C_121, COMP_LOOP_C_122, COMP_LOOP_C_123, COMP_LOOP_C_124,
      COMP_LOOP_C_125, COMP_LOOP_C_126, COMP_LOOP_C_127, COMP_LOOP_C_128, COMP_LOOP_C_129,
      COMP_LOOP_C_130, COMP_LOOP_C_131, COMP_LOOP_C_132, COMP_LOOP_C_133, COMP_LOOP_C_134,
      COMP_LOOP_C_135, COMP_LOOP_C_136, COMP_LOOP_C_137, COMP_LOOP_C_138, COMP_LOOP_C_139,
      COMP_LOOP_C_140, COMP_LOOP_C_141, COMP_LOOP_C_142, COMP_LOOP_C_143, COMP_LOOP_C_144,
      COMP_LOOP_C_145, COMP_LOOP_C_146, COMP_LOOP_C_147, COMP_LOOP_C_148, COMP_LOOP_C_149,
      COMP_LOOP_C_150, COMP_LOOP_C_151, COMP_LOOP_4_modExp_dev_1_while_C_0, COMP_LOOP_4_modExp_dev_1_while_C_1,
      COMP_LOOP_4_modExp_dev_1_while_C_2, COMP_LOOP_4_modExp_dev_1_while_C_3, COMP_LOOP_4_modExp_dev_1_while_C_4,
      COMP_LOOP_4_modExp_dev_1_while_C_5, COMP_LOOP_4_modExp_dev_1_while_C_6, COMP_LOOP_4_modExp_dev_1_while_C_7,
      COMP_LOOP_4_modExp_dev_1_while_C_8, COMP_LOOP_4_modExp_dev_1_while_C_9, COMP_LOOP_4_modExp_dev_1_while_C_10,
      COMP_LOOP_4_modExp_dev_1_while_C_11, COMP_LOOP_C_152, COMP_LOOP_C_153, COMP_LOOP_C_154,
      COMP_LOOP_C_155, COMP_LOOP_C_156, COMP_LOOP_C_157, COMP_LOOP_C_158, COMP_LOOP_C_159,
      COMP_LOOP_C_160, COMP_LOOP_C_161, COMP_LOOP_C_162, COMP_LOOP_C_163, COMP_LOOP_C_164,
      COMP_LOOP_C_165, COMP_LOOP_C_166, COMP_LOOP_C_167, COMP_LOOP_C_168, COMP_LOOP_C_169,
      COMP_LOOP_C_170, COMP_LOOP_C_171, COMP_LOOP_C_172, COMP_LOOP_C_173, COMP_LOOP_C_174,
      COMP_LOOP_C_175, COMP_LOOP_C_176, COMP_LOOP_C_177, COMP_LOOP_C_178, COMP_LOOP_C_179,
      COMP_LOOP_C_180, COMP_LOOP_C_181, COMP_LOOP_C_182, COMP_LOOP_C_183, COMP_LOOP_C_184,
      COMP_LOOP_C_185, COMP_LOOP_C_186, COMP_LOOP_C_187, COMP_LOOP_C_188, COMP_LOOP_C_189,
      COMP_LOOP_C_190, COMP_LOOP_C_191, COMP_LOOP_C_192, COMP_LOOP_C_193, COMP_LOOP_C_194,
      COMP_LOOP_C_195, COMP_LOOP_C_196, COMP_LOOP_5_modExp_dev_1_while_C_0, COMP_LOOP_5_modExp_dev_1_while_C_1,
      COMP_LOOP_5_modExp_dev_1_while_C_2, COMP_LOOP_5_modExp_dev_1_while_C_3, COMP_LOOP_5_modExp_dev_1_while_C_4,
      COMP_LOOP_5_modExp_dev_1_while_C_5, COMP_LOOP_5_modExp_dev_1_while_C_6, COMP_LOOP_5_modExp_dev_1_while_C_7,
      COMP_LOOP_5_modExp_dev_1_while_C_8, COMP_LOOP_5_modExp_dev_1_while_C_9, COMP_LOOP_5_modExp_dev_1_while_C_10,
      COMP_LOOP_5_modExp_dev_1_while_C_11, COMP_LOOP_C_197, COMP_LOOP_C_198, COMP_LOOP_C_199,
      COMP_LOOP_C_200, COMP_LOOP_C_201, COMP_LOOP_C_202, COMP_LOOP_C_203, COMP_LOOP_C_204,
      COMP_LOOP_C_205, COMP_LOOP_C_206, COMP_LOOP_C_207, COMP_LOOP_C_208, COMP_LOOP_C_209,
      COMP_LOOP_C_210, COMP_LOOP_C_211, COMP_LOOP_C_212, COMP_LOOP_C_213, COMP_LOOP_C_214,
      COMP_LOOP_C_215, COMP_LOOP_C_216, COMP_LOOP_C_217, COMP_LOOP_C_218, COMP_LOOP_C_219,
      COMP_LOOP_C_220, COMP_LOOP_C_221, COMP_LOOP_C_222, COMP_LOOP_C_223, COMP_LOOP_C_224,
      COMP_LOOP_C_225, COMP_LOOP_C_226, COMP_LOOP_C_227, COMP_LOOP_C_228, COMP_LOOP_C_229,
      COMP_LOOP_C_230, COMP_LOOP_C_231, COMP_LOOP_C_232, COMP_LOOP_C_233, COMP_LOOP_C_234,
      COMP_LOOP_C_235, COMP_LOOP_C_236, COMP_LOOP_C_237, COMP_LOOP_C_238, COMP_LOOP_C_239,
      COMP_LOOP_C_240, COMP_LOOP_C_241, COMP_LOOP_6_modExp_dev_1_while_C_0, COMP_LOOP_6_modExp_dev_1_while_C_1,
      COMP_LOOP_6_modExp_dev_1_while_C_2, COMP_LOOP_6_modExp_dev_1_while_C_3, COMP_LOOP_6_modExp_dev_1_while_C_4,
      COMP_LOOP_6_modExp_dev_1_while_C_5, COMP_LOOP_6_modExp_dev_1_while_C_6, COMP_LOOP_6_modExp_dev_1_while_C_7,
      COMP_LOOP_6_modExp_dev_1_while_C_8, COMP_LOOP_6_modExp_dev_1_while_C_9, COMP_LOOP_6_modExp_dev_1_while_C_10,
      COMP_LOOP_6_modExp_dev_1_while_C_11, COMP_LOOP_C_242, COMP_LOOP_C_243, COMP_LOOP_C_244,
      COMP_LOOP_C_245, COMP_LOOP_C_246, COMP_LOOP_C_247, COMP_LOOP_C_248, COMP_LOOP_C_249,
      COMP_LOOP_C_250, COMP_LOOP_C_251, COMP_LOOP_C_252, COMP_LOOP_C_253, COMP_LOOP_C_254,
      COMP_LOOP_C_255, COMP_LOOP_C_256, COMP_LOOP_C_257, COMP_LOOP_C_258, COMP_LOOP_C_259,
      COMP_LOOP_C_260, COMP_LOOP_C_261, COMP_LOOP_C_262, COMP_LOOP_C_263, COMP_LOOP_C_264,
      COMP_LOOP_C_265, COMP_LOOP_C_266, COMP_LOOP_C_267, COMP_LOOP_C_268, COMP_LOOP_C_269,
      COMP_LOOP_C_270, COMP_LOOP_C_271, COMP_LOOP_C_272, COMP_LOOP_C_273, COMP_LOOP_C_274,
      COMP_LOOP_C_275, COMP_LOOP_C_276, COMP_LOOP_C_277, COMP_LOOP_C_278, COMP_LOOP_C_279,
      COMP_LOOP_C_280, COMP_LOOP_C_281, COMP_LOOP_C_282, COMP_LOOP_C_283, COMP_LOOP_C_284,
      COMP_LOOP_C_285, COMP_LOOP_C_286, COMP_LOOP_7_modExp_dev_1_while_C_0, COMP_LOOP_7_modExp_dev_1_while_C_1,
      COMP_LOOP_7_modExp_dev_1_while_C_2, COMP_LOOP_7_modExp_dev_1_while_C_3, COMP_LOOP_7_modExp_dev_1_while_C_4,
      COMP_LOOP_7_modExp_dev_1_while_C_5, COMP_LOOP_7_modExp_dev_1_while_C_6, COMP_LOOP_7_modExp_dev_1_while_C_7,
      COMP_LOOP_7_modExp_dev_1_while_C_8, COMP_LOOP_7_modExp_dev_1_while_C_9, COMP_LOOP_7_modExp_dev_1_while_C_10,
      COMP_LOOP_7_modExp_dev_1_while_C_11, COMP_LOOP_C_287, COMP_LOOP_C_288, COMP_LOOP_C_289,
      COMP_LOOP_C_290, COMP_LOOP_C_291, COMP_LOOP_C_292, COMP_LOOP_C_293, COMP_LOOP_C_294,
      COMP_LOOP_C_295, COMP_LOOP_C_296, COMP_LOOP_C_297, COMP_LOOP_C_298, COMP_LOOP_C_299,
      COMP_LOOP_C_300, COMP_LOOP_C_301, COMP_LOOP_C_302, COMP_LOOP_C_303, COMP_LOOP_C_304,
      COMP_LOOP_C_305, COMP_LOOP_C_306, COMP_LOOP_C_307, COMP_LOOP_C_308, COMP_LOOP_C_309,
      COMP_LOOP_C_310, COMP_LOOP_C_311, COMP_LOOP_C_312, COMP_LOOP_C_313, COMP_LOOP_C_314,
      COMP_LOOP_C_315, COMP_LOOP_C_316, COMP_LOOP_C_317, COMP_LOOP_C_318, COMP_LOOP_C_319,
      COMP_LOOP_C_320, COMP_LOOP_C_321, COMP_LOOP_C_322, COMP_LOOP_C_323, COMP_LOOP_C_324,
      COMP_LOOP_C_325, COMP_LOOP_C_326, COMP_LOOP_C_327, COMP_LOOP_C_328, COMP_LOOP_C_329,
      COMP_LOOP_C_330, COMP_LOOP_C_331, COMP_LOOP_8_modExp_dev_1_while_C_0, COMP_LOOP_8_modExp_dev_1_while_C_1,
      COMP_LOOP_8_modExp_dev_1_while_C_2, COMP_LOOP_8_modExp_dev_1_while_C_3, COMP_LOOP_8_modExp_dev_1_while_C_4,
      COMP_LOOP_8_modExp_dev_1_while_C_5, COMP_LOOP_8_modExp_dev_1_while_C_6, COMP_LOOP_8_modExp_dev_1_while_C_7,
      COMP_LOOP_8_modExp_dev_1_while_C_8, COMP_LOOP_8_modExp_dev_1_while_C_9, COMP_LOOP_8_modExp_dev_1_while_C_10,
      COMP_LOOP_8_modExp_dev_1_while_C_11, COMP_LOOP_C_332, COMP_LOOP_C_333, COMP_LOOP_C_334,
      COMP_LOOP_C_335, COMP_LOOP_C_336, COMP_LOOP_C_337, COMP_LOOP_C_338, COMP_LOOP_C_339,
      COMP_LOOP_C_340, COMP_LOOP_C_341, COMP_LOOP_C_342, COMP_LOOP_C_343, COMP_LOOP_C_344,
      COMP_LOOP_C_345, COMP_LOOP_C_346, COMP_LOOP_C_347, COMP_LOOP_C_348, COMP_LOOP_C_349,
      COMP_LOOP_C_350, COMP_LOOP_C_351, COMP_LOOP_C_352, COMP_LOOP_C_353, COMP_LOOP_C_354,
      COMP_LOOP_C_355, COMP_LOOP_C_356, COMP_LOOP_C_357, COMP_LOOP_C_358, COMP_LOOP_C_359,
      COMP_LOOP_C_360, COMP_LOOP_C_361, COMP_LOOP_C_362, COMP_LOOP_C_363, COMP_LOOP_C_364,
      COMP_LOOP_C_365, COMP_LOOP_C_366, COMP_LOOP_C_367, COMP_LOOP_C_368, COMP_LOOP_C_369,
      COMP_LOOP_C_370, COMP_LOOP_C_371, COMP_LOOP_C_372, COMP_LOOP_C_373, COMP_LOOP_C_374,
      COMP_LOOP_C_375, COMP_LOOP_C_376, COMP_LOOP_9_modExp_dev_1_while_C_0, COMP_LOOP_9_modExp_dev_1_while_C_1,
      COMP_LOOP_9_modExp_dev_1_while_C_2, COMP_LOOP_9_modExp_dev_1_while_C_3, COMP_LOOP_9_modExp_dev_1_while_C_4,
      COMP_LOOP_9_modExp_dev_1_while_C_5, COMP_LOOP_9_modExp_dev_1_while_C_6, COMP_LOOP_9_modExp_dev_1_while_C_7,
      COMP_LOOP_9_modExp_dev_1_while_C_8, COMP_LOOP_9_modExp_dev_1_while_C_9, COMP_LOOP_9_modExp_dev_1_while_C_10,
      COMP_LOOP_9_modExp_dev_1_while_C_11, COMP_LOOP_C_377, COMP_LOOP_C_378, COMP_LOOP_C_379,
      COMP_LOOP_C_380, COMP_LOOP_C_381, COMP_LOOP_C_382, COMP_LOOP_C_383, COMP_LOOP_C_384,
      COMP_LOOP_C_385, COMP_LOOP_C_386, COMP_LOOP_C_387, COMP_LOOP_C_388, COMP_LOOP_C_389,
      COMP_LOOP_C_390, COMP_LOOP_C_391, COMP_LOOP_C_392, COMP_LOOP_C_393, COMP_LOOP_C_394,
      COMP_LOOP_C_395, COMP_LOOP_C_396, COMP_LOOP_C_397, COMP_LOOP_C_398, COMP_LOOP_C_399,
      COMP_LOOP_C_400, COMP_LOOP_C_401, COMP_LOOP_C_402, COMP_LOOP_C_403, COMP_LOOP_C_404,
      COMP_LOOP_C_405, COMP_LOOP_C_406, COMP_LOOP_C_407, COMP_LOOP_C_408, COMP_LOOP_C_409,
      COMP_LOOP_C_410, COMP_LOOP_C_411, COMP_LOOP_C_412, COMP_LOOP_C_413, COMP_LOOP_C_414,
      COMP_LOOP_C_415, COMP_LOOP_C_416, COMP_LOOP_C_417, COMP_LOOP_C_418, COMP_LOOP_C_419,
      COMP_LOOP_C_420, COMP_LOOP_C_421, COMP_LOOP_10_modExp_dev_1_while_C_0, COMP_LOOP_10_modExp_dev_1_while_C_1,
      COMP_LOOP_10_modExp_dev_1_while_C_2, COMP_LOOP_10_modExp_dev_1_while_C_3, COMP_LOOP_10_modExp_dev_1_while_C_4,
      COMP_LOOP_10_modExp_dev_1_while_C_5, COMP_LOOP_10_modExp_dev_1_while_C_6, COMP_LOOP_10_modExp_dev_1_while_C_7,
      COMP_LOOP_10_modExp_dev_1_while_C_8, COMP_LOOP_10_modExp_dev_1_while_C_9, COMP_LOOP_10_modExp_dev_1_while_C_10,
      COMP_LOOP_10_modExp_dev_1_while_C_11, COMP_LOOP_C_422, COMP_LOOP_C_423, COMP_LOOP_C_424,
      COMP_LOOP_C_425, COMP_LOOP_C_426, COMP_LOOP_C_427, COMP_LOOP_C_428, COMP_LOOP_C_429,
      COMP_LOOP_C_430, COMP_LOOP_C_431, COMP_LOOP_C_432, COMP_LOOP_C_433, COMP_LOOP_C_434,
      COMP_LOOP_C_435, COMP_LOOP_C_436, COMP_LOOP_C_437, COMP_LOOP_C_438, COMP_LOOP_C_439,
      COMP_LOOP_C_440, COMP_LOOP_C_441, COMP_LOOP_C_442, COMP_LOOP_C_443, COMP_LOOP_C_444,
      COMP_LOOP_C_445, COMP_LOOP_C_446, COMP_LOOP_C_447, COMP_LOOP_C_448, COMP_LOOP_C_449,
      COMP_LOOP_C_450, COMP_LOOP_C_451, COMP_LOOP_C_452, COMP_LOOP_C_453, COMP_LOOP_C_454,
      COMP_LOOP_C_455, COMP_LOOP_C_456, COMP_LOOP_C_457, COMP_LOOP_C_458, COMP_LOOP_C_459,
      COMP_LOOP_C_460, COMP_LOOP_C_461, COMP_LOOP_C_462, COMP_LOOP_C_463, COMP_LOOP_C_464,
      COMP_LOOP_C_465, COMP_LOOP_C_466, COMP_LOOP_11_modExp_dev_1_while_C_0, COMP_LOOP_11_modExp_dev_1_while_C_1,
      COMP_LOOP_11_modExp_dev_1_while_C_2, COMP_LOOP_11_modExp_dev_1_while_C_3, COMP_LOOP_11_modExp_dev_1_while_C_4,
      COMP_LOOP_11_modExp_dev_1_while_C_5, COMP_LOOP_11_modExp_dev_1_while_C_6, COMP_LOOP_11_modExp_dev_1_while_C_7,
      COMP_LOOP_11_modExp_dev_1_while_C_8, COMP_LOOP_11_modExp_dev_1_while_C_9, COMP_LOOP_11_modExp_dev_1_while_C_10,
      COMP_LOOP_11_modExp_dev_1_while_C_11, COMP_LOOP_C_467, COMP_LOOP_C_468, COMP_LOOP_C_469,
      COMP_LOOP_C_470, COMP_LOOP_C_471, COMP_LOOP_C_472, COMP_LOOP_C_473, COMP_LOOP_C_474,
      COMP_LOOP_C_475, COMP_LOOP_C_476, COMP_LOOP_C_477, COMP_LOOP_C_478, COMP_LOOP_C_479,
      COMP_LOOP_C_480, COMP_LOOP_C_481, COMP_LOOP_C_482, COMP_LOOP_C_483, COMP_LOOP_C_484,
      COMP_LOOP_C_485, COMP_LOOP_C_486, COMP_LOOP_C_487, COMP_LOOP_C_488, COMP_LOOP_C_489,
      COMP_LOOP_C_490, COMP_LOOP_C_491, COMP_LOOP_C_492, COMP_LOOP_C_493, COMP_LOOP_C_494,
      COMP_LOOP_C_495, COMP_LOOP_C_496, COMP_LOOP_C_497, COMP_LOOP_C_498, COMP_LOOP_C_499,
      COMP_LOOP_C_500, COMP_LOOP_C_501, COMP_LOOP_C_502, COMP_LOOP_C_503, COMP_LOOP_C_504,
      COMP_LOOP_C_505, COMP_LOOP_C_506, COMP_LOOP_C_507, COMP_LOOP_C_508, COMP_LOOP_C_509,
      COMP_LOOP_C_510, COMP_LOOP_C_511, COMP_LOOP_12_modExp_dev_1_while_C_0, COMP_LOOP_12_modExp_dev_1_while_C_1,
      COMP_LOOP_12_modExp_dev_1_while_C_2, COMP_LOOP_12_modExp_dev_1_while_C_3, COMP_LOOP_12_modExp_dev_1_while_C_4,
      COMP_LOOP_12_modExp_dev_1_while_C_5, COMP_LOOP_12_modExp_dev_1_while_C_6, COMP_LOOP_12_modExp_dev_1_while_C_7,
      COMP_LOOP_12_modExp_dev_1_while_C_8, COMP_LOOP_12_modExp_dev_1_while_C_9, COMP_LOOP_12_modExp_dev_1_while_C_10,
      COMP_LOOP_12_modExp_dev_1_while_C_11, COMP_LOOP_C_512, COMP_LOOP_C_513, COMP_LOOP_C_514,
      COMP_LOOP_C_515, COMP_LOOP_C_516, COMP_LOOP_C_517, COMP_LOOP_C_518, COMP_LOOP_C_519,
      COMP_LOOP_C_520, COMP_LOOP_C_521, COMP_LOOP_C_522, COMP_LOOP_C_523, COMP_LOOP_C_524,
      COMP_LOOP_C_525, COMP_LOOP_C_526, COMP_LOOP_C_527, COMP_LOOP_C_528, COMP_LOOP_C_529,
      COMP_LOOP_C_530, COMP_LOOP_C_531, COMP_LOOP_C_532, COMP_LOOP_C_533, COMP_LOOP_C_534,
      COMP_LOOP_C_535, COMP_LOOP_C_536, COMP_LOOP_C_537, COMP_LOOP_C_538, COMP_LOOP_C_539,
      COMP_LOOP_C_540, COMP_LOOP_C_541, COMP_LOOP_C_542, COMP_LOOP_C_543, COMP_LOOP_C_544,
      COMP_LOOP_C_545, COMP_LOOP_C_546, COMP_LOOP_C_547, COMP_LOOP_C_548, COMP_LOOP_C_549,
      COMP_LOOP_C_550, COMP_LOOP_C_551, COMP_LOOP_C_552, COMP_LOOP_C_553, COMP_LOOP_C_554,
      COMP_LOOP_C_555, COMP_LOOP_C_556, COMP_LOOP_13_modExp_dev_1_while_C_0, COMP_LOOP_13_modExp_dev_1_while_C_1,
      COMP_LOOP_13_modExp_dev_1_while_C_2, COMP_LOOP_13_modExp_dev_1_while_C_3, COMP_LOOP_13_modExp_dev_1_while_C_4,
      COMP_LOOP_13_modExp_dev_1_while_C_5, COMP_LOOP_13_modExp_dev_1_while_C_6, COMP_LOOP_13_modExp_dev_1_while_C_7,
      COMP_LOOP_13_modExp_dev_1_while_C_8, COMP_LOOP_13_modExp_dev_1_while_C_9, COMP_LOOP_13_modExp_dev_1_while_C_10,
      COMP_LOOP_13_modExp_dev_1_while_C_11, COMP_LOOP_C_557, COMP_LOOP_C_558, COMP_LOOP_C_559,
      COMP_LOOP_C_560, COMP_LOOP_C_561, COMP_LOOP_C_562, COMP_LOOP_C_563, COMP_LOOP_C_564,
      COMP_LOOP_C_565, COMP_LOOP_C_566, COMP_LOOP_C_567, COMP_LOOP_C_568, COMP_LOOP_C_569,
      COMP_LOOP_C_570, COMP_LOOP_C_571, COMP_LOOP_C_572, COMP_LOOP_C_573, COMP_LOOP_C_574,
      COMP_LOOP_C_575, COMP_LOOP_C_576, COMP_LOOP_C_577, COMP_LOOP_C_578, COMP_LOOP_C_579,
      COMP_LOOP_C_580, COMP_LOOP_C_581, COMP_LOOP_C_582, COMP_LOOP_C_583, COMP_LOOP_C_584,
      COMP_LOOP_C_585, COMP_LOOP_C_586, COMP_LOOP_C_587, COMP_LOOP_C_588, COMP_LOOP_C_589,
      COMP_LOOP_C_590, COMP_LOOP_C_591, COMP_LOOP_C_592, COMP_LOOP_C_593, COMP_LOOP_C_594,
      COMP_LOOP_C_595, COMP_LOOP_C_596, COMP_LOOP_C_597, COMP_LOOP_C_598, COMP_LOOP_C_599,
      COMP_LOOP_C_600, COMP_LOOP_C_601, COMP_LOOP_14_modExp_dev_1_while_C_0, COMP_LOOP_14_modExp_dev_1_while_C_1,
      COMP_LOOP_14_modExp_dev_1_while_C_2, COMP_LOOP_14_modExp_dev_1_while_C_3, COMP_LOOP_14_modExp_dev_1_while_C_4,
      COMP_LOOP_14_modExp_dev_1_while_C_5, COMP_LOOP_14_modExp_dev_1_while_C_6, COMP_LOOP_14_modExp_dev_1_while_C_7,
      COMP_LOOP_14_modExp_dev_1_while_C_8, COMP_LOOP_14_modExp_dev_1_while_C_9, COMP_LOOP_14_modExp_dev_1_while_C_10,
      COMP_LOOP_14_modExp_dev_1_while_C_11, COMP_LOOP_C_602, COMP_LOOP_C_603, COMP_LOOP_C_604,
      COMP_LOOP_C_605, COMP_LOOP_C_606, COMP_LOOP_C_607, COMP_LOOP_C_608, COMP_LOOP_C_609,
      COMP_LOOP_C_610, COMP_LOOP_C_611, COMP_LOOP_C_612, COMP_LOOP_C_613, COMP_LOOP_C_614,
      COMP_LOOP_C_615, COMP_LOOP_C_616, COMP_LOOP_C_617, COMP_LOOP_C_618, COMP_LOOP_C_619,
      COMP_LOOP_C_620, COMP_LOOP_C_621, COMP_LOOP_C_622, COMP_LOOP_C_623, COMP_LOOP_C_624,
      COMP_LOOP_C_625, COMP_LOOP_C_626, COMP_LOOP_C_627, COMP_LOOP_C_628, COMP_LOOP_C_629,
      COMP_LOOP_C_630, COMP_LOOP_C_631, COMP_LOOP_C_632, COMP_LOOP_C_633, COMP_LOOP_C_634,
      COMP_LOOP_C_635, COMP_LOOP_C_636, COMP_LOOP_C_637, COMP_LOOP_C_638, COMP_LOOP_C_639,
      COMP_LOOP_C_640, COMP_LOOP_C_641, COMP_LOOP_C_642, COMP_LOOP_C_643, COMP_LOOP_C_644,
      COMP_LOOP_C_645, COMP_LOOP_C_646, COMP_LOOP_15_modExp_dev_1_while_C_0, COMP_LOOP_15_modExp_dev_1_while_C_1,
      COMP_LOOP_15_modExp_dev_1_while_C_2, COMP_LOOP_15_modExp_dev_1_while_C_3, COMP_LOOP_15_modExp_dev_1_while_C_4,
      COMP_LOOP_15_modExp_dev_1_while_C_5, COMP_LOOP_15_modExp_dev_1_while_C_6, COMP_LOOP_15_modExp_dev_1_while_C_7,
      COMP_LOOP_15_modExp_dev_1_while_C_8, COMP_LOOP_15_modExp_dev_1_while_C_9, COMP_LOOP_15_modExp_dev_1_while_C_10,
      COMP_LOOP_15_modExp_dev_1_while_C_11, COMP_LOOP_C_647, COMP_LOOP_C_648, COMP_LOOP_C_649,
      COMP_LOOP_C_650, COMP_LOOP_C_651, COMP_LOOP_C_652, COMP_LOOP_C_653, COMP_LOOP_C_654,
      COMP_LOOP_C_655, COMP_LOOP_C_656, COMP_LOOP_C_657, COMP_LOOP_C_658, COMP_LOOP_C_659,
      COMP_LOOP_C_660, COMP_LOOP_C_661, COMP_LOOP_C_662, COMP_LOOP_C_663, COMP_LOOP_C_664,
      COMP_LOOP_C_665, COMP_LOOP_C_666, COMP_LOOP_C_667, COMP_LOOP_C_668, COMP_LOOP_C_669,
      COMP_LOOP_C_670, COMP_LOOP_C_671, COMP_LOOP_C_672, COMP_LOOP_C_673, COMP_LOOP_C_674,
      COMP_LOOP_C_675, COMP_LOOP_C_676, COMP_LOOP_C_677, COMP_LOOP_C_678, COMP_LOOP_C_679,
      COMP_LOOP_C_680, COMP_LOOP_C_681, COMP_LOOP_C_682, COMP_LOOP_C_683, COMP_LOOP_C_684,
      COMP_LOOP_C_685, COMP_LOOP_C_686, COMP_LOOP_C_687, COMP_LOOP_C_688, COMP_LOOP_C_689,
      COMP_LOOP_C_690, COMP_LOOP_C_691, COMP_LOOP_16_modExp_dev_1_while_C_0, COMP_LOOP_16_modExp_dev_1_while_C_1,
      COMP_LOOP_16_modExp_dev_1_while_C_2, COMP_LOOP_16_modExp_dev_1_while_C_3, COMP_LOOP_16_modExp_dev_1_while_C_4,
      COMP_LOOP_16_modExp_dev_1_while_C_5, COMP_LOOP_16_modExp_dev_1_while_C_6, COMP_LOOP_16_modExp_dev_1_while_C_7,
      COMP_LOOP_16_modExp_dev_1_while_C_8, COMP_LOOP_16_modExp_dev_1_while_C_9, COMP_LOOP_16_modExp_dev_1_while_C_10,
      COMP_LOOP_16_modExp_dev_1_while_C_11, COMP_LOOP_C_692, COMP_LOOP_C_693, COMP_LOOP_C_694,
      COMP_LOOP_C_695, COMP_LOOP_C_696, COMP_LOOP_C_697, COMP_LOOP_C_698, COMP_LOOP_C_699,
      COMP_LOOP_C_700, COMP_LOOP_C_701, COMP_LOOP_C_702, COMP_LOOP_C_703, COMP_LOOP_C_704,
      COMP_LOOP_C_705, COMP_LOOP_C_706, COMP_LOOP_C_707, COMP_LOOP_C_708, COMP_LOOP_C_709,
      COMP_LOOP_C_710, COMP_LOOP_C_711, COMP_LOOP_C_712, COMP_LOOP_C_713, COMP_LOOP_C_714,
      COMP_LOOP_C_715, COMP_LOOP_C_716, COMP_LOOP_C_717, COMP_LOOP_C_718, COMP_LOOP_C_719,
      COMP_LOOP_C_720, STAGE_VEC_LOOP_C_1, STAGE_MAIN_LOOP_C_4, main_C_1);

  SIGNAL state_var : inPlaceNTT_DIF_core_core_fsm_1_ST;
  SIGNAL state_var_NS : inPlaceNTT_DIF_core_core_fsm_1_ST;

BEGIN
  inPlaceNTT_DIF_core_core_fsm_1 : PROCESS (STAGE_MAIN_LOOP_C_3_tr0, modExp_dev_while_C_11_tr0,
      STAGE_VEC_LOOP_C_0_tr0, COMP_LOOP_C_16_tr0, COMP_LOOP_1_modExp_dev_1_while_C_11_tr0,
      COMP_LOOP_C_45_tr0, COMP_LOOP_2_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_90_tr0,
      COMP_LOOP_3_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_135_tr0, COMP_LOOP_4_modExp_dev_1_while_C_11_tr0,
      COMP_LOOP_C_180_tr0, COMP_LOOP_5_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_225_tr0,
      COMP_LOOP_6_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_270_tr0, COMP_LOOP_7_modExp_dev_1_while_C_11_tr0,
      COMP_LOOP_C_315_tr0, COMP_LOOP_8_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_360_tr0,
      COMP_LOOP_9_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_405_tr0, COMP_LOOP_10_modExp_dev_1_while_C_11_tr0,
      COMP_LOOP_C_450_tr0, COMP_LOOP_11_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_495_tr0,
      COMP_LOOP_12_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_540_tr0, COMP_LOOP_13_modExp_dev_1_while_C_11_tr0,
      COMP_LOOP_C_585_tr0, COMP_LOOP_14_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_630_tr0,
      COMP_LOOP_15_modExp_dev_1_while_C_11_tr0, COMP_LOOP_C_675_tr0, COMP_LOOP_16_modExp_dev_1_while_C_11_tr0,
      COMP_LOOP_C_720_tr0, STAGE_VEC_LOOP_C_1_tr0, STAGE_MAIN_LOOP_C_4_tr0, state_var)
  BEGIN
    CASE state_var IS
      WHEN STAGE_MAIN_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000001");
        state_var_NS <= STAGE_MAIN_LOOP_C_1;
      WHEN STAGE_MAIN_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000010");
        state_var_NS <= STAGE_MAIN_LOOP_C_2;
      WHEN STAGE_MAIN_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000011");
        state_var_NS <= STAGE_MAIN_LOOP_C_3;
      WHEN STAGE_MAIN_LOOP_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000100");
        IF ( STAGE_MAIN_LOOP_C_3_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_0;
        ELSE
          state_var_NS <= modExp_dev_while_C_0;
        END IF;
      WHEN modExp_dev_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000101");
        state_var_NS <= modExp_dev_while_C_1;
      WHEN modExp_dev_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000110");
        state_var_NS <= modExp_dev_while_C_2;
      WHEN modExp_dev_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000111");
        state_var_NS <= modExp_dev_while_C_3;
      WHEN modExp_dev_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001000");
        state_var_NS <= modExp_dev_while_C_4;
      WHEN modExp_dev_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001001");
        state_var_NS <= modExp_dev_while_C_5;
      WHEN modExp_dev_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001010");
        state_var_NS <= modExp_dev_while_C_6;
      WHEN modExp_dev_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001011");
        state_var_NS <= modExp_dev_while_C_7;
      WHEN modExp_dev_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001100");
        state_var_NS <= modExp_dev_while_C_8;
      WHEN modExp_dev_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001101");
        state_var_NS <= modExp_dev_while_C_9;
      WHEN modExp_dev_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001110");
        state_var_NS <= modExp_dev_while_C_10;
      WHEN modExp_dev_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001111");
        state_var_NS <= modExp_dev_while_C_11;
      WHEN modExp_dev_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010000");
        IF ( modExp_dev_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_0;
        ELSE
          state_var_NS <= modExp_dev_while_C_0;
        END IF;
      WHEN STAGE_VEC_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010001");
        IF ( STAGE_VEC_LOOP_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN COMP_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010010");
        state_var_NS <= COMP_LOOP_C_1;
      WHEN COMP_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010011");
        state_var_NS <= COMP_LOOP_C_2;
      WHEN COMP_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010100");
        state_var_NS <= COMP_LOOP_C_3;
      WHEN COMP_LOOP_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010101");
        state_var_NS <= COMP_LOOP_C_4;
      WHEN COMP_LOOP_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010110");
        state_var_NS <= COMP_LOOP_C_5;
      WHEN COMP_LOOP_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010111");
        state_var_NS <= COMP_LOOP_C_6;
      WHEN COMP_LOOP_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011000");
        state_var_NS <= COMP_LOOP_C_7;
      WHEN COMP_LOOP_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011001");
        state_var_NS <= COMP_LOOP_C_8;
      WHEN COMP_LOOP_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011010");
        state_var_NS <= COMP_LOOP_C_9;
      WHEN COMP_LOOP_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011011");
        state_var_NS <= COMP_LOOP_C_10;
      WHEN COMP_LOOP_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011100");
        state_var_NS <= COMP_LOOP_C_11;
      WHEN COMP_LOOP_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011101");
        state_var_NS <= COMP_LOOP_C_12;
      WHEN COMP_LOOP_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011110");
        state_var_NS <= COMP_LOOP_C_13;
      WHEN COMP_LOOP_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011111");
        state_var_NS <= COMP_LOOP_C_14;
      WHEN COMP_LOOP_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100000");
        state_var_NS <= COMP_LOOP_C_15;
      WHEN COMP_LOOP_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100001");
        state_var_NS <= COMP_LOOP_C_16;
      WHEN COMP_LOOP_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100010");
        IF ( COMP_LOOP_C_16_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_17;
        ELSE
          state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100011");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100100");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100101");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100110");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100111");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101000");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101001");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101010");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101011");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101100");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101101");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101110");
        IF ( COMP_LOOP_1_modExp_dev_1_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_17;
        ELSE
          state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101111");
        state_var_NS <= COMP_LOOP_C_18;
      WHEN COMP_LOOP_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110000");
        state_var_NS <= COMP_LOOP_C_19;
      WHEN COMP_LOOP_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110001");
        state_var_NS <= COMP_LOOP_C_20;
      WHEN COMP_LOOP_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110010");
        state_var_NS <= COMP_LOOP_C_21;
      WHEN COMP_LOOP_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110011");
        state_var_NS <= COMP_LOOP_C_22;
      WHEN COMP_LOOP_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110100");
        state_var_NS <= COMP_LOOP_C_23;
      WHEN COMP_LOOP_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110101");
        state_var_NS <= COMP_LOOP_C_24;
      WHEN COMP_LOOP_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110110");
        state_var_NS <= COMP_LOOP_C_25;
      WHEN COMP_LOOP_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110111");
        state_var_NS <= COMP_LOOP_C_26;
      WHEN COMP_LOOP_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111000");
        state_var_NS <= COMP_LOOP_C_27;
      WHEN COMP_LOOP_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111001");
        state_var_NS <= COMP_LOOP_C_28;
      WHEN COMP_LOOP_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111010");
        state_var_NS <= COMP_LOOP_C_29;
      WHEN COMP_LOOP_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111011");
        state_var_NS <= COMP_LOOP_C_30;
      WHEN COMP_LOOP_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111100");
        state_var_NS <= COMP_LOOP_C_31;
      WHEN COMP_LOOP_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111101");
        state_var_NS <= COMP_LOOP_C_32;
      WHEN COMP_LOOP_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111110");
        state_var_NS <= COMP_LOOP_C_33;
      WHEN COMP_LOOP_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111111");
        state_var_NS <= COMP_LOOP_C_34;
      WHEN COMP_LOOP_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000000");
        state_var_NS <= COMP_LOOP_C_35;
      WHEN COMP_LOOP_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000001");
        state_var_NS <= COMP_LOOP_C_36;
      WHEN COMP_LOOP_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000010");
        state_var_NS <= COMP_LOOP_C_37;
      WHEN COMP_LOOP_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000011");
        state_var_NS <= COMP_LOOP_C_38;
      WHEN COMP_LOOP_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000100");
        state_var_NS <= COMP_LOOP_C_39;
      WHEN COMP_LOOP_C_39 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000101");
        state_var_NS <= COMP_LOOP_C_40;
      WHEN COMP_LOOP_C_40 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000110");
        state_var_NS <= COMP_LOOP_C_41;
      WHEN COMP_LOOP_C_41 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000111");
        state_var_NS <= COMP_LOOP_C_42;
      WHEN COMP_LOOP_C_42 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001000");
        state_var_NS <= COMP_LOOP_C_43;
      WHEN COMP_LOOP_C_43 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001001");
        state_var_NS <= COMP_LOOP_C_44;
      WHEN COMP_LOOP_C_44 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001010");
        state_var_NS <= COMP_LOOP_C_45;
      WHEN COMP_LOOP_C_45 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001011");
        IF ( COMP_LOOP_C_45_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_46;
        END IF;
      WHEN COMP_LOOP_C_46 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001100");
        state_var_NS <= COMP_LOOP_C_47;
      WHEN COMP_LOOP_C_47 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001101");
        state_var_NS <= COMP_LOOP_C_48;
      WHEN COMP_LOOP_C_48 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001110");
        state_var_NS <= COMP_LOOP_C_49;
      WHEN COMP_LOOP_C_49 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001111");
        state_var_NS <= COMP_LOOP_C_50;
      WHEN COMP_LOOP_C_50 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010000");
        state_var_NS <= COMP_LOOP_C_51;
      WHEN COMP_LOOP_C_51 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010001");
        state_var_NS <= COMP_LOOP_C_52;
      WHEN COMP_LOOP_C_52 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010010");
        state_var_NS <= COMP_LOOP_C_53;
      WHEN COMP_LOOP_C_53 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010011");
        state_var_NS <= COMP_LOOP_C_54;
      WHEN COMP_LOOP_C_54 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010100");
        state_var_NS <= COMP_LOOP_C_55;
      WHEN COMP_LOOP_C_55 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010101");
        state_var_NS <= COMP_LOOP_C_56;
      WHEN COMP_LOOP_C_56 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010110");
        state_var_NS <= COMP_LOOP_C_57;
      WHEN COMP_LOOP_C_57 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010111");
        state_var_NS <= COMP_LOOP_C_58;
      WHEN COMP_LOOP_C_58 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011000");
        state_var_NS <= COMP_LOOP_C_59;
      WHEN COMP_LOOP_C_59 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011001");
        state_var_NS <= COMP_LOOP_C_60;
      WHEN COMP_LOOP_C_60 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011010");
        state_var_NS <= COMP_LOOP_C_61;
      WHEN COMP_LOOP_C_61 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011011");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011100");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011101");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011110");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011111");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100000");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100001");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100010");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100011");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100100");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100101");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100110");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100111");
        IF ( COMP_LOOP_2_modExp_dev_1_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_62;
        ELSE
          state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_62 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101000");
        state_var_NS <= COMP_LOOP_C_63;
      WHEN COMP_LOOP_C_63 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101001");
        state_var_NS <= COMP_LOOP_C_64;
      WHEN COMP_LOOP_C_64 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101010");
        state_var_NS <= COMP_LOOP_C_65;
      WHEN COMP_LOOP_C_65 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101011");
        state_var_NS <= COMP_LOOP_C_66;
      WHEN COMP_LOOP_C_66 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101100");
        state_var_NS <= COMP_LOOP_C_67;
      WHEN COMP_LOOP_C_67 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101101");
        state_var_NS <= COMP_LOOP_C_68;
      WHEN COMP_LOOP_C_68 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101110");
        state_var_NS <= COMP_LOOP_C_69;
      WHEN COMP_LOOP_C_69 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101111");
        state_var_NS <= COMP_LOOP_C_70;
      WHEN COMP_LOOP_C_70 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110000");
        state_var_NS <= COMP_LOOP_C_71;
      WHEN COMP_LOOP_C_71 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110001");
        state_var_NS <= COMP_LOOP_C_72;
      WHEN COMP_LOOP_C_72 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110010");
        state_var_NS <= COMP_LOOP_C_73;
      WHEN COMP_LOOP_C_73 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110011");
        state_var_NS <= COMP_LOOP_C_74;
      WHEN COMP_LOOP_C_74 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110100");
        state_var_NS <= COMP_LOOP_C_75;
      WHEN COMP_LOOP_C_75 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110101");
        state_var_NS <= COMP_LOOP_C_76;
      WHEN COMP_LOOP_C_76 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110110");
        state_var_NS <= COMP_LOOP_C_77;
      WHEN COMP_LOOP_C_77 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110111");
        state_var_NS <= COMP_LOOP_C_78;
      WHEN COMP_LOOP_C_78 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111000");
        state_var_NS <= COMP_LOOP_C_79;
      WHEN COMP_LOOP_C_79 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111001");
        state_var_NS <= COMP_LOOP_C_80;
      WHEN COMP_LOOP_C_80 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111010");
        state_var_NS <= COMP_LOOP_C_81;
      WHEN COMP_LOOP_C_81 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111011");
        state_var_NS <= COMP_LOOP_C_82;
      WHEN COMP_LOOP_C_82 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111100");
        state_var_NS <= COMP_LOOP_C_83;
      WHEN COMP_LOOP_C_83 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111101");
        state_var_NS <= COMP_LOOP_C_84;
      WHEN COMP_LOOP_C_84 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111110");
        state_var_NS <= COMP_LOOP_C_85;
      WHEN COMP_LOOP_C_85 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111111");
        state_var_NS <= COMP_LOOP_C_86;
      WHEN COMP_LOOP_C_86 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000000");
        state_var_NS <= COMP_LOOP_C_87;
      WHEN COMP_LOOP_C_87 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000001");
        state_var_NS <= COMP_LOOP_C_88;
      WHEN COMP_LOOP_C_88 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000010");
        state_var_NS <= COMP_LOOP_C_89;
      WHEN COMP_LOOP_C_89 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000011");
        state_var_NS <= COMP_LOOP_C_90;
      WHEN COMP_LOOP_C_90 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000100");
        IF ( COMP_LOOP_C_90_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_91;
        END IF;
      WHEN COMP_LOOP_C_91 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000101");
        state_var_NS <= COMP_LOOP_C_92;
      WHEN COMP_LOOP_C_92 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000110");
        state_var_NS <= COMP_LOOP_C_93;
      WHEN COMP_LOOP_C_93 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000111");
        state_var_NS <= COMP_LOOP_C_94;
      WHEN COMP_LOOP_C_94 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001000");
        state_var_NS <= COMP_LOOP_C_95;
      WHEN COMP_LOOP_C_95 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001001");
        state_var_NS <= COMP_LOOP_C_96;
      WHEN COMP_LOOP_C_96 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001010");
        state_var_NS <= COMP_LOOP_C_97;
      WHEN COMP_LOOP_C_97 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001011");
        state_var_NS <= COMP_LOOP_C_98;
      WHEN COMP_LOOP_C_98 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001100");
        state_var_NS <= COMP_LOOP_C_99;
      WHEN COMP_LOOP_C_99 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001101");
        state_var_NS <= COMP_LOOP_C_100;
      WHEN COMP_LOOP_C_100 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001110");
        state_var_NS <= COMP_LOOP_C_101;
      WHEN COMP_LOOP_C_101 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001111");
        state_var_NS <= COMP_LOOP_C_102;
      WHEN COMP_LOOP_C_102 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010000");
        state_var_NS <= COMP_LOOP_C_103;
      WHEN COMP_LOOP_C_103 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010001");
        state_var_NS <= COMP_LOOP_C_104;
      WHEN COMP_LOOP_C_104 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010010");
        state_var_NS <= COMP_LOOP_C_105;
      WHEN COMP_LOOP_C_105 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010011");
        state_var_NS <= COMP_LOOP_C_106;
      WHEN COMP_LOOP_C_106 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010100");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010101");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010110");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010111");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011000");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011001");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011010");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011011");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011100");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011101");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011110");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011111");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100000");
        IF ( COMP_LOOP_3_modExp_dev_1_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_107;
        ELSE
          state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_107 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100001");
        state_var_NS <= COMP_LOOP_C_108;
      WHEN COMP_LOOP_C_108 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100010");
        state_var_NS <= COMP_LOOP_C_109;
      WHEN COMP_LOOP_C_109 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100011");
        state_var_NS <= COMP_LOOP_C_110;
      WHEN COMP_LOOP_C_110 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100100");
        state_var_NS <= COMP_LOOP_C_111;
      WHEN COMP_LOOP_C_111 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100101");
        state_var_NS <= COMP_LOOP_C_112;
      WHEN COMP_LOOP_C_112 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100110");
        state_var_NS <= COMP_LOOP_C_113;
      WHEN COMP_LOOP_C_113 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100111");
        state_var_NS <= COMP_LOOP_C_114;
      WHEN COMP_LOOP_C_114 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101000");
        state_var_NS <= COMP_LOOP_C_115;
      WHEN COMP_LOOP_C_115 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101001");
        state_var_NS <= COMP_LOOP_C_116;
      WHEN COMP_LOOP_C_116 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101010");
        state_var_NS <= COMP_LOOP_C_117;
      WHEN COMP_LOOP_C_117 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101011");
        state_var_NS <= COMP_LOOP_C_118;
      WHEN COMP_LOOP_C_118 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101100");
        state_var_NS <= COMP_LOOP_C_119;
      WHEN COMP_LOOP_C_119 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101101");
        state_var_NS <= COMP_LOOP_C_120;
      WHEN COMP_LOOP_C_120 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101110");
        state_var_NS <= COMP_LOOP_C_121;
      WHEN COMP_LOOP_C_121 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101111");
        state_var_NS <= COMP_LOOP_C_122;
      WHEN COMP_LOOP_C_122 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110000");
        state_var_NS <= COMP_LOOP_C_123;
      WHEN COMP_LOOP_C_123 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110001");
        state_var_NS <= COMP_LOOP_C_124;
      WHEN COMP_LOOP_C_124 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110010");
        state_var_NS <= COMP_LOOP_C_125;
      WHEN COMP_LOOP_C_125 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110011");
        state_var_NS <= COMP_LOOP_C_126;
      WHEN COMP_LOOP_C_126 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110100");
        state_var_NS <= COMP_LOOP_C_127;
      WHEN COMP_LOOP_C_127 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110101");
        state_var_NS <= COMP_LOOP_C_128;
      WHEN COMP_LOOP_C_128 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110110");
        state_var_NS <= COMP_LOOP_C_129;
      WHEN COMP_LOOP_C_129 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110111");
        state_var_NS <= COMP_LOOP_C_130;
      WHEN COMP_LOOP_C_130 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111000");
        state_var_NS <= COMP_LOOP_C_131;
      WHEN COMP_LOOP_C_131 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111001");
        state_var_NS <= COMP_LOOP_C_132;
      WHEN COMP_LOOP_C_132 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111010");
        state_var_NS <= COMP_LOOP_C_133;
      WHEN COMP_LOOP_C_133 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111011");
        state_var_NS <= COMP_LOOP_C_134;
      WHEN COMP_LOOP_C_134 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111100");
        state_var_NS <= COMP_LOOP_C_135;
      WHEN COMP_LOOP_C_135 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111101");
        IF ( COMP_LOOP_C_135_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_136;
        END IF;
      WHEN COMP_LOOP_C_136 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111110");
        state_var_NS <= COMP_LOOP_C_137;
      WHEN COMP_LOOP_C_137 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111111");
        state_var_NS <= COMP_LOOP_C_138;
      WHEN COMP_LOOP_C_138 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000000");
        state_var_NS <= COMP_LOOP_C_139;
      WHEN COMP_LOOP_C_139 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000001");
        state_var_NS <= COMP_LOOP_C_140;
      WHEN COMP_LOOP_C_140 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000010");
        state_var_NS <= COMP_LOOP_C_141;
      WHEN COMP_LOOP_C_141 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000011");
        state_var_NS <= COMP_LOOP_C_142;
      WHEN COMP_LOOP_C_142 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000100");
        state_var_NS <= COMP_LOOP_C_143;
      WHEN COMP_LOOP_C_143 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000101");
        state_var_NS <= COMP_LOOP_C_144;
      WHEN COMP_LOOP_C_144 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000110");
        state_var_NS <= COMP_LOOP_C_145;
      WHEN COMP_LOOP_C_145 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000111");
        state_var_NS <= COMP_LOOP_C_146;
      WHEN COMP_LOOP_C_146 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001000");
        state_var_NS <= COMP_LOOP_C_147;
      WHEN COMP_LOOP_C_147 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001001");
        state_var_NS <= COMP_LOOP_C_148;
      WHEN COMP_LOOP_C_148 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001010");
        state_var_NS <= COMP_LOOP_C_149;
      WHEN COMP_LOOP_C_149 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001011");
        state_var_NS <= COMP_LOOP_C_150;
      WHEN COMP_LOOP_C_150 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001100");
        state_var_NS <= COMP_LOOP_C_151;
      WHEN COMP_LOOP_C_151 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001101");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001110");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001111");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010000");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010001");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010010");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010011");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010100");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010101");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010110");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010111");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011000");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011001");
        IF ( COMP_LOOP_4_modExp_dev_1_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_152;
        ELSE
          state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_152 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011010");
        state_var_NS <= COMP_LOOP_C_153;
      WHEN COMP_LOOP_C_153 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011011");
        state_var_NS <= COMP_LOOP_C_154;
      WHEN COMP_LOOP_C_154 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011100");
        state_var_NS <= COMP_LOOP_C_155;
      WHEN COMP_LOOP_C_155 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011101");
        state_var_NS <= COMP_LOOP_C_156;
      WHEN COMP_LOOP_C_156 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011110");
        state_var_NS <= COMP_LOOP_C_157;
      WHEN COMP_LOOP_C_157 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011111");
        state_var_NS <= COMP_LOOP_C_158;
      WHEN COMP_LOOP_C_158 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100000");
        state_var_NS <= COMP_LOOP_C_159;
      WHEN COMP_LOOP_C_159 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100001");
        state_var_NS <= COMP_LOOP_C_160;
      WHEN COMP_LOOP_C_160 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100010");
        state_var_NS <= COMP_LOOP_C_161;
      WHEN COMP_LOOP_C_161 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100011");
        state_var_NS <= COMP_LOOP_C_162;
      WHEN COMP_LOOP_C_162 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100100");
        state_var_NS <= COMP_LOOP_C_163;
      WHEN COMP_LOOP_C_163 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100101");
        state_var_NS <= COMP_LOOP_C_164;
      WHEN COMP_LOOP_C_164 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100110");
        state_var_NS <= COMP_LOOP_C_165;
      WHEN COMP_LOOP_C_165 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100111");
        state_var_NS <= COMP_LOOP_C_166;
      WHEN COMP_LOOP_C_166 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101000");
        state_var_NS <= COMP_LOOP_C_167;
      WHEN COMP_LOOP_C_167 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101001");
        state_var_NS <= COMP_LOOP_C_168;
      WHEN COMP_LOOP_C_168 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101010");
        state_var_NS <= COMP_LOOP_C_169;
      WHEN COMP_LOOP_C_169 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101011");
        state_var_NS <= COMP_LOOP_C_170;
      WHEN COMP_LOOP_C_170 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101100");
        state_var_NS <= COMP_LOOP_C_171;
      WHEN COMP_LOOP_C_171 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101101");
        state_var_NS <= COMP_LOOP_C_172;
      WHEN COMP_LOOP_C_172 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101110");
        state_var_NS <= COMP_LOOP_C_173;
      WHEN COMP_LOOP_C_173 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101111");
        state_var_NS <= COMP_LOOP_C_174;
      WHEN COMP_LOOP_C_174 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110000");
        state_var_NS <= COMP_LOOP_C_175;
      WHEN COMP_LOOP_C_175 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110001");
        state_var_NS <= COMP_LOOP_C_176;
      WHEN COMP_LOOP_C_176 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110010");
        state_var_NS <= COMP_LOOP_C_177;
      WHEN COMP_LOOP_C_177 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110011");
        state_var_NS <= COMP_LOOP_C_178;
      WHEN COMP_LOOP_C_178 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110100");
        state_var_NS <= COMP_LOOP_C_179;
      WHEN COMP_LOOP_C_179 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110101");
        state_var_NS <= COMP_LOOP_C_180;
      WHEN COMP_LOOP_C_180 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110110");
        IF ( COMP_LOOP_C_180_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_181;
        END IF;
      WHEN COMP_LOOP_C_181 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110111");
        state_var_NS <= COMP_LOOP_C_182;
      WHEN COMP_LOOP_C_182 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111000");
        state_var_NS <= COMP_LOOP_C_183;
      WHEN COMP_LOOP_C_183 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111001");
        state_var_NS <= COMP_LOOP_C_184;
      WHEN COMP_LOOP_C_184 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111010");
        state_var_NS <= COMP_LOOP_C_185;
      WHEN COMP_LOOP_C_185 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111011");
        state_var_NS <= COMP_LOOP_C_186;
      WHEN COMP_LOOP_C_186 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111100");
        state_var_NS <= COMP_LOOP_C_187;
      WHEN COMP_LOOP_C_187 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111101");
        state_var_NS <= COMP_LOOP_C_188;
      WHEN COMP_LOOP_C_188 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111110");
        state_var_NS <= COMP_LOOP_C_189;
      WHEN COMP_LOOP_C_189 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111111");
        state_var_NS <= COMP_LOOP_C_190;
      WHEN COMP_LOOP_C_190 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000000");
        state_var_NS <= COMP_LOOP_C_191;
      WHEN COMP_LOOP_C_191 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000001");
        state_var_NS <= COMP_LOOP_C_192;
      WHEN COMP_LOOP_C_192 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000010");
        state_var_NS <= COMP_LOOP_C_193;
      WHEN COMP_LOOP_C_193 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000011");
        state_var_NS <= COMP_LOOP_C_194;
      WHEN COMP_LOOP_C_194 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000100");
        state_var_NS <= COMP_LOOP_C_195;
      WHEN COMP_LOOP_C_195 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000101");
        state_var_NS <= COMP_LOOP_C_196;
      WHEN COMP_LOOP_C_196 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000110");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000111");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001000");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001001");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001010");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001011");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001100");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001101");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001110");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001111");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010000");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010001");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010010");
        IF ( COMP_LOOP_5_modExp_dev_1_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_197;
        ELSE
          state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_197 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010011");
        state_var_NS <= COMP_LOOP_C_198;
      WHEN COMP_LOOP_C_198 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010100");
        state_var_NS <= COMP_LOOP_C_199;
      WHEN COMP_LOOP_C_199 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010101");
        state_var_NS <= COMP_LOOP_C_200;
      WHEN COMP_LOOP_C_200 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010110");
        state_var_NS <= COMP_LOOP_C_201;
      WHEN COMP_LOOP_C_201 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010111");
        state_var_NS <= COMP_LOOP_C_202;
      WHEN COMP_LOOP_C_202 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011000");
        state_var_NS <= COMP_LOOP_C_203;
      WHEN COMP_LOOP_C_203 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011001");
        state_var_NS <= COMP_LOOP_C_204;
      WHEN COMP_LOOP_C_204 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011010");
        state_var_NS <= COMP_LOOP_C_205;
      WHEN COMP_LOOP_C_205 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011011");
        state_var_NS <= COMP_LOOP_C_206;
      WHEN COMP_LOOP_C_206 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011100");
        state_var_NS <= COMP_LOOP_C_207;
      WHEN COMP_LOOP_C_207 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011101");
        state_var_NS <= COMP_LOOP_C_208;
      WHEN COMP_LOOP_C_208 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011110");
        state_var_NS <= COMP_LOOP_C_209;
      WHEN COMP_LOOP_C_209 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011111");
        state_var_NS <= COMP_LOOP_C_210;
      WHEN COMP_LOOP_C_210 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100000");
        state_var_NS <= COMP_LOOP_C_211;
      WHEN COMP_LOOP_C_211 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100001");
        state_var_NS <= COMP_LOOP_C_212;
      WHEN COMP_LOOP_C_212 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100010");
        state_var_NS <= COMP_LOOP_C_213;
      WHEN COMP_LOOP_C_213 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100011");
        state_var_NS <= COMP_LOOP_C_214;
      WHEN COMP_LOOP_C_214 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100100");
        state_var_NS <= COMP_LOOP_C_215;
      WHEN COMP_LOOP_C_215 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100101");
        state_var_NS <= COMP_LOOP_C_216;
      WHEN COMP_LOOP_C_216 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100110");
        state_var_NS <= COMP_LOOP_C_217;
      WHEN COMP_LOOP_C_217 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100111");
        state_var_NS <= COMP_LOOP_C_218;
      WHEN COMP_LOOP_C_218 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101000");
        state_var_NS <= COMP_LOOP_C_219;
      WHEN COMP_LOOP_C_219 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101001");
        state_var_NS <= COMP_LOOP_C_220;
      WHEN COMP_LOOP_C_220 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101010");
        state_var_NS <= COMP_LOOP_C_221;
      WHEN COMP_LOOP_C_221 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101011");
        state_var_NS <= COMP_LOOP_C_222;
      WHEN COMP_LOOP_C_222 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101100");
        state_var_NS <= COMP_LOOP_C_223;
      WHEN COMP_LOOP_C_223 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101101");
        state_var_NS <= COMP_LOOP_C_224;
      WHEN COMP_LOOP_C_224 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101110");
        state_var_NS <= COMP_LOOP_C_225;
      WHEN COMP_LOOP_C_225 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101111");
        IF ( COMP_LOOP_C_225_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_226;
        END IF;
      WHEN COMP_LOOP_C_226 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110000");
        state_var_NS <= COMP_LOOP_C_227;
      WHEN COMP_LOOP_C_227 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110001");
        state_var_NS <= COMP_LOOP_C_228;
      WHEN COMP_LOOP_C_228 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110010");
        state_var_NS <= COMP_LOOP_C_229;
      WHEN COMP_LOOP_C_229 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110011");
        state_var_NS <= COMP_LOOP_C_230;
      WHEN COMP_LOOP_C_230 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110100");
        state_var_NS <= COMP_LOOP_C_231;
      WHEN COMP_LOOP_C_231 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110101");
        state_var_NS <= COMP_LOOP_C_232;
      WHEN COMP_LOOP_C_232 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110110");
        state_var_NS <= COMP_LOOP_C_233;
      WHEN COMP_LOOP_C_233 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110111");
        state_var_NS <= COMP_LOOP_C_234;
      WHEN COMP_LOOP_C_234 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111000");
        state_var_NS <= COMP_LOOP_C_235;
      WHEN COMP_LOOP_C_235 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111001");
        state_var_NS <= COMP_LOOP_C_236;
      WHEN COMP_LOOP_C_236 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111010");
        state_var_NS <= COMP_LOOP_C_237;
      WHEN COMP_LOOP_C_237 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111011");
        state_var_NS <= COMP_LOOP_C_238;
      WHEN COMP_LOOP_C_238 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111100");
        state_var_NS <= COMP_LOOP_C_239;
      WHEN COMP_LOOP_C_239 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111101");
        state_var_NS <= COMP_LOOP_C_240;
      WHEN COMP_LOOP_C_240 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111110");
        state_var_NS <= COMP_LOOP_C_241;
      WHEN COMP_LOOP_C_241 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111111");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000000");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000001");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000010");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000011");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000100");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000101");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000110");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000111");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001000");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001001");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001010");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001011");
        IF ( COMP_LOOP_6_modExp_dev_1_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_242;
        ELSE
          state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_242 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001100");
        state_var_NS <= COMP_LOOP_C_243;
      WHEN COMP_LOOP_C_243 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001101");
        state_var_NS <= COMP_LOOP_C_244;
      WHEN COMP_LOOP_C_244 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001110");
        state_var_NS <= COMP_LOOP_C_245;
      WHEN COMP_LOOP_C_245 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001111");
        state_var_NS <= COMP_LOOP_C_246;
      WHEN COMP_LOOP_C_246 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010000");
        state_var_NS <= COMP_LOOP_C_247;
      WHEN COMP_LOOP_C_247 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010001");
        state_var_NS <= COMP_LOOP_C_248;
      WHEN COMP_LOOP_C_248 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010010");
        state_var_NS <= COMP_LOOP_C_249;
      WHEN COMP_LOOP_C_249 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010011");
        state_var_NS <= COMP_LOOP_C_250;
      WHEN COMP_LOOP_C_250 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010100");
        state_var_NS <= COMP_LOOP_C_251;
      WHEN COMP_LOOP_C_251 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010101");
        state_var_NS <= COMP_LOOP_C_252;
      WHEN COMP_LOOP_C_252 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010110");
        state_var_NS <= COMP_LOOP_C_253;
      WHEN COMP_LOOP_C_253 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010111");
        state_var_NS <= COMP_LOOP_C_254;
      WHEN COMP_LOOP_C_254 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011000");
        state_var_NS <= COMP_LOOP_C_255;
      WHEN COMP_LOOP_C_255 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011001");
        state_var_NS <= COMP_LOOP_C_256;
      WHEN COMP_LOOP_C_256 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011010");
        state_var_NS <= COMP_LOOP_C_257;
      WHEN COMP_LOOP_C_257 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011011");
        state_var_NS <= COMP_LOOP_C_258;
      WHEN COMP_LOOP_C_258 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011100");
        state_var_NS <= COMP_LOOP_C_259;
      WHEN COMP_LOOP_C_259 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011101");
        state_var_NS <= COMP_LOOP_C_260;
      WHEN COMP_LOOP_C_260 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011110");
        state_var_NS <= COMP_LOOP_C_261;
      WHEN COMP_LOOP_C_261 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011111");
        state_var_NS <= COMP_LOOP_C_262;
      WHEN COMP_LOOP_C_262 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100000");
        state_var_NS <= COMP_LOOP_C_263;
      WHEN COMP_LOOP_C_263 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100001");
        state_var_NS <= COMP_LOOP_C_264;
      WHEN COMP_LOOP_C_264 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100010");
        state_var_NS <= COMP_LOOP_C_265;
      WHEN COMP_LOOP_C_265 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100011");
        state_var_NS <= COMP_LOOP_C_266;
      WHEN COMP_LOOP_C_266 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100100");
        state_var_NS <= COMP_LOOP_C_267;
      WHEN COMP_LOOP_C_267 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100101");
        state_var_NS <= COMP_LOOP_C_268;
      WHEN COMP_LOOP_C_268 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100110");
        state_var_NS <= COMP_LOOP_C_269;
      WHEN COMP_LOOP_C_269 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100111");
        state_var_NS <= COMP_LOOP_C_270;
      WHEN COMP_LOOP_C_270 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101000");
        IF ( COMP_LOOP_C_270_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_271;
        END IF;
      WHEN COMP_LOOP_C_271 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101001");
        state_var_NS <= COMP_LOOP_C_272;
      WHEN COMP_LOOP_C_272 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101010");
        state_var_NS <= COMP_LOOP_C_273;
      WHEN COMP_LOOP_C_273 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101011");
        state_var_NS <= COMP_LOOP_C_274;
      WHEN COMP_LOOP_C_274 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101100");
        state_var_NS <= COMP_LOOP_C_275;
      WHEN COMP_LOOP_C_275 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101101");
        state_var_NS <= COMP_LOOP_C_276;
      WHEN COMP_LOOP_C_276 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101110");
        state_var_NS <= COMP_LOOP_C_277;
      WHEN COMP_LOOP_C_277 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101111");
        state_var_NS <= COMP_LOOP_C_278;
      WHEN COMP_LOOP_C_278 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110000");
        state_var_NS <= COMP_LOOP_C_279;
      WHEN COMP_LOOP_C_279 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110001");
        state_var_NS <= COMP_LOOP_C_280;
      WHEN COMP_LOOP_C_280 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110010");
        state_var_NS <= COMP_LOOP_C_281;
      WHEN COMP_LOOP_C_281 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110011");
        state_var_NS <= COMP_LOOP_C_282;
      WHEN COMP_LOOP_C_282 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110100");
        state_var_NS <= COMP_LOOP_C_283;
      WHEN COMP_LOOP_C_283 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110101");
        state_var_NS <= COMP_LOOP_C_284;
      WHEN COMP_LOOP_C_284 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110110");
        state_var_NS <= COMP_LOOP_C_285;
      WHEN COMP_LOOP_C_285 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110111");
        state_var_NS <= COMP_LOOP_C_286;
      WHEN COMP_LOOP_C_286 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111000");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111001");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111010");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111011");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111100");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111101");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111110");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111111");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000000");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000001");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000010");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000011");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000100");
        IF ( COMP_LOOP_7_modExp_dev_1_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_287;
        ELSE
          state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_287 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000101");
        state_var_NS <= COMP_LOOP_C_288;
      WHEN COMP_LOOP_C_288 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000110");
        state_var_NS <= COMP_LOOP_C_289;
      WHEN COMP_LOOP_C_289 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000111");
        state_var_NS <= COMP_LOOP_C_290;
      WHEN COMP_LOOP_C_290 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001000");
        state_var_NS <= COMP_LOOP_C_291;
      WHEN COMP_LOOP_C_291 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001001");
        state_var_NS <= COMP_LOOP_C_292;
      WHEN COMP_LOOP_C_292 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001010");
        state_var_NS <= COMP_LOOP_C_293;
      WHEN COMP_LOOP_C_293 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001011");
        state_var_NS <= COMP_LOOP_C_294;
      WHEN COMP_LOOP_C_294 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001100");
        state_var_NS <= COMP_LOOP_C_295;
      WHEN COMP_LOOP_C_295 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001101");
        state_var_NS <= COMP_LOOP_C_296;
      WHEN COMP_LOOP_C_296 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001110");
        state_var_NS <= COMP_LOOP_C_297;
      WHEN COMP_LOOP_C_297 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001111");
        state_var_NS <= COMP_LOOP_C_298;
      WHEN COMP_LOOP_C_298 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010000");
        state_var_NS <= COMP_LOOP_C_299;
      WHEN COMP_LOOP_C_299 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010001");
        state_var_NS <= COMP_LOOP_C_300;
      WHEN COMP_LOOP_C_300 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010010");
        state_var_NS <= COMP_LOOP_C_301;
      WHEN COMP_LOOP_C_301 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010011");
        state_var_NS <= COMP_LOOP_C_302;
      WHEN COMP_LOOP_C_302 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010100");
        state_var_NS <= COMP_LOOP_C_303;
      WHEN COMP_LOOP_C_303 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010101");
        state_var_NS <= COMP_LOOP_C_304;
      WHEN COMP_LOOP_C_304 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010110");
        state_var_NS <= COMP_LOOP_C_305;
      WHEN COMP_LOOP_C_305 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010111");
        state_var_NS <= COMP_LOOP_C_306;
      WHEN COMP_LOOP_C_306 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011000");
        state_var_NS <= COMP_LOOP_C_307;
      WHEN COMP_LOOP_C_307 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011001");
        state_var_NS <= COMP_LOOP_C_308;
      WHEN COMP_LOOP_C_308 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011010");
        state_var_NS <= COMP_LOOP_C_309;
      WHEN COMP_LOOP_C_309 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011011");
        state_var_NS <= COMP_LOOP_C_310;
      WHEN COMP_LOOP_C_310 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011100");
        state_var_NS <= COMP_LOOP_C_311;
      WHEN COMP_LOOP_C_311 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011101");
        state_var_NS <= COMP_LOOP_C_312;
      WHEN COMP_LOOP_C_312 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011110");
        state_var_NS <= COMP_LOOP_C_313;
      WHEN COMP_LOOP_C_313 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011111");
        state_var_NS <= COMP_LOOP_C_314;
      WHEN COMP_LOOP_C_314 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100000");
        state_var_NS <= COMP_LOOP_C_315;
      WHEN COMP_LOOP_C_315 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100001");
        IF ( COMP_LOOP_C_315_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_316;
        END IF;
      WHEN COMP_LOOP_C_316 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100010");
        state_var_NS <= COMP_LOOP_C_317;
      WHEN COMP_LOOP_C_317 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100011");
        state_var_NS <= COMP_LOOP_C_318;
      WHEN COMP_LOOP_C_318 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100100");
        state_var_NS <= COMP_LOOP_C_319;
      WHEN COMP_LOOP_C_319 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100101");
        state_var_NS <= COMP_LOOP_C_320;
      WHEN COMP_LOOP_C_320 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100110");
        state_var_NS <= COMP_LOOP_C_321;
      WHEN COMP_LOOP_C_321 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100111");
        state_var_NS <= COMP_LOOP_C_322;
      WHEN COMP_LOOP_C_322 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101000");
        state_var_NS <= COMP_LOOP_C_323;
      WHEN COMP_LOOP_C_323 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101001");
        state_var_NS <= COMP_LOOP_C_324;
      WHEN COMP_LOOP_C_324 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101010");
        state_var_NS <= COMP_LOOP_C_325;
      WHEN COMP_LOOP_C_325 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101011");
        state_var_NS <= COMP_LOOP_C_326;
      WHEN COMP_LOOP_C_326 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101100");
        state_var_NS <= COMP_LOOP_C_327;
      WHEN COMP_LOOP_C_327 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101101");
        state_var_NS <= COMP_LOOP_C_328;
      WHEN COMP_LOOP_C_328 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101110");
        state_var_NS <= COMP_LOOP_C_329;
      WHEN COMP_LOOP_C_329 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101111");
        state_var_NS <= COMP_LOOP_C_330;
      WHEN COMP_LOOP_C_330 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110000");
        state_var_NS <= COMP_LOOP_C_331;
      WHEN COMP_LOOP_C_331 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110001");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110010");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110011");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110100");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110101");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110110");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110111");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111000");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111001");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111010");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111011");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111100");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111101");
        IF ( COMP_LOOP_8_modExp_dev_1_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_332;
        ELSE
          state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_332 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111110");
        state_var_NS <= COMP_LOOP_C_333;
      WHEN COMP_LOOP_C_333 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111111");
        state_var_NS <= COMP_LOOP_C_334;
      WHEN COMP_LOOP_C_334 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000000");
        state_var_NS <= COMP_LOOP_C_335;
      WHEN COMP_LOOP_C_335 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000001");
        state_var_NS <= COMP_LOOP_C_336;
      WHEN COMP_LOOP_C_336 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000010");
        state_var_NS <= COMP_LOOP_C_337;
      WHEN COMP_LOOP_C_337 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000011");
        state_var_NS <= COMP_LOOP_C_338;
      WHEN COMP_LOOP_C_338 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000100");
        state_var_NS <= COMP_LOOP_C_339;
      WHEN COMP_LOOP_C_339 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000101");
        state_var_NS <= COMP_LOOP_C_340;
      WHEN COMP_LOOP_C_340 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000110");
        state_var_NS <= COMP_LOOP_C_341;
      WHEN COMP_LOOP_C_341 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000111");
        state_var_NS <= COMP_LOOP_C_342;
      WHEN COMP_LOOP_C_342 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001000");
        state_var_NS <= COMP_LOOP_C_343;
      WHEN COMP_LOOP_C_343 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001001");
        state_var_NS <= COMP_LOOP_C_344;
      WHEN COMP_LOOP_C_344 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001010");
        state_var_NS <= COMP_LOOP_C_345;
      WHEN COMP_LOOP_C_345 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001011");
        state_var_NS <= COMP_LOOP_C_346;
      WHEN COMP_LOOP_C_346 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001100");
        state_var_NS <= COMP_LOOP_C_347;
      WHEN COMP_LOOP_C_347 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001101");
        state_var_NS <= COMP_LOOP_C_348;
      WHEN COMP_LOOP_C_348 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001110");
        state_var_NS <= COMP_LOOP_C_349;
      WHEN COMP_LOOP_C_349 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001111");
        state_var_NS <= COMP_LOOP_C_350;
      WHEN COMP_LOOP_C_350 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010000");
        state_var_NS <= COMP_LOOP_C_351;
      WHEN COMP_LOOP_C_351 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010001");
        state_var_NS <= COMP_LOOP_C_352;
      WHEN COMP_LOOP_C_352 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010010");
        state_var_NS <= COMP_LOOP_C_353;
      WHEN COMP_LOOP_C_353 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010011");
        state_var_NS <= COMP_LOOP_C_354;
      WHEN COMP_LOOP_C_354 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010100");
        state_var_NS <= COMP_LOOP_C_355;
      WHEN COMP_LOOP_C_355 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010101");
        state_var_NS <= COMP_LOOP_C_356;
      WHEN COMP_LOOP_C_356 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010110");
        state_var_NS <= COMP_LOOP_C_357;
      WHEN COMP_LOOP_C_357 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010111");
        state_var_NS <= COMP_LOOP_C_358;
      WHEN COMP_LOOP_C_358 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011000");
        state_var_NS <= COMP_LOOP_C_359;
      WHEN COMP_LOOP_C_359 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011001");
        state_var_NS <= COMP_LOOP_C_360;
      WHEN COMP_LOOP_C_360 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011010");
        IF ( COMP_LOOP_C_360_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_361;
        END IF;
      WHEN COMP_LOOP_C_361 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011011");
        state_var_NS <= COMP_LOOP_C_362;
      WHEN COMP_LOOP_C_362 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011100");
        state_var_NS <= COMP_LOOP_C_363;
      WHEN COMP_LOOP_C_363 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011101");
        state_var_NS <= COMP_LOOP_C_364;
      WHEN COMP_LOOP_C_364 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011110");
        state_var_NS <= COMP_LOOP_C_365;
      WHEN COMP_LOOP_C_365 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011111");
        state_var_NS <= COMP_LOOP_C_366;
      WHEN COMP_LOOP_C_366 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100000");
        state_var_NS <= COMP_LOOP_C_367;
      WHEN COMP_LOOP_C_367 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100001");
        state_var_NS <= COMP_LOOP_C_368;
      WHEN COMP_LOOP_C_368 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100010");
        state_var_NS <= COMP_LOOP_C_369;
      WHEN COMP_LOOP_C_369 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100011");
        state_var_NS <= COMP_LOOP_C_370;
      WHEN COMP_LOOP_C_370 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100100");
        state_var_NS <= COMP_LOOP_C_371;
      WHEN COMP_LOOP_C_371 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100101");
        state_var_NS <= COMP_LOOP_C_372;
      WHEN COMP_LOOP_C_372 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100110");
        state_var_NS <= COMP_LOOP_C_373;
      WHEN COMP_LOOP_C_373 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100111");
        state_var_NS <= COMP_LOOP_C_374;
      WHEN COMP_LOOP_C_374 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101000");
        state_var_NS <= COMP_LOOP_C_375;
      WHEN COMP_LOOP_C_375 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101001");
        state_var_NS <= COMP_LOOP_C_376;
      WHEN COMP_LOOP_C_376 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101010");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101011");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101100");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101101");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101110");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101111");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110000");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110001");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110010");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110011");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110100");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110101");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110110");
        IF ( COMP_LOOP_9_modExp_dev_1_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_377;
        ELSE
          state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_377 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110111");
        state_var_NS <= COMP_LOOP_C_378;
      WHEN COMP_LOOP_C_378 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111000");
        state_var_NS <= COMP_LOOP_C_379;
      WHEN COMP_LOOP_C_379 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111001");
        state_var_NS <= COMP_LOOP_C_380;
      WHEN COMP_LOOP_C_380 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111010");
        state_var_NS <= COMP_LOOP_C_381;
      WHEN COMP_LOOP_C_381 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111011");
        state_var_NS <= COMP_LOOP_C_382;
      WHEN COMP_LOOP_C_382 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111100");
        state_var_NS <= COMP_LOOP_C_383;
      WHEN COMP_LOOP_C_383 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111101");
        state_var_NS <= COMP_LOOP_C_384;
      WHEN COMP_LOOP_C_384 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111110");
        state_var_NS <= COMP_LOOP_C_385;
      WHEN COMP_LOOP_C_385 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111111");
        state_var_NS <= COMP_LOOP_C_386;
      WHEN COMP_LOOP_C_386 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000000");
        state_var_NS <= COMP_LOOP_C_387;
      WHEN COMP_LOOP_C_387 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000001");
        state_var_NS <= COMP_LOOP_C_388;
      WHEN COMP_LOOP_C_388 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000010");
        state_var_NS <= COMP_LOOP_C_389;
      WHEN COMP_LOOP_C_389 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000011");
        state_var_NS <= COMP_LOOP_C_390;
      WHEN COMP_LOOP_C_390 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000100");
        state_var_NS <= COMP_LOOP_C_391;
      WHEN COMP_LOOP_C_391 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000101");
        state_var_NS <= COMP_LOOP_C_392;
      WHEN COMP_LOOP_C_392 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000110");
        state_var_NS <= COMP_LOOP_C_393;
      WHEN COMP_LOOP_C_393 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000111");
        state_var_NS <= COMP_LOOP_C_394;
      WHEN COMP_LOOP_C_394 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001000");
        state_var_NS <= COMP_LOOP_C_395;
      WHEN COMP_LOOP_C_395 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001001");
        state_var_NS <= COMP_LOOP_C_396;
      WHEN COMP_LOOP_C_396 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001010");
        state_var_NS <= COMP_LOOP_C_397;
      WHEN COMP_LOOP_C_397 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001011");
        state_var_NS <= COMP_LOOP_C_398;
      WHEN COMP_LOOP_C_398 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001100");
        state_var_NS <= COMP_LOOP_C_399;
      WHEN COMP_LOOP_C_399 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001101");
        state_var_NS <= COMP_LOOP_C_400;
      WHEN COMP_LOOP_C_400 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001110");
        state_var_NS <= COMP_LOOP_C_401;
      WHEN COMP_LOOP_C_401 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001111");
        state_var_NS <= COMP_LOOP_C_402;
      WHEN COMP_LOOP_C_402 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010000");
        state_var_NS <= COMP_LOOP_C_403;
      WHEN COMP_LOOP_C_403 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010001");
        state_var_NS <= COMP_LOOP_C_404;
      WHEN COMP_LOOP_C_404 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010010");
        state_var_NS <= COMP_LOOP_C_405;
      WHEN COMP_LOOP_C_405 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010011");
        IF ( COMP_LOOP_C_405_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_406;
        END IF;
      WHEN COMP_LOOP_C_406 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010100");
        state_var_NS <= COMP_LOOP_C_407;
      WHEN COMP_LOOP_C_407 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010101");
        state_var_NS <= COMP_LOOP_C_408;
      WHEN COMP_LOOP_C_408 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010110");
        state_var_NS <= COMP_LOOP_C_409;
      WHEN COMP_LOOP_C_409 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010111");
        state_var_NS <= COMP_LOOP_C_410;
      WHEN COMP_LOOP_C_410 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011000");
        state_var_NS <= COMP_LOOP_C_411;
      WHEN COMP_LOOP_C_411 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011001");
        state_var_NS <= COMP_LOOP_C_412;
      WHEN COMP_LOOP_C_412 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011010");
        state_var_NS <= COMP_LOOP_C_413;
      WHEN COMP_LOOP_C_413 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011011");
        state_var_NS <= COMP_LOOP_C_414;
      WHEN COMP_LOOP_C_414 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011100");
        state_var_NS <= COMP_LOOP_C_415;
      WHEN COMP_LOOP_C_415 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011101");
        state_var_NS <= COMP_LOOP_C_416;
      WHEN COMP_LOOP_C_416 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011110");
        state_var_NS <= COMP_LOOP_C_417;
      WHEN COMP_LOOP_C_417 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011111");
        state_var_NS <= COMP_LOOP_C_418;
      WHEN COMP_LOOP_C_418 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100000");
        state_var_NS <= COMP_LOOP_C_419;
      WHEN COMP_LOOP_C_419 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100001");
        state_var_NS <= COMP_LOOP_C_420;
      WHEN COMP_LOOP_C_420 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100010");
        state_var_NS <= COMP_LOOP_C_421;
      WHEN COMP_LOOP_C_421 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100011");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100100");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100101");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100110");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100111");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101000");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101001");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101010");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101011");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101100");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101101");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101110");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101111");
        IF ( COMP_LOOP_10_modExp_dev_1_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_422;
        ELSE
          state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_422 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110000");
        state_var_NS <= COMP_LOOP_C_423;
      WHEN COMP_LOOP_C_423 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110001");
        state_var_NS <= COMP_LOOP_C_424;
      WHEN COMP_LOOP_C_424 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110010");
        state_var_NS <= COMP_LOOP_C_425;
      WHEN COMP_LOOP_C_425 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110011");
        state_var_NS <= COMP_LOOP_C_426;
      WHEN COMP_LOOP_C_426 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110100");
        state_var_NS <= COMP_LOOP_C_427;
      WHEN COMP_LOOP_C_427 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110101");
        state_var_NS <= COMP_LOOP_C_428;
      WHEN COMP_LOOP_C_428 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110110");
        state_var_NS <= COMP_LOOP_C_429;
      WHEN COMP_LOOP_C_429 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110111");
        state_var_NS <= COMP_LOOP_C_430;
      WHEN COMP_LOOP_C_430 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111000");
        state_var_NS <= COMP_LOOP_C_431;
      WHEN COMP_LOOP_C_431 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111001");
        state_var_NS <= COMP_LOOP_C_432;
      WHEN COMP_LOOP_C_432 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111010");
        state_var_NS <= COMP_LOOP_C_433;
      WHEN COMP_LOOP_C_433 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111011");
        state_var_NS <= COMP_LOOP_C_434;
      WHEN COMP_LOOP_C_434 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111100");
        state_var_NS <= COMP_LOOP_C_435;
      WHEN COMP_LOOP_C_435 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111101");
        state_var_NS <= COMP_LOOP_C_436;
      WHEN COMP_LOOP_C_436 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111110");
        state_var_NS <= COMP_LOOP_C_437;
      WHEN COMP_LOOP_C_437 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111111");
        state_var_NS <= COMP_LOOP_C_438;
      WHEN COMP_LOOP_C_438 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000000");
        state_var_NS <= COMP_LOOP_C_439;
      WHEN COMP_LOOP_C_439 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000001");
        state_var_NS <= COMP_LOOP_C_440;
      WHEN COMP_LOOP_C_440 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000010");
        state_var_NS <= COMP_LOOP_C_441;
      WHEN COMP_LOOP_C_441 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000011");
        state_var_NS <= COMP_LOOP_C_442;
      WHEN COMP_LOOP_C_442 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000100");
        state_var_NS <= COMP_LOOP_C_443;
      WHEN COMP_LOOP_C_443 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000101");
        state_var_NS <= COMP_LOOP_C_444;
      WHEN COMP_LOOP_C_444 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000110");
        state_var_NS <= COMP_LOOP_C_445;
      WHEN COMP_LOOP_C_445 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000111");
        state_var_NS <= COMP_LOOP_C_446;
      WHEN COMP_LOOP_C_446 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001000");
        state_var_NS <= COMP_LOOP_C_447;
      WHEN COMP_LOOP_C_447 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001001");
        state_var_NS <= COMP_LOOP_C_448;
      WHEN COMP_LOOP_C_448 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001010");
        state_var_NS <= COMP_LOOP_C_449;
      WHEN COMP_LOOP_C_449 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001011");
        state_var_NS <= COMP_LOOP_C_450;
      WHEN COMP_LOOP_C_450 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001100");
        IF ( COMP_LOOP_C_450_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_451;
        END IF;
      WHEN COMP_LOOP_C_451 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001101");
        state_var_NS <= COMP_LOOP_C_452;
      WHEN COMP_LOOP_C_452 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001110");
        state_var_NS <= COMP_LOOP_C_453;
      WHEN COMP_LOOP_C_453 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001111");
        state_var_NS <= COMP_LOOP_C_454;
      WHEN COMP_LOOP_C_454 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010000");
        state_var_NS <= COMP_LOOP_C_455;
      WHEN COMP_LOOP_C_455 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010001");
        state_var_NS <= COMP_LOOP_C_456;
      WHEN COMP_LOOP_C_456 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010010");
        state_var_NS <= COMP_LOOP_C_457;
      WHEN COMP_LOOP_C_457 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010011");
        state_var_NS <= COMP_LOOP_C_458;
      WHEN COMP_LOOP_C_458 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010100");
        state_var_NS <= COMP_LOOP_C_459;
      WHEN COMP_LOOP_C_459 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010101");
        state_var_NS <= COMP_LOOP_C_460;
      WHEN COMP_LOOP_C_460 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010110");
        state_var_NS <= COMP_LOOP_C_461;
      WHEN COMP_LOOP_C_461 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010111");
        state_var_NS <= COMP_LOOP_C_462;
      WHEN COMP_LOOP_C_462 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011000");
        state_var_NS <= COMP_LOOP_C_463;
      WHEN COMP_LOOP_C_463 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011001");
        state_var_NS <= COMP_LOOP_C_464;
      WHEN COMP_LOOP_C_464 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011010");
        state_var_NS <= COMP_LOOP_C_465;
      WHEN COMP_LOOP_C_465 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011011");
        state_var_NS <= COMP_LOOP_C_466;
      WHEN COMP_LOOP_C_466 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011100");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011101");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011110");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011111");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100000");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100001");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100010");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100011");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100100");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100101");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100110");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100111");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101000");
        IF ( COMP_LOOP_11_modExp_dev_1_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_467;
        ELSE
          state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_467 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101001");
        state_var_NS <= COMP_LOOP_C_468;
      WHEN COMP_LOOP_C_468 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101010");
        state_var_NS <= COMP_LOOP_C_469;
      WHEN COMP_LOOP_C_469 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101011");
        state_var_NS <= COMP_LOOP_C_470;
      WHEN COMP_LOOP_C_470 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101100");
        state_var_NS <= COMP_LOOP_C_471;
      WHEN COMP_LOOP_C_471 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101101");
        state_var_NS <= COMP_LOOP_C_472;
      WHEN COMP_LOOP_C_472 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101110");
        state_var_NS <= COMP_LOOP_C_473;
      WHEN COMP_LOOP_C_473 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101111");
        state_var_NS <= COMP_LOOP_C_474;
      WHEN COMP_LOOP_C_474 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110000");
        state_var_NS <= COMP_LOOP_C_475;
      WHEN COMP_LOOP_C_475 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110001");
        state_var_NS <= COMP_LOOP_C_476;
      WHEN COMP_LOOP_C_476 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110010");
        state_var_NS <= COMP_LOOP_C_477;
      WHEN COMP_LOOP_C_477 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110011");
        state_var_NS <= COMP_LOOP_C_478;
      WHEN COMP_LOOP_C_478 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110100");
        state_var_NS <= COMP_LOOP_C_479;
      WHEN COMP_LOOP_C_479 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110101");
        state_var_NS <= COMP_LOOP_C_480;
      WHEN COMP_LOOP_C_480 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110110");
        state_var_NS <= COMP_LOOP_C_481;
      WHEN COMP_LOOP_C_481 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110111");
        state_var_NS <= COMP_LOOP_C_482;
      WHEN COMP_LOOP_C_482 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111000");
        state_var_NS <= COMP_LOOP_C_483;
      WHEN COMP_LOOP_C_483 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111001");
        state_var_NS <= COMP_LOOP_C_484;
      WHEN COMP_LOOP_C_484 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111010");
        state_var_NS <= COMP_LOOP_C_485;
      WHEN COMP_LOOP_C_485 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111011");
        state_var_NS <= COMP_LOOP_C_486;
      WHEN COMP_LOOP_C_486 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111100");
        state_var_NS <= COMP_LOOP_C_487;
      WHEN COMP_LOOP_C_487 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111101");
        state_var_NS <= COMP_LOOP_C_488;
      WHEN COMP_LOOP_C_488 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111110");
        state_var_NS <= COMP_LOOP_C_489;
      WHEN COMP_LOOP_C_489 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111111");
        state_var_NS <= COMP_LOOP_C_490;
      WHEN COMP_LOOP_C_490 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000000");
        state_var_NS <= COMP_LOOP_C_491;
      WHEN COMP_LOOP_C_491 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000001");
        state_var_NS <= COMP_LOOP_C_492;
      WHEN COMP_LOOP_C_492 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000010");
        state_var_NS <= COMP_LOOP_C_493;
      WHEN COMP_LOOP_C_493 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000011");
        state_var_NS <= COMP_LOOP_C_494;
      WHEN COMP_LOOP_C_494 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000100");
        state_var_NS <= COMP_LOOP_C_495;
      WHEN COMP_LOOP_C_495 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000101");
        IF ( COMP_LOOP_C_495_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_496;
        END IF;
      WHEN COMP_LOOP_C_496 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000110");
        state_var_NS <= COMP_LOOP_C_497;
      WHEN COMP_LOOP_C_497 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000111");
        state_var_NS <= COMP_LOOP_C_498;
      WHEN COMP_LOOP_C_498 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001000");
        state_var_NS <= COMP_LOOP_C_499;
      WHEN COMP_LOOP_C_499 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001001");
        state_var_NS <= COMP_LOOP_C_500;
      WHEN COMP_LOOP_C_500 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001010");
        state_var_NS <= COMP_LOOP_C_501;
      WHEN COMP_LOOP_C_501 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001011");
        state_var_NS <= COMP_LOOP_C_502;
      WHEN COMP_LOOP_C_502 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001100");
        state_var_NS <= COMP_LOOP_C_503;
      WHEN COMP_LOOP_C_503 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001101");
        state_var_NS <= COMP_LOOP_C_504;
      WHEN COMP_LOOP_C_504 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001110");
        state_var_NS <= COMP_LOOP_C_505;
      WHEN COMP_LOOP_C_505 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001111");
        state_var_NS <= COMP_LOOP_C_506;
      WHEN COMP_LOOP_C_506 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010000");
        state_var_NS <= COMP_LOOP_C_507;
      WHEN COMP_LOOP_C_507 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010001");
        state_var_NS <= COMP_LOOP_C_508;
      WHEN COMP_LOOP_C_508 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010010");
        state_var_NS <= COMP_LOOP_C_509;
      WHEN COMP_LOOP_C_509 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010011");
        state_var_NS <= COMP_LOOP_C_510;
      WHEN COMP_LOOP_C_510 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010100");
        state_var_NS <= COMP_LOOP_C_511;
      WHEN COMP_LOOP_C_511 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010101");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010110");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010111");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011000");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011001");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011010");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011011");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011100");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011101");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011110");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011111");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100000");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100001");
        IF ( COMP_LOOP_12_modExp_dev_1_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_512;
        ELSE
          state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_512 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100010");
        state_var_NS <= COMP_LOOP_C_513;
      WHEN COMP_LOOP_C_513 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100011");
        state_var_NS <= COMP_LOOP_C_514;
      WHEN COMP_LOOP_C_514 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100100");
        state_var_NS <= COMP_LOOP_C_515;
      WHEN COMP_LOOP_C_515 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100101");
        state_var_NS <= COMP_LOOP_C_516;
      WHEN COMP_LOOP_C_516 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100110");
        state_var_NS <= COMP_LOOP_C_517;
      WHEN COMP_LOOP_C_517 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100111");
        state_var_NS <= COMP_LOOP_C_518;
      WHEN COMP_LOOP_C_518 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101000");
        state_var_NS <= COMP_LOOP_C_519;
      WHEN COMP_LOOP_C_519 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101001");
        state_var_NS <= COMP_LOOP_C_520;
      WHEN COMP_LOOP_C_520 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101010");
        state_var_NS <= COMP_LOOP_C_521;
      WHEN COMP_LOOP_C_521 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101011");
        state_var_NS <= COMP_LOOP_C_522;
      WHEN COMP_LOOP_C_522 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101100");
        state_var_NS <= COMP_LOOP_C_523;
      WHEN COMP_LOOP_C_523 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101101");
        state_var_NS <= COMP_LOOP_C_524;
      WHEN COMP_LOOP_C_524 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101110");
        state_var_NS <= COMP_LOOP_C_525;
      WHEN COMP_LOOP_C_525 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101111");
        state_var_NS <= COMP_LOOP_C_526;
      WHEN COMP_LOOP_C_526 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110000");
        state_var_NS <= COMP_LOOP_C_527;
      WHEN COMP_LOOP_C_527 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110001");
        state_var_NS <= COMP_LOOP_C_528;
      WHEN COMP_LOOP_C_528 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110010");
        state_var_NS <= COMP_LOOP_C_529;
      WHEN COMP_LOOP_C_529 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110011");
        state_var_NS <= COMP_LOOP_C_530;
      WHEN COMP_LOOP_C_530 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110100");
        state_var_NS <= COMP_LOOP_C_531;
      WHEN COMP_LOOP_C_531 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110101");
        state_var_NS <= COMP_LOOP_C_532;
      WHEN COMP_LOOP_C_532 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110110");
        state_var_NS <= COMP_LOOP_C_533;
      WHEN COMP_LOOP_C_533 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110111");
        state_var_NS <= COMP_LOOP_C_534;
      WHEN COMP_LOOP_C_534 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111000");
        state_var_NS <= COMP_LOOP_C_535;
      WHEN COMP_LOOP_C_535 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111001");
        state_var_NS <= COMP_LOOP_C_536;
      WHEN COMP_LOOP_C_536 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111010");
        state_var_NS <= COMP_LOOP_C_537;
      WHEN COMP_LOOP_C_537 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111011");
        state_var_NS <= COMP_LOOP_C_538;
      WHEN COMP_LOOP_C_538 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111100");
        state_var_NS <= COMP_LOOP_C_539;
      WHEN COMP_LOOP_C_539 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111101");
        state_var_NS <= COMP_LOOP_C_540;
      WHEN COMP_LOOP_C_540 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111110");
        IF ( COMP_LOOP_C_540_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_541;
        END IF;
      WHEN COMP_LOOP_C_541 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111111");
        state_var_NS <= COMP_LOOP_C_542;
      WHEN COMP_LOOP_C_542 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000000");
        state_var_NS <= COMP_LOOP_C_543;
      WHEN COMP_LOOP_C_543 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000001");
        state_var_NS <= COMP_LOOP_C_544;
      WHEN COMP_LOOP_C_544 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000010");
        state_var_NS <= COMP_LOOP_C_545;
      WHEN COMP_LOOP_C_545 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000011");
        state_var_NS <= COMP_LOOP_C_546;
      WHEN COMP_LOOP_C_546 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000100");
        state_var_NS <= COMP_LOOP_C_547;
      WHEN COMP_LOOP_C_547 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000101");
        state_var_NS <= COMP_LOOP_C_548;
      WHEN COMP_LOOP_C_548 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000110");
        state_var_NS <= COMP_LOOP_C_549;
      WHEN COMP_LOOP_C_549 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000111");
        state_var_NS <= COMP_LOOP_C_550;
      WHEN COMP_LOOP_C_550 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001000");
        state_var_NS <= COMP_LOOP_C_551;
      WHEN COMP_LOOP_C_551 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001001");
        state_var_NS <= COMP_LOOP_C_552;
      WHEN COMP_LOOP_C_552 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001010");
        state_var_NS <= COMP_LOOP_C_553;
      WHEN COMP_LOOP_C_553 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001011");
        state_var_NS <= COMP_LOOP_C_554;
      WHEN COMP_LOOP_C_554 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001100");
        state_var_NS <= COMP_LOOP_C_555;
      WHEN COMP_LOOP_C_555 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001101");
        state_var_NS <= COMP_LOOP_C_556;
      WHEN COMP_LOOP_C_556 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001110");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001111");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010000");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010001");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010010");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010011");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010100");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010101");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010110");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010111");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011000");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011001");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011010");
        IF ( COMP_LOOP_13_modExp_dev_1_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_557;
        ELSE
          state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_557 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011011");
        state_var_NS <= COMP_LOOP_C_558;
      WHEN COMP_LOOP_C_558 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011100");
        state_var_NS <= COMP_LOOP_C_559;
      WHEN COMP_LOOP_C_559 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011101");
        state_var_NS <= COMP_LOOP_C_560;
      WHEN COMP_LOOP_C_560 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011110");
        state_var_NS <= COMP_LOOP_C_561;
      WHEN COMP_LOOP_C_561 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011111");
        state_var_NS <= COMP_LOOP_C_562;
      WHEN COMP_LOOP_C_562 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100000");
        state_var_NS <= COMP_LOOP_C_563;
      WHEN COMP_LOOP_C_563 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100001");
        state_var_NS <= COMP_LOOP_C_564;
      WHEN COMP_LOOP_C_564 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100010");
        state_var_NS <= COMP_LOOP_C_565;
      WHEN COMP_LOOP_C_565 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100011");
        state_var_NS <= COMP_LOOP_C_566;
      WHEN COMP_LOOP_C_566 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100100");
        state_var_NS <= COMP_LOOP_C_567;
      WHEN COMP_LOOP_C_567 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100101");
        state_var_NS <= COMP_LOOP_C_568;
      WHEN COMP_LOOP_C_568 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100110");
        state_var_NS <= COMP_LOOP_C_569;
      WHEN COMP_LOOP_C_569 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100111");
        state_var_NS <= COMP_LOOP_C_570;
      WHEN COMP_LOOP_C_570 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101000");
        state_var_NS <= COMP_LOOP_C_571;
      WHEN COMP_LOOP_C_571 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101001");
        state_var_NS <= COMP_LOOP_C_572;
      WHEN COMP_LOOP_C_572 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101010");
        state_var_NS <= COMP_LOOP_C_573;
      WHEN COMP_LOOP_C_573 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101011");
        state_var_NS <= COMP_LOOP_C_574;
      WHEN COMP_LOOP_C_574 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101100");
        state_var_NS <= COMP_LOOP_C_575;
      WHEN COMP_LOOP_C_575 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101101");
        state_var_NS <= COMP_LOOP_C_576;
      WHEN COMP_LOOP_C_576 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101110");
        state_var_NS <= COMP_LOOP_C_577;
      WHEN COMP_LOOP_C_577 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101111");
        state_var_NS <= COMP_LOOP_C_578;
      WHEN COMP_LOOP_C_578 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110000");
        state_var_NS <= COMP_LOOP_C_579;
      WHEN COMP_LOOP_C_579 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110001");
        state_var_NS <= COMP_LOOP_C_580;
      WHEN COMP_LOOP_C_580 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110010");
        state_var_NS <= COMP_LOOP_C_581;
      WHEN COMP_LOOP_C_581 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110011");
        state_var_NS <= COMP_LOOP_C_582;
      WHEN COMP_LOOP_C_582 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110100");
        state_var_NS <= COMP_LOOP_C_583;
      WHEN COMP_LOOP_C_583 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110101");
        state_var_NS <= COMP_LOOP_C_584;
      WHEN COMP_LOOP_C_584 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110110");
        state_var_NS <= COMP_LOOP_C_585;
      WHEN COMP_LOOP_C_585 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110111");
        IF ( COMP_LOOP_C_585_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_586;
        END IF;
      WHEN COMP_LOOP_C_586 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111000");
        state_var_NS <= COMP_LOOP_C_587;
      WHEN COMP_LOOP_C_587 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111001");
        state_var_NS <= COMP_LOOP_C_588;
      WHEN COMP_LOOP_C_588 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111010");
        state_var_NS <= COMP_LOOP_C_589;
      WHEN COMP_LOOP_C_589 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111011");
        state_var_NS <= COMP_LOOP_C_590;
      WHEN COMP_LOOP_C_590 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111100");
        state_var_NS <= COMP_LOOP_C_591;
      WHEN COMP_LOOP_C_591 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111101");
        state_var_NS <= COMP_LOOP_C_592;
      WHEN COMP_LOOP_C_592 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111110");
        state_var_NS <= COMP_LOOP_C_593;
      WHEN COMP_LOOP_C_593 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111111");
        state_var_NS <= COMP_LOOP_C_594;
      WHEN COMP_LOOP_C_594 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000000");
        state_var_NS <= COMP_LOOP_C_595;
      WHEN COMP_LOOP_C_595 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000001");
        state_var_NS <= COMP_LOOP_C_596;
      WHEN COMP_LOOP_C_596 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000010");
        state_var_NS <= COMP_LOOP_C_597;
      WHEN COMP_LOOP_C_597 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000011");
        state_var_NS <= COMP_LOOP_C_598;
      WHEN COMP_LOOP_C_598 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000100");
        state_var_NS <= COMP_LOOP_C_599;
      WHEN COMP_LOOP_C_599 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000101");
        state_var_NS <= COMP_LOOP_C_600;
      WHEN COMP_LOOP_C_600 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000110");
        state_var_NS <= COMP_LOOP_C_601;
      WHEN COMP_LOOP_C_601 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000111");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100001000");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100001001");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100001010");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100001011");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100001100");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100001101");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100001110");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100001111");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100010000");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100010001");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100010010");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100010011");
        IF ( COMP_LOOP_14_modExp_dev_1_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_602;
        ELSE
          state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_602 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100010100");
        state_var_NS <= COMP_LOOP_C_603;
      WHEN COMP_LOOP_C_603 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100010101");
        state_var_NS <= COMP_LOOP_C_604;
      WHEN COMP_LOOP_C_604 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100010110");
        state_var_NS <= COMP_LOOP_C_605;
      WHEN COMP_LOOP_C_605 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100010111");
        state_var_NS <= COMP_LOOP_C_606;
      WHEN COMP_LOOP_C_606 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100011000");
        state_var_NS <= COMP_LOOP_C_607;
      WHEN COMP_LOOP_C_607 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100011001");
        state_var_NS <= COMP_LOOP_C_608;
      WHEN COMP_LOOP_C_608 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100011010");
        state_var_NS <= COMP_LOOP_C_609;
      WHEN COMP_LOOP_C_609 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100011011");
        state_var_NS <= COMP_LOOP_C_610;
      WHEN COMP_LOOP_C_610 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100011100");
        state_var_NS <= COMP_LOOP_C_611;
      WHEN COMP_LOOP_C_611 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100011101");
        state_var_NS <= COMP_LOOP_C_612;
      WHEN COMP_LOOP_C_612 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100011110");
        state_var_NS <= COMP_LOOP_C_613;
      WHEN COMP_LOOP_C_613 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100011111");
        state_var_NS <= COMP_LOOP_C_614;
      WHEN COMP_LOOP_C_614 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100100000");
        state_var_NS <= COMP_LOOP_C_615;
      WHEN COMP_LOOP_C_615 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100100001");
        state_var_NS <= COMP_LOOP_C_616;
      WHEN COMP_LOOP_C_616 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100100010");
        state_var_NS <= COMP_LOOP_C_617;
      WHEN COMP_LOOP_C_617 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100100011");
        state_var_NS <= COMP_LOOP_C_618;
      WHEN COMP_LOOP_C_618 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100100100");
        state_var_NS <= COMP_LOOP_C_619;
      WHEN COMP_LOOP_C_619 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100100101");
        state_var_NS <= COMP_LOOP_C_620;
      WHEN COMP_LOOP_C_620 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100100110");
        state_var_NS <= COMP_LOOP_C_621;
      WHEN COMP_LOOP_C_621 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100100111");
        state_var_NS <= COMP_LOOP_C_622;
      WHEN COMP_LOOP_C_622 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100101000");
        state_var_NS <= COMP_LOOP_C_623;
      WHEN COMP_LOOP_C_623 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100101001");
        state_var_NS <= COMP_LOOP_C_624;
      WHEN COMP_LOOP_C_624 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100101010");
        state_var_NS <= COMP_LOOP_C_625;
      WHEN COMP_LOOP_C_625 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100101011");
        state_var_NS <= COMP_LOOP_C_626;
      WHEN COMP_LOOP_C_626 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100101100");
        state_var_NS <= COMP_LOOP_C_627;
      WHEN COMP_LOOP_C_627 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100101101");
        state_var_NS <= COMP_LOOP_C_628;
      WHEN COMP_LOOP_C_628 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100101110");
        state_var_NS <= COMP_LOOP_C_629;
      WHEN COMP_LOOP_C_629 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100101111");
        state_var_NS <= COMP_LOOP_C_630;
      WHEN COMP_LOOP_C_630 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100110000");
        IF ( COMP_LOOP_C_630_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_631;
        END IF;
      WHEN COMP_LOOP_C_631 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100110001");
        state_var_NS <= COMP_LOOP_C_632;
      WHEN COMP_LOOP_C_632 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100110010");
        state_var_NS <= COMP_LOOP_C_633;
      WHEN COMP_LOOP_C_633 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100110011");
        state_var_NS <= COMP_LOOP_C_634;
      WHEN COMP_LOOP_C_634 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100110100");
        state_var_NS <= COMP_LOOP_C_635;
      WHEN COMP_LOOP_C_635 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100110101");
        state_var_NS <= COMP_LOOP_C_636;
      WHEN COMP_LOOP_C_636 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100110110");
        state_var_NS <= COMP_LOOP_C_637;
      WHEN COMP_LOOP_C_637 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100110111");
        state_var_NS <= COMP_LOOP_C_638;
      WHEN COMP_LOOP_C_638 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100111000");
        state_var_NS <= COMP_LOOP_C_639;
      WHEN COMP_LOOP_C_639 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100111001");
        state_var_NS <= COMP_LOOP_C_640;
      WHEN COMP_LOOP_C_640 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100111010");
        state_var_NS <= COMP_LOOP_C_641;
      WHEN COMP_LOOP_C_641 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100111011");
        state_var_NS <= COMP_LOOP_C_642;
      WHEN COMP_LOOP_C_642 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100111100");
        state_var_NS <= COMP_LOOP_C_643;
      WHEN COMP_LOOP_C_643 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100111101");
        state_var_NS <= COMP_LOOP_C_644;
      WHEN COMP_LOOP_C_644 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100111110");
        state_var_NS <= COMP_LOOP_C_645;
      WHEN COMP_LOOP_C_645 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100111111");
        state_var_NS <= COMP_LOOP_C_646;
      WHEN COMP_LOOP_C_646 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101000000");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101000001");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101000010");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101000011");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101000100");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101000101");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101000110");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101000111");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101001000");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101001001");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101001010");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101001011");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101001100");
        IF ( COMP_LOOP_15_modExp_dev_1_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_647;
        ELSE
          state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_647 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101001101");
        state_var_NS <= COMP_LOOP_C_648;
      WHEN COMP_LOOP_C_648 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101001110");
        state_var_NS <= COMP_LOOP_C_649;
      WHEN COMP_LOOP_C_649 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101001111");
        state_var_NS <= COMP_LOOP_C_650;
      WHEN COMP_LOOP_C_650 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101010000");
        state_var_NS <= COMP_LOOP_C_651;
      WHEN COMP_LOOP_C_651 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101010001");
        state_var_NS <= COMP_LOOP_C_652;
      WHEN COMP_LOOP_C_652 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101010010");
        state_var_NS <= COMP_LOOP_C_653;
      WHEN COMP_LOOP_C_653 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101010011");
        state_var_NS <= COMP_LOOP_C_654;
      WHEN COMP_LOOP_C_654 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101010100");
        state_var_NS <= COMP_LOOP_C_655;
      WHEN COMP_LOOP_C_655 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101010101");
        state_var_NS <= COMP_LOOP_C_656;
      WHEN COMP_LOOP_C_656 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101010110");
        state_var_NS <= COMP_LOOP_C_657;
      WHEN COMP_LOOP_C_657 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101010111");
        state_var_NS <= COMP_LOOP_C_658;
      WHEN COMP_LOOP_C_658 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101011000");
        state_var_NS <= COMP_LOOP_C_659;
      WHEN COMP_LOOP_C_659 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101011001");
        state_var_NS <= COMP_LOOP_C_660;
      WHEN COMP_LOOP_C_660 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101011010");
        state_var_NS <= COMP_LOOP_C_661;
      WHEN COMP_LOOP_C_661 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101011011");
        state_var_NS <= COMP_LOOP_C_662;
      WHEN COMP_LOOP_C_662 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101011100");
        state_var_NS <= COMP_LOOP_C_663;
      WHEN COMP_LOOP_C_663 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101011101");
        state_var_NS <= COMP_LOOP_C_664;
      WHEN COMP_LOOP_C_664 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101011110");
        state_var_NS <= COMP_LOOP_C_665;
      WHEN COMP_LOOP_C_665 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101011111");
        state_var_NS <= COMP_LOOP_C_666;
      WHEN COMP_LOOP_C_666 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101100000");
        state_var_NS <= COMP_LOOP_C_667;
      WHEN COMP_LOOP_C_667 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101100001");
        state_var_NS <= COMP_LOOP_C_668;
      WHEN COMP_LOOP_C_668 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101100010");
        state_var_NS <= COMP_LOOP_C_669;
      WHEN COMP_LOOP_C_669 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101100011");
        state_var_NS <= COMP_LOOP_C_670;
      WHEN COMP_LOOP_C_670 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101100100");
        state_var_NS <= COMP_LOOP_C_671;
      WHEN COMP_LOOP_C_671 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101100101");
        state_var_NS <= COMP_LOOP_C_672;
      WHEN COMP_LOOP_C_672 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101100110");
        state_var_NS <= COMP_LOOP_C_673;
      WHEN COMP_LOOP_C_673 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101100111");
        state_var_NS <= COMP_LOOP_C_674;
      WHEN COMP_LOOP_C_674 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101101000");
        state_var_NS <= COMP_LOOP_C_675;
      WHEN COMP_LOOP_C_675 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101101001");
        IF ( COMP_LOOP_C_675_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_676;
        END IF;
      WHEN COMP_LOOP_C_676 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101101010");
        state_var_NS <= COMP_LOOP_C_677;
      WHEN COMP_LOOP_C_677 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101101011");
        state_var_NS <= COMP_LOOP_C_678;
      WHEN COMP_LOOP_C_678 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101101100");
        state_var_NS <= COMP_LOOP_C_679;
      WHEN COMP_LOOP_C_679 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101101101");
        state_var_NS <= COMP_LOOP_C_680;
      WHEN COMP_LOOP_C_680 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101101110");
        state_var_NS <= COMP_LOOP_C_681;
      WHEN COMP_LOOP_C_681 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101101111");
        state_var_NS <= COMP_LOOP_C_682;
      WHEN COMP_LOOP_C_682 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101110000");
        state_var_NS <= COMP_LOOP_C_683;
      WHEN COMP_LOOP_C_683 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101110001");
        state_var_NS <= COMP_LOOP_C_684;
      WHEN COMP_LOOP_C_684 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101110010");
        state_var_NS <= COMP_LOOP_C_685;
      WHEN COMP_LOOP_C_685 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101110011");
        state_var_NS <= COMP_LOOP_C_686;
      WHEN COMP_LOOP_C_686 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101110100");
        state_var_NS <= COMP_LOOP_C_687;
      WHEN COMP_LOOP_C_687 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101110101");
        state_var_NS <= COMP_LOOP_C_688;
      WHEN COMP_LOOP_C_688 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101110110");
        state_var_NS <= COMP_LOOP_C_689;
      WHEN COMP_LOOP_C_689 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101110111");
        state_var_NS <= COMP_LOOP_C_690;
      WHEN COMP_LOOP_C_690 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101111000");
        state_var_NS <= COMP_LOOP_C_691;
      WHEN COMP_LOOP_C_691 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101111001");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101111010");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101111011");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101111100");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101111101");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101111110");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1101111111");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110000000");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110000001");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110000010");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110000011");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110000100");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110000101");
        IF ( COMP_LOOP_16_modExp_dev_1_while_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_692;
        ELSE
          state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_692 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110000110");
        state_var_NS <= COMP_LOOP_C_693;
      WHEN COMP_LOOP_C_693 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110000111");
        state_var_NS <= COMP_LOOP_C_694;
      WHEN COMP_LOOP_C_694 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110001000");
        state_var_NS <= COMP_LOOP_C_695;
      WHEN COMP_LOOP_C_695 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110001001");
        state_var_NS <= COMP_LOOP_C_696;
      WHEN COMP_LOOP_C_696 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110001010");
        state_var_NS <= COMP_LOOP_C_697;
      WHEN COMP_LOOP_C_697 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110001011");
        state_var_NS <= COMP_LOOP_C_698;
      WHEN COMP_LOOP_C_698 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110001100");
        state_var_NS <= COMP_LOOP_C_699;
      WHEN COMP_LOOP_C_699 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110001101");
        state_var_NS <= COMP_LOOP_C_700;
      WHEN COMP_LOOP_C_700 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110001110");
        state_var_NS <= COMP_LOOP_C_701;
      WHEN COMP_LOOP_C_701 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110001111");
        state_var_NS <= COMP_LOOP_C_702;
      WHEN COMP_LOOP_C_702 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110010000");
        state_var_NS <= COMP_LOOP_C_703;
      WHEN COMP_LOOP_C_703 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110010001");
        state_var_NS <= COMP_LOOP_C_704;
      WHEN COMP_LOOP_C_704 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110010010");
        state_var_NS <= COMP_LOOP_C_705;
      WHEN COMP_LOOP_C_705 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110010011");
        state_var_NS <= COMP_LOOP_C_706;
      WHEN COMP_LOOP_C_706 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110010100");
        state_var_NS <= COMP_LOOP_C_707;
      WHEN COMP_LOOP_C_707 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110010101");
        state_var_NS <= COMP_LOOP_C_708;
      WHEN COMP_LOOP_C_708 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110010110");
        state_var_NS <= COMP_LOOP_C_709;
      WHEN COMP_LOOP_C_709 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110010111");
        state_var_NS <= COMP_LOOP_C_710;
      WHEN COMP_LOOP_C_710 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110011000");
        state_var_NS <= COMP_LOOP_C_711;
      WHEN COMP_LOOP_C_711 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110011001");
        state_var_NS <= COMP_LOOP_C_712;
      WHEN COMP_LOOP_C_712 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110011010");
        state_var_NS <= COMP_LOOP_C_713;
      WHEN COMP_LOOP_C_713 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110011011");
        state_var_NS <= COMP_LOOP_C_714;
      WHEN COMP_LOOP_C_714 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110011100");
        state_var_NS <= COMP_LOOP_C_715;
      WHEN COMP_LOOP_C_715 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110011101");
        state_var_NS <= COMP_LOOP_C_716;
      WHEN COMP_LOOP_C_716 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110011110");
        state_var_NS <= COMP_LOOP_C_717;
      WHEN COMP_LOOP_C_717 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110011111");
        state_var_NS <= COMP_LOOP_C_718;
      WHEN COMP_LOOP_C_718 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110100000");
        state_var_NS <= COMP_LOOP_C_719;
      WHEN COMP_LOOP_C_719 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110100001");
        state_var_NS <= COMP_LOOP_C_720;
      WHEN COMP_LOOP_C_720 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110100010");
        IF ( COMP_LOOP_C_720_tr0 = '1' ) THEN
          state_var_NS <= STAGE_VEC_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN STAGE_VEC_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110100011");
        IF ( STAGE_VEC_LOOP_C_1_tr0 = '1' ) THEN
          state_var_NS <= STAGE_MAIN_LOOP_C_4;
        ELSE
          state_var_NS <= STAGE_VEC_LOOP_C_0;
        END IF;
      WHEN STAGE_MAIN_LOOP_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110100100");
        IF ( STAGE_MAIN_LOOP_C_4_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSE
          state_var_NS <= STAGE_MAIN_LOOP_C_0;
        END IF;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1110100101");
        state_var_NS <= main_C_0;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000");
        state_var_NS <= STAGE_MAIN_LOOP_C_0;
    END CASE;
  END PROCESS inPlaceNTT_DIF_core_core_fsm_1;

  inPlaceNTT_DIF_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        state_var <= state_var_NS;
      END IF;
    END IF;
  END PROCESS inPlaceNTT_DIF_core_core_fsm_1_REG;

END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_core_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_core_wait_dp IS
  PORT(
    ensig_cgo_iro : IN STD_LOGIC;
    ensig_cgo : IN STD_LOGIC;
    COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_core_wait_dp;

ARCHITECTURE v7 OF inPlaceNTT_DIF_core_wait_dp IS
  -- Default Constants

BEGIN
  COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en <= ensig_cgo OR ensig_cgo_iro;
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC;
    vec_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_0_i_adra_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_1_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_2_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_3_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_4_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_5_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_6_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_7_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_8_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_9_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_10_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_11_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_12_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_13_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_14_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_15_i_wea_d_pff : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_core;

ARCHITECTURE v7 OF inPlaceNTT_DIF_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL p_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL r_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_return_rsc_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en : STD_LOGIC;
  SIGNAL modExp_dev_while_rem_cmp_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modExp_dev_while_rem_cmp_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_MAIN_LOOP_div_cmp_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_MAIN_LOOP_div_cmp_b : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL STAGE_MAIN_LOOP_div_cmp_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL fsm_output : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_1_operator_64_false_acc_tmp : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL or_tmp : STD_LOGIC;
  SIGNAL nor_tmp_1 : STD_LOGIC;
  SIGNAL nor_tmp_3 : STD_LOGIC;
  SIGNAL and_dcpl : STD_LOGIC;
  SIGNAL and_dcpl_5 : STD_LOGIC;
  SIGNAL or_tmp_33 : STD_LOGIC;
  SIGNAL mux_tmp_79 : STD_LOGIC;
  SIGNAL nor_tmp_87 : STD_LOGIC;
  SIGNAL mux_tmp_302 : STD_LOGIC;
  SIGNAL or_tmp_235 : STD_LOGIC;
  SIGNAL nor_tmp_130 : STD_LOGIC;
  SIGNAL and_tmp_11 : STD_LOGIC;
  SIGNAL and_dcpl_44 : STD_LOGIC;
  SIGNAL and_dcpl_70 : STD_LOGIC;
  SIGNAL not_tmp_266 : STD_LOGIC;
  SIGNAL and_dcpl_91 : STD_LOGIC;
  SIGNAL and_dcpl_92 : STD_LOGIC;
  SIGNAL and_dcpl_93 : STD_LOGIC;
  SIGNAL and_dcpl_94 : STD_LOGIC;
  SIGNAL and_dcpl_95 : STD_LOGIC;
  SIGNAL and_dcpl_96 : STD_LOGIC;
  SIGNAL and_dcpl_97 : STD_LOGIC;
  SIGNAL and_dcpl_98 : STD_LOGIC;
  SIGNAL or_tmp_546 : STD_LOGIC;
  SIGNAL and_dcpl_105 : STD_LOGIC;
  SIGNAL and_dcpl_106 : STD_LOGIC;
  SIGNAL and_dcpl_109 : STD_LOGIC;
  SIGNAL xor_dcpl : STD_LOGIC;
  SIGNAL and_dcpl_113 : STD_LOGIC;
  SIGNAL not_tmp_280 : STD_LOGIC;
  SIGNAL and_dcpl_125 : STD_LOGIC;
  SIGNAL and_dcpl_131 : STD_LOGIC;
  SIGNAL and_dcpl_135 : STD_LOGIC;
  SIGNAL and_dcpl_143 : STD_LOGIC;
  SIGNAL and_dcpl_146 : STD_LOGIC;
  SIGNAL and_dcpl_147 : STD_LOGIC;
  SIGNAL and_dcpl_158 : STD_LOGIC;
  SIGNAL and_dcpl_159 : STD_LOGIC;
  SIGNAL not_tmp_292 : STD_LOGIC;
  SIGNAL and_dcpl_176 : STD_LOGIC;
  SIGNAL and_dcpl_192 : STD_LOGIC;
  SIGNAL and_dcpl_199 : STD_LOGIC;
  SIGNAL or_tmp_591 : STD_LOGIC;
  SIGNAL and_dcpl_225 : STD_LOGIC;
  SIGNAL not_tmp_311 : STD_LOGIC;
  SIGNAL not_tmp_312 : STD_LOGIC;
  SIGNAL nand_tmp_16 : STD_LOGIC;
  SIGNAL or_tmp_669 : STD_LOGIC;
  SIGNAL nand_tmp_19 : STD_LOGIC;
  SIGNAL not_tmp_322 : STD_LOGIC;
  SIGNAL nand_tmp_22 : STD_LOGIC;
  SIGNAL nand_tmp_28 : STD_LOGIC;
  SIGNAL nand_tmp_34 : STD_LOGIC;
  SIGNAL nand_tmp_40 : STD_LOGIC;
  SIGNAL nand_tmp_46 : STD_LOGIC;
  SIGNAL nand_tmp_52 : STD_LOGIC;
  SIGNAL nand_tmp_58 : STD_LOGIC;
  SIGNAL nand_tmp_64 : STD_LOGIC;
  SIGNAL nand_tmp_70 : STD_LOGIC;
  SIGNAL nand_tmp_76 : STD_LOGIC;
  SIGNAL nand_tmp_82 : STD_LOGIC;
  SIGNAL nand_tmp_88 : STD_LOGIC;
  SIGNAL nand_tmp_94 : STD_LOGIC;
  SIGNAL nand_tmp_100 : STD_LOGIC;
  SIGNAL nand_tmp_106 : STD_LOGIC;
  SIGNAL or_tmp_2322 : STD_LOGIC;
  SIGNAL mux_tmp_2110 : STD_LOGIC;
  SIGNAL mux_tmp_2111 : STD_LOGIC;
  SIGNAL mux_tmp_2112 : STD_LOGIC;
  SIGNAL mux_tmp_2113 : STD_LOGIC;
  SIGNAL or_tmp_2324 : STD_LOGIC;
  SIGNAL mux_tmp_2114 : STD_LOGIC;
  SIGNAL mux_tmp_2118 : STD_LOGIC;
  SIGNAL mux_tmp_2124 : STD_LOGIC;
  SIGNAL mux_tmp_2127 : STD_LOGIC;
  SIGNAL mux_tmp_2129 : STD_LOGIC;
  SIGNAL mux_tmp_2130 : STD_LOGIC;
  SIGNAL mux_tmp_2131 : STD_LOGIC;
  SIGNAL mux_tmp_2132 : STD_LOGIC;
  SIGNAL mux_tmp_2135 : STD_LOGIC;
  SIGNAL mux_tmp_2139 : STD_LOGIC;
  SIGNAL mux_tmp_2142 : STD_LOGIC;
  SIGNAL nor_tmp_357 : STD_LOGIC;
  SIGNAL mux_tmp_2161 : STD_LOGIC;
  SIGNAL and_dcpl_239 : STD_LOGIC;
  SIGNAL and_dcpl_240 : STD_LOGIC;
  SIGNAL or_tmp_2348 : STD_LOGIC;
  SIGNAL or_tmp_2352 : STD_LOGIC;
  SIGNAL or_tmp_2355 : STD_LOGIC;
  SIGNAL and_dcpl_241 : STD_LOGIC;
  SIGNAL and_dcpl_242 : STD_LOGIC;
  SIGNAL and_dcpl_243 : STD_LOGIC;
  SIGNAL and_dcpl_244 : STD_LOGIC;
  SIGNAL and_dcpl_245 : STD_LOGIC;
  SIGNAL and_dcpl_246 : STD_LOGIC;
  SIGNAL and_dcpl_248 : STD_LOGIC;
  SIGNAL and_dcpl_249 : STD_LOGIC;
  SIGNAL and_dcpl_251 : STD_LOGIC;
  SIGNAL and_dcpl_252 : STD_LOGIC;
  SIGNAL and_dcpl_253 : STD_LOGIC;
  SIGNAL and_dcpl_254 : STD_LOGIC;
  SIGNAL and_dcpl_255 : STD_LOGIC;
  SIGNAL and_dcpl_256 : STD_LOGIC;
  SIGNAL and_dcpl_257 : STD_LOGIC;
  SIGNAL and_dcpl_258 : STD_LOGIC;
  SIGNAL and_dcpl_259 : STD_LOGIC;
  SIGNAL and_dcpl_260 : STD_LOGIC;
  SIGNAL and_dcpl_261 : STD_LOGIC;
  SIGNAL and_dcpl_262 : STD_LOGIC;
  SIGNAL and_dcpl_263 : STD_LOGIC;
  SIGNAL and_dcpl_264 : STD_LOGIC;
  SIGNAL and_dcpl_265 : STD_LOGIC;
  SIGNAL and_dcpl_266 : STD_LOGIC;
  SIGNAL and_dcpl_267 : STD_LOGIC;
  SIGNAL and_dcpl_268 : STD_LOGIC;
  SIGNAL and_dcpl_269 : STD_LOGIC;
  SIGNAL and_dcpl_270 : STD_LOGIC;
  SIGNAL and_dcpl_271 : STD_LOGIC;
  SIGNAL and_dcpl_273 : STD_LOGIC;
  SIGNAL and_dcpl_275 : STD_LOGIC;
  SIGNAL and_dcpl_276 : STD_LOGIC;
  SIGNAL and_dcpl_278 : STD_LOGIC;
  SIGNAL and_dcpl_279 : STD_LOGIC;
  SIGNAL and_dcpl_280 : STD_LOGIC;
  SIGNAL and_dcpl_282 : STD_LOGIC;
  SIGNAL and_dcpl_283 : STD_LOGIC;
  SIGNAL and_dcpl_284 : STD_LOGIC;
  SIGNAL and_dcpl_285 : STD_LOGIC;
  SIGNAL and_dcpl_286 : STD_LOGIC;
  SIGNAL and_dcpl_287 : STD_LOGIC;
  SIGNAL and_dcpl_288 : STD_LOGIC;
  SIGNAL and_dcpl_289 : STD_LOGIC;
  SIGNAL or_tmp_2368 : STD_LOGIC;
  SIGNAL mux_tmp_2215 : STD_LOGIC;
  SIGNAL mux_tmp_2216 : STD_LOGIC;
  SIGNAL or_tmp_2373 : STD_LOGIC;
  SIGNAL or_tmp_2381 : STD_LOGIC;
  SIGNAL mux_tmp_2223 : STD_LOGIC;
  SIGNAL mux_tmp_2226 : STD_LOGIC;
  SIGNAL and_dcpl_290 : STD_LOGIC;
  SIGNAL or_tmp_2391 : STD_LOGIC;
  SIGNAL or_tmp_2393 : STD_LOGIC;
  SIGNAL or_tmp_2395 : STD_LOGIC;
  SIGNAL mux_tmp_2244 : STD_LOGIC;
  SIGNAL or_tmp_2401 : STD_LOGIC;
  SIGNAL or_tmp_2402 : STD_LOGIC;
  SIGNAL mux_tmp_2247 : STD_LOGIC;
  SIGNAL or_tmp_2406 : STD_LOGIC;
  SIGNAL mux_tmp_2250 : STD_LOGIC;
  SIGNAL not_tmp_572 : STD_LOGIC;
  SIGNAL or_tmp_2409 : STD_LOGIC;
  SIGNAL mux_tmp_2276 : STD_LOGIC;
  SIGNAL and_dcpl_293 : STD_LOGIC;
  SIGNAL and_dcpl_294 : STD_LOGIC;
  SIGNAL and_dcpl_295 : STD_LOGIC;
  SIGNAL or_tmp_2439 : STD_LOGIC;
  SIGNAL and_tmp_24 : STD_LOGIC;
  SIGNAL nor_tmp_388 : STD_LOGIC;
  SIGNAL or_tmp_2447 : STD_LOGIC;
  SIGNAL or_tmp_2451 : STD_LOGIC;
  SIGNAL not_tmp_597 : STD_LOGIC;
  SIGNAL mux_tmp_2377 : STD_LOGIC;
  SIGNAL or_tmp_2548 : STD_LOGIC;
  SIGNAL or_tmp_2549 : STD_LOGIC;
  SIGNAL mux_tmp_2380 : STD_LOGIC;
  SIGNAL nor_tmp_399 : STD_LOGIC;
  SIGNAL mux_tmp_2381 : STD_LOGIC;
  SIGNAL mux_tmp_2382 : STD_LOGIC;
  SIGNAL not_tmp_617 : STD_LOGIC;
  SIGNAL mux_tmp_2389 : STD_LOGIC;
  SIGNAL or_tmp_2551 : STD_LOGIC;
  SIGNAL or_tmp_2552 : STD_LOGIC;
  SIGNAL mux_tmp_2400 : STD_LOGIC;
  SIGNAL nor_tmp_403 : STD_LOGIC;
  SIGNAL and_dcpl_307 : STD_LOGIC;
  SIGNAL and_dcpl_311 : STD_LOGIC;
  SIGNAL and_dcpl_313 : STD_LOGIC;
  SIGNAL and_dcpl_317 : STD_LOGIC;
  SIGNAL and_dcpl_319 : STD_LOGIC;
  SIGNAL and_dcpl_321 : STD_LOGIC;
  SIGNAL and_dcpl_323 : STD_LOGIC;
  SIGNAL and_dcpl_329 : STD_LOGIC;
  SIGNAL and_dcpl_331 : STD_LOGIC;
  SIGNAL and_dcpl_345 : STD_LOGIC;
  SIGNAL and_dcpl_346 : STD_LOGIC;
  SIGNAL mux_tmp_2449 : STD_LOGIC;
  SIGNAL mux_tmp_2450 : STD_LOGIC;
  SIGNAL or_dcpl_72 : STD_LOGIC;
  SIGNAL mux_tmp_2457 : STD_LOGIC;
  SIGNAL mux_tmp_2458 : STD_LOGIC;
  SIGNAL mux_tmp_2459 : STD_LOGIC;
  SIGNAL or_tmp_2585 : STD_LOGIC;
  SIGNAL mux_tmp_2461 : STD_LOGIC;
  SIGNAL mux_tmp_2462 : STD_LOGIC;
  SIGNAL mux_tmp_2467 : STD_LOGIC;
  SIGNAL mux_tmp_2468 : STD_LOGIC;
  SIGNAL or_tmp_2587 : STD_LOGIC;
  SIGNAL mux_tmp_2469 : STD_LOGIC;
  SIGNAL mux_tmp_2470 : STD_LOGIC;
  SIGNAL or_tmp_2588 : STD_LOGIC;
  SIGNAL mux_tmp_2474 : STD_LOGIC;
  SIGNAL nand_tmp_140 : STD_LOGIC;
  SIGNAL nor_tmp_417 : STD_LOGIC;
  SIGNAL mux_tmp_2529 : STD_LOGIC;
  SIGNAL not_tmp_662 : STD_LOGIC;
  SIGNAL mux_tmp_2538 : STD_LOGIC;
  SIGNAL not_tmp_664 : STD_LOGIC;
  SIGNAL and_dcpl_354 : STD_LOGIC;
  SIGNAL and_dcpl_357 : STD_LOGIC;
  SIGNAL and_dcpl_359 : STD_LOGIC;
  SIGNAL nor_tmp_427 : STD_LOGIC;
  SIGNAL and_dcpl_361 : STD_LOGIC;
  SIGNAL mux_tmp_2574 : STD_LOGIC;
  SIGNAL or_tmp_2638 : STD_LOGIC;
  SIGNAL mux_tmp_2583 : STD_LOGIC;
  SIGNAL and_dcpl_364 : STD_LOGIC;
  SIGNAL and_dcpl_367 : STD_LOGIC;
  SIGNAL and_dcpl_370 : STD_LOGIC;
  SIGNAL not_tmp_696 : STD_LOGIC;
  SIGNAL not_tmp_698 : STD_LOGIC;
  SIGNAL and_dcpl_372 : STD_LOGIC;
  SIGNAL mux_tmp_2612 : STD_LOGIC;
  SIGNAL not_tmp_703 : STD_LOGIC;
  SIGNAL mux_tmp_2614 : STD_LOGIC;
  SIGNAL not_tmp_706 : STD_LOGIC;
  SIGNAL or_tmp_2668 : STD_LOGIC;
  SIGNAL and_tmp_32 : STD_LOGIC;
  SIGNAL mux_tmp_2625 : STD_LOGIC;
  SIGNAL mux_tmp_2626 : STD_LOGIC;
  SIGNAL nor_tmp_459 : STD_LOGIC;
  SIGNAL mux_tmp_2653 : STD_LOGIC;
  SIGNAL nor_tmp_463 : STD_LOGIC;
  SIGNAL nor_tmp_467 : STD_LOGIC;
  SIGNAL mux_tmp_2666 : STD_LOGIC;
  SIGNAL not_tmp_729 : STD_LOGIC;
  SIGNAL mux_tmp_2689 : STD_LOGIC;
  SIGNAL mux_tmp_2713 : STD_LOGIC;
  SIGNAL mux_tmp_2714 : STD_LOGIC;
  SIGNAL mux_tmp_2720 : STD_LOGIC;
  SIGNAL or_tmp_2733 : STD_LOGIC;
  SIGNAL or_tmp_2734 : STD_LOGIC;
  SIGNAL mux_tmp_2721 : STD_LOGIC;
  SIGNAL or_tmp_2735 : STD_LOGIC;
  SIGNAL or_tmp_2736 : STD_LOGIC;
  SIGNAL mux_tmp_2724 : STD_LOGIC;
  SIGNAL nand_tmp_148 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm : STD_LOGIC;
  SIGNAL operator_64_false_1_slc_operator_64_false_1_acc_5_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_8_psp_sva_1 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_k_9_4_sva_4_0 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_cse_4_sva_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL STAGE_VEC_LOOP_j_sva_9_0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_slc_operator_64_false_acc_1_60_itm : STD_LOGIC;
  SIGNAL operator_64_false_acc_cse_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_12_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_12_psp_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_7_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_2_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_8_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_psp_sva : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_4_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_13_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_14_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_11_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_10_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_9_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_6_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_8_psp_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_13_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_cse_12_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_11_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_cse_8_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_7_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_3_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_cse_4_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_cse_14_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_9_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_cse_10_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_cse_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_15_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_cse_6_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_5_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_cse_2_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_1_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL STAGE_MAIN_LOOP_lshift_psp_1_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_cse_2_sva_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_2_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_3_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_4_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_5_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_6_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_7_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_8_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_9_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_10_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_11_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_12_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_13_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_14_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_15_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL operator_64_false_acc_cse_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL and_332_m1c : STD_LOGIC;
  SIGNAL and_334_m1c : STD_LOGIC;
  SIGNAL and_335_m1c : STD_LOGIC;
  SIGNAL and_338_m1c : STD_LOGIC;
  SIGNAL and_340_m1c : STD_LOGIC;
  SIGNAL and_342_m1c : STD_LOGIC;
  SIGNAL and_344_m1c : STD_LOGIC;
  SIGNAL and_346_m1c : STD_LOGIC;
  SIGNAL and_348_m1c : STD_LOGIC;
  SIGNAL and_350_m1c : STD_LOGIC;
  SIGNAL and_351_m1c : STD_LOGIC;
  SIGNAL and_352_m1c : STD_LOGIC;
  SIGNAL and_354_m1c : STD_LOGIC;
  SIGNAL and_356_m1c : STD_LOGIC;
  SIGNAL and_358_m1c : STD_LOGIC;
  SIGNAL nand_437_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_triosy_0_15_obj_ld_cse : STD_LOGIC;
  SIGNAL reg_ensig_cgo_cse : STD_LOGIC;
  SIGNAL nor_368_cse : STD_LOGIC;
  SIGNAL and_516_cse : STD_LOGIC;
  SIGNAL and_515_cse : STD_LOGIC;
  SIGNAL reg_COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat_cse : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL or_602_cse : STD_LOGIC;
  SIGNAL or_2500_cse : STD_LOGIC;
  SIGNAL or_2700_cse : STD_LOGIC;
  SIGNAL or_598_cse : STD_LOGIC;
  SIGNAL and_697_cse : STD_LOGIC;
  SIGNAL and_711_cse : STD_LOGIC;
  SIGNAL or_111_cse : STD_LOGIC;
  SIGNAL and_581_cse : STD_LOGIC;
  SIGNAL or_307_cse : STD_LOGIC;
  SIGNAL or_165_cse : STD_LOGIC;
  SIGNAL nor_813_cse : STD_LOGIC;
  SIGNAL or_420_cse : STD_LOGIC;
  SIGNAL and_459_cse : STD_LOGIC;
  SIGNAL and_623_cse : STD_LOGIC;
  SIGNAL and_679_cse : STD_LOGIC;
  SIGNAL or_2733_cse : STD_LOGIC;
  SIGNAL and_756_cse : STD_LOGIC;
  SIGNAL nor_936_cse : STD_LOGIC;
  SIGNAL and_475_cse : STD_LOGIC;
  SIGNAL and_613_cse : STD_LOGIC;
  SIGNAL nor_832_cse : STD_LOGIC;
  SIGNAL nand_442_cse : STD_LOGIC;
  SIGNAL or_694_cse : STD_LOGIC;
  SIGNAL or_803_cse : STD_LOGIC;
  SIGNAL or_909_cse : STD_LOGIC;
  SIGNAL or_1018_cse : STD_LOGIC;
  SIGNAL or_1124_cse : STD_LOGIC;
  SIGNAL or_1233_cse : STD_LOGIC;
  SIGNAL or_1339_cse : STD_LOGIC;
  SIGNAL or_1448_cse : STD_LOGIC;
  SIGNAL nand_169_cse : STD_LOGIC;
  SIGNAL nand_445_cse : STD_LOGIC;
  SIGNAL mux_2252_cse : STD_LOGIC;
  SIGNAL or_2573_cse : STD_LOGIC;
  SIGNAL or_204_cse : STD_LOGIC;
  SIGNAL mux_156_cse : STD_LOGIC;
  SIGNAL nor_510_cse : STD_LOGIC;
  SIGNAL mux_494_cse : STD_LOGIC;
  SIGNAL nor_569_cse : STD_LOGIC;
  SIGNAL nor_497_cse : STD_LOGIC;
  SIGNAL mux_2374_cse : STD_LOGIC;
  SIGNAL or_2549_cse : STD_LOGIC;
  SIGNAL nor_558_cse : STD_LOGIC;
  SIGNAL mux_792_cse : STD_LOGIC;
  SIGNAL mux_79_cse : STD_LOGIC;
  SIGNAL mux_1112_cse : STD_LOGIC;
  SIGNAL mux_1031_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_244_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_62_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_185_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_64_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_65_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_66_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_6_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_68_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_69_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_70_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_72_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_12_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_13_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_14_itm : STD_LOGIC;
  SIGNAL tmp_1_lpi_4_dfm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_10_lpi_4_dfm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_10_modExp_dev_1_while_mul_mut : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_5_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_51_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_52_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_77_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_54_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_79_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_80_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_81_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_57_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_83_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_84_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_85_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_86_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_87_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_88_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_89_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_9_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_91_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_92_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_137_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_94_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_139_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_140_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_141_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_97_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_143_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_144_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_145_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_146_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_147_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_148_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_149_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_13_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_131_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_132_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_197_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_134_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_199_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_200_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_201_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_137_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_203_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_204_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_205_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_206_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_207_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_208_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_209_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_17_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_171_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_172_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_257_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_174_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_259_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_260_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_261_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_177_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_263_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_264_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_265_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_266_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_267_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_268_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_269_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_21_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_211_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_212_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_317_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_214_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_319_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_320_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_321_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_217_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_323_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_324_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_325_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_326_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_327_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_328_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_329_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_25_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_251_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_252_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_377_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_254_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_379_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_380_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_381_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_257_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_383_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_384_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_385_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_386_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_387_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_388_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_389_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_29_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_291_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_292_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_437_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_294_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_439_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_440_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_441_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_297_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_443_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_444_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_445_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_446_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_447_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_448_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_449_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_33_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_331_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_332_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_497_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_334_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_499_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_500_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_501_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_337_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_503_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_504_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_505_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_506_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_507_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_508_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_509_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_37_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_371_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_372_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_557_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_374_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_559_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_560_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_561_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_377_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_563_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_564_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_565_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_566_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_567_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_568_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_569_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_41_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_411_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_412_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_617_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_414_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_619_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_620_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_621_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_417_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_623_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_624_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_625_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_626_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_627_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_628_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_629_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_45_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_451_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_452_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_677_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_454_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_679_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_680_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_681_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_457_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_683_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_684_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_685_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_686_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_687_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_688_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_689_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_49_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_491_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_492_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_737_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_494_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_739_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_740_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_741_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_497_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_743_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_744_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_745_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_746_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_747_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_748_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_749_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_53_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_531_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_532_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_797_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_534_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_799_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_800_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_801_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_537_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_803_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_804_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_805_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_806_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_807_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_808_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_809_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_57_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_571_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_572_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_857_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_574_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_859_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_860_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_861_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_577_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_863_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_864_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_865_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_866_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_867_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_868_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_869_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_61_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_611_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_612_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_917_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_614_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_919_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_920_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_921_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_617_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_923_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_924_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_925_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_926_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_927_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_928_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_929_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_psp_sva : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL p_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mux_2240_itm : STD_LOGIC;
  SIGNAL mux_2232_itm : STD_LOGIC;
  SIGNAL mux_2336_itm : STD_LOGIC;
  SIGNAL mux_2586_itm : STD_LOGIC;
  SIGNAL mux_2688_itm : STD_LOGIC;
  SIGNAL mux_2703_itm : STD_LOGIC;
  SIGNAL mux_2715_itm : STD_LOGIC;
  SIGNAL mux_2727_itm : STD_LOGIC;
  SIGNAL mux_2734_itm : STD_LOGIC;
  SIGNAL mux_2745_itm : STD_LOGIC;
  SIGNAL or_tmp_2740 : STD_LOGIC;
  SIGNAL or_tmp_2743 : STD_LOGIC;
  SIGNAL mux_tmp_2749 : STD_LOGIC;
  SIGNAL nand_tmp_150 : STD_LOGIC;
  SIGNAL and_dcpl_402 : STD_LOGIC;
  SIGNAL z_out : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL and_dcpl_418 : STD_LOGIC;
  SIGNAL z_out_1 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL and_dcpl_419 : STD_LOGIC;
  SIGNAL and_dcpl_421 : STD_LOGIC;
  SIGNAL and_dcpl_423 : STD_LOGIC;
  SIGNAL and_dcpl_424 : STD_LOGIC;
  SIGNAL and_dcpl_427 : STD_LOGIC;
  SIGNAL and_dcpl_429 : STD_LOGIC;
  SIGNAL and_dcpl_431 : STD_LOGIC;
  SIGNAL and_dcpl_432 : STD_LOGIC;
  SIGNAL and_dcpl_433 : STD_LOGIC;
  SIGNAL and_dcpl_434 : STD_LOGIC;
  SIGNAL and_dcpl_435 : STD_LOGIC;
  SIGNAL and_dcpl_436 : STD_LOGIC;
  SIGNAL and_dcpl_437 : STD_LOGIC;
  SIGNAL and_dcpl_439 : STD_LOGIC;
  SIGNAL and_dcpl_440 : STD_LOGIC;
  SIGNAL and_dcpl_441 : STD_LOGIC;
  SIGNAL and_dcpl_442 : STD_LOGIC;
  SIGNAL and_dcpl_444 : STD_LOGIC;
  SIGNAL and_dcpl_445 : STD_LOGIC;
  SIGNAL and_dcpl_449 : STD_LOGIC;
  SIGNAL and_dcpl_451 : STD_LOGIC;
  SIGNAL and_dcpl_452 : STD_LOGIC;
  SIGNAL and_dcpl_453 : STD_LOGIC;
  SIGNAL and_dcpl_454 : STD_LOGIC;
  SIGNAL and_dcpl_456 : STD_LOGIC;
  SIGNAL and_dcpl_457 : STD_LOGIC;
  SIGNAL and_dcpl_458 : STD_LOGIC;
  SIGNAL and_dcpl_462 : STD_LOGIC;
  SIGNAL and_dcpl_464 : STD_LOGIC;
  SIGNAL and_dcpl_465 : STD_LOGIC;
  SIGNAL and_dcpl_466 : STD_LOGIC;
  SIGNAL and_dcpl_468 : STD_LOGIC;
  SIGNAL and_dcpl_469 : STD_LOGIC;
  SIGNAL and_dcpl_470 : STD_LOGIC;
  SIGNAL and_dcpl_471 : STD_LOGIC;
  SIGNAL and_dcpl_474 : STD_LOGIC;
  SIGNAL and_dcpl_476 : STD_LOGIC;
  SIGNAL and_dcpl_478 : STD_LOGIC;
  SIGNAL and_dcpl_481 : STD_LOGIC;
  SIGNAL and_dcpl_483 : STD_LOGIC;
  SIGNAL and_dcpl_484 : STD_LOGIC;
  SIGNAL and_dcpl_487 : STD_LOGIC;
  SIGNAL and_dcpl_489 : STD_LOGIC;
  SIGNAL and_dcpl_490 : STD_LOGIC;
  SIGNAL and_dcpl_491 : STD_LOGIC;
  SIGNAL and_dcpl_493 : STD_LOGIC;
  SIGNAL and_dcpl_495 : STD_LOGIC;
  SIGNAL and_dcpl_496 : STD_LOGIC;
  SIGNAL and_dcpl_498 : STD_LOGIC;
  SIGNAL z_out_2 : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL and_dcpl_505 : STD_LOGIC;
  SIGNAL and_dcpl_507 : STD_LOGIC;
  SIGNAL and_dcpl_508 : STD_LOGIC;
  SIGNAL and_dcpl_509 : STD_LOGIC;
  SIGNAL and_dcpl_510 : STD_LOGIC;
  SIGNAL and_dcpl_511 : STD_LOGIC;
  SIGNAL and_dcpl_523 : STD_LOGIC;
  SIGNAL and_dcpl_525 : STD_LOGIC;
  SIGNAL and_dcpl_530 : STD_LOGIC;
  SIGNAL and_dcpl_534 : STD_LOGIC;
  SIGNAL and_dcpl_543 : STD_LOGIC;
  SIGNAL and_dcpl_544 : STD_LOGIC;
  SIGNAL z_out_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL and_dcpl_582 : STD_LOGIC;
  SIGNAL and_dcpl_584 : STD_LOGIC;
  SIGNAL and_dcpl_589 : STD_LOGIC;
  SIGNAL and_dcpl_593 : STD_LOGIC;
  SIGNAL and_dcpl_599 : STD_LOGIC;
  SIGNAL and_dcpl_621 : STD_LOGIC;
  SIGNAL z_out_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL r_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_MAIN_LOOP_acc_1_psp_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL modExp_dev_result_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_1_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_12_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_14_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_19_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_20_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_21_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_17_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_23_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_24_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_25_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_26_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_27_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_28_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_29_itm : STD_LOGIC;
  SIGNAL modExp_dev_exp_1_sva_63_9 : STD_LOGIC_VECTOR (54 DOWNTO 0);
  SIGNAL modExp_dev_exp_1_sva_8_4 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL STAGE_MAIN_LOOP_lshift_psp_1_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_10_modExp_dev_1_while_mul_mut_mx0c4 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_modExp_dev_1_while_mul_mut_mx0c5 : STD_LOGIC;
  SIGNAL STAGE_VEC_LOOP_j_sva_9_0_mx0c1 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c3 :
      STD_LOGIC;
  SIGNAL COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c4 :
      STD_LOGIC;
  SIGNAL COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c5 :
      STD_LOGIC;
  SIGNAL COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c6 :
      STD_LOGIC;
  SIGNAL COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c7 :
      STD_LOGIC;
  SIGNAL COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c8 :
      STD_LOGIC;
  SIGNAL COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c9 :
      STD_LOGIC;
  SIGNAL COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c10 :
      STD_LOGIC;
  SIGNAL COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c11 :
      STD_LOGIC;
  SIGNAL COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c12 :
      STD_LOGIC;
  SIGNAL COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c13 :
      STD_LOGIC;
  SIGNAL operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c1 : STD_LOGIC;
  SIGNAL operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c2 : STD_LOGIC;
  SIGNAL operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c3 : STD_LOGIC;
  SIGNAL operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c4 : STD_LOGIC;
  SIGNAL tmp_1_lpi_4_dfm_mx0c0 : STD_LOGIC;
  SIGNAL and_330_rgt : STD_LOGIC;
  SIGNAL or_2938_cse : STD_LOGIC;
  SIGNAL nor_554_cse : STD_LOGIC;
  SIGNAL or_2955_cse : STD_LOGIC;
  SIGNAL mux_2332_cse : STD_LOGIC;
  SIGNAL mux_2326_cse : STD_LOGIC;
  SIGNAL or_2929_cse : STD_LOGIC;
  SIGNAL mux_2829_cse : STD_LOGIC;
  SIGNAL nand_176_cse : STD_LOGIC;
  SIGNAL mux_2830_cse : STD_LOGIC;
  SIGNAL and_920_cse : STD_LOGIC;
  SIGNAL and_936_cse : STD_LOGIC;
  SIGNAL and_945_cse : STD_LOGIC;
  SIGNAL and_950_cse : STD_LOGIC;
  SIGNAL and_953_cse : STD_LOGIC;
  SIGNAL and_957_cse : STD_LOGIC;
  SIGNAL and_964_cse : STD_LOGIC;
  SIGNAL and_966_cse : STD_LOGIC;
  SIGNAL and_973_cse : STD_LOGIC;
  SIGNAL and_975_cse : STD_LOGIC;
  SIGNAL and_978_cse : STD_LOGIC;
  SIGNAL mux_2835_cse : STD_LOGIC;
  SIGNAL or_2960_cse : STD_LOGIC;
  SIGNAL and_925_cse : STD_LOGIC;
  SIGNAL and_940_cse : STD_LOGIC;
  SIGNAL and_960_cse : STD_LOGIC;
  SIGNAL and_970_cse : STD_LOGIC;
  SIGNAL mux_tmp_2812 : STD_LOGIC;
  SIGNAL mux_tmp_2813 : STD_LOGIC;
  SIGNAL mux_tmp_2815 : STD_LOGIC;
  SIGNAL mux_tmp_2823 : STD_LOGIC;
  SIGNAL mux_tmp_2824 : STD_LOGIC;
  SIGNAL nand_490_cse : STD_LOGIC;
  SIGNAL nor_1040_cse : STD_LOGIC;
  SIGNAL or_3018_cse : STD_LOGIC;
  SIGNAL nor_1039_cse : STD_LOGIC;
  SIGNAL and_694_cse : STD_LOGIC;
  SIGNAL mux_2797_itm : STD_LOGIC;
  SIGNAL mux_2545_itm : STD_LOGIC;
  SIGNAL mux_2863_itm : STD_LOGIC;
  SIGNAL operator_64_false_or_120_itm : STD_LOGIC;
  SIGNAL operator_64_false_or_121_cse : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_or_1_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_slc_acc_3_12_1_slc : STD_LOGIC_VECTOR (11 DOWNTO 0);

  SIGNAL mux_2239_nl : STD_LOGIC;
  SIGNAL mux_2238_nl : STD_LOGIC;
  SIGNAL mux_2237_nl : STD_LOGIC;
  SIGNAL mux_2236_nl : STD_LOGIC;
  SIGNAL mux_2235_nl : STD_LOGIC;
  SIGNAL mux_2234_nl : STD_LOGIC;
  SIGNAL mux_2233_nl : STD_LOGIC;
  SIGNAL mux_2231_nl : STD_LOGIC;
  SIGNAL mux_2230_nl : STD_LOGIC;
  SIGNAL mux_2229_nl : STD_LOGIC;
  SIGNAL mux_2228_nl : STD_LOGIC;
  SIGNAL mux_2227_nl : STD_LOGIC;
  SIGNAL mux_2226_nl : STD_LOGIC;
  SIGNAL mux_2225_nl : STD_LOGIC;
  SIGNAL mux_2224_nl : STD_LOGIC;
  SIGNAL mux_2223_nl : STD_LOGIC;
  SIGNAL mux_2222_nl : STD_LOGIC;
  SIGNAL mux_2221_nl : STD_LOGIC;
  SIGNAL mux_2220_nl : STD_LOGIC;
  SIGNAL mux_2219_nl : STD_LOGIC;
  SIGNAL mux_2218_nl : STD_LOGIC;
  SIGNAL mux_2217_nl : STD_LOGIC;
  SIGNAL mux_2216_nl : STD_LOGIC;
  SIGNAL mux_2215_nl : STD_LOGIC;
  SIGNAL mux_2214_nl : STD_LOGIC;
  SIGNAL mux_2213_nl : STD_LOGIC;
  SIGNAL mux_2211_nl : STD_LOGIC;
  SIGNAL mux_2210_nl : STD_LOGIC;
  SIGNAL mux_2209_nl : STD_LOGIC;
  SIGNAL mux_2208_nl : STD_LOGIC;
  SIGNAL or_2841_nl : STD_LOGIC;
  SIGNAL mux_2207_nl : STD_LOGIC;
  SIGNAL mux_2206_nl : STD_LOGIC;
  SIGNAL mux_2205_nl : STD_LOGIC;
  SIGNAL mux_2204_nl : STD_LOGIC;
  SIGNAL mux_2203_nl : STD_LOGIC;
  SIGNAL mux_2202_nl : STD_LOGIC;
  SIGNAL mux_2201_nl : STD_LOGIC;
  SIGNAL mux_2200_nl : STD_LOGIC;
  SIGNAL or_2392_nl : STD_LOGIC;
  SIGNAL mux_2199_nl : STD_LOGIC;
  SIGNAL mux_2198_nl : STD_LOGIC;
  SIGNAL mux_2197_nl : STD_LOGIC;
  SIGNAL mux_2196_nl : STD_LOGIC;
  SIGNAL mux_2195_nl : STD_LOGIC;
  SIGNAL mux_2194_nl : STD_LOGIC;
  SIGNAL mux_2192_nl : STD_LOGIC;
  SIGNAL mux_2191_nl : STD_LOGIC;
  SIGNAL mux_2189_nl : STD_LOGIC;
  SIGNAL mux_2188_nl : STD_LOGIC;
  SIGNAL mux_2187_nl : STD_LOGIC;
  SIGNAL mux_2185_nl : STD_LOGIC;
  SIGNAL mux_2184_nl : STD_LOGIC;
  SIGNAL mux_2179_nl : STD_LOGIC;
  SIGNAL mux_2173_nl : STD_LOGIC;
  SIGNAL mux_2172_nl : STD_LOGIC;
  SIGNAL mux_2171_nl : STD_LOGIC;
  SIGNAL mux_2170_nl : STD_LOGIC;
  SIGNAL mux_2168_nl : STD_LOGIC;
  SIGNAL mux_2167_nl : STD_LOGIC;
  SIGNAL mux_2166_nl : STD_LOGIC;
  SIGNAL mux_2323_nl : STD_LOGIC;
  SIGNAL mux_2322_nl : STD_LOGIC;
  SIGNAL mux_2321_nl : STD_LOGIC;
  SIGNAL mux_2320_nl : STD_LOGIC;
  SIGNAL mux_2319_nl : STD_LOGIC;
  SIGNAL mux_2318_nl : STD_LOGIC;
  SIGNAL or_2479_nl : STD_LOGIC;
  SIGNAL mux_2317_nl : STD_LOGIC;
  SIGNAL mux_2316_nl : STD_LOGIC;
  SIGNAL mux_2315_nl : STD_LOGIC;
  SIGNAL mux_2314_nl : STD_LOGIC;
  SIGNAL nand_177_nl : STD_LOGIC;
  SIGNAL mux_2313_nl : STD_LOGIC;
  SIGNAL or_2477_nl : STD_LOGIC;
  SIGNAL mux_2312_nl : STD_LOGIC;
  SIGNAL mux_2311_nl : STD_LOGIC;
  SIGNAL mux_2310_nl : STD_LOGIC;
  SIGNAL or_2476_nl : STD_LOGIC;
  SIGNAL mux_2309_nl : STD_LOGIC;
  SIGNAL nand_178_nl : STD_LOGIC;
  SIGNAL mux_2308_nl : STD_LOGIC;
  SIGNAL mux_2307_nl : STD_LOGIC;
  SIGNAL mux_2306_nl : STD_LOGIC;
  SIGNAL mux_2305_nl : STD_LOGIC;
  SIGNAL mux_2304_nl : STD_LOGIC;
  SIGNAL mux_2303_nl : STD_LOGIC;
  SIGNAL mux_2302_nl : STD_LOGIC;
  SIGNAL mux_2300_nl : STD_LOGIC;
  SIGNAL mux_2299_nl : STD_LOGIC;
  SIGNAL or_2468_nl : STD_LOGIC;
  SIGNAL mux_2297_nl : STD_LOGIC;
  SIGNAL mux_2296_nl : STD_LOGIC;
  SIGNAL or_2461_nl : STD_LOGIC;
  SIGNAL mux_2294_nl : STD_LOGIC;
  SIGNAL mux_2293_nl : STD_LOGIC;
  SIGNAL mux_2292_nl : STD_LOGIC;
  SIGNAL or_2455_nl : STD_LOGIC;
  SIGNAL mux_2339_nl : STD_LOGIC;
  SIGNAL mux_2338_nl : STD_LOGIC;
  SIGNAL mux_2337_nl : STD_LOGIC;
  SIGNAL nor_549_nl : STD_LOGIC;
  SIGNAL and_511_nl : STD_LOGIC;
  SIGNAL and_512_nl : STD_LOGIC;
  SIGNAL and_513_nl : STD_LOGIC;
  SIGNAL mux_1016_nl : STD_LOGIC;
  SIGNAL nor_548_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_2_nl : STD_LOGIC;
  SIGNAL mux_2427_nl : STD_LOGIC;
  SIGNAL nor_524_nl : STD_LOGIC;
  SIGNAL and_331_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_2_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_3_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_4_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_5_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_6_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_7_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_8_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_9_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_11_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_12_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_13_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_14_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_15_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_16_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_17_nl : STD_LOGIC;
  SIGNAL mux_2475_nl : STD_LOGIC;
  SIGNAL mux_2474_nl : STD_LOGIC;
  SIGNAL mux_2473_nl : STD_LOGIC;
  SIGNAL mux_2472_nl : STD_LOGIC;
  SIGNAL mux_2471_nl : STD_LOGIC;
  SIGNAL mux_2470_nl : STD_LOGIC;
  SIGNAL or_2623_nl : STD_LOGIC;
  SIGNAL mux_2469_nl : STD_LOGIC;
  SIGNAL or_2622_nl : STD_LOGIC;
  SIGNAL mux_2468_nl : STD_LOGIC;
  SIGNAL mux_2467_nl : STD_LOGIC;
  SIGNAL mux_2466_nl : STD_LOGIC;
  SIGNAL mux_2465_nl : STD_LOGIC;
  SIGNAL mux_2464_nl : STD_LOGIC;
  SIGNAL mux_2463_nl : STD_LOGIC;
  SIGNAL mux_2462_nl : STD_LOGIC;
  SIGNAL mux_2461_nl : STD_LOGIC;
  SIGNAL mux_2460_nl : STD_LOGIC;
  SIGNAL mux_2459_nl : STD_LOGIC;
  SIGNAL mux_2458_nl : STD_LOGIC;
  SIGNAL or_2621_nl : STD_LOGIC;
  SIGNAL mux_2457_nl : STD_LOGIC;
  SIGNAL mux_2456_nl : STD_LOGIC;
  SIGNAL mux_2455_nl : STD_LOGIC;
  SIGNAL mux_2454_nl : STD_LOGIC;
  SIGNAL mux_2453_nl : STD_LOGIC;
  SIGNAL mux_2452_nl : STD_LOGIC;
  SIGNAL mux_2450_nl : STD_LOGIC;
  SIGNAL mux_2449_nl : STD_LOGIC;
  SIGNAL mux_2448_nl : STD_LOGIC;
  SIGNAL mux_2447_nl : STD_LOGIC;
  SIGNAL mux_2446_nl : STD_LOGIC;
  SIGNAL mux_2445_nl : STD_LOGIC;
  SIGNAL mux_2444_nl : STD_LOGIC;
  SIGNAL mux_2443_nl : STD_LOGIC;
  SIGNAL mux_2442_nl : STD_LOGIC;
  SIGNAL mux_2441_nl : STD_LOGIC;
  SIGNAL mux_2437_nl : STD_LOGIC;
  SIGNAL mux_2436_nl : STD_LOGIC;
  SIGNAL mux_2435_nl : STD_LOGIC;
  SIGNAL mux_2434_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_17_nl : STD_LOGIC;
  SIGNAL modExp_dev_while_or_nl : STD_LOGIC;
  SIGNAL modExp_dev_while_or_1_nl : STD_LOGIC;
  SIGNAL nand_486_nl : STD_LOGIC;
  SIGNAL mux_2864_nl : STD_LOGIC;
  SIGNAL nor_nl : STD_LOGIC;
  SIGNAL nor_1038_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_2_nl_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL operator_64_false_and_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL operator_64_false_mux1h_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL and_421_nl : STD_LOGIC;
  SIGNAL and_422_nl : STD_LOGIC;
  SIGNAL and_423_nl : STD_LOGIC;
  SIGNAL and_424_nl : STD_LOGIC;
  SIGNAL and_425_nl : STD_LOGIC;
  SIGNAL and_426_nl : STD_LOGIC;
  SIGNAL and_427_nl : STD_LOGIC;
  SIGNAL and_428_nl : STD_LOGIC;
  SIGNAL and_429_nl : STD_LOGIC;
  SIGNAL and_430_nl : STD_LOGIC;
  SIGNAL and_431_nl : STD_LOGIC;
  SIGNAL and_432_nl : STD_LOGIC;
  SIGNAL and_433_nl : STD_LOGIC;
  SIGNAL and_434_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nand_nl : STD_LOGIC;
  SIGNAL and_435_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_acc_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL mux_2590_nl : STD_LOGIC;
  SIGNAL or_2696_nl : STD_LOGIC;
  SIGNAL mux_2587_nl : STD_LOGIC;
  SIGNAL mux_2592_nl : STD_LOGIC;
  SIGNAL mux_2591_nl : STD_LOGIC;
  SIGNAL or_2699_nl : STD_LOGIC;
  SIGNAL mux_2599_nl : STD_LOGIC;
  SIGNAL mux_2598_nl : STD_LOGIC;
  SIGNAL mux_2597_nl : STD_LOGIC;
  SIGNAL mux_2596_nl : STD_LOGIC;
  SIGNAL mux_2594_nl : STD_LOGIC;
  SIGNAL mux_2593_nl : STD_LOGIC;
  SIGNAL mux_2601_nl : STD_LOGIC;
  SIGNAL mux_2600_nl : STD_LOGIC;
  SIGNAL or_2701_nl : STD_LOGIC;
  SIGNAL mux_2612_nl : STD_LOGIC;
  SIGNAL mux_2611_nl : STD_LOGIC;
  SIGNAL and_485_nl : STD_LOGIC;
  SIGNAL mux_2616_nl : STD_LOGIC;
  SIGNAL or_2824_nl : STD_LOGIC;
  SIGNAL mux_2615_nl : STD_LOGIC;
  SIGNAL mux_2614_nl : STD_LOGIC;
  SIGNAL or_2825_nl : STD_LOGIC;
  SIGNAL nand_161_nl : STD_LOGIC;
  SIGNAL nand_162_nl : STD_LOGIC;
  SIGNAL mux_2621_nl : STD_LOGIC;
  SIGNAL or_2707_nl : STD_LOGIC;
  SIGNAL mux_2620_nl : STD_LOGIC;
  SIGNAL mux_2619_nl : STD_LOGIC;
  SIGNAL and_482_nl : STD_LOGIC;
  SIGNAL mux_2624_nl : STD_LOGIC;
  SIGNAL or_2708_nl : STD_LOGIC;
  SIGNAL mux_2623_nl : STD_LOGIC;
  SIGNAL and_480_nl : STD_LOGIC;
  SIGNAL mux_2633_nl : STD_LOGIC;
  SIGNAL mux_2632_nl : STD_LOGIC;
  SIGNAL mux_2631_nl : STD_LOGIC;
  SIGNAL mux_2630_nl : STD_LOGIC;
  SIGNAL mux_2629_nl : STD_LOGIC;
  SIGNAL mux_2628_nl : STD_LOGIC;
  SIGNAL mux_2627_nl : STD_LOGIC;
  SIGNAL mux_2626_nl : STD_LOGIC;
  SIGNAL mux_2640_nl : STD_LOGIC;
  SIGNAL mux_2639_nl : STD_LOGIC;
  SIGNAL mux_2638_nl : STD_LOGIC;
  SIGNAL mux_2637_nl : STD_LOGIC;
  SIGNAL nor_511_nl : STD_LOGIC;
  SIGNAL and_473_nl : STD_LOGIC;
  SIGNAL mux_2641_nl : STD_LOGIC;
  SIGNAL and_393_nl : STD_LOGIC;
  SIGNAL mux_2645_nl : STD_LOGIC;
  SIGNAL and_397_nl : STD_LOGIC;
  SIGNAL mux_2649_nl : STD_LOGIC;
  SIGNAL mux_2648_nl : STD_LOGIC;
  SIGNAL mux_2647_nl : STD_LOGIC;
  SIGNAL mux_2646_nl : STD_LOGIC;
  SIGNAL nor_937_nl : STD_LOGIC;
  SIGNAL and_754_nl : STD_LOGIC;
  SIGNAL and_755_nl : STD_LOGIC;
  SIGNAL mux_2657_nl : STD_LOGIC;
  SIGNAL mux_2656_nl : STD_LOGIC;
  SIGNAL mux_2655_nl : STD_LOGIC;
  SIGNAL or_196_nl : STD_LOGIC;
  SIGNAL mux_2654_nl : STD_LOGIC;
  SIGNAL mux_2653_nl : STD_LOGIC;
  SIGNAL or_2651_nl : STD_LOGIC;
  SIGNAL or_2732_nl : STD_LOGIC;
  SIGNAL mux_2670_nl : STD_LOGIC;
  SIGNAL mux_2669_nl : STD_LOGIC;
  SIGNAL mux_2668_nl : STD_LOGIC;
  SIGNAL mux_2667_nl : STD_LOGIC;
  SIGNAL mux_2666_nl : STD_LOGIC;
  SIGNAL mux_2681_nl : STD_LOGIC;
  SIGNAL mux_2680_nl : STD_LOGIC;
  SIGNAL mux_2679_nl : STD_LOGIC;
  SIGNAL mux_2678_nl : STD_LOGIC;
  SIGNAL or_2743_nl : STD_LOGIC;
  SIGNAL or_2748_nl : STD_LOGIC;
  SIGNAL mux_2692_nl : STD_LOGIC;
  SIGNAL mux_2691_nl : STD_LOGIC;
  SIGNAL nor_503_nl : STD_LOGIC;
  SIGNAL mux_2690_nl : STD_LOGIC;
  SIGNAL nor_504_nl : STD_LOGIC;
  SIGNAL and_409_nl : STD_LOGIC;
  SIGNAL mux_2708_nl : STD_LOGIC;
  SIGNAL mux_2707_nl : STD_LOGIC;
  SIGNAL mux_2706_nl : STD_LOGIC;
  SIGNAL nor_500_nl : STD_LOGIC;
  SIGNAL and_452_nl : STD_LOGIC;
  SIGNAL mux_2705_nl : STD_LOGIC;
  SIGNAL or_2755_nl : STD_LOGIC;
  SIGNAL mux_2713_nl : STD_LOGIC;
  SIGNAL mux_2712_nl : STD_LOGIC;
  SIGNAL mux_2711_nl : STD_LOGIC;
  SIGNAL nor_498_nl : STD_LOGIC;
  SIGNAL mux_2710_nl : STD_LOGIC;
  SIGNAL nor_499_nl : STD_LOGIC;
  SIGNAL and_410_nl : STD_LOGIC;
  SIGNAL mux_2722_nl : STD_LOGIC;
  SIGNAL mux_2721_nl : STD_LOGIC;
  SIGNAL mux_2720_nl : STD_LOGIC;
  SIGNAL mux_2719_nl : STD_LOGIC;
  SIGNAL mux_2718_nl : STD_LOGIC;
  SIGNAL and_636_nl : STD_LOGIC;
  SIGNAL mux_2730_nl : STD_LOGIC;
  SIGNAL mux_2729_nl : STD_LOGIC;
  SIGNAL or_2814_nl : STD_LOGIC;
  SIGNAL mux_2728_nl : STD_LOGIC;
  SIGNAL or_2815_nl : STD_LOGIC;
  SIGNAL nand_156_nl : STD_LOGIC;
  SIGNAL mux_2733_nl : STD_LOGIC;
  SIGNAL mux_2732_nl : STD_LOGIC;
  SIGNAL or_2812_nl : STD_LOGIC;
  SIGNAL mux_2731_nl : STD_LOGIC;
  SIGNAL or_411_nl : STD_LOGIC;
  SIGNAL or_2777_nl : STD_LOGIC;
  SIGNAL nand_154_nl : STD_LOGIC;
  SIGNAL and_413_nl : STD_LOGIC;
  SIGNAL and_414_nl : STD_LOGIC;
  SIGNAL mux_2736_nl : STD_LOGIC;
  SIGNAL or_2891_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_11_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_35_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_18_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_19_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_20_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_21_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_22_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_23_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_24_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_25_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_26_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_27_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_28_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_29_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_30_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_31_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_32_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_33_nl : STD_LOGIC;
  SIGNAL not_7089_nl : STD_LOGIC;
  SIGNAL mux_2893_nl : STD_LOGIC;
  SIGNAL mux_2892_nl : STD_LOGIC;
  SIGNAL nand_nl : STD_LOGIC;
  SIGNAL mux_2891_nl : STD_LOGIC;
  SIGNAL mux_2890_nl : STD_LOGIC;
  SIGNAL nor_1035_nl : STD_LOGIC;
  SIGNAL mux_2889_nl : STD_LOGIC;
  SIGNAL mux_2896_nl : STD_LOGIC;
  SIGNAL or_3019_nl : STD_LOGIC;
  SIGNAL mux_2888_nl : STD_LOGIC;
  SIGNAL mux_2887_nl : STD_LOGIC;
  SIGNAL mux_2895_nl : STD_LOGIC;
  SIGNAL mux_2885_nl : STD_LOGIC;
  SIGNAL or_3017_nl : STD_LOGIC;
  SIGNAL mux_2884_nl : STD_LOGIC;
  SIGNAL mux_2883_nl : STD_LOGIC;
  SIGNAL mux_2882_nl : STD_LOGIC;
  SIGNAL mux_2881_nl : STD_LOGIC;
  SIGNAL mux_2880_nl : STD_LOGIC;
  SIGNAL mux_2879_nl : STD_LOGIC;
  SIGNAL mux_2878_nl : STD_LOGIC;
  SIGNAL mux_2875_nl : STD_LOGIC;
  SIGNAL mux_2874_nl : STD_LOGIC;
  SIGNAL or_3011_nl : STD_LOGIC;
  SIGNAL mux_2873_nl : STD_LOGIC;
  SIGNAL or_3008_nl : STD_LOGIC;
  SIGNAL mux_2872_nl : STD_LOGIC;
  SIGNAL mux_2871_nl : STD_LOGIC;
  SIGNAL mux_2870_nl : STD_LOGIC;
  SIGNAL mux_2869_nl : STD_LOGIC;
  SIGNAL or_3006_nl : STD_LOGIC;
  SIGNAL mux_2867_nl : STD_LOGIC;
  SIGNAL or_3005_nl : STD_LOGIC;
  SIGNAL or_3004_nl : STD_LOGIC;
  SIGNAL or_424_nl : STD_LOGIC;
  SIGNAL or_444_nl : STD_LOGIC;
  SIGNAL or_533_nl : STD_LOGIC;
  SIGNAL mux_1049_nl : STD_LOGIC;
  SIGNAL mux_1048_nl : STD_LOGIC;
  SIGNAL or_2836_nl : STD_LOGIC;
  SIGNAL nand_389_nl : STD_LOGIC;
  SIGNAL nand_390_nl : STD_LOGIC;
  SIGNAL nand_391_nl : STD_LOGIC;
  SIGNAL nor_809_nl : STD_LOGIC;
  SIGNAL nor_810_nl : STD_LOGIC;
  SIGNAL and_741_nl : STD_LOGIC;
  SIGNAL nor_797_nl : STD_LOGIC;
  SIGNAL mux_1085_nl : STD_LOGIC;
  SIGNAL nor_775_nl : STD_LOGIC;
  SIGNAL nor_776_nl : STD_LOGIC;
  SIGNAL mux_1111_nl : STD_LOGIC;
  SIGNAL or_735_nl : STD_LOGIC;
  SIGNAL mux_1153_nl : STD_LOGIC;
  SIGNAL nor_763_nl : STD_LOGIC;
  SIGNAL nor_764_nl : STD_LOGIC;
  SIGNAL mux_1221_nl : STD_LOGIC;
  SIGNAL nor_751_nl : STD_LOGIC;
  SIGNAL nor_752_nl : STD_LOGIC;
  SIGNAL mux_1289_nl : STD_LOGIC;
  SIGNAL nor_739_nl : STD_LOGIC;
  SIGNAL nor_740_nl : STD_LOGIC;
  SIGNAL mux_1357_nl : STD_LOGIC;
  SIGNAL nor_727_nl : STD_LOGIC;
  SIGNAL nor_728_nl : STD_LOGIC;
  SIGNAL mux_1425_nl : STD_LOGIC;
  SIGNAL nor_715_nl : STD_LOGIC;
  SIGNAL nor_716_nl : STD_LOGIC;
  SIGNAL mux_1493_nl : STD_LOGIC;
  SIGNAL nor_703_nl : STD_LOGIC;
  SIGNAL nor_704_nl : STD_LOGIC;
  SIGNAL mux_1561_nl : STD_LOGIC;
  SIGNAL nor_691_nl : STD_LOGIC;
  SIGNAL nor_692_nl : STD_LOGIC;
  SIGNAL mux_1629_nl : STD_LOGIC;
  SIGNAL nor_679_nl : STD_LOGIC;
  SIGNAL nor_680_nl : STD_LOGIC;
  SIGNAL mux_1697_nl : STD_LOGIC;
  SIGNAL nor_667_nl : STD_LOGIC;
  SIGNAL nor_668_nl : STD_LOGIC;
  SIGNAL mux_1765_nl : STD_LOGIC;
  SIGNAL nor_655_nl : STD_LOGIC;
  SIGNAL nor_656_nl : STD_LOGIC;
  SIGNAL mux_1833_nl : STD_LOGIC;
  SIGNAL nor_643_nl : STD_LOGIC;
  SIGNAL nor_644_nl : STD_LOGIC;
  SIGNAL mux_1901_nl : STD_LOGIC;
  SIGNAL nor_631_nl : STD_LOGIC;
  SIGNAL nor_632_nl : STD_LOGIC;
  SIGNAL mux_1969_nl : STD_LOGIC;
  SIGNAL nor_619_nl : STD_LOGIC;
  SIGNAL nor_620_nl : STD_LOGIC;
  SIGNAL mux_2037_nl : STD_LOGIC;
  SIGNAL nor_607_nl : STD_LOGIC;
  SIGNAL nor_608_nl : STD_LOGIC;
  SIGNAL mux_2105_nl : STD_LOGIC;
  SIGNAL nor_595_nl : STD_LOGIC;
  SIGNAL nor_596_nl : STD_LOGIC;
  SIGNAL or_2390_nl : STD_LOGIC;
  SIGNAL mux_2174_nl : STD_LOGIC;
  SIGNAL mux_2177_nl : STD_LOGIC;
  SIGNAL mux_2176_nl : STD_LOGIC;
  SIGNAL or_2412_nl : STD_LOGIC;
  SIGNAL or_2411_nl : STD_LOGIC;
  SIGNAL or_2634_nl : STD_LOGIC;
  SIGNAL or_2431_nl : STD_LOGIC;
  SIGNAL nand_180_nl : STD_LOGIC;
  SIGNAL or_2464_nl : STD_LOGIC;
  SIGNAL or_2462_nl : STD_LOGIC;
  SIGNAL nor_552_nl : STD_LOGIC;
  SIGNAL or_2486_nl : STD_LOGIC;
  SIGNAL or_2484_nl : STD_LOGIC;
  SIGNAL nor_550_nl : STD_LOGIC;
  SIGNAL nor_551_nl : STD_LOGIC;
  SIGNAL mux_2335_nl : STD_LOGIC;
  SIGNAL or_2498_nl : STD_LOGIC;
  SIGNAL mux_2334_nl : STD_LOGIC;
  SIGNAL or_2497_nl : STD_LOGIC;
  SIGNAL or_2495_nl : STD_LOGIC;
  SIGNAL mux_2333_nl : STD_LOGIC;
  SIGNAL nand_120_nl : STD_LOGIC;
  SIGNAL or_2492_nl : STD_LOGIC;
  SIGNAL mux_2331_nl : STD_LOGIC;
  SIGNAL or_2491_nl : STD_LOGIC;
  SIGNAL mux_2330_nl : STD_LOGIC;
  SIGNAL mux_2329_nl : STD_LOGIC;
  SIGNAL mux_2328_nl : STD_LOGIC;
  SIGNAL or_2489_nl : STD_LOGIC;
  SIGNAL or_2488_nl : STD_LOGIC;
  SIGNAL mux_2325_nl : STD_LOGIC;
  SIGNAL nand_175_nl : STD_LOGIC;
  SIGNAL mux_2324_nl : STD_LOGIC;
  SIGNAL or_2482_nl : STD_LOGIC;
  SIGNAL or_2480_nl : STD_LOGIC;
  SIGNAL mux_2358_nl : STD_LOGIC;
  SIGNAL mux_2357_nl : STD_LOGIC;
  SIGNAL nor_541_nl : STD_LOGIC;
  SIGNAL nor_542_nl : STD_LOGIC;
  SIGNAL mux_2356_nl : STD_LOGIC;
  SIGNAL and_506_nl : STD_LOGIC;
  SIGNAL mux_2355_nl : STD_LOGIC;
  SIGNAL or_2521_nl : STD_LOGIC;
  SIGNAL mux_2354_nl : STD_LOGIC;
  SIGNAL nor_825_nl : STD_LOGIC;
  SIGNAL nor_544_nl : STD_LOGIC;
  SIGNAL mux_2353_nl : STD_LOGIC;
  SIGNAL or_2518_nl : STD_LOGIC;
  SIGNAL mux_2352_nl : STD_LOGIC;
  SIGNAL mux_2351_nl : STD_LOGIC;
  SIGNAL nor_545_nl : STD_LOGIC;
  SIGNAL mux_2350_nl : STD_LOGIC;
  SIGNAL or_2831_nl : STD_LOGIC;
  SIGNAL and_507_nl : STD_LOGIC;
  SIGNAL mux_2348_nl : STD_LOGIC;
  SIGNAL or_2510_nl : STD_LOGIC;
  SIGNAL and_508_nl : STD_LOGIC;
  SIGNAL mux_2347_nl : STD_LOGIC;
  SIGNAL nor_546_nl : STD_LOGIC;
  SIGNAL nor_547_nl : STD_LOGIC;
  SIGNAL or_2555_nl : STD_LOGIC;
  SIGNAL nand_420_nl : STD_LOGIC;
  SIGNAL or_2612_nl : STD_LOGIC;
  SIGNAL mux_2439_nl : STD_LOGIC;
  SIGNAL mux_2438_nl : STD_LOGIC;
  SIGNAL mux_2511_nl : STD_LOGIC;
  SIGNAL mux_2507_nl : STD_LOGIC;
  SIGNAL nand_137_nl : STD_LOGIC;
  SIGNAL mux_2524_nl : STD_LOGIC;
  SIGNAL mux_2531_nl : STD_LOGIC;
  SIGNAL and_494_nl : STD_LOGIC;
  SIGNAL nor_516_nl : STD_LOGIC;
  SIGNAL and_489_nl : STD_LOGIC;
  SIGNAL mux_2585_nl : STD_LOGIC;
  SIGNAL mux_2584_nl : STD_LOGIC;
  SIGNAL mux_2583_nl : STD_LOGIC;
  SIGNAL mux_2582_nl : STD_LOGIC;
  SIGNAL mux_2581_nl : STD_LOGIC;
  SIGNAL mux_2610_nl : STD_LOGIC;
  SIGNAL mux_2609_nl : STD_LOGIC;
  SIGNAL mux_2608_nl : STD_LOGIC;
  SIGNAL mux_2607_nl : STD_LOGIC;
  SIGNAL mux_2606_nl : STD_LOGIC;
  SIGNAL or_2877_nl : STD_LOGIC;
  SIGNAL mux_2605_nl : STD_LOGIC;
  SIGNAL mux_2604_nl : STD_LOGIC;
  SIGNAL mux_2603_nl : STD_LOGIC;
  SIGNAL mux_2602_nl : STD_LOGIC;
  SIGNAL or_2604_nl : STD_LOGIC;
  SIGNAL mux_2613_nl : STD_LOGIC;
  SIGNAL mux_2618_nl : STD_LOGIC;
  SIGNAL mux_2617_nl : STD_LOGIC;
  SIGNAL and_483_nl : STD_LOGIC;
  SIGNAL mux_2622_nl : STD_LOGIC;
  SIGNAL nor_871_nl : STD_LOGIC;
  SIGNAL and_684_nl : STD_LOGIC;
  SIGNAL mux_2636_nl : STD_LOGIC;
  SIGNAL or_2712_nl : STD_LOGIC;
  SIGNAL mux_2635_nl : STD_LOGIC;
  SIGNAL mux_2644_nl : STD_LOGIC;
  SIGNAL nor_940_nl : STD_LOGIC;
  SIGNAL mux_2643_nl : STD_LOGIC;
  SIGNAL or_2719_nl : STD_LOGIC;
  SIGNAL or_2900_nl : STD_LOGIC;
  SIGNAL mux_2642_nl : STD_LOGIC;
  SIGNAL and_395_nl : STD_LOGIC;
  SIGNAL mux_2651_nl : STD_LOGIC;
  SIGNAL and_400_nl : STD_LOGIC;
  SIGNAL mux_2650_nl : STD_LOGIC;
  SIGNAL mux_2661_nl : STD_LOGIC;
  SIGNAL and_403_nl : STD_LOGIC;
  SIGNAL mux_2660_nl : STD_LOGIC;
  SIGNAL mux_2659_nl : STD_LOGIC;
  SIGNAL mux_2664_nl : STD_LOGIC;
  SIGNAL mux_2674_nl : STD_LOGIC;
  SIGNAL or_2740_nl : STD_LOGIC;
  SIGNAL mux_2673_nl : STD_LOGIC;
  SIGNAL or_2737_nl : STD_LOGIC;
  SIGNAL mux_2672_nl : STD_LOGIC;
  SIGNAL or_2735_nl : STD_LOGIC;
  SIGNAL mux_2687_nl : STD_LOGIC;
  SIGNAL mux_2686_nl : STD_LOGIC;
  SIGNAL mux_2685_nl : STD_LOGIC;
  SIGNAL or_2747_nl : STD_LOGIC;
  SIGNAL mux_2684_nl : STD_LOGIC;
  SIGNAL and_461_nl : STD_LOGIC;
  SIGNAL mux_2702_nl : STD_LOGIC;
  SIGNAL mux_2701_nl : STD_LOGIC;
  SIGNAL mux_2700_nl : STD_LOGIC;
  SIGNAL mux_2699_nl : STD_LOGIC;
  SIGNAL mux_2698_nl : STD_LOGIC;
  SIGNAL mux_2697_nl : STD_LOGIC;
  SIGNAL mux_2696_nl : STD_LOGIC;
  SIGNAL mux_2695_nl : STD_LOGIC;
  SIGNAL or_2762_nl : STD_LOGIC;
  SIGNAL mux_2726_nl : STD_LOGIC;
  SIGNAL mux_2725_nl : STD_LOGIC;
  SIGNAL mux_2724_nl : STD_LOGIC;
  SIGNAL nor_494_nl : STD_LOGIC;
  SIGNAL and_444_nl : STD_LOGIC;
  SIGNAL and_445_nl : STD_LOGIC;
  SIGNAL and_412_nl : STD_LOGIC;
  SIGNAL mux_2739_nl : STD_LOGIC;
  SIGNAL mux_2744_nl : STD_LOGIC;
  SIGNAL mux_2743_nl : STD_LOGIC;
  SIGNAL mux_2742_nl : STD_LOGIC;
  SIGNAL mux_2741_nl : STD_LOGIC;
  SIGNAL nor_490_nl : STD_LOGIC;
  SIGNAL mux_2763_nl : STD_LOGIC;
  SIGNAL mux_2762_nl : STD_LOGIC;
  SIGNAL nand_145_nl : STD_LOGIC;
  SIGNAL mux_2783_nl : STD_LOGIC;
  SIGNAL mux_2782_nl : STD_LOGIC;
  SIGNAL mux_2796_nl : STD_LOGIC;
  SIGNAL mux_2795_nl : STD_LOGIC;
  SIGNAL mux_2794_nl : STD_LOGIC;
  SIGNAL mux_2793_nl : STD_LOGIC;
  SIGNAL mux_2792_nl : STD_LOGIC;
  SIGNAL mux_2791_nl : STD_LOGIC;
  SIGNAL mux_2790_nl : STD_LOGIC;
  SIGNAL mux_2789_nl : STD_LOGIC;
  SIGNAL mux_2788_nl : STD_LOGIC;
  SIGNAL mux_2787_nl : STD_LOGIC;
  SIGNAL mux_2786_nl : STD_LOGIC;
  SIGNAL mux_2785_nl : STD_LOGIC;
  SIGNAL mux_2784_nl : STD_LOGIC;
  SIGNAL mux_2781_nl : STD_LOGIC;
  SIGNAL nand_147_nl : STD_LOGIC;
  SIGNAL mux_2780_nl : STD_LOGIC;
  SIGNAL mux_2779_nl : STD_LOGIC;
  SIGNAL mux_2778_nl : STD_LOGIC;
  SIGNAL mux_2777_nl : STD_LOGIC;
  SIGNAL mux_2776_nl : STD_LOGIC;
  SIGNAL nand_146_nl : STD_LOGIC;
  SIGNAL mux_2774_nl : STD_LOGIC;
  SIGNAL mux_2773_nl : STD_LOGIC;
  SIGNAL mux_2770_nl : STD_LOGIC;
  SIGNAL mux_2769_nl : STD_LOGIC;
  SIGNAL mux_2768_nl : STD_LOGIC;
  SIGNAL nor_489_nl : STD_LOGIC;
  SIGNAL mux_2767_nl : STD_LOGIC;
  SIGNAL mux_2371_nl : STD_LOGIC;
  SIGNAL mux_2370_nl : STD_LOGIC;
  SIGNAL and_504_nl : STD_LOGIC;
  SIGNAL nor_534_nl : STD_LOGIC;
  SIGNAL mux_2369_nl : STD_LOGIC;
  SIGNAL or_2547_nl : STD_LOGIC;
  SIGNAL nand_126_nl : STD_LOGIC;
  SIGNAL and_505_nl : STD_LOGIC;
  SIGNAL mux_2367_nl : STD_LOGIC;
  SIGNAL nor_535_nl : STD_LOGIC;
  SIGNAL nor_536_nl : STD_LOGIC;
  SIGNAL mux_2366_nl : STD_LOGIC;
  SIGNAL nor_537_nl : STD_LOGIC;
  SIGNAL mux_2365_nl : STD_LOGIC;
  SIGNAL or_2539_nl : STD_LOGIC;
  SIGNAL mux_2364_nl : STD_LOGIC;
  SIGNAL mux_2362_nl : STD_LOGIC;
  SIGNAL nor_538_nl : STD_LOGIC;
  SIGNAL mux_2361_nl : STD_LOGIC;
  SIGNAL or_2531_nl : STD_LOGIC;
  SIGNAL or_2530_nl : STD_LOGIC;
  SIGNAL mux_2360_nl : STD_LOGIC;
  SIGNAL nor_539_nl : STD_LOGIC;
  SIGNAL nor_540_nl : STD_LOGIC;
  SIGNAL mux_2385_nl : STD_LOGIC;
  SIGNAL mux_2384_nl : STD_LOGIC;
  SIGNAL nor_525_nl : STD_LOGIC;
  SIGNAL mux_2383_nl : STD_LOGIC;
  SIGNAL mux_2382_nl : STD_LOGIC;
  SIGNAL or_2571_nl : STD_LOGIC;
  SIGNAL or_2625_nl : STD_LOGIC;
  SIGNAL nand_172_nl : STD_LOGIC;
  SIGNAL and_501_nl : STD_LOGIC;
  SIGNAL mux_2381_nl : STD_LOGIC;
  SIGNAL nor_526_nl : STD_LOGIC;
  SIGNAL nor_527_nl : STD_LOGIC;
  SIGNAL mux_2380_nl : STD_LOGIC;
  SIGNAL nor_528_nl : STD_LOGIC;
  SIGNAL and_502_nl : STD_LOGIC;
  SIGNAL mux_2379_nl : STD_LOGIC;
  SIGNAL or_2560_nl : STD_LOGIC;
  SIGNAL mux_2378_nl : STD_LOGIC;
  SIGNAL mux_2377_nl : STD_LOGIC;
  SIGNAL and_503_nl : STD_LOGIC;
  SIGNAL mux_2376_nl : STD_LOGIC;
  SIGNAL nor_529_nl : STD_LOGIC;
  SIGNAL nor_530_nl : STD_LOGIC;
  SIGNAL mux_2375_nl : STD_LOGIC;
  SIGNAL nor_532_nl : STD_LOGIC;
  SIGNAL nor_533_nl : STD_LOGIC;
  SIGNAL mux_2373_nl : STD_LOGIC;
  SIGNAL or_2550_nl : STD_LOGIC;
  SIGNAL mux_2544_nl : STD_LOGIC;
  SIGNAL mux_2543_nl : STD_LOGIC;
  SIGNAL mux_2542_nl : STD_LOGIC;
  SIGNAL mux_2541_nl : STD_LOGIC;
  SIGNAL or_2664_nl : STD_LOGIC;
  SIGNAL mux_2540_nl : STD_LOGIC;
  SIGNAL mux_2539_nl : STD_LOGIC;
  SIGNAL mux_2538_nl : STD_LOGIC;
  SIGNAL mux_2537_nl : STD_LOGIC;
  SIGNAL mux_2536_nl : STD_LOGIC;
  SIGNAL mux_2535_nl : STD_LOGIC;
  SIGNAL mux_2534_nl : STD_LOGIC;
  SIGNAL mux_2533_nl : STD_LOGIC;
  SIGNAL mux_2532_nl : STD_LOGIC;
  SIGNAL mux_2530_nl : STD_LOGIC;
  SIGNAL nand_139_nl : STD_LOGIC;
  SIGNAL mux_2529_nl : STD_LOGIC;
  SIGNAL mux_2528_nl : STD_LOGIC;
  SIGNAL mux_2527_nl : STD_LOGIC;
  SIGNAL mux_2526_nl : STD_LOGIC;
  SIGNAL nand_138_nl : STD_LOGIC;
  SIGNAL mux_2523_nl : STD_LOGIC;
  SIGNAL mux_2522_nl : STD_LOGIC;
  SIGNAL mux_2517_nl : STD_LOGIC;
  SIGNAL mux_2516_nl : STD_LOGIC;
  SIGNAL mux_2515_nl : STD_LOGIC;
  SIGNAL nor_520_nl : STD_LOGIC;
  SIGNAL mux_2514_nl : STD_LOGIC;
  SIGNAL and_125_nl : STD_LOGIC;
  SIGNAL mux_1051_nl : STD_LOGIC;
  SIGNAL or_508_nl : STD_LOGIC;
  SIGNAL and_132_nl : STD_LOGIC;
  SIGNAL and_136_nl : STD_LOGIC;
  SIGNAL and_139_nl : STD_LOGIC;
  SIGNAL mux_1052_nl : STD_LOGIC;
  SIGNAL nor_811_nl : STD_LOGIC;
  SIGNAL nor_812_nl : STD_LOGIC;
  SIGNAL and_144_nl : STD_LOGIC;
  SIGNAL and_149_nl : STD_LOGIC;
  SIGNAL mux_1054_nl : STD_LOGIC;
  SIGNAL and_556_nl : STD_LOGIC;
  SIGNAL nor_808_nl : STD_LOGIC;
  SIGNAL and_151_nl : STD_LOGIC;
  SIGNAL mux_1055_nl : STD_LOGIC;
  SIGNAL nor_806_nl : STD_LOGIC;
  SIGNAL nor_807_nl : STD_LOGIC;
  SIGNAL and_156_nl : STD_LOGIC;
  SIGNAL mux_1056_nl : STD_LOGIC;
  SIGNAL nor_804_nl : STD_LOGIC;
  SIGNAL nor_805_nl : STD_LOGIC;
  SIGNAL and_159_nl : STD_LOGIC;
  SIGNAL mux_1057_nl : STD_LOGIC;
  SIGNAL nor_802_nl : STD_LOGIC;
  SIGNAL nor_803_nl : STD_LOGIC;
  SIGNAL and_163_nl : STD_LOGIC;
  SIGNAL mux_1058_nl : STD_LOGIC;
  SIGNAL and_555_nl : STD_LOGIC;
  SIGNAL nor_801_nl : STD_LOGIC;
  SIGNAL and_171_nl : STD_LOGIC;
  SIGNAL and_175_nl : STD_LOGIC;
  SIGNAL mux_1059_nl : STD_LOGIC;
  SIGNAL nor_799_nl : STD_LOGIC;
  SIGNAL nor_800_nl : STD_LOGIC;
  SIGNAL and_179_nl : STD_LOGIC;
  SIGNAL mux_1060_nl : STD_LOGIC;
  SIGNAL nor_798_nl : STD_LOGIC;
  SIGNAL and_554_nl : STD_LOGIC;
  SIGNAL and_184_nl : STD_LOGIC;
  SIGNAL and_188_nl : STD_LOGIC;
  SIGNAL and_191_nl : STD_LOGIC;
  SIGNAL mux_1062_nl : STD_LOGIC;
  SIGNAL nor_795_nl : STD_LOGIC;
  SIGNAL nor_796_nl : STD_LOGIC;
  SIGNAL and_196_nl : STD_LOGIC;
  SIGNAL mux_1063_nl : STD_LOGIC;
  SIGNAL nor_793_nl : STD_LOGIC;
  SIGNAL nor_794_nl : STD_LOGIC;
  SIGNAL and_200_nl : STD_LOGIC;
  SIGNAL mux_1064_nl : STD_LOGIC;
  SIGNAL and_552_nl : STD_LOGIC;
  SIGNAL nor_792_nl : STD_LOGIC;
  SIGNAL and_205_nl : STD_LOGIC;
  SIGNAL mux_1065_nl : STD_LOGIC;
  SIGNAL nor_790_nl : STD_LOGIC;
  SIGNAL nor_791_nl : STD_LOGIC;
  SIGNAL and_208_nl : STD_LOGIC;
  SIGNAL mux_1066_nl : STD_LOGIC;
  SIGNAL nor_788_nl : STD_LOGIC;
  SIGNAL nor_789_nl : STD_LOGIC;
  SIGNAL and_213_nl : STD_LOGIC;
  SIGNAL and_218_nl : STD_LOGIC;
  SIGNAL and_223_nl : STD_LOGIC;
  SIGNAL and_227_nl : STD_LOGIC;
  SIGNAL mux_1067_nl : STD_LOGIC;
  SIGNAL nor_786_nl : STD_LOGIC;
  SIGNAL and_762_nl : STD_LOGIC;
  SIGNAL and_231_nl : STD_LOGIC;
  SIGNAL mux_1068_nl : STD_LOGIC;
  SIGNAL and_551_nl : STD_LOGIC;
  SIGNAL nor_785_nl : STD_LOGIC;
  SIGNAL and_234_nl : STD_LOGIC;
  SIGNAL mux_1069_nl : STD_LOGIC;
  SIGNAL and_237_nl : STD_LOGIC;
  SIGNAL mux_1070_nl : STD_LOGIC;
  SIGNAL and_550_nl : STD_LOGIC;
  SIGNAL nor_784_nl : STD_LOGIC;
  SIGNAL and_240_nl : STD_LOGIC;
  SIGNAL mux_1071_nl : STD_LOGIC;
  SIGNAL nor_782_nl : STD_LOGIC;
  SIGNAL nor_783_nl : STD_LOGIC;
  SIGNAL and_245_nl : STD_LOGIC;
  SIGNAL mux_1072_nl : STD_LOGIC;
  SIGNAL nor_781_nl : STD_LOGIC;
  SIGNAL and_549_nl : STD_LOGIC;
  SIGNAL and_249_nl : STD_LOGIC;
  SIGNAL mux_1073_nl : STD_LOGIC;
  SIGNAL nor_779_nl : STD_LOGIC;
  SIGNAL nor_780_nl : STD_LOGIC;
  SIGNAL and_250_nl : STD_LOGIC;
  SIGNAL and_254_nl : STD_LOGIC;
  SIGNAL mux_1074_nl : STD_LOGIC;
  SIGNAL nor_777_nl : STD_LOGIC;
  SIGNAL nor_778_nl : STD_LOGIC;
  SIGNAL mux_1107_nl : STD_LOGIC;
  SIGNAL mux_1106_nl : STD_LOGIC;
  SIGNAL mux_1105_nl : STD_LOGIC;
  SIGNAL nand_18_nl : STD_LOGIC;
  SIGNAL mux_1104_nl : STD_LOGIC;
  SIGNAL mux_1103_nl : STD_LOGIC;
  SIGNAL nor_765_nl : STD_LOGIC;
  SIGNAL nor_766_nl : STD_LOGIC;
  SIGNAL mux_1102_nl : STD_LOGIC;
  SIGNAL nor_767_nl : STD_LOGIC;
  SIGNAL nor_768_nl : STD_LOGIC;
  SIGNAL mux_1101_nl : STD_LOGIC;
  SIGNAL nand_17_nl : STD_LOGIC;
  SIGNAL mux_1100_nl : STD_LOGIC;
  SIGNAL nor_769_nl : STD_LOGIC;
  SIGNAL nor_770_nl : STD_LOGIC;
  SIGNAL mux_1099_nl : STD_LOGIC;
  SIGNAL mux_1098_nl : STD_LOGIC;
  SIGNAL or_711_nl : STD_LOGIC;
  SIGNAL or_709_nl : STD_LOGIC;
  SIGNAL or_708_nl : STD_LOGIC;
  SIGNAL mux_1097_nl : STD_LOGIC;
  SIGNAL or_707_nl : STD_LOGIC;
  SIGNAL mux_1096_nl : STD_LOGIC;
  SIGNAL mux_1095_nl : STD_LOGIC;
  SIGNAL or_706_nl : STD_LOGIC;
  SIGNAL or_705_nl : STD_LOGIC;
  SIGNAL mux_1094_nl : STD_LOGIC;
  SIGNAL or_703_nl : STD_LOGIC;
  SIGNAL or_701_nl : STD_LOGIC;
  SIGNAL mux_1093_nl : STD_LOGIC;
  SIGNAL or_699_nl : STD_LOGIC;
  SIGNAL mux_1092_nl : STD_LOGIC;
  SIGNAL or_698_nl : STD_LOGIC;
  SIGNAL or_697_nl : STD_LOGIC;
  SIGNAL or_696_nl : STD_LOGIC;
  SIGNAL mux_1091_nl : STD_LOGIC;
  SIGNAL mux_1090_nl : STD_LOGIC;
  SIGNAL mux_1089_nl : STD_LOGIC;
  SIGNAL mux_1088_nl : STD_LOGIC;
  SIGNAL mux_1087_nl : STD_LOGIC;
  SIGNAL or_692_nl : STD_LOGIC;
  SIGNAL mux_1086_nl : STD_LOGIC;
  SIGNAL or_691_nl : STD_LOGIC;
  SIGNAL nand_15_nl : STD_LOGIC;
  SIGNAL mux_1084_nl : STD_LOGIC;
  SIGNAL mux_1083_nl : STD_LOGIC;
  SIGNAL nor_771_nl : STD_LOGIC;
  SIGNAL nor_772_nl : STD_LOGIC;
  SIGNAL mux_1082_nl : STD_LOGIC;
  SIGNAL nor_773_nl : STD_LOGIC;
  SIGNAL nor_774_nl : STD_LOGIC;
  SIGNAL mux_1081_nl : STD_LOGIC;
  SIGNAL mux_1080_nl : STD_LOGIC;
  SIGNAL mux_1079_nl : STD_LOGIC;
  SIGNAL or_680_nl : STD_LOGIC;
  SIGNAL mux_1078_nl : STD_LOGIC;
  SIGNAL or_678_nl : STD_LOGIC;
  SIGNAL or_676_nl : STD_LOGIC;
  SIGNAL or_675_nl : STD_LOGIC;
  SIGNAL mux_1077_nl : STD_LOGIC;
  SIGNAL or_674_nl : STD_LOGIC;
  SIGNAL or_673_nl : STD_LOGIC;
  SIGNAL or_672_nl : STD_LOGIC;
  SIGNAL mux_1076_nl : STD_LOGIC;
  SIGNAL mux_1075_nl : STD_LOGIC;
  SIGNAL or_671_nl : STD_LOGIC;
  SIGNAL or_670_nl : STD_LOGIC;
  SIGNAL or_668_nl : STD_LOGIC;
  SIGNAL mux_1142_nl : STD_LOGIC;
  SIGNAL mux_1141_nl : STD_LOGIC;
  SIGNAL mux_1140_nl : STD_LOGIC;
  SIGNAL mux_1139_nl : STD_LOGIC;
  SIGNAL or_775_nl : STD_LOGIC;
  SIGNAL mux_1138_nl : STD_LOGIC;
  SIGNAL or_773_nl : STD_LOGIC;
  SIGNAL mux_1137_nl : STD_LOGIC;
  SIGNAL or_772_nl : STD_LOGIC;
  SIGNAL or_771_nl : STD_LOGIC;
  SIGNAL mux_1136_nl : STD_LOGIC;
  SIGNAL mux_1135_nl : STD_LOGIC;
  SIGNAL mux_1134_nl : STD_LOGIC;
  SIGNAL or_770_nl : STD_LOGIC;
  SIGNAL or_768_nl : STD_LOGIC;
  SIGNAL or_766_nl : STD_LOGIC;
  SIGNAL or_764_nl : STD_LOGIC;
  SIGNAL mux_1133_nl : STD_LOGIC;
  SIGNAL mux_1132_nl : STD_LOGIC;
  SIGNAL mux_1131_nl : STD_LOGIC;
  SIGNAL mux_1130_nl : STD_LOGIC;
  SIGNAL or_763_nl : STD_LOGIC;
  SIGNAL or_762_nl : STD_LOGIC;
  SIGNAL or_761_nl : STD_LOGIC;
  SIGNAL or_760_nl : STD_LOGIC;
  SIGNAL mux_1129_nl : STD_LOGIC;
  SIGNAL mux_1128_nl : STD_LOGIC;
  SIGNAL or_758_nl : STD_LOGIC;
  SIGNAL mux_1127_nl : STD_LOGIC;
  SIGNAL or_757_nl : STD_LOGIC;
  SIGNAL or_756_nl : STD_LOGIC;
  SIGNAL or_755_nl : STD_LOGIC;
  SIGNAL mux_1126_nl : STD_LOGIC;
  SIGNAL mux_1125_nl : STD_LOGIC;
  SIGNAL mux_1124_nl : STD_LOGIC;
  SIGNAL mux_1123_nl : STD_LOGIC;
  SIGNAL mux_1122_nl : STD_LOGIC;
  SIGNAL or_754_nl : STD_LOGIC;
  SIGNAL or_752_nl : STD_LOGIC;
  SIGNAL or_750_nl : STD_LOGIC;
  SIGNAL nand_20_nl : STD_LOGIC;
  SIGNAL mux_1121_nl : STD_LOGIC;
  SIGNAL mux_1120_nl : STD_LOGIC;
  SIGNAL mux_1119_nl : STD_LOGIC;
  SIGNAL or_748_nl : STD_LOGIC;
  SIGNAL or_747_nl : STD_LOGIC;
  SIGNAL or_745_nl : STD_LOGIC;
  SIGNAL or_744_nl : STD_LOGIC;
  SIGNAL mux_1118_nl : STD_LOGIC;
  SIGNAL mux_1117_nl : STD_LOGIC;
  SIGNAL or_742_nl : STD_LOGIC;
  SIGNAL or_740_nl : STD_LOGIC;
  SIGNAL mux_1116_nl : STD_LOGIC;
  SIGNAL or_739_nl : STD_LOGIC;
  SIGNAL mux_1115_nl : STD_LOGIC;
  SIGNAL or_737_nl : STD_LOGIC;
  SIGNAL mux_1114_nl : STD_LOGIC;
  SIGNAL mux_1113_nl : STD_LOGIC;
  SIGNAL or_730_nl : STD_LOGIC;
  SIGNAL or_729_nl : STD_LOGIC;
  SIGNAL or_727_nl : STD_LOGIC;
  SIGNAL or_726_nl : STD_LOGIC;
  SIGNAL mux_1110_nl : STD_LOGIC;
  SIGNAL or_725_nl : STD_LOGIC;
  SIGNAL mux_1109_nl : STD_LOGIC;
  SIGNAL or_724_nl : STD_LOGIC;
  SIGNAL mux_1108_nl : STD_LOGIC;
  SIGNAL or_723_nl : STD_LOGIC;
  SIGNAL or_722_nl : STD_LOGIC;
  SIGNAL mux_1175_nl : STD_LOGIC;
  SIGNAL mux_1174_nl : STD_LOGIC;
  SIGNAL mux_1173_nl : STD_LOGIC;
  SIGNAL nand_24_nl : STD_LOGIC;
  SIGNAL mux_1172_nl : STD_LOGIC;
  SIGNAL mux_1171_nl : STD_LOGIC;
  SIGNAL nor_753_nl : STD_LOGIC;
  SIGNAL nor_754_nl : STD_LOGIC;
  SIGNAL mux_1170_nl : STD_LOGIC;
  SIGNAL nor_755_nl : STD_LOGIC;
  SIGNAL nor_756_nl : STD_LOGIC;
  SIGNAL mux_1169_nl : STD_LOGIC;
  SIGNAL nand_23_nl : STD_LOGIC;
  SIGNAL mux_1168_nl : STD_LOGIC;
  SIGNAL nor_757_nl : STD_LOGIC;
  SIGNAL nor_758_nl : STD_LOGIC;
  SIGNAL mux_1167_nl : STD_LOGIC;
  SIGNAL mux_1166_nl : STD_LOGIC;
  SIGNAL or_820_nl : STD_LOGIC;
  SIGNAL or_818_nl : STD_LOGIC;
  SIGNAL or_817_nl : STD_LOGIC;
  SIGNAL mux_1165_nl : STD_LOGIC;
  SIGNAL or_816_nl : STD_LOGIC;
  SIGNAL mux_1164_nl : STD_LOGIC;
  SIGNAL mux_1163_nl : STD_LOGIC;
  SIGNAL or_815_nl : STD_LOGIC;
  SIGNAL or_814_nl : STD_LOGIC;
  SIGNAL mux_1162_nl : STD_LOGIC;
  SIGNAL or_812_nl : STD_LOGIC;
  SIGNAL or_810_nl : STD_LOGIC;
  SIGNAL mux_1161_nl : STD_LOGIC;
  SIGNAL or_808_nl : STD_LOGIC;
  SIGNAL mux_1160_nl : STD_LOGIC;
  SIGNAL or_807_nl : STD_LOGIC;
  SIGNAL or_806_nl : STD_LOGIC;
  SIGNAL or_805_nl : STD_LOGIC;
  SIGNAL mux_1159_nl : STD_LOGIC;
  SIGNAL mux_1158_nl : STD_LOGIC;
  SIGNAL mux_1157_nl : STD_LOGIC;
  SIGNAL mux_1156_nl : STD_LOGIC;
  SIGNAL mux_1155_nl : STD_LOGIC;
  SIGNAL or_801_nl : STD_LOGIC;
  SIGNAL mux_1154_nl : STD_LOGIC;
  SIGNAL or_800_nl : STD_LOGIC;
  SIGNAL nand_21_nl : STD_LOGIC;
  SIGNAL mux_1152_nl : STD_LOGIC;
  SIGNAL mux_1151_nl : STD_LOGIC;
  SIGNAL nor_759_nl : STD_LOGIC;
  SIGNAL nor_760_nl : STD_LOGIC;
  SIGNAL mux_1150_nl : STD_LOGIC;
  SIGNAL nor_761_nl : STD_LOGIC;
  SIGNAL nor_762_nl : STD_LOGIC;
  SIGNAL mux_1149_nl : STD_LOGIC;
  SIGNAL mux_1148_nl : STD_LOGIC;
  SIGNAL mux_1147_nl : STD_LOGIC;
  SIGNAL or_789_nl : STD_LOGIC;
  SIGNAL mux_1146_nl : STD_LOGIC;
  SIGNAL or_787_nl : STD_LOGIC;
  SIGNAL or_785_nl : STD_LOGIC;
  SIGNAL or_784_nl : STD_LOGIC;
  SIGNAL mux_1145_nl : STD_LOGIC;
  SIGNAL or_783_nl : STD_LOGIC;
  SIGNAL or_782_nl : STD_LOGIC;
  SIGNAL or_781_nl : STD_LOGIC;
  SIGNAL mux_1144_nl : STD_LOGIC;
  SIGNAL mux_1143_nl : STD_LOGIC;
  SIGNAL or_780_nl : STD_LOGIC;
  SIGNAL or_779_nl : STD_LOGIC;
  SIGNAL or_777_nl : STD_LOGIC;
  SIGNAL mux_1210_nl : STD_LOGIC;
  SIGNAL mux_1209_nl : STD_LOGIC;
  SIGNAL mux_1208_nl : STD_LOGIC;
  SIGNAL mux_1207_nl : STD_LOGIC;
  SIGNAL or_881_nl : STD_LOGIC;
  SIGNAL mux_1206_nl : STD_LOGIC;
  SIGNAL or_879_nl : STD_LOGIC;
  SIGNAL mux_1205_nl : STD_LOGIC;
  SIGNAL or_878_nl : STD_LOGIC;
  SIGNAL or_877_nl : STD_LOGIC;
  SIGNAL mux_1204_nl : STD_LOGIC;
  SIGNAL mux_1203_nl : STD_LOGIC;
  SIGNAL mux_1202_nl : STD_LOGIC;
  SIGNAL or_876_nl : STD_LOGIC;
  SIGNAL or_874_nl : STD_LOGIC;
  SIGNAL or_872_nl : STD_LOGIC;
  SIGNAL or_870_nl : STD_LOGIC;
  SIGNAL mux_1201_nl : STD_LOGIC;
  SIGNAL mux_1200_nl : STD_LOGIC;
  SIGNAL mux_1199_nl : STD_LOGIC;
  SIGNAL mux_1198_nl : STD_LOGIC;
  SIGNAL or_869_nl : STD_LOGIC;
  SIGNAL or_868_nl : STD_LOGIC;
  SIGNAL or_867_nl : STD_LOGIC;
  SIGNAL or_866_nl : STD_LOGIC;
  SIGNAL mux_1197_nl : STD_LOGIC;
  SIGNAL mux_1196_nl : STD_LOGIC;
  SIGNAL or_864_nl : STD_LOGIC;
  SIGNAL mux_1195_nl : STD_LOGIC;
  SIGNAL or_863_nl : STD_LOGIC;
  SIGNAL or_862_nl : STD_LOGIC;
  SIGNAL or_861_nl : STD_LOGIC;
  SIGNAL mux_1194_nl : STD_LOGIC;
  SIGNAL mux_1193_nl : STD_LOGIC;
  SIGNAL mux_1192_nl : STD_LOGIC;
  SIGNAL mux_1191_nl : STD_LOGIC;
  SIGNAL mux_1190_nl : STD_LOGIC;
  SIGNAL or_860_nl : STD_LOGIC;
  SIGNAL or_858_nl : STD_LOGIC;
  SIGNAL or_856_nl : STD_LOGIC;
  SIGNAL nand_26_nl : STD_LOGIC;
  SIGNAL mux_1189_nl : STD_LOGIC;
  SIGNAL mux_1188_nl : STD_LOGIC;
  SIGNAL or_854_nl : STD_LOGIC;
  SIGNAL mux_1187_nl : STD_LOGIC;
  SIGNAL or_852_nl : STD_LOGIC;
  SIGNAL nor_277_nl : STD_LOGIC;
  SIGNAL or_851_nl : STD_LOGIC;
  SIGNAL mux_1186_nl : STD_LOGIC;
  SIGNAL mux_1185_nl : STD_LOGIC;
  SIGNAL or_849_nl : STD_LOGIC;
  SIGNAL or_847_nl : STD_LOGIC;
  SIGNAL mux_1184_nl : STD_LOGIC;
  SIGNAL or_846_nl : STD_LOGIC;
  SIGNAL mux_1183_nl : STD_LOGIC;
  SIGNAL or_844_nl : STD_LOGIC;
  SIGNAL mux_1182_nl : STD_LOGIC;
  SIGNAL or_842_nl : STD_LOGIC;
  SIGNAL mux_1181_nl : STD_LOGIC;
  SIGNAL nor_275_nl : STD_LOGIC;
  SIGNAL nor_274_nl : STD_LOGIC;
  SIGNAL or_835_nl : STD_LOGIC;
  SIGNAL mux_1178_nl : STD_LOGIC;
  SIGNAL or_834_nl : STD_LOGIC;
  SIGNAL mux_1177_nl : STD_LOGIC;
  SIGNAL or_833_nl : STD_LOGIC;
  SIGNAL mux_1176_nl : STD_LOGIC;
  SIGNAL or_832_nl : STD_LOGIC;
  SIGNAL or_831_nl : STD_LOGIC;
  SIGNAL mux_1243_nl : STD_LOGIC;
  SIGNAL mux_1242_nl : STD_LOGIC;
  SIGNAL mux_1241_nl : STD_LOGIC;
  SIGNAL nand_30_nl : STD_LOGIC;
  SIGNAL mux_1240_nl : STD_LOGIC;
  SIGNAL mux_1239_nl : STD_LOGIC;
  SIGNAL nor_741_nl : STD_LOGIC;
  SIGNAL nor_742_nl : STD_LOGIC;
  SIGNAL mux_1238_nl : STD_LOGIC;
  SIGNAL nor_743_nl : STD_LOGIC;
  SIGNAL nor_744_nl : STD_LOGIC;
  SIGNAL mux_1237_nl : STD_LOGIC;
  SIGNAL nand_29_nl : STD_LOGIC;
  SIGNAL mux_1236_nl : STD_LOGIC;
  SIGNAL nor_745_nl : STD_LOGIC;
  SIGNAL nor_746_nl : STD_LOGIC;
  SIGNAL mux_1235_nl : STD_LOGIC;
  SIGNAL mux_1234_nl : STD_LOGIC;
  SIGNAL or_926_nl : STD_LOGIC;
  SIGNAL or_924_nl : STD_LOGIC;
  SIGNAL or_923_nl : STD_LOGIC;
  SIGNAL mux_1233_nl : STD_LOGIC;
  SIGNAL or_922_nl : STD_LOGIC;
  SIGNAL mux_1232_nl : STD_LOGIC;
  SIGNAL mux_1231_nl : STD_LOGIC;
  SIGNAL or_921_nl : STD_LOGIC;
  SIGNAL or_920_nl : STD_LOGIC;
  SIGNAL mux_1230_nl : STD_LOGIC;
  SIGNAL or_918_nl : STD_LOGIC;
  SIGNAL or_916_nl : STD_LOGIC;
  SIGNAL mux_1229_nl : STD_LOGIC;
  SIGNAL or_914_nl : STD_LOGIC;
  SIGNAL mux_1228_nl : STD_LOGIC;
  SIGNAL or_913_nl : STD_LOGIC;
  SIGNAL or_912_nl : STD_LOGIC;
  SIGNAL or_911_nl : STD_LOGIC;
  SIGNAL mux_1227_nl : STD_LOGIC;
  SIGNAL mux_1226_nl : STD_LOGIC;
  SIGNAL mux_1225_nl : STD_LOGIC;
  SIGNAL mux_1224_nl : STD_LOGIC;
  SIGNAL mux_1223_nl : STD_LOGIC;
  SIGNAL or_907_nl : STD_LOGIC;
  SIGNAL mux_1222_nl : STD_LOGIC;
  SIGNAL or_906_nl : STD_LOGIC;
  SIGNAL nand_27_nl : STD_LOGIC;
  SIGNAL mux_1220_nl : STD_LOGIC;
  SIGNAL mux_1219_nl : STD_LOGIC;
  SIGNAL nor_747_nl : STD_LOGIC;
  SIGNAL nor_748_nl : STD_LOGIC;
  SIGNAL mux_1218_nl : STD_LOGIC;
  SIGNAL nor_749_nl : STD_LOGIC;
  SIGNAL nor_750_nl : STD_LOGIC;
  SIGNAL mux_1217_nl : STD_LOGIC;
  SIGNAL mux_1216_nl : STD_LOGIC;
  SIGNAL mux_1215_nl : STD_LOGIC;
  SIGNAL or_895_nl : STD_LOGIC;
  SIGNAL mux_1214_nl : STD_LOGIC;
  SIGNAL or_893_nl : STD_LOGIC;
  SIGNAL or_891_nl : STD_LOGIC;
  SIGNAL or_890_nl : STD_LOGIC;
  SIGNAL mux_1213_nl : STD_LOGIC;
  SIGNAL or_889_nl : STD_LOGIC;
  SIGNAL or_888_nl : STD_LOGIC;
  SIGNAL or_887_nl : STD_LOGIC;
  SIGNAL mux_1212_nl : STD_LOGIC;
  SIGNAL mux_1211_nl : STD_LOGIC;
  SIGNAL or_886_nl : STD_LOGIC;
  SIGNAL or_885_nl : STD_LOGIC;
  SIGNAL or_883_nl : STD_LOGIC;
  SIGNAL mux_1278_nl : STD_LOGIC;
  SIGNAL mux_1277_nl : STD_LOGIC;
  SIGNAL mux_1276_nl : STD_LOGIC;
  SIGNAL mux_1275_nl : STD_LOGIC;
  SIGNAL or_990_nl : STD_LOGIC;
  SIGNAL mux_1274_nl : STD_LOGIC;
  SIGNAL or_988_nl : STD_LOGIC;
  SIGNAL mux_1273_nl : STD_LOGIC;
  SIGNAL or_987_nl : STD_LOGIC;
  SIGNAL or_986_nl : STD_LOGIC;
  SIGNAL mux_1272_nl : STD_LOGIC;
  SIGNAL mux_1271_nl : STD_LOGIC;
  SIGNAL mux_1270_nl : STD_LOGIC;
  SIGNAL or_985_nl : STD_LOGIC;
  SIGNAL or_983_nl : STD_LOGIC;
  SIGNAL or_981_nl : STD_LOGIC;
  SIGNAL or_979_nl : STD_LOGIC;
  SIGNAL mux_1269_nl : STD_LOGIC;
  SIGNAL mux_1268_nl : STD_LOGIC;
  SIGNAL mux_1267_nl : STD_LOGIC;
  SIGNAL mux_1266_nl : STD_LOGIC;
  SIGNAL or_978_nl : STD_LOGIC;
  SIGNAL or_977_nl : STD_LOGIC;
  SIGNAL or_976_nl : STD_LOGIC;
  SIGNAL or_975_nl : STD_LOGIC;
  SIGNAL mux_1265_nl : STD_LOGIC;
  SIGNAL mux_1264_nl : STD_LOGIC;
  SIGNAL or_973_nl : STD_LOGIC;
  SIGNAL mux_1263_nl : STD_LOGIC;
  SIGNAL or_972_nl : STD_LOGIC;
  SIGNAL or_971_nl : STD_LOGIC;
  SIGNAL or_970_nl : STD_LOGIC;
  SIGNAL mux_1262_nl : STD_LOGIC;
  SIGNAL mux_1261_nl : STD_LOGIC;
  SIGNAL mux_1260_nl : STD_LOGIC;
  SIGNAL mux_1259_nl : STD_LOGIC;
  SIGNAL mux_1258_nl : STD_LOGIC;
  SIGNAL or_969_nl : STD_LOGIC;
  SIGNAL or_967_nl : STD_LOGIC;
  SIGNAL or_965_nl : STD_LOGIC;
  SIGNAL nand_32_nl : STD_LOGIC;
  SIGNAL mux_1257_nl : STD_LOGIC;
  SIGNAL mux_1256_nl : STD_LOGIC;
  SIGNAL mux_1255_nl : STD_LOGIC;
  SIGNAL or_963_nl : STD_LOGIC;
  SIGNAL or_962_nl : STD_LOGIC;
  SIGNAL or_960_nl : STD_LOGIC;
  SIGNAL or_959_nl : STD_LOGIC;
  SIGNAL mux_1254_nl : STD_LOGIC;
  SIGNAL mux_1253_nl : STD_LOGIC;
  SIGNAL or_957_nl : STD_LOGIC;
  SIGNAL or_955_nl : STD_LOGIC;
  SIGNAL mux_1252_nl : STD_LOGIC;
  SIGNAL or_954_nl : STD_LOGIC;
  SIGNAL mux_1251_nl : STD_LOGIC;
  SIGNAL or_952_nl : STD_LOGIC;
  SIGNAL mux_1250_nl : STD_LOGIC;
  SIGNAL mux_1249_nl : STD_LOGIC;
  SIGNAL or_945_nl : STD_LOGIC;
  SIGNAL or_944_nl : STD_LOGIC;
  SIGNAL or_942_nl : STD_LOGIC;
  SIGNAL or_941_nl : STD_LOGIC;
  SIGNAL mux_1246_nl : STD_LOGIC;
  SIGNAL or_940_nl : STD_LOGIC;
  SIGNAL mux_1245_nl : STD_LOGIC;
  SIGNAL or_939_nl : STD_LOGIC;
  SIGNAL mux_1244_nl : STD_LOGIC;
  SIGNAL or_938_nl : STD_LOGIC;
  SIGNAL or_937_nl : STD_LOGIC;
  SIGNAL mux_1311_nl : STD_LOGIC;
  SIGNAL mux_1310_nl : STD_LOGIC;
  SIGNAL mux_1309_nl : STD_LOGIC;
  SIGNAL nand_36_nl : STD_LOGIC;
  SIGNAL mux_1308_nl : STD_LOGIC;
  SIGNAL mux_1307_nl : STD_LOGIC;
  SIGNAL nor_729_nl : STD_LOGIC;
  SIGNAL nor_730_nl : STD_LOGIC;
  SIGNAL mux_1306_nl : STD_LOGIC;
  SIGNAL nor_731_nl : STD_LOGIC;
  SIGNAL nor_732_nl : STD_LOGIC;
  SIGNAL mux_1305_nl : STD_LOGIC;
  SIGNAL nand_35_nl : STD_LOGIC;
  SIGNAL mux_1304_nl : STD_LOGIC;
  SIGNAL nor_733_nl : STD_LOGIC;
  SIGNAL nor_734_nl : STD_LOGIC;
  SIGNAL mux_1303_nl : STD_LOGIC;
  SIGNAL mux_1302_nl : STD_LOGIC;
  SIGNAL or_1035_nl : STD_LOGIC;
  SIGNAL or_1033_nl : STD_LOGIC;
  SIGNAL or_1032_nl : STD_LOGIC;
  SIGNAL mux_1301_nl : STD_LOGIC;
  SIGNAL or_1031_nl : STD_LOGIC;
  SIGNAL mux_1300_nl : STD_LOGIC;
  SIGNAL mux_1299_nl : STD_LOGIC;
  SIGNAL or_1030_nl : STD_LOGIC;
  SIGNAL or_1029_nl : STD_LOGIC;
  SIGNAL mux_1298_nl : STD_LOGIC;
  SIGNAL or_1027_nl : STD_LOGIC;
  SIGNAL or_1025_nl : STD_LOGIC;
  SIGNAL mux_1297_nl : STD_LOGIC;
  SIGNAL or_1023_nl : STD_LOGIC;
  SIGNAL mux_1296_nl : STD_LOGIC;
  SIGNAL or_1022_nl : STD_LOGIC;
  SIGNAL or_1021_nl : STD_LOGIC;
  SIGNAL or_1020_nl : STD_LOGIC;
  SIGNAL mux_1295_nl : STD_LOGIC;
  SIGNAL mux_1294_nl : STD_LOGIC;
  SIGNAL mux_1293_nl : STD_LOGIC;
  SIGNAL mux_1292_nl : STD_LOGIC;
  SIGNAL mux_1291_nl : STD_LOGIC;
  SIGNAL or_1016_nl : STD_LOGIC;
  SIGNAL mux_1290_nl : STD_LOGIC;
  SIGNAL or_1015_nl : STD_LOGIC;
  SIGNAL nand_33_nl : STD_LOGIC;
  SIGNAL mux_1288_nl : STD_LOGIC;
  SIGNAL mux_1287_nl : STD_LOGIC;
  SIGNAL nor_735_nl : STD_LOGIC;
  SIGNAL nor_736_nl : STD_LOGIC;
  SIGNAL mux_1286_nl : STD_LOGIC;
  SIGNAL nor_737_nl : STD_LOGIC;
  SIGNAL nor_738_nl : STD_LOGIC;
  SIGNAL mux_1285_nl : STD_LOGIC;
  SIGNAL mux_1284_nl : STD_LOGIC;
  SIGNAL mux_1283_nl : STD_LOGIC;
  SIGNAL or_1004_nl : STD_LOGIC;
  SIGNAL mux_1282_nl : STD_LOGIC;
  SIGNAL or_1002_nl : STD_LOGIC;
  SIGNAL or_1000_nl : STD_LOGIC;
  SIGNAL or_999_nl : STD_LOGIC;
  SIGNAL mux_1281_nl : STD_LOGIC;
  SIGNAL or_998_nl : STD_LOGIC;
  SIGNAL or_997_nl : STD_LOGIC;
  SIGNAL or_996_nl : STD_LOGIC;
  SIGNAL mux_1280_nl : STD_LOGIC;
  SIGNAL mux_1279_nl : STD_LOGIC;
  SIGNAL or_995_nl : STD_LOGIC;
  SIGNAL or_994_nl : STD_LOGIC;
  SIGNAL or_992_nl : STD_LOGIC;
  SIGNAL mux_1346_nl : STD_LOGIC;
  SIGNAL mux_1345_nl : STD_LOGIC;
  SIGNAL mux_1344_nl : STD_LOGIC;
  SIGNAL mux_1343_nl : STD_LOGIC;
  SIGNAL or_1096_nl : STD_LOGIC;
  SIGNAL mux_1342_nl : STD_LOGIC;
  SIGNAL or_1094_nl : STD_LOGIC;
  SIGNAL mux_1341_nl : STD_LOGIC;
  SIGNAL or_1093_nl : STD_LOGIC;
  SIGNAL or_1092_nl : STD_LOGIC;
  SIGNAL mux_1340_nl : STD_LOGIC;
  SIGNAL mux_1339_nl : STD_LOGIC;
  SIGNAL mux_1338_nl : STD_LOGIC;
  SIGNAL or_1091_nl : STD_LOGIC;
  SIGNAL or_1089_nl : STD_LOGIC;
  SIGNAL or_1087_nl : STD_LOGIC;
  SIGNAL or_1085_nl : STD_LOGIC;
  SIGNAL mux_1337_nl : STD_LOGIC;
  SIGNAL mux_1336_nl : STD_LOGIC;
  SIGNAL mux_1335_nl : STD_LOGIC;
  SIGNAL mux_1334_nl : STD_LOGIC;
  SIGNAL or_1084_nl : STD_LOGIC;
  SIGNAL or_1083_nl : STD_LOGIC;
  SIGNAL or_1082_nl : STD_LOGIC;
  SIGNAL or_1081_nl : STD_LOGIC;
  SIGNAL mux_1333_nl : STD_LOGIC;
  SIGNAL mux_1332_nl : STD_LOGIC;
  SIGNAL nand_357_nl : STD_LOGIC;
  SIGNAL mux_1331_nl : STD_LOGIC;
  SIGNAL or_1078_nl : STD_LOGIC;
  SIGNAL or_1077_nl : STD_LOGIC;
  SIGNAL or_1076_nl : STD_LOGIC;
  SIGNAL mux_1330_nl : STD_LOGIC;
  SIGNAL mux_1329_nl : STD_LOGIC;
  SIGNAL mux_1328_nl : STD_LOGIC;
  SIGNAL mux_1327_nl : STD_LOGIC;
  SIGNAL mux_1326_nl : STD_LOGIC;
  SIGNAL or_1075_nl : STD_LOGIC;
  SIGNAL or_1073_nl : STD_LOGIC;
  SIGNAL or_1071_nl : STD_LOGIC;
  SIGNAL nand_38_nl : STD_LOGIC;
  SIGNAL mux_1325_nl : STD_LOGIC;
  SIGNAL mux_1324_nl : STD_LOGIC;
  SIGNAL or_1069_nl : STD_LOGIC;
  SIGNAL mux_1323_nl : STD_LOGIC;
  SIGNAL or_1067_nl : STD_LOGIC;
  SIGNAL nor_288_nl : STD_LOGIC;
  SIGNAL or_1066_nl : STD_LOGIC;
  SIGNAL mux_1322_nl : STD_LOGIC;
  SIGNAL mux_1321_nl : STD_LOGIC;
  SIGNAL or_1064_nl : STD_LOGIC;
  SIGNAL or_1062_nl : STD_LOGIC;
  SIGNAL mux_1320_nl : STD_LOGIC;
  SIGNAL or_1061_nl : STD_LOGIC;
  SIGNAL mux_1319_nl : STD_LOGIC;
  SIGNAL or_1059_nl : STD_LOGIC;
  SIGNAL mux_1318_nl : STD_LOGIC;
  SIGNAL or_1057_nl : STD_LOGIC;
  SIGNAL mux_1317_nl : STD_LOGIC;
  SIGNAL nor_286_nl : STD_LOGIC;
  SIGNAL nor_285_nl : STD_LOGIC;
  SIGNAL or_1050_nl : STD_LOGIC;
  SIGNAL mux_1314_nl : STD_LOGIC;
  SIGNAL or_1049_nl : STD_LOGIC;
  SIGNAL mux_1313_nl : STD_LOGIC;
  SIGNAL or_1048_nl : STD_LOGIC;
  SIGNAL mux_1312_nl : STD_LOGIC;
  SIGNAL or_1047_nl : STD_LOGIC;
  SIGNAL or_1046_nl : STD_LOGIC;
  SIGNAL mux_1379_nl : STD_LOGIC;
  SIGNAL mux_1378_nl : STD_LOGIC;
  SIGNAL mux_1377_nl : STD_LOGIC;
  SIGNAL nand_42_nl : STD_LOGIC;
  SIGNAL mux_1376_nl : STD_LOGIC;
  SIGNAL mux_1375_nl : STD_LOGIC;
  SIGNAL nor_717_nl : STD_LOGIC;
  SIGNAL nor_718_nl : STD_LOGIC;
  SIGNAL mux_1374_nl : STD_LOGIC;
  SIGNAL nor_719_nl : STD_LOGIC;
  SIGNAL nor_720_nl : STD_LOGIC;
  SIGNAL mux_1373_nl : STD_LOGIC;
  SIGNAL nand_41_nl : STD_LOGIC;
  SIGNAL mux_1372_nl : STD_LOGIC;
  SIGNAL nor_721_nl : STD_LOGIC;
  SIGNAL nor_722_nl : STD_LOGIC;
  SIGNAL mux_1371_nl : STD_LOGIC;
  SIGNAL mux_1370_nl : STD_LOGIC;
  SIGNAL or_1141_nl : STD_LOGIC;
  SIGNAL or_1139_nl : STD_LOGIC;
  SIGNAL or_1138_nl : STD_LOGIC;
  SIGNAL mux_1369_nl : STD_LOGIC;
  SIGNAL or_1137_nl : STD_LOGIC;
  SIGNAL mux_1368_nl : STD_LOGIC;
  SIGNAL mux_1367_nl : STD_LOGIC;
  SIGNAL or_1136_nl : STD_LOGIC;
  SIGNAL or_1135_nl : STD_LOGIC;
  SIGNAL mux_1366_nl : STD_LOGIC;
  SIGNAL or_1133_nl : STD_LOGIC;
  SIGNAL or_1131_nl : STD_LOGIC;
  SIGNAL mux_1365_nl : STD_LOGIC;
  SIGNAL or_1129_nl : STD_LOGIC;
  SIGNAL mux_1364_nl : STD_LOGIC;
  SIGNAL or_1128_nl : STD_LOGIC;
  SIGNAL or_1127_nl : STD_LOGIC;
  SIGNAL or_1126_nl : STD_LOGIC;
  SIGNAL mux_1363_nl : STD_LOGIC;
  SIGNAL mux_1362_nl : STD_LOGIC;
  SIGNAL mux_1361_nl : STD_LOGIC;
  SIGNAL mux_1360_nl : STD_LOGIC;
  SIGNAL mux_1359_nl : STD_LOGIC;
  SIGNAL or_1122_nl : STD_LOGIC;
  SIGNAL mux_1358_nl : STD_LOGIC;
  SIGNAL or_1121_nl : STD_LOGIC;
  SIGNAL nand_39_nl : STD_LOGIC;
  SIGNAL mux_1356_nl : STD_LOGIC;
  SIGNAL mux_1355_nl : STD_LOGIC;
  SIGNAL nor_723_nl : STD_LOGIC;
  SIGNAL nor_724_nl : STD_LOGIC;
  SIGNAL mux_1354_nl : STD_LOGIC;
  SIGNAL nor_725_nl : STD_LOGIC;
  SIGNAL nor_726_nl : STD_LOGIC;
  SIGNAL mux_1353_nl : STD_LOGIC;
  SIGNAL mux_1352_nl : STD_LOGIC;
  SIGNAL mux_1351_nl : STD_LOGIC;
  SIGNAL or_1110_nl : STD_LOGIC;
  SIGNAL mux_1350_nl : STD_LOGIC;
  SIGNAL or_1108_nl : STD_LOGIC;
  SIGNAL or_1106_nl : STD_LOGIC;
  SIGNAL or_1105_nl : STD_LOGIC;
  SIGNAL mux_1349_nl : STD_LOGIC;
  SIGNAL or_1104_nl : STD_LOGIC;
  SIGNAL or_1103_nl : STD_LOGIC;
  SIGNAL or_1102_nl : STD_LOGIC;
  SIGNAL mux_1348_nl : STD_LOGIC;
  SIGNAL mux_1347_nl : STD_LOGIC;
  SIGNAL or_1101_nl : STD_LOGIC;
  SIGNAL or_1100_nl : STD_LOGIC;
  SIGNAL or_1098_nl : STD_LOGIC;
  SIGNAL mux_1414_nl : STD_LOGIC;
  SIGNAL mux_1413_nl : STD_LOGIC;
  SIGNAL mux_1412_nl : STD_LOGIC;
  SIGNAL mux_1411_nl : STD_LOGIC;
  SIGNAL or_1205_nl : STD_LOGIC;
  SIGNAL mux_1410_nl : STD_LOGIC;
  SIGNAL or_1203_nl : STD_LOGIC;
  SIGNAL mux_1409_nl : STD_LOGIC;
  SIGNAL or_1202_nl : STD_LOGIC;
  SIGNAL or_1201_nl : STD_LOGIC;
  SIGNAL mux_1408_nl : STD_LOGIC;
  SIGNAL mux_1407_nl : STD_LOGIC;
  SIGNAL mux_1406_nl : STD_LOGIC;
  SIGNAL or_1200_nl : STD_LOGIC;
  SIGNAL or_1198_nl : STD_LOGIC;
  SIGNAL or_1196_nl : STD_LOGIC;
  SIGNAL or_1194_nl : STD_LOGIC;
  SIGNAL mux_1405_nl : STD_LOGIC;
  SIGNAL mux_1404_nl : STD_LOGIC;
  SIGNAL mux_1403_nl : STD_LOGIC;
  SIGNAL mux_1402_nl : STD_LOGIC;
  SIGNAL or_1193_nl : STD_LOGIC;
  SIGNAL or_1192_nl : STD_LOGIC;
  SIGNAL or_1191_nl : STD_LOGIC;
  SIGNAL or_1190_nl : STD_LOGIC;
  SIGNAL mux_1401_nl : STD_LOGIC;
  SIGNAL mux_1400_nl : STD_LOGIC;
  SIGNAL or_1188_nl : STD_LOGIC;
  SIGNAL mux_1399_nl : STD_LOGIC;
  SIGNAL or_1187_nl : STD_LOGIC;
  SIGNAL or_1186_nl : STD_LOGIC;
  SIGNAL or_1185_nl : STD_LOGIC;
  SIGNAL mux_1398_nl : STD_LOGIC;
  SIGNAL mux_1397_nl : STD_LOGIC;
  SIGNAL mux_1396_nl : STD_LOGIC;
  SIGNAL mux_1395_nl : STD_LOGIC;
  SIGNAL mux_1394_nl : STD_LOGIC;
  SIGNAL or_1184_nl : STD_LOGIC;
  SIGNAL or_1182_nl : STD_LOGIC;
  SIGNAL or_1180_nl : STD_LOGIC;
  SIGNAL nand_44_nl : STD_LOGIC;
  SIGNAL mux_1393_nl : STD_LOGIC;
  SIGNAL mux_1392_nl : STD_LOGIC;
  SIGNAL mux_1391_nl : STD_LOGIC;
  SIGNAL or_1178_nl : STD_LOGIC;
  SIGNAL or_1177_nl : STD_LOGIC;
  SIGNAL or_1175_nl : STD_LOGIC;
  SIGNAL or_1174_nl : STD_LOGIC;
  SIGNAL mux_1390_nl : STD_LOGIC;
  SIGNAL mux_1389_nl : STD_LOGIC;
  SIGNAL or_1172_nl : STD_LOGIC;
  SIGNAL or_1170_nl : STD_LOGIC;
  SIGNAL mux_1388_nl : STD_LOGIC;
  SIGNAL or_1169_nl : STD_LOGIC;
  SIGNAL mux_1387_nl : STD_LOGIC;
  SIGNAL or_1167_nl : STD_LOGIC;
  SIGNAL mux_1386_nl : STD_LOGIC;
  SIGNAL mux_1385_nl : STD_LOGIC;
  SIGNAL or_1160_nl : STD_LOGIC;
  SIGNAL or_1159_nl : STD_LOGIC;
  SIGNAL or_1157_nl : STD_LOGIC;
  SIGNAL or_1156_nl : STD_LOGIC;
  SIGNAL mux_1382_nl : STD_LOGIC;
  SIGNAL or_1155_nl : STD_LOGIC;
  SIGNAL mux_1381_nl : STD_LOGIC;
  SIGNAL or_1154_nl : STD_LOGIC;
  SIGNAL mux_1380_nl : STD_LOGIC;
  SIGNAL or_1153_nl : STD_LOGIC;
  SIGNAL or_1152_nl : STD_LOGIC;
  SIGNAL mux_1447_nl : STD_LOGIC;
  SIGNAL mux_1446_nl : STD_LOGIC;
  SIGNAL mux_1445_nl : STD_LOGIC;
  SIGNAL nand_48_nl : STD_LOGIC;
  SIGNAL mux_1444_nl : STD_LOGIC;
  SIGNAL mux_1443_nl : STD_LOGIC;
  SIGNAL nor_705_nl : STD_LOGIC;
  SIGNAL nor_706_nl : STD_LOGIC;
  SIGNAL mux_1442_nl : STD_LOGIC;
  SIGNAL nor_707_nl : STD_LOGIC;
  SIGNAL nor_708_nl : STD_LOGIC;
  SIGNAL mux_1441_nl : STD_LOGIC;
  SIGNAL nand_47_nl : STD_LOGIC;
  SIGNAL mux_1440_nl : STD_LOGIC;
  SIGNAL nor_709_nl : STD_LOGIC;
  SIGNAL nor_710_nl : STD_LOGIC;
  SIGNAL mux_1439_nl : STD_LOGIC;
  SIGNAL mux_1438_nl : STD_LOGIC;
  SIGNAL or_1250_nl : STD_LOGIC;
  SIGNAL or_1248_nl : STD_LOGIC;
  SIGNAL or_1247_nl : STD_LOGIC;
  SIGNAL mux_1437_nl : STD_LOGIC;
  SIGNAL or_1246_nl : STD_LOGIC;
  SIGNAL mux_1436_nl : STD_LOGIC;
  SIGNAL mux_1435_nl : STD_LOGIC;
  SIGNAL or_1245_nl : STD_LOGIC;
  SIGNAL or_1244_nl : STD_LOGIC;
  SIGNAL mux_1434_nl : STD_LOGIC;
  SIGNAL or_1242_nl : STD_LOGIC;
  SIGNAL or_1240_nl : STD_LOGIC;
  SIGNAL mux_1433_nl : STD_LOGIC;
  SIGNAL or_1238_nl : STD_LOGIC;
  SIGNAL mux_1432_nl : STD_LOGIC;
  SIGNAL or_1237_nl : STD_LOGIC;
  SIGNAL or_1236_nl : STD_LOGIC;
  SIGNAL or_1235_nl : STD_LOGIC;
  SIGNAL mux_1431_nl : STD_LOGIC;
  SIGNAL mux_1430_nl : STD_LOGIC;
  SIGNAL mux_1429_nl : STD_LOGIC;
  SIGNAL mux_1428_nl : STD_LOGIC;
  SIGNAL mux_1427_nl : STD_LOGIC;
  SIGNAL or_1231_nl : STD_LOGIC;
  SIGNAL mux_1426_nl : STD_LOGIC;
  SIGNAL or_1230_nl : STD_LOGIC;
  SIGNAL nand_45_nl : STD_LOGIC;
  SIGNAL mux_1424_nl : STD_LOGIC;
  SIGNAL mux_1423_nl : STD_LOGIC;
  SIGNAL nor_711_nl : STD_LOGIC;
  SIGNAL nor_712_nl : STD_LOGIC;
  SIGNAL mux_1422_nl : STD_LOGIC;
  SIGNAL nor_713_nl : STD_LOGIC;
  SIGNAL nor_714_nl : STD_LOGIC;
  SIGNAL mux_1421_nl : STD_LOGIC;
  SIGNAL mux_1420_nl : STD_LOGIC;
  SIGNAL mux_1419_nl : STD_LOGIC;
  SIGNAL or_1219_nl : STD_LOGIC;
  SIGNAL mux_1418_nl : STD_LOGIC;
  SIGNAL or_1217_nl : STD_LOGIC;
  SIGNAL or_1215_nl : STD_LOGIC;
  SIGNAL or_1214_nl : STD_LOGIC;
  SIGNAL mux_1417_nl : STD_LOGIC;
  SIGNAL or_1213_nl : STD_LOGIC;
  SIGNAL or_1212_nl : STD_LOGIC;
  SIGNAL or_1211_nl : STD_LOGIC;
  SIGNAL mux_1416_nl : STD_LOGIC;
  SIGNAL mux_1415_nl : STD_LOGIC;
  SIGNAL or_1210_nl : STD_LOGIC;
  SIGNAL or_1209_nl : STD_LOGIC;
  SIGNAL or_1207_nl : STD_LOGIC;
  SIGNAL mux_1482_nl : STD_LOGIC;
  SIGNAL mux_1481_nl : STD_LOGIC;
  SIGNAL mux_1480_nl : STD_LOGIC;
  SIGNAL mux_1479_nl : STD_LOGIC;
  SIGNAL or_1311_nl : STD_LOGIC;
  SIGNAL mux_1478_nl : STD_LOGIC;
  SIGNAL or_1309_nl : STD_LOGIC;
  SIGNAL mux_1477_nl : STD_LOGIC;
  SIGNAL or_1308_nl : STD_LOGIC;
  SIGNAL or_1307_nl : STD_LOGIC;
  SIGNAL mux_1476_nl : STD_LOGIC;
  SIGNAL mux_1475_nl : STD_LOGIC;
  SIGNAL mux_1474_nl : STD_LOGIC;
  SIGNAL or_1306_nl : STD_LOGIC;
  SIGNAL or_1304_nl : STD_LOGIC;
  SIGNAL or_1302_nl : STD_LOGIC;
  SIGNAL or_1300_nl : STD_LOGIC;
  SIGNAL mux_1473_nl : STD_LOGIC;
  SIGNAL mux_1472_nl : STD_LOGIC;
  SIGNAL mux_1471_nl : STD_LOGIC;
  SIGNAL mux_1470_nl : STD_LOGIC;
  SIGNAL or_1299_nl : STD_LOGIC;
  SIGNAL or_1298_nl : STD_LOGIC;
  SIGNAL or_1297_nl : STD_LOGIC;
  SIGNAL or_1296_nl : STD_LOGIC;
  SIGNAL mux_1469_nl : STD_LOGIC;
  SIGNAL mux_1468_nl : STD_LOGIC;
  SIGNAL nand_346_nl : STD_LOGIC;
  SIGNAL mux_1467_nl : STD_LOGIC;
  SIGNAL or_1293_nl : STD_LOGIC;
  SIGNAL or_1292_nl : STD_LOGIC;
  SIGNAL or_1291_nl : STD_LOGIC;
  SIGNAL mux_1466_nl : STD_LOGIC;
  SIGNAL mux_1465_nl : STD_LOGIC;
  SIGNAL mux_1464_nl : STD_LOGIC;
  SIGNAL mux_1463_nl : STD_LOGIC;
  SIGNAL mux_1462_nl : STD_LOGIC;
  SIGNAL or_1290_nl : STD_LOGIC;
  SIGNAL or_1288_nl : STD_LOGIC;
  SIGNAL or_1286_nl : STD_LOGIC;
  SIGNAL nand_50_nl : STD_LOGIC;
  SIGNAL mux_1461_nl : STD_LOGIC;
  SIGNAL mux_1460_nl : STD_LOGIC;
  SIGNAL or_1284_nl : STD_LOGIC;
  SIGNAL mux_1459_nl : STD_LOGIC;
  SIGNAL or_1282_nl : STD_LOGIC;
  SIGNAL nor_299_nl : STD_LOGIC;
  SIGNAL or_1281_nl : STD_LOGIC;
  SIGNAL mux_1458_nl : STD_LOGIC;
  SIGNAL mux_1457_nl : STD_LOGIC;
  SIGNAL or_1279_nl : STD_LOGIC;
  SIGNAL or_1277_nl : STD_LOGIC;
  SIGNAL mux_1456_nl : STD_LOGIC;
  SIGNAL or_1276_nl : STD_LOGIC;
  SIGNAL mux_1455_nl : STD_LOGIC;
  SIGNAL or_1274_nl : STD_LOGIC;
  SIGNAL mux_1454_nl : STD_LOGIC;
  SIGNAL or_1272_nl : STD_LOGIC;
  SIGNAL mux_1453_nl : STD_LOGIC;
  SIGNAL nor_297_nl : STD_LOGIC;
  SIGNAL nor_296_nl : STD_LOGIC;
  SIGNAL or_1265_nl : STD_LOGIC;
  SIGNAL mux_1450_nl : STD_LOGIC;
  SIGNAL or_1264_nl : STD_LOGIC;
  SIGNAL mux_1449_nl : STD_LOGIC;
  SIGNAL or_1263_nl : STD_LOGIC;
  SIGNAL mux_1448_nl : STD_LOGIC;
  SIGNAL or_1262_nl : STD_LOGIC;
  SIGNAL or_1261_nl : STD_LOGIC;
  SIGNAL mux_1515_nl : STD_LOGIC;
  SIGNAL mux_1514_nl : STD_LOGIC;
  SIGNAL mux_1513_nl : STD_LOGIC;
  SIGNAL nand_54_nl : STD_LOGIC;
  SIGNAL mux_1512_nl : STD_LOGIC;
  SIGNAL mux_1511_nl : STD_LOGIC;
  SIGNAL nor_693_nl : STD_LOGIC;
  SIGNAL nor_694_nl : STD_LOGIC;
  SIGNAL mux_1510_nl : STD_LOGIC;
  SIGNAL nor_695_nl : STD_LOGIC;
  SIGNAL nor_696_nl : STD_LOGIC;
  SIGNAL mux_1509_nl : STD_LOGIC;
  SIGNAL nand_53_nl : STD_LOGIC;
  SIGNAL mux_1508_nl : STD_LOGIC;
  SIGNAL nor_697_nl : STD_LOGIC;
  SIGNAL nor_698_nl : STD_LOGIC;
  SIGNAL mux_1507_nl : STD_LOGIC;
  SIGNAL mux_1506_nl : STD_LOGIC;
  SIGNAL or_1356_nl : STD_LOGIC;
  SIGNAL or_1354_nl : STD_LOGIC;
  SIGNAL or_1353_nl : STD_LOGIC;
  SIGNAL mux_1505_nl : STD_LOGIC;
  SIGNAL or_1352_nl : STD_LOGIC;
  SIGNAL mux_1504_nl : STD_LOGIC;
  SIGNAL mux_1503_nl : STD_LOGIC;
  SIGNAL or_1351_nl : STD_LOGIC;
  SIGNAL or_1350_nl : STD_LOGIC;
  SIGNAL mux_1502_nl : STD_LOGIC;
  SIGNAL or_1348_nl : STD_LOGIC;
  SIGNAL or_1346_nl : STD_LOGIC;
  SIGNAL mux_1501_nl : STD_LOGIC;
  SIGNAL or_1344_nl : STD_LOGIC;
  SIGNAL mux_1500_nl : STD_LOGIC;
  SIGNAL or_1343_nl : STD_LOGIC;
  SIGNAL or_1342_nl : STD_LOGIC;
  SIGNAL or_1341_nl : STD_LOGIC;
  SIGNAL mux_1499_nl : STD_LOGIC;
  SIGNAL mux_1498_nl : STD_LOGIC;
  SIGNAL mux_1497_nl : STD_LOGIC;
  SIGNAL mux_1496_nl : STD_LOGIC;
  SIGNAL mux_1495_nl : STD_LOGIC;
  SIGNAL or_1337_nl : STD_LOGIC;
  SIGNAL mux_1494_nl : STD_LOGIC;
  SIGNAL or_1336_nl : STD_LOGIC;
  SIGNAL nand_51_nl : STD_LOGIC;
  SIGNAL mux_1492_nl : STD_LOGIC;
  SIGNAL mux_1491_nl : STD_LOGIC;
  SIGNAL nor_699_nl : STD_LOGIC;
  SIGNAL nor_700_nl : STD_LOGIC;
  SIGNAL mux_1490_nl : STD_LOGIC;
  SIGNAL nor_701_nl : STD_LOGIC;
  SIGNAL nor_702_nl : STD_LOGIC;
  SIGNAL mux_1489_nl : STD_LOGIC;
  SIGNAL mux_1488_nl : STD_LOGIC;
  SIGNAL mux_1487_nl : STD_LOGIC;
  SIGNAL or_1325_nl : STD_LOGIC;
  SIGNAL mux_1486_nl : STD_LOGIC;
  SIGNAL or_1323_nl : STD_LOGIC;
  SIGNAL or_1321_nl : STD_LOGIC;
  SIGNAL or_1320_nl : STD_LOGIC;
  SIGNAL mux_1485_nl : STD_LOGIC;
  SIGNAL or_1319_nl : STD_LOGIC;
  SIGNAL or_1318_nl : STD_LOGIC;
  SIGNAL or_1317_nl : STD_LOGIC;
  SIGNAL mux_1484_nl : STD_LOGIC;
  SIGNAL mux_1483_nl : STD_LOGIC;
  SIGNAL or_1316_nl : STD_LOGIC;
  SIGNAL or_1315_nl : STD_LOGIC;
  SIGNAL or_1313_nl : STD_LOGIC;
  SIGNAL mux_1550_nl : STD_LOGIC;
  SIGNAL mux_1549_nl : STD_LOGIC;
  SIGNAL mux_1548_nl : STD_LOGIC;
  SIGNAL mux_1547_nl : STD_LOGIC;
  SIGNAL or_1420_nl : STD_LOGIC;
  SIGNAL mux_1546_nl : STD_LOGIC;
  SIGNAL or_1418_nl : STD_LOGIC;
  SIGNAL mux_1545_nl : STD_LOGIC;
  SIGNAL or_1417_nl : STD_LOGIC;
  SIGNAL or_1416_nl : STD_LOGIC;
  SIGNAL mux_1544_nl : STD_LOGIC;
  SIGNAL mux_1543_nl : STD_LOGIC;
  SIGNAL mux_1542_nl : STD_LOGIC;
  SIGNAL or_1415_nl : STD_LOGIC;
  SIGNAL or_1413_nl : STD_LOGIC;
  SIGNAL or_1411_nl : STD_LOGIC;
  SIGNAL or_1409_nl : STD_LOGIC;
  SIGNAL mux_1541_nl : STD_LOGIC;
  SIGNAL mux_1540_nl : STD_LOGIC;
  SIGNAL mux_1539_nl : STD_LOGIC;
  SIGNAL mux_1538_nl : STD_LOGIC;
  SIGNAL or_1408_nl : STD_LOGIC;
  SIGNAL or_1407_nl : STD_LOGIC;
  SIGNAL or_1406_nl : STD_LOGIC;
  SIGNAL or_1405_nl : STD_LOGIC;
  SIGNAL mux_1537_nl : STD_LOGIC;
  SIGNAL mux_1536_nl : STD_LOGIC;
  SIGNAL nand_340_nl : STD_LOGIC;
  SIGNAL mux_1535_nl : STD_LOGIC;
  SIGNAL or_1402_nl : STD_LOGIC;
  SIGNAL or_1401_nl : STD_LOGIC;
  SIGNAL or_1400_nl : STD_LOGIC;
  SIGNAL mux_1534_nl : STD_LOGIC;
  SIGNAL mux_1533_nl : STD_LOGIC;
  SIGNAL mux_1532_nl : STD_LOGIC;
  SIGNAL mux_1531_nl : STD_LOGIC;
  SIGNAL mux_1530_nl : STD_LOGIC;
  SIGNAL or_1399_nl : STD_LOGIC;
  SIGNAL or_1397_nl : STD_LOGIC;
  SIGNAL or_1395_nl : STD_LOGIC;
  SIGNAL nand_56_nl : STD_LOGIC;
  SIGNAL mux_1529_nl : STD_LOGIC;
  SIGNAL mux_1528_nl : STD_LOGIC;
  SIGNAL mux_1527_nl : STD_LOGIC;
  SIGNAL or_1393_nl : STD_LOGIC;
  SIGNAL or_1392_nl : STD_LOGIC;
  SIGNAL or_1390_nl : STD_LOGIC;
  SIGNAL or_1389_nl : STD_LOGIC;
  SIGNAL mux_1526_nl : STD_LOGIC;
  SIGNAL mux_1525_nl : STD_LOGIC;
  SIGNAL or_1387_nl : STD_LOGIC;
  SIGNAL or_1385_nl : STD_LOGIC;
  SIGNAL mux_1524_nl : STD_LOGIC;
  SIGNAL or_1384_nl : STD_LOGIC;
  SIGNAL mux_1523_nl : STD_LOGIC;
  SIGNAL or_1382_nl : STD_LOGIC;
  SIGNAL mux_1522_nl : STD_LOGIC;
  SIGNAL mux_1521_nl : STD_LOGIC;
  SIGNAL or_1375_nl : STD_LOGIC;
  SIGNAL or_1374_nl : STD_LOGIC;
  SIGNAL or_1372_nl : STD_LOGIC;
  SIGNAL or_1371_nl : STD_LOGIC;
  SIGNAL mux_1518_nl : STD_LOGIC;
  SIGNAL or_1370_nl : STD_LOGIC;
  SIGNAL mux_1517_nl : STD_LOGIC;
  SIGNAL or_1369_nl : STD_LOGIC;
  SIGNAL mux_1516_nl : STD_LOGIC;
  SIGNAL or_1368_nl : STD_LOGIC;
  SIGNAL or_1367_nl : STD_LOGIC;
  SIGNAL mux_1583_nl : STD_LOGIC;
  SIGNAL mux_1582_nl : STD_LOGIC;
  SIGNAL mux_1581_nl : STD_LOGIC;
  SIGNAL nand_60_nl : STD_LOGIC;
  SIGNAL mux_1580_nl : STD_LOGIC;
  SIGNAL mux_1579_nl : STD_LOGIC;
  SIGNAL nor_681_nl : STD_LOGIC;
  SIGNAL nor_682_nl : STD_LOGIC;
  SIGNAL mux_1578_nl : STD_LOGIC;
  SIGNAL and_773_nl : STD_LOGIC;
  SIGNAL and_779_nl : STD_LOGIC;
  SIGNAL mux_1577_nl : STD_LOGIC;
  SIGNAL nand_59_nl : STD_LOGIC;
  SIGNAL mux_1576_nl : STD_LOGIC;
  SIGNAL nor_685_nl : STD_LOGIC;
  SIGNAL nor_686_nl : STD_LOGIC;
  SIGNAL mux_1575_nl : STD_LOGIC;
  SIGNAL mux_1574_nl : STD_LOGIC;
  SIGNAL or_1465_nl : STD_LOGIC;
  SIGNAL or_1463_nl : STD_LOGIC;
  SIGNAL or_1462_nl : STD_LOGIC;
  SIGNAL mux_1573_nl : STD_LOGIC;
  SIGNAL or_1461_nl : STD_LOGIC;
  SIGNAL mux_1572_nl : STD_LOGIC;
  SIGNAL mux_1571_nl : STD_LOGIC;
  SIGNAL nand_331_nl : STD_LOGIC;
  SIGNAL nand_472_nl : STD_LOGIC;
  SIGNAL mux_1570_nl : STD_LOGIC;
  SIGNAL or_1457_nl : STD_LOGIC;
  SIGNAL or_1455_nl : STD_LOGIC;
  SIGNAL mux_1569_nl : STD_LOGIC;
  SIGNAL or_1453_nl : STD_LOGIC;
  SIGNAL mux_1568_nl : STD_LOGIC;
  SIGNAL or_1452_nl : STD_LOGIC;
  SIGNAL or_1451_nl : STD_LOGIC;
  SIGNAL or_1450_nl : STD_LOGIC;
  SIGNAL mux_1567_nl : STD_LOGIC;
  SIGNAL mux_1566_nl : STD_LOGIC;
  SIGNAL mux_1565_nl : STD_LOGIC;
  SIGNAL mux_1564_nl : STD_LOGIC;
  SIGNAL mux_1563_nl : STD_LOGIC;
  SIGNAL or_1446_nl : STD_LOGIC;
  SIGNAL mux_1562_nl : STD_LOGIC;
  SIGNAL or_1445_nl : STD_LOGIC;
  SIGNAL nand_57_nl : STD_LOGIC;
  SIGNAL mux_1560_nl : STD_LOGIC;
  SIGNAL mux_1559_nl : STD_LOGIC;
  SIGNAL nor_687_nl : STD_LOGIC;
  SIGNAL nor_688_nl : STD_LOGIC;
  SIGNAL mux_1558_nl : STD_LOGIC;
  SIGNAL and_789_nl : STD_LOGIC;
  SIGNAL and_790_nl : STD_LOGIC;
  SIGNAL mux_1557_nl : STD_LOGIC;
  SIGNAL mux_1556_nl : STD_LOGIC;
  SIGNAL mux_1555_nl : STD_LOGIC;
  SIGNAL or_1434_nl : STD_LOGIC;
  SIGNAL mux_1554_nl : STD_LOGIC;
  SIGNAL or_1432_nl : STD_LOGIC;
  SIGNAL or_1430_nl : STD_LOGIC;
  SIGNAL or_1429_nl : STD_LOGIC;
  SIGNAL mux_1553_nl : STD_LOGIC;
  SIGNAL or_1428_nl : STD_LOGIC;
  SIGNAL or_1427_nl : STD_LOGIC;
  SIGNAL or_1426_nl : STD_LOGIC;
  SIGNAL mux_1552_nl : STD_LOGIC;
  SIGNAL mux_1551_nl : STD_LOGIC;
  SIGNAL nand_336_nl : STD_LOGIC;
  SIGNAL nand_453_nl : STD_LOGIC;
  SIGNAL or_1422_nl : STD_LOGIC;
  SIGNAL mux_1618_nl : STD_LOGIC;
  SIGNAL mux_1617_nl : STD_LOGIC;
  SIGNAL mux_1616_nl : STD_LOGIC;
  SIGNAL mux_1615_nl : STD_LOGIC;
  SIGNAL or_1526_nl : STD_LOGIC;
  SIGNAL mux_1614_nl : STD_LOGIC;
  SIGNAL nand_317_nl : STD_LOGIC;
  SIGNAL mux_1613_nl : STD_LOGIC;
  SIGNAL or_1523_nl : STD_LOGIC;
  SIGNAL or_1522_nl : STD_LOGIC;
  SIGNAL mux_1612_nl : STD_LOGIC;
  SIGNAL mux_1611_nl : STD_LOGIC;
  SIGNAL mux_1610_nl : STD_LOGIC;
  SIGNAL or_1521_nl : STD_LOGIC;
  SIGNAL or_1519_nl : STD_LOGIC;
  SIGNAL or_1517_nl : STD_LOGIC;
  SIGNAL or_1515_nl : STD_LOGIC;
  SIGNAL mux_1609_nl : STD_LOGIC;
  SIGNAL mux_1608_nl : STD_LOGIC;
  SIGNAL mux_1607_nl : STD_LOGIC;
  SIGNAL mux_1606_nl : STD_LOGIC;
  SIGNAL nand_318_nl : STD_LOGIC;
  SIGNAL nand_319_nl : STD_LOGIC;
  SIGNAL or_1512_nl : STD_LOGIC;
  SIGNAL or_1511_nl : STD_LOGIC;
  SIGNAL mux_1605_nl : STD_LOGIC;
  SIGNAL mux_1604_nl : STD_LOGIC;
  SIGNAL nand_320_nl : STD_LOGIC;
  SIGNAL mux_1603_nl : STD_LOGIC;
  SIGNAL or_1508_nl : STD_LOGIC;
  SIGNAL or_1507_nl : STD_LOGIC;
  SIGNAL or_1506_nl : STD_LOGIC;
  SIGNAL mux_1602_nl : STD_LOGIC;
  SIGNAL mux_1601_nl : STD_LOGIC;
  SIGNAL mux_1600_nl : STD_LOGIC;
  SIGNAL mux_1599_nl : STD_LOGIC;
  SIGNAL mux_1598_nl : STD_LOGIC;
  SIGNAL or_1505_nl : STD_LOGIC;
  SIGNAL or_1503_nl : STD_LOGIC;
  SIGNAL or_1501_nl : STD_LOGIC;
  SIGNAL nand_62_nl : STD_LOGIC;
  SIGNAL mux_1597_nl : STD_LOGIC;
  SIGNAL mux_1596_nl : STD_LOGIC;
  SIGNAL nand_467_nl : STD_LOGIC;
  SIGNAL mux_1595_nl : STD_LOGIC;
  SIGNAL nand_323_nl : STD_LOGIC;
  SIGNAL and_546_nl : STD_LOGIC;
  SIGNAL nand_463_nl : STD_LOGIC;
  SIGNAL mux_1594_nl : STD_LOGIC;
  SIGNAL mux_1593_nl : STD_LOGIC;
  SIGNAL or_1494_nl : STD_LOGIC;
  SIGNAL or_1492_nl : STD_LOGIC;
  SIGNAL mux_1592_nl : STD_LOGIC;
  SIGNAL or_1491_nl : STD_LOGIC;
  SIGNAL mux_1591_nl : STD_LOGIC;
  SIGNAL or_1489_nl : STD_LOGIC;
  SIGNAL mux_1590_nl : STD_LOGIC;
  SIGNAL or_1487_nl : STD_LOGIC;
  SIGNAL mux_1589_nl : STD_LOGIC;
  SIGNAL and_547_nl : STD_LOGIC;
  SIGNAL and_548_nl : STD_LOGIC;
  SIGNAL or_1480_nl : STD_LOGIC;
  SIGNAL mux_1586_nl : STD_LOGIC;
  SIGNAL or_1479_nl : STD_LOGIC;
  SIGNAL mux_1585_nl : STD_LOGIC;
  SIGNAL or_1478_nl : STD_LOGIC;
  SIGNAL mux_1584_nl : STD_LOGIC;
  SIGNAL or_1477_nl : STD_LOGIC;
  SIGNAL or_1476_nl : STD_LOGIC;
  SIGNAL mux_1651_nl : STD_LOGIC;
  SIGNAL mux_1650_nl : STD_LOGIC;
  SIGNAL mux_1649_nl : STD_LOGIC;
  SIGNAL nand_66_nl : STD_LOGIC;
  SIGNAL mux_1648_nl : STD_LOGIC;
  SIGNAL mux_1647_nl : STD_LOGIC;
  SIGNAL nor_669_nl : STD_LOGIC;
  SIGNAL nor_670_nl : STD_LOGIC;
  SIGNAL mux_1646_nl : STD_LOGIC;
  SIGNAL nor_671_nl : STD_LOGIC;
  SIGNAL nor_672_nl : STD_LOGIC;
  SIGNAL mux_1645_nl : STD_LOGIC;
  SIGNAL nand_65_nl : STD_LOGIC;
  SIGNAL mux_1644_nl : STD_LOGIC;
  SIGNAL nor_673_nl : STD_LOGIC;
  SIGNAL nor_674_nl : STD_LOGIC;
  SIGNAL mux_1643_nl : STD_LOGIC;
  SIGNAL mux_1642_nl : STD_LOGIC;
  SIGNAL or_1571_nl : STD_LOGIC;
  SIGNAL or_1569_nl : STD_LOGIC;
  SIGNAL or_1568_nl : STD_LOGIC;
  SIGNAL mux_1641_nl : STD_LOGIC;
  SIGNAL or_1567_nl : STD_LOGIC;
  SIGNAL mux_1640_nl : STD_LOGIC;
  SIGNAL mux_1639_nl : STD_LOGIC;
  SIGNAL or_1566_nl : STD_LOGIC;
  SIGNAL or_1565_nl : STD_LOGIC;
  SIGNAL mux_1638_nl : STD_LOGIC;
  SIGNAL or_1563_nl : STD_LOGIC;
  SIGNAL or_1561_nl : STD_LOGIC;
  SIGNAL mux_1637_nl : STD_LOGIC;
  SIGNAL or_1559_nl : STD_LOGIC;
  SIGNAL mux_1636_nl : STD_LOGIC;
  SIGNAL or_1558_nl : STD_LOGIC;
  SIGNAL or_1557_nl : STD_LOGIC;
  SIGNAL or_1556_nl : STD_LOGIC;
  SIGNAL mux_1635_nl : STD_LOGIC;
  SIGNAL mux_1634_nl : STD_LOGIC;
  SIGNAL mux_1633_nl : STD_LOGIC;
  SIGNAL mux_1632_nl : STD_LOGIC;
  SIGNAL or_1554_nl : STD_LOGIC;
  SIGNAL mux_1631_nl : STD_LOGIC;
  SIGNAL mux_1630_nl : STD_LOGIC;
  SIGNAL or_1551_nl : STD_LOGIC;
  SIGNAL nand_63_nl : STD_LOGIC;
  SIGNAL mux_1628_nl : STD_LOGIC;
  SIGNAL mux_1627_nl : STD_LOGIC;
  SIGNAL nor_675_nl : STD_LOGIC;
  SIGNAL nor_676_nl : STD_LOGIC;
  SIGNAL mux_1626_nl : STD_LOGIC;
  SIGNAL nor_677_nl : STD_LOGIC;
  SIGNAL nor_678_nl : STD_LOGIC;
  SIGNAL mux_1625_nl : STD_LOGIC;
  SIGNAL mux_1624_nl : STD_LOGIC;
  SIGNAL mux_1623_nl : STD_LOGIC;
  SIGNAL or_1540_nl : STD_LOGIC;
  SIGNAL mux_1622_nl : STD_LOGIC;
  SIGNAL or_1538_nl : STD_LOGIC;
  SIGNAL or_1536_nl : STD_LOGIC;
  SIGNAL or_1535_nl : STD_LOGIC;
  SIGNAL mux_1621_nl : STD_LOGIC;
  SIGNAL or_1534_nl : STD_LOGIC;
  SIGNAL or_1533_nl : STD_LOGIC;
  SIGNAL or_1532_nl : STD_LOGIC;
  SIGNAL mux_1620_nl : STD_LOGIC;
  SIGNAL mux_1619_nl : STD_LOGIC;
  SIGNAL or_1531_nl : STD_LOGIC;
  SIGNAL or_1530_nl : STD_LOGIC;
  SIGNAL or_1528_nl : STD_LOGIC;
  SIGNAL mux_1686_nl : STD_LOGIC;
  SIGNAL mux_1685_nl : STD_LOGIC;
  SIGNAL mux_1684_nl : STD_LOGIC;
  SIGNAL mux_1683_nl : STD_LOGIC;
  SIGNAL or_1635_nl : STD_LOGIC;
  SIGNAL mux_1682_nl : STD_LOGIC;
  SIGNAL or_1633_nl : STD_LOGIC;
  SIGNAL mux_1681_nl : STD_LOGIC;
  SIGNAL or_1632_nl : STD_LOGIC;
  SIGNAL or_1631_nl : STD_LOGIC;
  SIGNAL mux_1680_nl : STD_LOGIC;
  SIGNAL mux_1679_nl : STD_LOGIC;
  SIGNAL mux_1678_nl : STD_LOGIC;
  SIGNAL or_1630_nl : STD_LOGIC;
  SIGNAL or_1628_nl : STD_LOGIC;
  SIGNAL or_1626_nl : STD_LOGIC;
  SIGNAL or_1624_nl : STD_LOGIC;
  SIGNAL mux_1677_nl : STD_LOGIC;
  SIGNAL mux_1676_nl : STD_LOGIC;
  SIGNAL mux_1675_nl : STD_LOGIC;
  SIGNAL mux_1674_nl : STD_LOGIC;
  SIGNAL or_1623_nl : STD_LOGIC;
  SIGNAL or_1622_nl : STD_LOGIC;
  SIGNAL or_1621_nl : STD_LOGIC;
  SIGNAL or_1620_nl : STD_LOGIC;
  SIGNAL mux_1673_nl : STD_LOGIC;
  SIGNAL mux_1672_nl : STD_LOGIC;
  SIGNAL or_1618_nl : STD_LOGIC;
  SIGNAL mux_1671_nl : STD_LOGIC;
  SIGNAL or_1617_nl : STD_LOGIC;
  SIGNAL or_1616_nl : STD_LOGIC;
  SIGNAL or_1615_nl : STD_LOGIC;
  SIGNAL mux_1670_nl : STD_LOGIC;
  SIGNAL mux_1669_nl : STD_LOGIC;
  SIGNAL mux_1668_nl : STD_LOGIC;
  SIGNAL mux_1667_nl : STD_LOGIC;
  SIGNAL mux_1666_nl : STD_LOGIC;
  SIGNAL or_1614_nl : STD_LOGIC;
  SIGNAL or_1612_nl : STD_LOGIC;
  SIGNAL or_1610_nl : STD_LOGIC;
  SIGNAL nand_68_nl : STD_LOGIC;
  SIGNAL mux_1665_nl : STD_LOGIC;
  SIGNAL mux_1664_nl : STD_LOGIC;
  SIGNAL mux_1663_nl : STD_LOGIC;
  SIGNAL or_1608_nl : STD_LOGIC;
  SIGNAL or_1607_nl : STD_LOGIC;
  SIGNAL or_1605_nl : STD_LOGIC;
  SIGNAL or_1604_nl : STD_LOGIC;
  SIGNAL mux_1662_nl : STD_LOGIC;
  SIGNAL mux_1661_nl : STD_LOGIC;
  SIGNAL or_1602_nl : STD_LOGIC;
  SIGNAL or_1600_nl : STD_LOGIC;
  SIGNAL mux_1660_nl : STD_LOGIC;
  SIGNAL or_1599_nl : STD_LOGIC;
  SIGNAL mux_1659_nl : STD_LOGIC;
  SIGNAL or_1597_nl : STD_LOGIC;
  SIGNAL mux_1658_nl : STD_LOGIC;
  SIGNAL mux_1657_nl : STD_LOGIC;
  SIGNAL or_1590_nl : STD_LOGIC;
  SIGNAL or_1589_nl : STD_LOGIC;
  SIGNAL or_1587_nl : STD_LOGIC;
  SIGNAL or_1586_nl : STD_LOGIC;
  SIGNAL mux_1654_nl : STD_LOGIC;
  SIGNAL or_1585_nl : STD_LOGIC;
  SIGNAL mux_1653_nl : STD_LOGIC;
  SIGNAL or_1584_nl : STD_LOGIC;
  SIGNAL mux_1652_nl : STD_LOGIC;
  SIGNAL or_1583_nl : STD_LOGIC;
  SIGNAL or_1582_nl : STD_LOGIC;
  SIGNAL mux_1719_nl : STD_LOGIC;
  SIGNAL mux_1718_nl : STD_LOGIC;
  SIGNAL mux_1717_nl : STD_LOGIC;
  SIGNAL nand_72_nl : STD_LOGIC;
  SIGNAL mux_1716_nl : STD_LOGIC;
  SIGNAL mux_1715_nl : STD_LOGIC;
  SIGNAL nor_657_nl : STD_LOGIC;
  SIGNAL nor_658_nl : STD_LOGIC;
  SIGNAL mux_1714_nl : STD_LOGIC;
  SIGNAL nor_659_nl : STD_LOGIC;
  SIGNAL nor_660_nl : STD_LOGIC;
  SIGNAL mux_1713_nl : STD_LOGIC;
  SIGNAL nand_71_nl : STD_LOGIC;
  SIGNAL mux_1712_nl : STD_LOGIC;
  SIGNAL nor_661_nl : STD_LOGIC;
  SIGNAL nor_662_nl : STD_LOGIC;
  SIGNAL mux_1711_nl : STD_LOGIC;
  SIGNAL mux_1710_nl : STD_LOGIC;
  SIGNAL or_1680_nl : STD_LOGIC;
  SIGNAL or_1678_nl : STD_LOGIC;
  SIGNAL or_1677_nl : STD_LOGIC;
  SIGNAL mux_1709_nl : STD_LOGIC;
  SIGNAL or_1676_nl : STD_LOGIC;
  SIGNAL mux_1708_nl : STD_LOGIC;
  SIGNAL mux_1707_nl : STD_LOGIC;
  SIGNAL or_1675_nl : STD_LOGIC;
  SIGNAL or_1674_nl : STD_LOGIC;
  SIGNAL mux_1706_nl : STD_LOGIC;
  SIGNAL or_1672_nl : STD_LOGIC;
  SIGNAL or_1670_nl : STD_LOGIC;
  SIGNAL mux_1705_nl : STD_LOGIC;
  SIGNAL or_1668_nl : STD_LOGIC;
  SIGNAL mux_1704_nl : STD_LOGIC;
  SIGNAL or_1667_nl : STD_LOGIC;
  SIGNAL or_1666_nl : STD_LOGIC;
  SIGNAL or_1665_nl : STD_LOGIC;
  SIGNAL mux_1703_nl : STD_LOGIC;
  SIGNAL mux_1702_nl : STD_LOGIC;
  SIGNAL mux_1701_nl : STD_LOGIC;
  SIGNAL mux_1700_nl : STD_LOGIC;
  SIGNAL or_1663_nl : STD_LOGIC;
  SIGNAL mux_1699_nl : STD_LOGIC;
  SIGNAL mux_1698_nl : STD_LOGIC;
  SIGNAL or_1660_nl : STD_LOGIC;
  SIGNAL nand_69_nl : STD_LOGIC;
  SIGNAL mux_1696_nl : STD_LOGIC;
  SIGNAL mux_1695_nl : STD_LOGIC;
  SIGNAL nor_663_nl : STD_LOGIC;
  SIGNAL nor_664_nl : STD_LOGIC;
  SIGNAL mux_1694_nl : STD_LOGIC;
  SIGNAL nor_665_nl : STD_LOGIC;
  SIGNAL nor_666_nl : STD_LOGIC;
  SIGNAL mux_1693_nl : STD_LOGIC;
  SIGNAL mux_1692_nl : STD_LOGIC;
  SIGNAL mux_1691_nl : STD_LOGIC;
  SIGNAL or_1649_nl : STD_LOGIC;
  SIGNAL mux_1690_nl : STD_LOGIC;
  SIGNAL or_1647_nl : STD_LOGIC;
  SIGNAL or_1645_nl : STD_LOGIC;
  SIGNAL or_1644_nl : STD_LOGIC;
  SIGNAL mux_1689_nl : STD_LOGIC;
  SIGNAL or_1643_nl : STD_LOGIC;
  SIGNAL or_1642_nl : STD_LOGIC;
  SIGNAL or_1641_nl : STD_LOGIC;
  SIGNAL mux_1688_nl : STD_LOGIC;
  SIGNAL mux_1687_nl : STD_LOGIC;
  SIGNAL or_1640_nl : STD_LOGIC;
  SIGNAL or_1639_nl : STD_LOGIC;
  SIGNAL or_1637_nl : STD_LOGIC;
  SIGNAL mux_1754_nl : STD_LOGIC;
  SIGNAL mux_1753_nl : STD_LOGIC;
  SIGNAL mux_1752_nl : STD_LOGIC;
  SIGNAL mux_1751_nl : STD_LOGIC;
  SIGNAL or_1741_nl : STD_LOGIC;
  SIGNAL mux_1750_nl : STD_LOGIC;
  SIGNAL or_1739_nl : STD_LOGIC;
  SIGNAL mux_1749_nl : STD_LOGIC;
  SIGNAL or_1738_nl : STD_LOGIC;
  SIGNAL or_1737_nl : STD_LOGIC;
  SIGNAL mux_1748_nl : STD_LOGIC;
  SIGNAL mux_1747_nl : STD_LOGIC;
  SIGNAL mux_1746_nl : STD_LOGIC;
  SIGNAL or_1736_nl : STD_LOGIC;
  SIGNAL or_1734_nl : STD_LOGIC;
  SIGNAL or_1732_nl : STD_LOGIC;
  SIGNAL or_1730_nl : STD_LOGIC;
  SIGNAL mux_1745_nl : STD_LOGIC;
  SIGNAL mux_1744_nl : STD_LOGIC;
  SIGNAL mux_1743_nl : STD_LOGIC;
  SIGNAL mux_1742_nl : STD_LOGIC;
  SIGNAL or_1729_nl : STD_LOGIC;
  SIGNAL or_1728_nl : STD_LOGIC;
  SIGNAL or_1727_nl : STD_LOGIC;
  SIGNAL or_1726_nl : STD_LOGIC;
  SIGNAL mux_1741_nl : STD_LOGIC;
  SIGNAL mux_1740_nl : STD_LOGIC;
  SIGNAL nand_306_nl : STD_LOGIC;
  SIGNAL mux_1739_nl : STD_LOGIC;
  SIGNAL or_1723_nl : STD_LOGIC;
  SIGNAL or_1722_nl : STD_LOGIC;
  SIGNAL or_1721_nl : STD_LOGIC;
  SIGNAL mux_1738_nl : STD_LOGIC;
  SIGNAL mux_1737_nl : STD_LOGIC;
  SIGNAL mux_1736_nl : STD_LOGIC;
  SIGNAL mux_1735_nl : STD_LOGIC;
  SIGNAL mux_1734_nl : STD_LOGIC;
  SIGNAL or_1720_nl : STD_LOGIC;
  SIGNAL or_1718_nl : STD_LOGIC;
  SIGNAL or_1716_nl : STD_LOGIC;
  SIGNAL nand_74_nl : STD_LOGIC;
  SIGNAL mux_1733_nl : STD_LOGIC;
  SIGNAL mux_1732_nl : STD_LOGIC;
  SIGNAL or_1714_nl : STD_LOGIC;
  SIGNAL mux_1731_nl : STD_LOGIC;
  SIGNAL or_1712_nl : STD_LOGIC;
  SIGNAL nor_321_nl : STD_LOGIC;
  SIGNAL or_1711_nl : STD_LOGIC;
  SIGNAL mux_1730_nl : STD_LOGIC;
  SIGNAL mux_1729_nl : STD_LOGIC;
  SIGNAL or_1709_nl : STD_LOGIC;
  SIGNAL or_1707_nl : STD_LOGIC;
  SIGNAL mux_1728_nl : STD_LOGIC;
  SIGNAL or_1706_nl : STD_LOGIC;
  SIGNAL mux_1727_nl : STD_LOGIC;
  SIGNAL or_1704_nl : STD_LOGIC;
  SIGNAL mux_1726_nl : STD_LOGIC;
  SIGNAL or_1702_nl : STD_LOGIC;
  SIGNAL mux_1725_nl : STD_LOGIC;
  SIGNAL nor_319_nl : STD_LOGIC;
  SIGNAL nor_318_nl : STD_LOGIC;
  SIGNAL or_1695_nl : STD_LOGIC;
  SIGNAL mux_1722_nl : STD_LOGIC;
  SIGNAL or_1694_nl : STD_LOGIC;
  SIGNAL mux_1721_nl : STD_LOGIC;
  SIGNAL or_1693_nl : STD_LOGIC;
  SIGNAL mux_1720_nl : STD_LOGIC;
  SIGNAL or_1692_nl : STD_LOGIC;
  SIGNAL or_1691_nl : STD_LOGIC;
  SIGNAL mux_1787_nl : STD_LOGIC;
  SIGNAL mux_1786_nl : STD_LOGIC;
  SIGNAL mux_1785_nl : STD_LOGIC;
  SIGNAL nand_78_nl : STD_LOGIC;
  SIGNAL mux_1784_nl : STD_LOGIC;
  SIGNAL mux_1783_nl : STD_LOGIC;
  SIGNAL nor_645_nl : STD_LOGIC;
  SIGNAL nor_646_nl : STD_LOGIC;
  SIGNAL mux_1782_nl : STD_LOGIC;
  SIGNAL nor_647_nl : STD_LOGIC;
  SIGNAL nor_648_nl : STD_LOGIC;
  SIGNAL mux_1781_nl : STD_LOGIC;
  SIGNAL nand_77_nl : STD_LOGIC;
  SIGNAL mux_1780_nl : STD_LOGIC;
  SIGNAL nor_649_nl : STD_LOGIC;
  SIGNAL nor_650_nl : STD_LOGIC;
  SIGNAL mux_1779_nl : STD_LOGIC;
  SIGNAL mux_1778_nl : STD_LOGIC;
  SIGNAL or_1786_nl : STD_LOGIC;
  SIGNAL or_1784_nl : STD_LOGIC;
  SIGNAL or_1783_nl : STD_LOGIC;
  SIGNAL mux_1777_nl : STD_LOGIC;
  SIGNAL or_1782_nl : STD_LOGIC;
  SIGNAL mux_1776_nl : STD_LOGIC;
  SIGNAL mux_1775_nl : STD_LOGIC;
  SIGNAL or_1781_nl : STD_LOGIC;
  SIGNAL or_1780_nl : STD_LOGIC;
  SIGNAL mux_1774_nl : STD_LOGIC;
  SIGNAL or_1778_nl : STD_LOGIC;
  SIGNAL or_1776_nl : STD_LOGIC;
  SIGNAL mux_1773_nl : STD_LOGIC;
  SIGNAL or_1774_nl : STD_LOGIC;
  SIGNAL mux_1772_nl : STD_LOGIC;
  SIGNAL or_1773_nl : STD_LOGIC;
  SIGNAL or_1772_nl : STD_LOGIC;
  SIGNAL or_1771_nl : STD_LOGIC;
  SIGNAL mux_1771_nl : STD_LOGIC;
  SIGNAL mux_1770_nl : STD_LOGIC;
  SIGNAL mux_1769_nl : STD_LOGIC;
  SIGNAL mux_1768_nl : STD_LOGIC;
  SIGNAL or_1769_nl : STD_LOGIC;
  SIGNAL mux_1767_nl : STD_LOGIC;
  SIGNAL mux_1766_nl : STD_LOGIC;
  SIGNAL or_1766_nl : STD_LOGIC;
  SIGNAL nand_75_nl : STD_LOGIC;
  SIGNAL mux_1764_nl : STD_LOGIC;
  SIGNAL mux_1763_nl : STD_LOGIC;
  SIGNAL nor_651_nl : STD_LOGIC;
  SIGNAL nor_652_nl : STD_LOGIC;
  SIGNAL mux_1762_nl : STD_LOGIC;
  SIGNAL nor_653_nl : STD_LOGIC;
  SIGNAL nor_654_nl : STD_LOGIC;
  SIGNAL mux_1761_nl : STD_LOGIC;
  SIGNAL mux_1760_nl : STD_LOGIC;
  SIGNAL mux_1759_nl : STD_LOGIC;
  SIGNAL or_1755_nl : STD_LOGIC;
  SIGNAL mux_1758_nl : STD_LOGIC;
  SIGNAL or_1753_nl : STD_LOGIC;
  SIGNAL or_1751_nl : STD_LOGIC;
  SIGNAL or_1750_nl : STD_LOGIC;
  SIGNAL mux_1757_nl : STD_LOGIC;
  SIGNAL or_1749_nl : STD_LOGIC;
  SIGNAL or_1748_nl : STD_LOGIC;
  SIGNAL or_1747_nl : STD_LOGIC;
  SIGNAL mux_1756_nl : STD_LOGIC;
  SIGNAL mux_1755_nl : STD_LOGIC;
  SIGNAL or_1746_nl : STD_LOGIC;
  SIGNAL or_1745_nl : STD_LOGIC;
  SIGNAL or_1743_nl : STD_LOGIC;
  SIGNAL mux_1822_nl : STD_LOGIC;
  SIGNAL mux_1821_nl : STD_LOGIC;
  SIGNAL mux_1820_nl : STD_LOGIC;
  SIGNAL mux_1819_nl : STD_LOGIC;
  SIGNAL or_1850_nl : STD_LOGIC;
  SIGNAL mux_1818_nl : STD_LOGIC;
  SIGNAL or_1848_nl : STD_LOGIC;
  SIGNAL mux_1817_nl : STD_LOGIC;
  SIGNAL or_1847_nl : STD_LOGIC;
  SIGNAL or_1846_nl : STD_LOGIC;
  SIGNAL mux_1816_nl : STD_LOGIC;
  SIGNAL mux_1815_nl : STD_LOGIC;
  SIGNAL mux_1814_nl : STD_LOGIC;
  SIGNAL or_1845_nl : STD_LOGIC;
  SIGNAL or_1843_nl : STD_LOGIC;
  SIGNAL or_1841_nl : STD_LOGIC;
  SIGNAL or_1839_nl : STD_LOGIC;
  SIGNAL mux_1813_nl : STD_LOGIC;
  SIGNAL mux_1812_nl : STD_LOGIC;
  SIGNAL mux_1811_nl : STD_LOGIC;
  SIGNAL mux_1810_nl : STD_LOGIC;
  SIGNAL or_1838_nl : STD_LOGIC;
  SIGNAL or_1837_nl : STD_LOGIC;
  SIGNAL or_1836_nl : STD_LOGIC;
  SIGNAL or_1835_nl : STD_LOGIC;
  SIGNAL mux_1809_nl : STD_LOGIC;
  SIGNAL mux_1808_nl : STD_LOGIC;
  SIGNAL nand_300_nl : STD_LOGIC;
  SIGNAL mux_1807_nl : STD_LOGIC;
  SIGNAL or_1832_nl : STD_LOGIC;
  SIGNAL or_1831_nl : STD_LOGIC;
  SIGNAL or_1830_nl : STD_LOGIC;
  SIGNAL mux_1806_nl : STD_LOGIC;
  SIGNAL mux_1805_nl : STD_LOGIC;
  SIGNAL mux_1804_nl : STD_LOGIC;
  SIGNAL mux_1803_nl : STD_LOGIC;
  SIGNAL mux_1802_nl : STD_LOGIC;
  SIGNAL or_1829_nl : STD_LOGIC;
  SIGNAL or_1827_nl : STD_LOGIC;
  SIGNAL or_1825_nl : STD_LOGIC;
  SIGNAL nand_80_nl : STD_LOGIC;
  SIGNAL mux_1801_nl : STD_LOGIC;
  SIGNAL mux_1800_nl : STD_LOGIC;
  SIGNAL mux_1799_nl : STD_LOGIC;
  SIGNAL or_1823_nl : STD_LOGIC;
  SIGNAL or_1822_nl : STD_LOGIC;
  SIGNAL or_1820_nl : STD_LOGIC;
  SIGNAL or_1819_nl : STD_LOGIC;
  SIGNAL mux_1798_nl : STD_LOGIC;
  SIGNAL mux_1797_nl : STD_LOGIC;
  SIGNAL or_1817_nl : STD_LOGIC;
  SIGNAL or_1815_nl : STD_LOGIC;
  SIGNAL mux_1796_nl : STD_LOGIC;
  SIGNAL or_1814_nl : STD_LOGIC;
  SIGNAL mux_1795_nl : STD_LOGIC;
  SIGNAL or_1812_nl : STD_LOGIC;
  SIGNAL mux_1794_nl : STD_LOGIC;
  SIGNAL mux_1793_nl : STD_LOGIC;
  SIGNAL or_1805_nl : STD_LOGIC;
  SIGNAL or_1804_nl : STD_LOGIC;
  SIGNAL or_1802_nl : STD_LOGIC;
  SIGNAL or_1801_nl : STD_LOGIC;
  SIGNAL mux_1790_nl : STD_LOGIC;
  SIGNAL or_1800_nl : STD_LOGIC;
  SIGNAL mux_1789_nl : STD_LOGIC;
  SIGNAL or_1799_nl : STD_LOGIC;
  SIGNAL mux_1788_nl : STD_LOGIC;
  SIGNAL or_1798_nl : STD_LOGIC;
  SIGNAL or_1797_nl : STD_LOGIC;
  SIGNAL mux_1855_nl : STD_LOGIC;
  SIGNAL mux_1854_nl : STD_LOGIC;
  SIGNAL mux_1853_nl : STD_LOGIC;
  SIGNAL nand_84_nl : STD_LOGIC;
  SIGNAL mux_1852_nl : STD_LOGIC;
  SIGNAL mux_1851_nl : STD_LOGIC;
  SIGNAL nor_633_nl : STD_LOGIC;
  SIGNAL nor_634_nl : STD_LOGIC;
  SIGNAL mux_1850_nl : STD_LOGIC;
  SIGNAL and_772_nl : STD_LOGIC;
  SIGNAL and_778_nl : STD_LOGIC;
  SIGNAL mux_1849_nl : STD_LOGIC;
  SIGNAL nand_83_nl : STD_LOGIC;
  SIGNAL mux_1848_nl : STD_LOGIC;
  SIGNAL nor_637_nl : STD_LOGIC;
  SIGNAL nor_638_nl : STD_LOGIC;
  SIGNAL mux_1847_nl : STD_LOGIC;
  SIGNAL mux_1846_nl : STD_LOGIC;
  SIGNAL or_1895_nl : STD_LOGIC;
  SIGNAL or_1893_nl : STD_LOGIC;
  SIGNAL or_1892_nl : STD_LOGIC;
  SIGNAL mux_1845_nl : STD_LOGIC;
  SIGNAL or_1891_nl : STD_LOGIC;
  SIGNAL mux_1844_nl : STD_LOGIC;
  SIGNAL mux_1843_nl : STD_LOGIC;
  SIGNAL nand_291_nl : STD_LOGIC;
  SIGNAL nand_471_nl : STD_LOGIC;
  SIGNAL mux_1842_nl : STD_LOGIC;
  SIGNAL or_1887_nl : STD_LOGIC;
  SIGNAL or_1885_nl : STD_LOGIC;
  SIGNAL mux_1841_nl : STD_LOGIC;
  SIGNAL or_1883_nl : STD_LOGIC;
  SIGNAL mux_1840_nl : STD_LOGIC;
  SIGNAL or_1882_nl : STD_LOGIC;
  SIGNAL or_1881_nl : STD_LOGIC;
  SIGNAL or_1880_nl : STD_LOGIC;
  SIGNAL mux_1839_nl : STD_LOGIC;
  SIGNAL mux_1838_nl : STD_LOGIC;
  SIGNAL mux_1837_nl : STD_LOGIC;
  SIGNAL mux_1836_nl : STD_LOGIC;
  SIGNAL or_1878_nl : STD_LOGIC;
  SIGNAL mux_1835_nl : STD_LOGIC;
  SIGNAL mux_1834_nl : STD_LOGIC;
  SIGNAL or_1875_nl : STD_LOGIC;
  SIGNAL nand_81_nl : STD_LOGIC;
  SIGNAL mux_1832_nl : STD_LOGIC;
  SIGNAL mux_1831_nl : STD_LOGIC;
  SIGNAL nor_639_nl : STD_LOGIC;
  SIGNAL nor_640_nl : STD_LOGIC;
  SIGNAL mux_1830_nl : STD_LOGIC;
  SIGNAL and_787_nl : STD_LOGIC;
  SIGNAL and_788_nl : STD_LOGIC;
  SIGNAL mux_1829_nl : STD_LOGIC;
  SIGNAL mux_1828_nl : STD_LOGIC;
  SIGNAL mux_1827_nl : STD_LOGIC;
  SIGNAL or_1864_nl : STD_LOGIC;
  SIGNAL mux_1826_nl : STD_LOGIC;
  SIGNAL or_1862_nl : STD_LOGIC;
  SIGNAL or_1860_nl : STD_LOGIC;
  SIGNAL or_1859_nl : STD_LOGIC;
  SIGNAL mux_1825_nl : STD_LOGIC;
  SIGNAL or_1858_nl : STD_LOGIC;
  SIGNAL or_1857_nl : STD_LOGIC;
  SIGNAL or_1856_nl : STD_LOGIC;
  SIGNAL mux_1824_nl : STD_LOGIC;
  SIGNAL mux_1823_nl : STD_LOGIC;
  SIGNAL nand_296_nl : STD_LOGIC;
  SIGNAL nand_452_nl : STD_LOGIC;
  SIGNAL or_1852_nl : STD_LOGIC;
  SIGNAL mux_1890_nl : STD_LOGIC;
  SIGNAL mux_1889_nl : STD_LOGIC;
  SIGNAL mux_1888_nl : STD_LOGIC;
  SIGNAL mux_1887_nl : STD_LOGIC;
  SIGNAL or_1956_nl : STD_LOGIC;
  SIGNAL mux_1886_nl : STD_LOGIC;
  SIGNAL nand_277_nl : STD_LOGIC;
  SIGNAL mux_1885_nl : STD_LOGIC;
  SIGNAL or_1953_nl : STD_LOGIC;
  SIGNAL or_1952_nl : STD_LOGIC;
  SIGNAL mux_1884_nl : STD_LOGIC;
  SIGNAL mux_1883_nl : STD_LOGIC;
  SIGNAL mux_1882_nl : STD_LOGIC;
  SIGNAL or_1951_nl : STD_LOGIC;
  SIGNAL or_1949_nl : STD_LOGIC;
  SIGNAL or_1947_nl : STD_LOGIC;
  SIGNAL or_1945_nl : STD_LOGIC;
  SIGNAL mux_1881_nl : STD_LOGIC;
  SIGNAL mux_1880_nl : STD_LOGIC;
  SIGNAL mux_1879_nl : STD_LOGIC;
  SIGNAL mux_1878_nl : STD_LOGIC;
  SIGNAL nand_278_nl : STD_LOGIC;
  SIGNAL nand_279_nl : STD_LOGIC;
  SIGNAL or_1942_nl : STD_LOGIC;
  SIGNAL or_1941_nl : STD_LOGIC;
  SIGNAL mux_1877_nl : STD_LOGIC;
  SIGNAL mux_1876_nl : STD_LOGIC;
  SIGNAL nand_280_nl : STD_LOGIC;
  SIGNAL mux_1875_nl : STD_LOGIC;
  SIGNAL or_1938_nl : STD_LOGIC;
  SIGNAL or_1937_nl : STD_LOGIC;
  SIGNAL or_1936_nl : STD_LOGIC;
  SIGNAL mux_1874_nl : STD_LOGIC;
  SIGNAL mux_1873_nl : STD_LOGIC;
  SIGNAL mux_1872_nl : STD_LOGIC;
  SIGNAL mux_1871_nl : STD_LOGIC;
  SIGNAL mux_1870_nl : STD_LOGIC;
  SIGNAL or_1935_nl : STD_LOGIC;
  SIGNAL or_1933_nl : STD_LOGIC;
  SIGNAL or_1931_nl : STD_LOGIC;
  SIGNAL nand_86_nl : STD_LOGIC;
  SIGNAL mux_1869_nl : STD_LOGIC;
  SIGNAL mux_1868_nl : STD_LOGIC;
  SIGNAL nand_466_nl : STD_LOGIC;
  SIGNAL mux_1867_nl : STD_LOGIC;
  SIGNAL nand_283_nl : STD_LOGIC;
  SIGNAL and_543_nl : STD_LOGIC;
  SIGNAL nand_462_nl : STD_LOGIC;
  SIGNAL mux_1866_nl : STD_LOGIC;
  SIGNAL mux_1865_nl : STD_LOGIC;
  SIGNAL or_1924_nl : STD_LOGIC;
  SIGNAL or_1922_nl : STD_LOGIC;
  SIGNAL mux_1864_nl : STD_LOGIC;
  SIGNAL or_1921_nl : STD_LOGIC;
  SIGNAL mux_1863_nl : STD_LOGIC;
  SIGNAL or_1919_nl : STD_LOGIC;
  SIGNAL mux_1862_nl : STD_LOGIC;
  SIGNAL or_1917_nl : STD_LOGIC;
  SIGNAL mux_1861_nl : STD_LOGIC;
  SIGNAL and_544_nl : STD_LOGIC;
  SIGNAL and_545_nl : STD_LOGIC;
  SIGNAL or_1910_nl : STD_LOGIC;
  SIGNAL mux_1858_nl : STD_LOGIC;
  SIGNAL or_1909_nl : STD_LOGIC;
  SIGNAL mux_1857_nl : STD_LOGIC;
  SIGNAL or_1908_nl : STD_LOGIC;
  SIGNAL mux_1856_nl : STD_LOGIC;
  SIGNAL or_1907_nl : STD_LOGIC;
  SIGNAL or_1906_nl : STD_LOGIC;
  SIGNAL mux_1923_nl : STD_LOGIC;
  SIGNAL mux_1922_nl : STD_LOGIC;
  SIGNAL mux_1921_nl : STD_LOGIC;
  SIGNAL nand_90_nl : STD_LOGIC;
  SIGNAL mux_1920_nl : STD_LOGIC;
  SIGNAL mux_1919_nl : STD_LOGIC;
  SIGNAL nor_621_nl : STD_LOGIC;
  SIGNAL nor_622_nl : STD_LOGIC;
  SIGNAL mux_1918_nl : STD_LOGIC;
  SIGNAL nor_623_nl : STD_LOGIC;
  SIGNAL nor_624_nl : STD_LOGIC;
  SIGNAL mux_1917_nl : STD_LOGIC;
  SIGNAL nand_89_nl : STD_LOGIC;
  SIGNAL mux_1916_nl : STD_LOGIC;
  SIGNAL nor_625_nl : STD_LOGIC;
  SIGNAL nor_626_nl : STD_LOGIC;
  SIGNAL mux_1915_nl : STD_LOGIC;
  SIGNAL mux_1914_nl : STD_LOGIC;
  SIGNAL or_2001_nl : STD_LOGIC;
  SIGNAL or_1999_nl : STD_LOGIC;
  SIGNAL or_1998_nl : STD_LOGIC;
  SIGNAL mux_1913_nl : STD_LOGIC;
  SIGNAL or_1997_nl : STD_LOGIC;
  SIGNAL mux_1912_nl : STD_LOGIC;
  SIGNAL mux_1911_nl : STD_LOGIC;
  SIGNAL or_1996_nl : STD_LOGIC;
  SIGNAL or_1995_nl : STD_LOGIC;
  SIGNAL mux_1910_nl : STD_LOGIC;
  SIGNAL or_1993_nl : STD_LOGIC;
  SIGNAL or_1991_nl : STD_LOGIC;
  SIGNAL mux_1909_nl : STD_LOGIC;
  SIGNAL or_1989_nl : STD_LOGIC;
  SIGNAL mux_1908_nl : STD_LOGIC;
  SIGNAL or_1988_nl : STD_LOGIC;
  SIGNAL or_1987_nl : STD_LOGIC;
  SIGNAL or_1986_nl : STD_LOGIC;
  SIGNAL mux_1907_nl : STD_LOGIC;
  SIGNAL mux_1906_nl : STD_LOGIC;
  SIGNAL mux_1905_nl : STD_LOGIC;
  SIGNAL mux_1904_nl : STD_LOGIC;
  SIGNAL or_1984_nl : STD_LOGIC;
  SIGNAL mux_1903_nl : STD_LOGIC;
  SIGNAL mux_1902_nl : STD_LOGIC;
  SIGNAL or_1981_nl : STD_LOGIC;
  SIGNAL nand_87_nl : STD_LOGIC;
  SIGNAL mux_1900_nl : STD_LOGIC;
  SIGNAL mux_1899_nl : STD_LOGIC;
  SIGNAL nor_627_nl : STD_LOGIC;
  SIGNAL nor_628_nl : STD_LOGIC;
  SIGNAL mux_1898_nl : STD_LOGIC;
  SIGNAL nor_629_nl : STD_LOGIC;
  SIGNAL nor_630_nl : STD_LOGIC;
  SIGNAL mux_1897_nl : STD_LOGIC;
  SIGNAL mux_1896_nl : STD_LOGIC;
  SIGNAL mux_1895_nl : STD_LOGIC;
  SIGNAL or_1970_nl : STD_LOGIC;
  SIGNAL mux_1894_nl : STD_LOGIC;
  SIGNAL or_1968_nl : STD_LOGIC;
  SIGNAL or_1966_nl : STD_LOGIC;
  SIGNAL or_1965_nl : STD_LOGIC;
  SIGNAL mux_1893_nl : STD_LOGIC;
  SIGNAL or_1964_nl : STD_LOGIC;
  SIGNAL or_1963_nl : STD_LOGIC;
  SIGNAL or_1962_nl : STD_LOGIC;
  SIGNAL mux_1892_nl : STD_LOGIC;
  SIGNAL mux_1891_nl : STD_LOGIC;
  SIGNAL or_1961_nl : STD_LOGIC;
  SIGNAL or_1960_nl : STD_LOGIC;
  SIGNAL or_1958_nl : STD_LOGIC;
  SIGNAL mux_1958_nl : STD_LOGIC;
  SIGNAL mux_1957_nl : STD_LOGIC;
  SIGNAL mux_1956_nl : STD_LOGIC;
  SIGNAL mux_1955_nl : STD_LOGIC;
  SIGNAL or_2065_nl : STD_LOGIC;
  SIGNAL mux_1954_nl : STD_LOGIC;
  SIGNAL or_2063_nl : STD_LOGIC;
  SIGNAL mux_1953_nl : STD_LOGIC;
  SIGNAL or_2062_nl : STD_LOGIC;
  SIGNAL or_2061_nl : STD_LOGIC;
  SIGNAL mux_1952_nl : STD_LOGIC;
  SIGNAL mux_1951_nl : STD_LOGIC;
  SIGNAL mux_1950_nl : STD_LOGIC;
  SIGNAL or_2060_nl : STD_LOGIC;
  SIGNAL or_2058_nl : STD_LOGIC;
  SIGNAL or_2056_nl : STD_LOGIC;
  SIGNAL or_2054_nl : STD_LOGIC;
  SIGNAL mux_1949_nl : STD_LOGIC;
  SIGNAL mux_1948_nl : STD_LOGIC;
  SIGNAL mux_1947_nl : STD_LOGIC;
  SIGNAL mux_1946_nl : STD_LOGIC;
  SIGNAL or_2053_nl : STD_LOGIC;
  SIGNAL or_2052_nl : STD_LOGIC;
  SIGNAL or_2051_nl : STD_LOGIC;
  SIGNAL or_2050_nl : STD_LOGIC;
  SIGNAL mux_1945_nl : STD_LOGIC;
  SIGNAL mux_1944_nl : STD_LOGIC;
  SIGNAL nand_271_nl : STD_LOGIC;
  SIGNAL mux_1943_nl : STD_LOGIC;
  SIGNAL or_2047_nl : STD_LOGIC;
  SIGNAL or_2046_nl : STD_LOGIC;
  SIGNAL or_2045_nl : STD_LOGIC;
  SIGNAL mux_1942_nl : STD_LOGIC;
  SIGNAL mux_1941_nl : STD_LOGIC;
  SIGNAL mux_1940_nl : STD_LOGIC;
  SIGNAL mux_1939_nl : STD_LOGIC;
  SIGNAL mux_1938_nl : STD_LOGIC;
  SIGNAL or_2044_nl : STD_LOGIC;
  SIGNAL or_2042_nl : STD_LOGIC;
  SIGNAL or_2040_nl : STD_LOGIC;
  SIGNAL nand_92_nl : STD_LOGIC;
  SIGNAL mux_1937_nl : STD_LOGIC;
  SIGNAL mux_1936_nl : STD_LOGIC;
  SIGNAL mux_1935_nl : STD_LOGIC;
  SIGNAL or_2038_nl : STD_LOGIC;
  SIGNAL or_2037_nl : STD_LOGIC;
  SIGNAL or_2035_nl : STD_LOGIC;
  SIGNAL or_2034_nl : STD_LOGIC;
  SIGNAL mux_1934_nl : STD_LOGIC;
  SIGNAL mux_1933_nl : STD_LOGIC;
  SIGNAL or_2032_nl : STD_LOGIC;
  SIGNAL or_2030_nl : STD_LOGIC;
  SIGNAL mux_1932_nl : STD_LOGIC;
  SIGNAL or_2029_nl : STD_LOGIC;
  SIGNAL mux_1931_nl : STD_LOGIC;
  SIGNAL or_2027_nl : STD_LOGIC;
  SIGNAL mux_1930_nl : STD_LOGIC;
  SIGNAL mux_1929_nl : STD_LOGIC;
  SIGNAL or_2020_nl : STD_LOGIC;
  SIGNAL or_2019_nl : STD_LOGIC;
  SIGNAL or_2017_nl : STD_LOGIC;
  SIGNAL or_2016_nl : STD_LOGIC;
  SIGNAL mux_1926_nl : STD_LOGIC;
  SIGNAL or_2015_nl : STD_LOGIC;
  SIGNAL mux_1925_nl : STD_LOGIC;
  SIGNAL or_2014_nl : STD_LOGIC;
  SIGNAL mux_1924_nl : STD_LOGIC;
  SIGNAL or_2013_nl : STD_LOGIC;
  SIGNAL or_2012_nl : STD_LOGIC;
  SIGNAL mux_1991_nl : STD_LOGIC;
  SIGNAL mux_1990_nl : STD_LOGIC;
  SIGNAL mux_1989_nl : STD_LOGIC;
  SIGNAL nand_96_nl : STD_LOGIC;
  SIGNAL mux_1988_nl : STD_LOGIC;
  SIGNAL mux_1987_nl : STD_LOGIC;
  SIGNAL nor_609_nl : STD_LOGIC;
  SIGNAL nor_610_nl : STD_LOGIC;
  SIGNAL mux_1986_nl : STD_LOGIC;
  SIGNAL and_771_nl : STD_LOGIC;
  SIGNAL and_777_nl : STD_LOGIC;
  SIGNAL mux_1985_nl : STD_LOGIC;
  SIGNAL nand_95_nl : STD_LOGIC;
  SIGNAL mux_1984_nl : STD_LOGIC;
  SIGNAL nor_613_nl : STD_LOGIC;
  SIGNAL nor_614_nl : STD_LOGIC;
  SIGNAL mux_1983_nl : STD_LOGIC;
  SIGNAL mux_1982_nl : STD_LOGIC;
  SIGNAL or_2110_nl : STD_LOGIC;
  SIGNAL or_2108_nl : STD_LOGIC;
  SIGNAL or_2107_nl : STD_LOGIC;
  SIGNAL mux_1981_nl : STD_LOGIC;
  SIGNAL or_2106_nl : STD_LOGIC;
  SIGNAL mux_1980_nl : STD_LOGIC;
  SIGNAL mux_1979_nl : STD_LOGIC;
  SIGNAL nand_262_nl : STD_LOGIC;
  SIGNAL nand_470_nl : STD_LOGIC;
  SIGNAL mux_1978_nl : STD_LOGIC;
  SIGNAL or_2102_nl : STD_LOGIC;
  SIGNAL or_2100_nl : STD_LOGIC;
  SIGNAL mux_1977_nl : STD_LOGIC;
  SIGNAL or_2098_nl : STD_LOGIC;
  SIGNAL mux_1976_nl : STD_LOGIC;
  SIGNAL or_2097_nl : STD_LOGIC;
  SIGNAL or_2096_nl : STD_LOGIC;
  SIGNAL or_2095_nl : STD_LOGIC;
  SIGNAL mux_1975_nl : STD_LOGIC;
  SIGNAL mux_1974_nl : STD_LOGIC;
  SIGNAL mux_1973_nl : STD_LOGIC;
  SIGNAL mux_1972_nl : STD_LOGIC;
  SIGNAL or_2093_nl : STD_LOGIC;
  SIGNAL mux_1971_nl : STD_LOGIC;
  SIGNAL mux_1970_nl : STD_LOGIC;
  SIGNAL or_2090_nl : STD_LOGIC;
  SIGNAL nand_93_nl : STD_LOGIC;
  SIGNAL mux_1968_nl : STD_LOGIC;
  SIGNAL mux_1967_nl : STD_LOGIC;
  SIGNAL nor_615_nl : STD_LOGIC;
  SIGNAL nor_616_nl : STD_LOGIC;
  SIGNAL mux_1966_nl : STD_LOGIC;
  SIGNAL and_785_nl : STD_LOGIC;
  SIGNAL and_786_nl : STD_LOGIC;
  SIGNAL mux_1965_nl : STD_LOGIC;
  SIGNAL mux_1964_nl : STD_LOGIC;
  SIGNAL mux_1963_nl : STD_LOGIC;
  SIGNAL or_2079_nl : STD_LOGIC;
  SIGNAL mux_1962_nl : STD_LOGIC;
  SIGNAL or_2077_nl : STD_LOGIC;
  SIGNAL or_2075_nl : STD_LOGIC;
  SIGNAL or_2074_nl : STD_LOGIC;
  SIGNAL mux_1961_nl : STD_LOGIC;
  SIGNAL or_2073_nl : STD_LOGIC;
  SIGNAL or_2072_nl : STD_LOGIC;
  SIGNAL or_2071_nl : STD_LOGIC;
  SIGNAL mux_1960_nl : STD_LOGIC;
  SIGNAL mux_1959_nl : STD_LOGIC;
  SIGNAL nand_267_nl : STD_LOGIC;
  SIGNAL nand_451_nl : STD_LOGIC;
  SIGNAL or_2067_nl : STD_LOGIC;
  SIGNAL mux_2026_nl : STD_LOGIC;
  SIGNAL mux_2025_nl : STD_LOGIC;
  SIGNAL mux_2024_nl : STD_LOGIC;
  SIGNAL mux_2023_nl : STD_LOGIC;
  SIGNAL or_2171_nl : STD_LOGIC;
  SIGNAL mux_2022_nl : STD_LOGIC;
  SIGNAL nand_248_nl : STD_LOGIC;
  SIGNAL mux_2021_nl : STD_LOGIC;
  SIGNAL or_2168_nl : STD_LOGIC;
  SIGNAL or_2167_nl : STD_LOGIC;
  SIGNAL mux_2020_nl : STD_LOGIC;
  SIGNAL mux_2019_nl : STD_LOGIC;
  SIGNAL mux_2018_nl : STD_LOGIC;
  SIGNAL or_2166_nl : STD_LOGIC;
  SIGNAL or_2164_nl : STD_LOGIC;
  SIGNAL or_2162_nl : STD_LOGIC;
  SIGNAL or_2160_nl : STD_LOGIC;
  SIGNAL mux_2017_nl : STD_LOGIC;
  SIGNAL mux_2016_nl : STD_LOGIC;
  SIGNAL mux_2015_nl : STD_LOGIC;
  SIGNAL mux_2014_nl : STD_LOGIC;
  SIGNAL nand_249_nl : STD_LOGIC;
  SIGNAL nand_250_nl : STD_LOGIC;
  SIGNAL or_2157_nl : STD_LOGIC;
  SIGNAL or_2156_nl : STD_LOGIC;
  SIGNAL mux_2013_nl : STD_LOGIC;
  SIGNAL mux_2012_nl : STD_LOGIC;
  SIGNAL nand_251_nl : STD_LOGIC;
  SIGNAL mux_2011_nl : STD_LOGIC;
  SIGNAL or_2153_nl : STD_LOGIC;
  SIGNAL or_2152_nl : STD_LOGIC;
  SIGNAL or_2151_nl : STD_LOGIC;
  SIGNAL mux_2010_nl : STD_LOGIC;
  SIGNAL mux_2009_nl : STD_LOGIC;
  SIGNAL mux_2008_nl : STD_LOGIC;
  SIGNAL mux_2007_nl : STD_LOGIC;
  SIGNAL mux_2006_nl : STD_LOGIC;
  SIGNAL or_2150_nl : STD_LOGIC;
  SIGNAL or_2148_nl : STD_LOGIC;
  SIGNAL or_2146_nl : STD_LOGIC;
  SIGNAL nand_98_nl : STD_LOGIC;
  SIGNAL mux_2005_nl : STD_LOGIC;
  SIGNAL mux_2004_nl : STD_LOGIC;
  SIGNAL nand_465_nl : STD_LOGIC;
  SIGNAL mux_2003_nl : STD_LOGIC;
  SIGNAL nand_254_nl : STD_LOGIC;
  SIGNAL and_540_nl : STD_LOGIC;
  SIGNAL nand_461_nl : STD_LOGIC;
  SIGNAL mux_2002_nl : STD_LOGIC;
  SIGNAL mux_2001_nl : STD_LOGIC;
  SIGNAL or_2139_nl : STD_LOGIC;
  SIGNAL or_2137_nl : STD_LOGIC;
  SIGNAL mux_2000_nl : STD_LOGIC;
  SIGNAL or_2136_nl : STD_LOGIC;
  SIGNAL mux_1999_nl : STD_LOGIC;
  SIGNAL or_2134_nl : STD_LOGIC;
  SIGNAL mux_1998_nl : STD_LOGIC;
  SIGNAL or_2132_nl : STD_LOGIC;
  SIGNAL mux_1997_nl : STD_LOGIC;
  SIGNAL and_541_nl : STD_LOGIC;
  SIGNAL and_542_nl : STD_LOGIC;
  SIGNAL or_2125_nl : STD_LOGIC;
  SIGNAL mux_1994_nl : STD_LOGIC;
  SIGNAL or_2124_nl : STD_LOGIC;
  SIGNAL mux_1993_nl : STD_LOGIC;
  SIGNAL or_2123_nl : STD_LOGIC;
  SIGNAL mux_1992_nl : STD_LOGIC;
  SIGNAL or_2122_nl : STD_LOGIC;
  SIGNAL or_2121_nl : STD_LOGIC;
  SIGNAL mux_2059_nl : STD_LOGIC;
  SIGNAL mux_2058_nl : STD_LOGIC;
  SIGNAL mux_2057_nl : STD_LOGIC;
  SIGNAL nand_102_nl : STD_LOGIC;
  SIGNAL mux_2056_nl : STD_LOGIC;
  SIGNAL mux_2055_nl : STD_LOGIC;
  SIGNAL nor_597_nl : STD_LOGIC;
  SIGNAL nor_598_nl : STD_LOGIC;
  SIGNAL mux_2054_nl : STD_LOGIC;
  SIGNAL and_770_nl : STD_LOGIC;
  SIGNAL and_776_nl : STD_LOGIC;
  SIGNAL mux_2053_nl : STD_LOGIC;
  SIGNAL nand_101_nl : STD_LOGIC;
  SIGNAL mux_2052_nl : STD_LOGIC;
  SIGNAL nor_601_nl : STD_LOGIC;
  SIGNAL nor_602_nl : STD_LOGIC;
  SIGNAL mux_2051_nl : STD_LOGIC;
  SIGNAL mux_2050_nl : STD_LOGIC;
  SIGNAL or_2216_nl : STD_LOGIC;
  SIGNAL or_2214_nl : STD_LOGIC;
  SIGNAL or_2213_nl : STD_LOGIC;
  SIGNAL mux_2049_nl : STD_LOGIC;
  SIGNAL or_2212_nl : STD_LOGIC;
  SIGNAL mux_2048_nl : STD_LOGIC;
  SIGNAL mux_2047_nl : STD_LOGIC;
  SIGNAL nand_239_nl : STD_LOGIC;
  SIGNAL nand_469_nl : STD_LOGIC;
  SIGNAL mux_2046_nl : STD_LOGIC;
  SIGNAL or_2208_nl : STD_LOGIC;
  SIGNAL or_2206_nl : STD_LOGIC;
  SIGNAL mux_2045_nl : STD_LOGIC;
  SIGNAL or_2204_nl : STD_LOGIC;
  SIGNAL mux_2044_nl : STD_LOGIC;
  SIGNAL or_2203_nl : STD_LOGIC;
  SIGNAL or_2202_nl : STD_LOGIC;
  SIGNAL or_2201_nl : STD_LOGIC;
  SIGNAL mux_2043_nl : STD_LOGIC;
  SIGNAL mux_2042_nl : STD_LOGIC;
  SIGNAL mux_2041_nl : STD_LOGIC;
  SIGNAL mux_2040_nl : STD_LOGIC;
  SIGNAL or_2199_nl : STD_LOGIC;
  SIGNAL mux_2039_nl : STD_LOGIC;
  SIGNAL mux_2038_nl : STD_LOGIC;
  SIGNAL or_2196_nl : STD_LOGIC;
  SIGNAL nand_99_nl : STD_LOGIC;
  SIGNAL mux_2036_nl : STD_LOGIC;
  SIGNAL mux_2035_nl : STD_LOGIC;
  SIGNAL nor_603_nl : STD_LOGIC;
  SIGNAL nor_604_nl : STD_LOGIC;
  SIGNAL mux_2034_nl : STD_LOGIC;
  SIGNAL and_783_nl : STD_LOGIC;
  SIGNAL and_784_nl : STD_LOGIC;
  SIGNAL mux_2033_nl : STD_LOGIC;
  SIGNAL mux_2032_nl : STD_LOGIC;
  SIGNAL mux_2031_nl : STD_LOGIC;
  SIGNAL or_2185_nl : STD_LOGIC;
  SIGNAL mux_2030_nl : STD_LOGIC;
  SIGNAL or_2183_nl : STD_LOGIC;
  SIGNAL or_2181_nl : STD_LOGIC;
  SIGNAL or_2180_nl : STD_LOGIC;
  SIGNAL mux_2029_nl : STD_LOGIC;
  SIGNAL or_2179_nl : STD_LOGIC;
  SIGNAL or_2178_nl : STD_LOGIC;
  SIGNAL or_2177_nl : STD_LOGIC;
  SIGNAL mux_2028_nl : STD_LOGIC;
  SIGNAL mux_2027_nl : STD_LOGIC;
  SIGNAL nand_244_nl : STD_LOGIC;
  SIGNAL nand_450_nl : STD_LOGIC;
  SIGNAL or_2173_nl : STD_LOGIC;
  SIGNAL mux_2094_nl : STD_LOGIC;
  SIGNAL mux_2093_nl : STD_LOGIC;
  SIGNAL mux_2092_nl : STD_LOGIC;
  SIGNAL mux_2091_nl : STD_LOGIC;
  SIGNAL or_2280_nl : STD_LOGIC;
  SIGNAL mux_2090_nl : STD_LOGIC;
  SIGNAL nand_222_nl : STD_LOGIC;
  SIGNAL mux_2089_nl : STD_LOGIC;
  SIGNAL or_2277_nl : STD_LOGIC;
  SIGNAL or_2276_nl : STD_LOGIC;
  SIGNAL mux_2088_nl : STD_LOGIC;
  SIGNAL mux_2087_nl : STD_LOGIC;
  SIGNAL mux_2086_nl : STD_LOGIC;
  SIGNAL or_2275_nl : STD_LOGIC;
  SIGNAL or_2273_nl : STD_LOGIC;
  SIGNAL or_2271_nl : STD_LOGIC;
  SIGNAL or_2269_nl : STD_LOGIC;
  SIGNAL mux_2085_nl : STD_LOGIC;
  SIGNAL mux_2084_nl : STD_LOGIC;
  SIGNAL mux_2083_nl : STD_LOGIC;
  SIGNAL mux_2082_nl : STD_LOGIC;
  SIGNAL nand_223_nl : STD_LOGIC;
  SIGNAL nand_224_nl : STD_LOGIC;
  SIGNAL or_2266_nl : STD_LOGIC;
  SIGNAL or_2265_nl : STD_LOGIC;
  SIGNAL mux_2081_nl : STD_LOGIC;
  SIGNAL mux_2080_nl : STD_LOGIC;
  SIGNAL nand_225_nl : STD_LOGIC;
  SIGNAL mux_2079_nl : STD_LOGIC;
  SIGNAL or_2262_nl : STD_LOGIC;
  SIGNAL or_2261_nl : STD_LOGIC;
  SIGNAL or_2260_nl : STD_LOGIC;
  SIGNAL mux_2078_nl : STD_LOGIC;
  SIGNAL mux_2077_nl : STD_LOGIC;
  SIGNAL mux_2076_nl : STD_LOGIC;
  SIGNAL mux_2075_nl : STD_LOGIC;
  SIGNAL mux_2074_nl : STD_LOGIC;
  SIGNAL or_2259_nl : STD_LOGIC;
  SIGNAL or_2257_nl : STD_LOGIC;
  SIGNAL or_2255_nl : STD_LOGIC;
  SIGNAL nand_104_nl : STD_LOGIC;
  SIGNAL mux_2073_nl : STD_LOGIC;
  SIGNAL mux_2072_nl : STD_LOGIC;
  SIGNAL mux_2071_nl : STD_LOGIC;
  SIGNAL nand_227_nl : STD_LOGIC;
  SIGNAL nand_464_nl : STD_LOGIC;
  SIGNAL nand_229_nl : STD_LOGIC;
  SIGNAL nand_460_nl : STD_LOGIC;
  SIGNAL mux_2070_nl : STD_LOGIC;
  SIGNAL mux_2069_nl : STD_LOGIC;
  SIGNAL or_2247_nl : STD_LOGIC;
  SIGNAL or_2245_nl : STD_LOGIC;
  SIGNAL mux_2068_nl : STD_LOGIC;
  SIGNAL or_2244_nl : STD_LOGIC;
  SIGNAL mux_2067_nl : STD_LOGIC;
  SIGNAL or_2242_nl : STD_LOGIC;
  SIGNAL mux_2066_nl : STD_LOGIC;
  SIGNAL mux_2065_nl : STD_LOGIC;
  SIGNAL nand_233_nl : STD_LOGIC;
  SIGNAL or_2234_nl : STD_LOGIC;
  SIGNAL nand_234_nl : STD_LOGIC;
  SIGNAL or_2231_nl : STD_LOGIC;
  SIGNAL mux_2062_nl : STD_LOGIC;
  SIGNAL or_2230_nl : STD_LOGIC;
  SIGNAL mux_2061_nl : STD_LOGIC;
  SIGNAL or_2229_nl : STD_LOGIC;
  SIGNAL mux_2060_nl : STD_LOGIC;
  SIGNAL or_2228_nl : STD_LOGIC;
  SIGNAL or_2227_nl : STD_LOGIC;
  SIGNAL mux_2127_nl : STD_LOGIC;
  SIGNAL mux_2126_nl : STD_LOGIC;
  SIGNAL mux_2125_nl : STD_LOGIC;
  SIGNAL nand_108_nl : STD_LOGIC;
  SIGNAL mux_2124_nl : STD_LOGIC;
  SIGNAL mux_2123_nl : STD_LOGIC;
  SIGNAL and_536_nl : STD_LOGIC;
  SIGNAL and_537_nl : STD_LOGIC;
  SIGNAL mux_2122_nl : STD_LOGIC;
  SIGNAL and_769_nl : STD_LOGIC;
  SIGNAL and_775_nl : STD_LOGIC;
  SIGNAL mux_2121_nl : STD_LOGIC;
  SIGNAL nand_107_nl : STD_LOGIC;
  SIGNAL mux_2120_nl : STD_LOGIC;
  SIGNAL nor_591_nl : STD_LOGIC;
  SIGNAL nor_592_nl : STD_LOGIC;
  SIGNAL mux_2119_nl : STD_LOGIC;
  SIGNAL mux_2118_nl : STD_LOGIC;
  SIGNAL or_2325_nl : STD_LOGIC;
  SIGNAL or_2323_nl : STD_LOGIC;
  SIGNAL or_2322_nl : STD_LOGIC;
  SIGNAL mux_2117_nl : STD_LOGIC;
  SIGNAL or_2321_nl : STD_LOGIC;
  SIGNAL mux_2116_nl : STD_LOGIC;
  SIGNAL mux_2115_nl : STD_LOGIC;
  SIGNAL nand_208_nl : STD_LOGIC;
  SIGNAL nand_468_nl : STD_LOGIC;
  SIGNAL mux_2114_nl : STD_LOGIC;
  SIGNAL or_2317_nl : STD_LOGIC;
  SIGNAL or_2315_nl : STD_LOGIC;
  SIGNAL mux_2113_nl : STD_LOGIC;
  SIGNAL or_2313_nl : STD_LOGIC;
  SIGNAL mux_2112_nl : STD_LOGIC;
  SIGNAL or_2312_nl : STD_LOGIC;
  SIGNAL or_2311_nl : STD_LOGIC;
  SIGNAL or_2310_nl : STD_LOGIC;
  SIGNAL mux_2111_nl : STD_LOGIC;
  SIGNAL mux_2110_nl : STD_LOGIC;
  SIGNAL mux_2109_nl : STD_LOGIC;
  SIGNAL mux_2108_nl : STD_LOGIC;
  SIGNAL or_2308_nl : STD_LOGIC;
  SIGNAL mux_2107_nl : STD_LOGIC;
  SIGNAL mux_2106_nl : STD_LOGIC;
  SIGNAL or_2305_nl : STD_LOGIC;
  SIGNAL nand_105_nl : STD_LOGIC;
  SIGNAL mux_2104_nl : STD_LOGIC;
  SIGNAL mux_2103_nl : STD_LOGIC;
  SIGNAL and_538_nl : STD_LOGIC;
  SIGNAL and_539_nl : STD_LOGIC;
  SIGNAL mux_2102_nl : STD_LOGIC;
  SIGNAL and_781_nl : STD_LOGIC;
  SIGNAL and_782_nl : STD_LOGIC;
  SIGNAL mux_2101_nl : STD_LOGIC;
  SIGNAL mux_2100_nl : STD_LOGIC;
  SIGNAL mux_2099_nl : STD_LOGIC;
  SIGNAL or_2294_nl : STD_LOGIC;
  SIGNAL mux_2098_nl : STD_LOGIC;
  SIGNAL or_2292_nl : STD_LOGIC;
  SIGNAL nand_215_nl : STD_LOGIC;
  SIGNAL or_2289_nl : STD_LOGIC;
  SIGNAL mux_2097_nl : STD_LOGIC;
  SIGNAL or_2288_nl : STD_LOGIC;
  SIGNAL or_2287_nl : STD_LOGIC;
  SIGNAL or_2286_nl : STD_LOGIC;
  SIGNAL mux_2096_nl : STD_LOGIC;
  SIGNAL mux_2095_nl : STD_LOGIC;
  SIGNAL nand_216_nl : STD_LOGIC;
  SIGNAL nand_449_nl : STD_LOGIC;
  SIGNAL or_2282_nl : STD_LOGIC;
  SIGNAL mux_2159_nl : STD_LOGIC;
  SIGNAL mux_2158_nl : STD_LOGIC;
  SIGNAL mux_2157_nl : STD_LOGIC;
  SIGNAL and_530_nl : STD_LOGIC;
  SIGNAL mux_2156_nl : STD_LOGIC;
  SIGNAL and_531_nl : STD_LOGIC;
  SIGNAL mux_2155_nl : STD_LOGIC;
  SIGNAL nor_570_nl : STD_LOGIC;
  SIGNAL nor_571_nl : STD_LOGIC;
  SIGNAL and_532_nl : STD_LOGIC;
  SIGNAL nor_572_nl : STD_LOGIC;
  SIGNAL mux_2154_nl : STD_LOGIC;
  SIGNAL mux_2153_nl : STD_LOGIC;
  SIGNAL nor_573_nl : STD_LOGIC;
  SIGNAL mux_2152_nl : STD_LOGIC;
  SIGNAL mux_2151_nl : STD_LOGIC;
  SIGNAL or_2835_nl : STD_LOGIC;
  SIGNAL nand_188_nl : STD_LOGIC;
  SIGNAL or_2377_nl : STD_LOGIC;
  SIGNAL mux_2150_nl : STD_LOGIC;
  SIGNAL mux_2149_nl : STD_LOGIC;
  SIGNAL and_533_nl : STD_LOGIC;
  SIGNAL mux_2148_nl : STD_LOGIC;
  SIGNAL and_766_nl : STD_LOGIC;
  SIGNAL and_767_nl : STD_LOGIC;
  SIGNAL nor_576_nl : STD_LOGIC;
  SIGNAL nor_577_nl : STD_LOGIC;
  SIGNAL mux_2147_nl : STD_LOGIC;
  SIGNAL nand_459_nl : STD_LOGIC;
  SIGNAL mux_2146_nl : STD_LOGIC;
  SIGNAL or_2365_nl : STD_LOGIC;
  SIGNAL mux_2145_nl : STD_LOGIC;
  SIGNAL nand_190_nl : STD_LOGIC;
  SIGNAL nand_191_nl : STD_LOGIC;
  SIGNAL mux_2144_nl : STD_LOGIC;
  SIGNAL mux_2143_nl : STD_LOGIC;
  SIGNAL mux_2142_nl : STD_LOGIC;
  SIGNAL nor_578_nl : STD_LOGIC;
  SIGNAL nor_579_nl : STD_LOGIC;
  SIGNAL mux_2141_nl : STD_LOGIC;
  SIGNAL mux_2140_nl : STD_LOGIC;
  SIGNAL nand_192_nl : STD_LOGIC;
  SIGNAL nand_193_nl : STD_LOGIC;
  SIGNAL or_2357_nl : STD_LOGIC;
  SIGNAL mux_2139_nl : STD_LOGIC;
  SIGNAL mux_2138_nl : STD_LOGIC;
  SIGNAL mux_2137_nl : STD_LOGIC;
  SIGNAL mux_2136_nl : STD_LOGIC;
  SIGNAL nor_580_nl : STD_LOGIC;
  SIGNAL nor_581_nl : STD_LOGIC;
  SIGNAL and_768_nl : STD_LOGIC;
  SIGNAL and_534_nl : STD_LOGIC;
  SIGNAL mux_2135_nl : STD_LOGIC;
  SIGNAL mux_2134_nl : STD_LOGIC;
  SIGNAL mux_2133_nl : STD_LOGIC;
  SIGNAL nand_448_nl : STD_LOGIC;
  SIGNAL nand_422_nl : STD_LOGIC;
  SIGNAL nand_197_nl : STD_LOGIC;
  SIGNAL or_2347_nl : STD_LOGIC;
  SIGNAL mux_2132_nl : STD_LOGIC;
  SIGNAL nor_583_nl : STD_LOGIC;
  SIGNAL mux_2131_nl : STD_LOGIC;
  SIGNAL nor_584_nl : STD_LOGIC;
  SIGNAL mux_2130_nl : STD_LOGIC;
  SIGNAL and_774_nl : STD_LOGIC;
  SIGNAL mux_2129_nl : STD_LOGIC;
  SIGNAL and_780_nl : STD_LOGIC;
  SIGNAL mux_2128_nl : STD_LOGIC;
  SIGNAL and_535_nl : STD_LOGIC;
  SIGNAL and_791_nl : STD_LOGIC;
  SIGNAL and_792_nl : STD_LOGIC;
  SIGNAL mux_2800_nl : STD_LOGIC;
  SIGNAL or_2913_nl : STD_LOGIC;
  SIGNAL mux_2799_nl : STD_LOGIC;
  SIGNAL or_2912_nl : STD_LOGIC;
  SIGNAL nand_481_nl : STD_LOGIC;
  SIGNAL mux_nl : STD_LOGIC;
  SIGNAL or_2999_nl : STD_LOGIC;
  SIGNAL or_2918_nl : STD_LOGIC;
  SIGNAL or_2917_nl : STD_LOGIC;
  SIGNAL mux_2834_nl : STD_LOGIC;
  SIGNAL mux_2833_nl : STD_LOGIC;
  SIGNAL nand_484_nl : STD_LOGIC;
  SIGNAL mux_2832_nl : STD_LOGIC;
  SIGNAL or_2958_nl : STD_LOGIC;
  SIGNAL mux_2828_nl : STD_LOGIC;
  SIGNAL or_2953_nl : STD_LOGIC;
  SIGNAL mux_2827_nl : STD_LOGIC;
  SIGNAL mux_2826_nl : STD_LOGIC;
  SIGNAL or_2952_nl : STD_LOGIC;
  SIGNAL or_2951_nl : STD_LOGIC;
  SIGNAL mux_2825_nl : STD_LOGIC;
  SIGNAL or_2950_nl : STD_LOGIC;
  SIGNAL or_2949_nl : STD_LOGIC;
  SIGNAL mux_2824_nl : STD_LOGIC;
  SIGNAL nand_479_nl : STD_LOGIC;
  SIGNAL mux_2823_nl : STD_LOGIC;
  SIGNAL mux_2822_nl : STD_LOGIC;
  SIGNAL or_2944_nl : STD_LOGIC;
  SIGNAL or_2943_nl : STD_LOGIC;
  SIGNAL or_2942_nl : STD_LOGIC;
  SIGNAL mux_2862_nl : STD_LOGIC;
  SIGNAL nand_477_nl : STD_LOGIC;
  SIGNAL mux_2861_nl : STD_LOGIC;
  SIGNAL mux_2860_nl : STD_LOGIC;
  SIGNAL or_2996_nl : STD_LOGIC;
  SIGNAL mux_2856_nl : STD_LOGIC;
  SIGNAL mux_2855_nl : STD_LOGIC;
  SIGNAL mux_2854_nl : STD_LOGIC;
  SIGNAL mux_2853_nl : STD_LOGIC;
  SIGNAL nand_476_nl : STD_LOGIC;
  SIGNAL or_2989_nl : STD_LOGIC;
  SIGNAL or_2987_nl : STD_LOGIC;
  SIGNAL or_2986_nl : STD_LOGIC;
  SIGNAL mux_2851_nl : STD_LOGIC;
  SIGNAL or_2984_nl : STD_LOGIC;
  SIGNAL nand_475_nl : STD_LOGIC;
  SIGNAL mux_2850_nl : STD_LOGIC;
  SIGNAL nor_1007_nl : STD_LOGIC;
  SIGNAL nor_1008_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux_291_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_mux1h_842_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mux_2897_nl : STD_LOGIC;
  SIGNAL mux_2898_nl : STD_LOGIC;
  SIGNAL mux_2899_nl : STD_LOGIC;
  SIGNAL or_3024_nl : STD_LOGIC;
  SIGNAL mux_2900_nl : STD_LOGIC;
  SIGNAL or_3025_nl : STD_LOGIC;
  SIGNAL mux_2901_nl : STD_LOGIC;
  SIGNAL nand_491_nl : STD_LOGIC;
  SIGNAL mux_2902_nl : STD_LOGIC;
  SIGNAL or_3026_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux_292_nl : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_mux_293_nl : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL acc_1_nl : STD_LOGIC_VECTOR (65 DOWNTO 0);
  SIGNAL operator_64_false_operator_64_false_or_58_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_130_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_58_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_131_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_59_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_132_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_60_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_133_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_61_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_134_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_62_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_135_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_63_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_136_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_64_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_137_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_65_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_138_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_66_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_139_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_67_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_140_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_68_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_141_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_69_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_142_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_70_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_143_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_71_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_144_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_72_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_145_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_73_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_146_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_74_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_147_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_75_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_148_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_76_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_149_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_77_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_150_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_78_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_151_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_79_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_152_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_80_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_153_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_81_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_154_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_82_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_155_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_83_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_156_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_84_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_157_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_85_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_158_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_86_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_159_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_87_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_160_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_88_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_161_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_89_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_162_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_90_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_163_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_91_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_164_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_92_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_165_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_93_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_166_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_94_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_167_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_95_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_168_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_96_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_169_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_97_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_170_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_98_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_171_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_99_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_172_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_100_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_173_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_101_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_174_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_102_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_175_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_103_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_176_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_104_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_177_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_105_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_178_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_106_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_179_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_107_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_180_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_108_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_181_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_109_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_182_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_110_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_183_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_111_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_184_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_112_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_185_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL operator_64_false_operator_64_false_nor_111_nl : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL operator_64_false_mux1h_62_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL operator_64_false_or_186_nl : STD_LOGIC;
  SIGNAL operator_64_false_mux1h_63_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL operator_64_false_or_187_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_188_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_or_59_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_189_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL operator_64_false_and_65_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL operator_64_false_operator_64_false_mux_113_nl : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL operator_64_false_nor_121_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_190_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL operator_64_false_and_66_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL operator_64_false_mux1h_64_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL operator_64_false_or_191_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_192_nl : STD_LOGIC;
  SIGNAL operator_64_false_nor_122_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_193_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_114_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_194_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_115_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_or_60_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_or_61_nl : STD_LOGIC;
  SIGNAL acc_2_nl : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_64_false_mux1h_3_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL operator_64_false_or_7_nl : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_nand_1_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_9_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL operator_64_false_mux1h_4_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL operator_64_false_or_10_nl : STD_LOGIC;
  SIGNAL operator_64_false_or_11_nl : STD_LOGIC;
  SIGNAL acc_3_nl : STD_LOGIC_VECTOR (12 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_3_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_4_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_and_451_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL not_7303_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_41_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_42_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL COMP_LOOP_mux1h_843_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL COMP_LOOP_or_43_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_992_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL COMP_LOOP_nor_626_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_993_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL COMP_LOOP_mux_294_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL COMP_LOOP_nor_627_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_452_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL COMP_LOOP_mux1h_844_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL not_7304_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_5_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_845_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_846_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_994_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_995_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_996_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_997_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_998_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_999_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1000_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1001_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1002_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1003_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1004_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1005_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1006_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1007_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1008_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_847_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1009_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1010_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1011_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1012_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1013_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1014_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1015_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1016_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1017_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1018_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1019_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1020_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1021_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1022_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1023_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_848_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_849_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1024_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1025_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1026_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1027_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1028_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1029_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1030_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1031_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1032_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1033_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1034_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1035_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1036_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1037_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1038_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_850_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_851_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_852_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_853_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1039_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1040_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1041_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1042_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1043_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1044_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1045_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1046_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1047_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1048_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1049_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1050_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1051_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1052_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1053_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_854_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_855_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_856_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_857_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_858_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_859_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_860_nl : STD_LOGIC;
  SIGNAL p_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL p_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL r_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL r_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT modulo_dev
    PORT (
      base_rsc_dat : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      m_rsc_dat : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      return_rsc_z : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      ccs_ccore_start_rsc_dat : IN STD_LOGIC;
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_srst : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_return_rsc_z_1 : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat : STD_LOGIC;

  SIGNAL modExp_dev_while_rem_cmp_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modExp_dev_while_rem_cmp_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modExp_dev_while_rem_cmp_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL STAGE_MAIN_LOOP_div_cmp_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_MAIN_LOOP_div_cmp_b_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL STAGE_MAIN_LOOP_div_cmp_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL STAGE_MAIN_LOOP_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL STAGE_MAIN_LOOP_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL STAGE_MAIN_LOOP_lshift_rg_z : STD_LOGIC_VECTOR (9 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_core_wait_dp
    PORT(
      ensig_cgo_iro : IN STD_LOGIC;
      ensig_cgo : IN STD_LOGIC;
      COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en : OUT STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_core_wait_dp_inst_ensig_cgo_iro : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      STAGE_MAIN_LOOP_C_3_tr0 : IN STD_LOGIC;
      modExp_dev_while_C_11_tr0 : IN STD_LOGIC;
      STAGE_VEC_LOOP_C_0_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_16_tr0 : IN STD_LOGIC;
      COMP_LOOP_1_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_45_tr0 : IN STD_LOGIC;
      COMP_LOOP_2_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_90_tr0 : IN STD_LOGIC;
      COMP_LOOP_3_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_135_tr0 : IN STD_LOGIC;
      COMP_LOOP_4_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_180_tr0 : IN STD_LOGIC;
      COMP_LOOP_5_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_225_tr0 : IN STD_LOGIC;
      COMP_LOOP_6_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_270_tr0 : IN STD_LOGIC;
      COMP_LOOP_7_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_315_tr0 : IN STD_LOGIC;
      COMP_LOOP_8_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_360_tr0 : IN STD_LOGIC;
      COMP_LOOP_9_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_405_tr0 : IN STD_LOGIC;
      COMP_LOOP_10_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_450_tr0 : IN STD_LOGIC;
      COMP_LOOP_11_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_495_tr0 : IN STD_LOGIC;
      COMP_LOOP_12_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_540_tr0 : IN STD_LOGIC;
      COMP_LOOP_13_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_585_tr0 : IN STD_LOGIC;
      COMP_LOOP_14_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_630_tr0 : IN STD_LOGIC;
      COMP_LOOP_15_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_675_tr0 : IN STD_LOGIC;
      COMP_LOOP_16_modExp_dev_1_while_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_720_tr0 : IN STD_LOGIC;
      STAGE_VEC_LOOP_C_1_tr0 : IN STD_LOGIC;
      STAGE_MAIN_LOOP_C_4_tr0 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (9 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_STAGE_MAIN_LOOP_C_3_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_STAGE_VEC_LOOP_C_0_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_16_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_45_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_90_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_135_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_180_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_225_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_270_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_315_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_360_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_405_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_450_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_495_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_540_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_585_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_630_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_675_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_STAGE_VEC_LOOP_C_1_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_STAGE_MAIN_LOOP_C_4_tr0 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_s_1_16_2(input_15 : STD_LOGIC;
  input_14 : STD_LOGIC;
  input_13 : STD_LOGIC;
  input_12 : STD_LOGIC;
  input_11 : STD_LOGIC;
  input_10 : STD_LOGIC;
  input_9 : STD_LOGIC;
  input_8 : STD_LOGIC;
  input_7 : STD_LOGIC;
  input_6 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(15 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
      tmp := sel(6);
      result := result or ( input_6 and tmp);
      tmp := sel(7);
      result := result or ( input_7 and tmp);
      tmp := sel(8);
      result := result or ( input_8 and tmp);
      tmp := sel(9);
      result := result or ( input_9 and tmp);
      tmp := sel(10);
      result := result or ( input_10 and tmp);
      tmp := sel(11);
      result := result or ( input_11 and tmp);
      tmp := sel(12);
      result := result or ( input_12 and tmp);
      tmp := sel(13);
      result := result or ( input_13 and tmp);
      tmp := sel(14);
      result := result or ( input_14 and tmp);
      tmp := sel(15);
      result := result or ( input_15 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_4_2(input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_2_4_2(input_3 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_3_2(input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_4_2(input_3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_16_2(input_15 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(15 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_16_2(input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(15 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_18_2(input_17 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(17 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_3_2(input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_4_2(input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_33_2(input_32 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_31 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_30 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_29 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_28 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_27 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_26 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_25 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_24 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_23 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_22 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_21 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_20 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(32 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
      tmp := (OTHERS=>sel( 20));
      result := result or ( input_20 and tmp);
      tmp := (OTHERS=>sel( 21));
      result := result or ( input_21 and tmp);
      tmp := (OTHERS=>sel( 22));
      result := result or ( input_22 and tmp);
      tmp := (OTHERS=>sel( 23));
      result := result or ( input_23 and tmp);
      tmp := (OTHERS=>sel( 24));
      result := result or ( input_24 and tmp);
      tmp := (OTHERS=>sel( 25));
      result := result or ( input_25 and tmp);
      tmp := (OTHERS=>sel( 26));
      result := result or ( input_26 and tmp);
      tmp := (OTHERS=>sel( 27));
      result := result or ( input_27 and tmp);
      tmp := (OTHERS=>sel( 28));
      result := result or ( input_28 and tmp);
      tmp := (OTHERS=>sel( 29));
      result := result or ( input_29 and tmp);
      tmp := (OTHERS=>sel( 30));
      result := result or ( input_30 and tmp);
      tmp := (OTHERS=>sel( 31));
      result := result or ( input_31 and tmp);
      tmp := (OTHERS=>sel( 32));
      result := result or ( input_32 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_3_2(input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_7_7_2(input_6 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_10_2_2(input_0 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(9 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_2_2_2(input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_3_2_2(input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_4_2_2(input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_55_2_2(input_0 : STD_LOGIC_VECTOR(54 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(54 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(54 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_64_2_2(input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_6_2_2(input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  p_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 5,
      width => 64
      )
    PORT MAP(
      dat => p_rsci_dat,
      idat => p_rsci_idat_1
    );
  p_rsci_dat <= p_rsc_dat;
  p_rsci_idat <= p_rsci_idat_1;

  r_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 6,
      width => 64
      )
    PORT MAP(
      dat => r_rsci_dat,
      idat => r_rsci_idat_1
    );
  r_rsci_dat <= r_rsc_dat;
  r_rsci_idat <= r_rsci_idat_1;

  vec_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_15_lz
    );
  vec_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_14_lz
    );
  vec_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_13_lz
    );
  vec_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_12_lz
    );
  vec_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_11_lz
    );
  vec_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_10_lz
    );
  vec_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_9_lz
    );
  vec_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_8_lz
    );
  vec_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_7_lz
    );
  vec_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_6_lz
    );
  vec_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_5_lz
    );
  vec_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_4_lz
    );
  vec_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_3_lz
    );
  vec_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_2_lz
    );
  vec_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_1_lz
    );
  vec_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_0_lz
    );
  p_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => p_rsc_triosy_lz
    );
  r_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => r_rsc_triosy_lz
    );
  COMP_LOOP_1_modulo_dev_cmp : modulo_dev
    PORT MAP(
      base_rsc_dat => COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat,
      m_rsc_dat => COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat,
      return_rsc_z => COMP_LOOP_1_modulo_dev_cmp_return_rsc_z_1,
      ccs_ccore_start_rsc_dat => COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat,
      ccs_ccore_clk => clk,
      ccs_ccore_srst => rst,
      ccs_ccore_en => COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en
    );
  COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat <= MUX_v_64_2_2(z_out_3, COMP_LOOP_10_modExp_dev_1_while_mul_mut,
      MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2((NOT((fsm_output(4)) OR (MUX_s_1_2_2((CONV_SL_1_1(fsm_output(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR nand_445_cse), (MUX_s_1_2_2(((NOT (fsm_output(0)))
      OR (NOT (fsm_output(2))) OR (fsm_output(8)) OR (fsm_output(5))), ((fsm_output(0))
      OR (fsm_output(2)) OR nand_445_cse), fsm_output(1))), fsm_output(9))))), ((fsm_output(4))
      AND (NOT (MUX_s_1_2_2(or_tmp_2355, (NOT((fsm_output(1)) AND (fsm_output(0))
      AND (fsm_output(2)) AND (NOT (fsm_output(8))) AND (fsm_output(5)))), fsm_output(9))))),
      fsm_output(6))), (MUX_s_1_2_2(((fsm_output(4)) AND (NOT (MUX_s_1_2_2(((fsm_output(1))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(2))) OR (fsm_output(8)) OR (NOT
      (fsm_output(5)))), or_tmp_2355, fsm_output(9))))), ((fsm_output(4)) AND (NOT
      (MUX_s_1_2_2(((NOT (fsm_output(1))) OR (fsm_output(0)) OR (fsm_output(2)) OR
      (NOT (fsm_output(8))) OR (fsm_output(5))), or_tmp_2352, fsm_output(9))))),
      fsm_output(6))), fsm_output(3))), (MUX_s_1_2_2((NOT((fsm_output(6)) OR (NOT
      (fsm_output(4))) OR (MUX_s_1_2_2(or_tmp_2352, or_tmp_2348, fsm_output(9))))),
      (MUX_s_1_2_2(nor_558_cse, (NOT((fsm_output(4)) OR (MUX_s_1_2_2(or_tmp_2348,
      ((fsm_output(1)) OR (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(8))
      OR (NOT (fsm_output(5)))), fsm_output(9))))), fsm_output(6))), fsm_output(3))),
      fsm_output(7)));
  COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat <= p_sva;
  COMP_LOOP_1_modulo_dev_cmp_return_rsc_z <= COMP_LOOP_1_modulo_dev_cmp_return_rsc_z_1;
  COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat <= NOT (MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2(((fsm_output(7))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (fsm_output(8)) OR (fsm_output(5))),
      or_2573_cse, fsm_output(1))), (MUX_s_1_2_2((NOT((fsm_output(4)) AND (NOT mux_2252_cse))),
      mux_tmp_2226, fsm_output(1))), fsm_output(9))), (MUX_s_1_2_2(or_tmp_2381, ((fsm_output(1))
      OR (NOT (fsm_output(7))) OR (fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(8))
      OR (fsm_output(5))), fsm_output(9))), fsm_output(6))), (MUX_s_1_2_2(mux_tmp_2223,
      (MUX_s_1_2_2((MUX_s_1_2_2((nor_368_cse OR mux_2252_cse), mux_tmp_2216, fsm_output(1))),
      ((NOT (fsm_output(1))) OR (fsm_output(7)) OR (fsm_output(4)) OR (NOT (fsm_output(2)))
      OR (fsm_output(8)) OR (fsm_output(5))), fsm_output(9))), fsm_output(6))), fsm_output(3))),
      (MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2(mux_tmp_2226, (MUX_s_1_2_2(((NOT
      (fsm_output(4))) OR (fsm_output(2)) OR (NOT (fsm_output(8))) OR (fsm_output(5))),
      mux_tmp_2215, fsm_output(7))), fsm_output(1))), (MUX_s_1_2_2(((fsm_output(7))
      OR (NOT (fsm_output(2))) OR (fsm_output(8)) OR (fsm_output(5))), or_2573_cse,
      fsm_output(1))), fsm_output(9))), mux_tmp_2223, fsm_output(6))), (MUX_s_1_2_2(((fsm_output(9))
      OR (MUX_s_1_2_2(((fsm_output(7)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2)))
      OR (fsm_output(8)) OR (NOT (fsm_output(5)))), (nor_368_cse OR (NOT (fsm_output(2)))
      OR (fsm_output(8)) OR (NOT (fsm_output(5)))), fsm_output(1)))), (MUX_s_1_2_2(((fsm_output(1))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (NOT (fsm_output(2))) OR (fsm_output(8))
      OR (fsm_output(5))), (MUX_s_1_2_2((MUX_s_1_2_2(or_tmp_2373, ((fsm_output(2))
      OR (fsm_output(8)) OR (NOT (fsm_output(5)))), fsm_output(7))), mux_tmp_2216,
      fsm_output(1))), fsm_output(9))), fsm_output(6))), fsm_output(3))), fsm_output(0)));

  modExp_dev_while_rem_cmp : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => modExp_dev_while_rem_cmp_a_1,
      b => modExp_dev_while_rem_cmp_b,
      z => modExp_dev_while_rem_cmp_z_1
    );
  modExp_dev_while_rem_cmp_a_1 <= modExp_dev_while_rem_cmp_a;
  modExp_dev_while_rem_cmp_b <= reg_COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat_cse;
  modExp_dev_while_rem_cmp_z <= modExp_dev_while_rem_cmp_z_1;

  STAGE_MAIN_LOOP_div_cmp : work.mgc_comps.mgc_div
    GENERIC MAP(
      width_a => 64,
      width_b => 10,
      signd => 0
      )
    PORT MAP(
      a => STAGE_MAIN_LOOP_div_cmp_a_1,
      b => STAGE_MAIN_LOOP_div_cmp_b_1,
      z => STAGE_MAIN_LOOP_div_cmp_z_1
    );
  STAGE_MAIN_LOOP_div_cmp_a_1 <= STAGE_MAIN_LOOP_div_cmp_a;
  STAGE_MAIN_LOOP_div_cmp_b_1 <= STAGE_MAIN_LOOP_div_cmp_b;
  STAGE_MAIN_LOOP_div_cmp_z <= STAGE_MAIN_LOOP_div_cmp_z_1;

  STAGE_MAIN_LOOP_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_l_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 0,
      width_s => 4,
      width_z => 10
      )
    PORT MAP(
      a => STAGE_MAIN_LOOP_lshift_rg_a,
      s => STAGE_MAIN_LOOP_lshift_rg_s,
      z => STAGE_MAIN_LOOP_lshift_rg_z
    );
  STAGE_MAIN_LOOP_lshift_rg_a(0) <= '1';
  STAGE_MAIN_LOOP_lshift_rg_s <= COMP_LOOP_slc_acc_3_12_1_slc(3 DOWNTO 0);
  STAGE_MAIN_LOOP_lshift_psp_1_sva_mx0w0 <= STAGE_MAIN_LOOP_lshift_rg_z;

  inPlaceNTT_DIF_core_wait_dp_inst : inPlaceNTT_DIF_core_wait_dp
    PORT MAP(
      ensig_cgo_iro => inPlaceNTT_DIF_core_wait_dp_inst_ensig_cgo_iro,
      ensig_cgo => reg_ensig_cgo_cse,
      COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en => COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en
    );
  inPlaceNTT_DIF_core_wait_dp_inst_ensig_cgo_iro <= NOT mux_2240_itm;

  inPlaceNTT_DIF_core_core_fsm_inst : inPlaceNTT_DIF_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      fsm_output => inPlaceNTT_DIF_core_core_fsm_inst_fsm_output,
      STAGE_MAIN_LOOP_C_3_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_STAGE_MAIN_LOOP_C_3_tr0,
      modExp_dev_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      STAGE_VEC_LOOP_C_0_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_STAGE_VEC_LOOP_C_0_tr0,
      COMP_LOOP_C_16_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_16_tr0,
      COMP_LOOP_1_modExp_dev_1_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      COMP_LOOP_C_45_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_45_tr0,
      COMP_LOOP_2_modExp_dev_1_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      COMP_LOOP_C_90_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_90_tr0,
      COMP_LOOP_3_modExp_dev_1_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      COMP_LOOP_C_135_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_135_tr0,
      COMP_LOOP_4_modExp_dev_1_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      COMP_LOOP_C_180_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_180_tr0,
      COMP_LOOP_5_modExp_dev_1_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      COMP_LOOP_C_225_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_225_tr0,
      COMP_LOOP_6_modExp_dev_1_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      COMP_LOOP_C_270_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_270_tr0,
      COMP_LOOP_7_modExp_dev_1_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      COMP_LOOP_C_315_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_315_tr0,
      COMP_LOOP_8_modExp_dev_1_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      COMP_LOOP_C_360_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_360_tr0,
      COMP_LOOP_9_modExp_dev_1_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      COMP_LOOP_C_405_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_405_tr0,
      COMP_LOOP_10_modExp_dev_1_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      COMP_LOOP_C_450_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_450_tr0,
      COMP_LOOP_11_modExp_dev_1_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      COMP_LOOP_C_495_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_495_tr0,
      COMP_LOOP_12_modExp_dev_1_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      COMP_LOOP_C_540_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_540_tr0,
      COMP_LOOP_13_modExp_dev_1_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      COMP_LOOP_C_585_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_585_tr0,
      COMP_LOOP_14_modExp_dev_1_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      COMP_LOOP_C_630_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_630_tr0,
      COMP_LOOP_15_modExp_dev_1_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      COMP_LOOP_C_675_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_675_tr0,
      COMP_LOOP_16_modExp_dev_1_while_C_11_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      COMP_LOOP_C_720_tr0 => COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm,
      STAGE_VEC_LOOP_C_1_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_STAGE_VEC_LOOP_C_1_tr0,
      STAGE_MAIN_LOOP_C_4_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_STAGE_MAIN_LOOP_C_4_tr0
    );
  fsm_output <= inPlaceNTT_DIF_core_core_fsm_inst_fsm_output;
  inPlaceNTT_DIF_core_core_fsm_inst_STAGE_MAIN_LOOP_C_3_tr0 <= NOT (z_out_2(64));
  inPlaceNTT_DIF_core_core_fsm_inst_STAGE_VEC_LOOP_C_0_tr0 <= NOT (z_out_2(63));
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_16_tr0 <= NOT operator_64_false_1_slc_operator_64_false_1_acc_5_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_45_tr0 <= NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_90_tr0 <= NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_135_tr0 <= NOT operator_64_false_slc_operator_64_false_acc_1_60_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_180_tr0 <= NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_225_tr0 <= NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_270_tr0 <= NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_315_tr0 <= NOT operator_64_false_slc_operator_64_false_acc_1_60_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_360_tr0 <= NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_405_tr0 <= NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_450_tr0 <= NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_495_tr0 <= NOT operator_64_false_slc_operator_64_false_acc_1_60_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_540_tr0 <= NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_585_tr0 <= NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_630_tr0 <= NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_675_tr0 <= NOT operator_64_false_slc_operator_64_false_acc_1_60_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_STAGE_VEC_LOOP_C_1_tr0 <= z_out_1(10);
  inPlaceNTT_DIF_core_core_fsm_inst_STAGE_MAIN_LOOP_C_4_tr0 <= z_out_2(4);

  nand_437_cse <= NOT(COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      AND (fsm_output(5)) AND (fsm_output(6)) AND (NOT (fsm_output(3))) AND (fsm_output(2)));
  mux_1112_cse <= MUX_s_1_2_2(or_tmp_669, nand_tmp_19, COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_2235_nl <= MUX_s_1_2_2(mux_2232_itm, (NOT mux_tmp_2129), fsm_output(4));
  mux_2233_nl <= MUX_s_1_2_2(mux_2232_itm, (NOT mux_tmp_2114), fsm_output(4));
  mux_2231_nl <= MUX_s_1_2_2(mux_tmp_2131, mux_tmp_2118, fsm_output(4));
  mux_2234_nl <= MUX_s_1_2_2(mux_2233_nl, mux_2231_nl, fsm_output(0));
  mux_2236_nl <= MUX_s_1_2_2(mux_2235_nl, mux_2234_nl, fsm_output(1));
  mux_2227_nl <= MUX_s_1_2_2(or_2733_cse, (NOT or_tmp_2324), fsm_output(9));
  mux_2228_nl <= MUX_s_1_2_2(mux_2227_nl, (fsm_output(8)), fsm_output(4));
  mux_2226_nl <= MUX_s_1_2_2(mux_tmp_2161, nor_tmp_357, fsm_output(4));
  mux_2229_nl <= MUX_s_1_2_2(mux_2228_nl, mux_2226_nl, fsm_output(0));
  mux_2224_nl <= MUX_s_1_2_2(mux_tmp_2112, and_679_cse, fsm_output(4));
  mux_2225_nl <= MUX_s_1_2_2(mux_2224_nl, mux_tmp_2139, fsm_output(0));
  mux_2230_nl <= MUX_s_1_2_2(mux_2229_nl, mux_2225_nl, fsm_output(1));
  mux_2237_nl <= MUX_s_1_2_2(mux_2236_nl, mux_2230_nl, fsm_output(5));
  mux_2223_nl <= MUX_s_1_2_2(mux_tmp_2142, mux_tmp_2139, fsm_output(5));
  mux_2238_nl <= MUX_s_1_2_2(mux_2237_nl, mux_2223_nl, fsm_output(6));
  mux_2221_nl <= MUX_s_1_2_2((NOT mux_tmp_2135), mux_tmp_2139, fsm_output(5));
  mux_2216_nl <= MUX_s_1_2_2(or_2733_cse, (fsm_output(7)), fsm_output(9));
  mux_2217_nl <= MUX_s_1_2_2(mux_tmp_2110, mux_2216_nl, fsm_output(4));
  mux_2218_nl <= MUX_s_1_2_2(mux_tmp_2142, mux_2217_nl, fsm_output(0));
  mux_2213_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), (fsm_output(8)), fsm_output(9));
  mux_2214_nl <= MUX_s_1_2_2(mux_2213_nl, mux_tmp_2161, fsm_output(4));
  mux_2211_nl <= MUX_s_1_2_2(or_tmp_2324, mux_tmp_2112, fsm_output(4));
  mux_2215_nl <= MUX_s_1_2_2(mux_2214_nl, mux_2211_nl, fsm_output(0));
  mux_2219_nl <= MUX_s_1_2_2(mux_2218_nl, mux_2215_nl, fsm_output(1));
  or_2841_nl <= (NOT (fsm_output(4))) OR (fsm_output(9));
  mux_2208_nl <= MUX_s_1_2_2((NOT or_tmp_2322), (fsm_output(8)), or_2841_nl);
  mux_2209_nl <= MUX_s_1_2_2(mux_tmp_2124, mux_2208_nl, fsm_output(0));
  mux_2206_nl <= MUX_s_1_2_2(nor_tmp_357, mux_tmp_2110, fsm_output(4));
  mux_2207_nl <= MUX_s_1_2_2(mux_2206_nl, mux_tmp_2111, fsm_output(0));
  mux_2210_nl <= MUX_s_1_2_2(mux_2209_nl, mux_2207_nl, fsm_output(1));
  mux_2220_nl <= MUX_s_1_2_2(mux_2219_nl, mux_2210_nl, fsm_output(5));
  mux_2222_nl <= MUX_s_1_2_2(mux_2221_nl, mux_2220_nl, fsm_output(6));
  mux_2239_nl <= MUX_s_1_2_2(mux_2238_nl, mux_2222_nl, fsm_output(3));
  or_2392_nl <= nor_569_cse OR (fsm_output(8));
  mux_2200_nl <= MUX_s_1_2_2((NOT or_tmp_2322), or_2392_nl, fsm_output(4));
  mux_2198_nl <= MUX_s_1_2_2(and_679_cse, (NOT (fsm_output(7))), fsm_output(9));
  mux_2199_nl <= MUX_s_1_2_2(mux_2198_nl, or_tmp_2324, fsm_output(4));
  mux_2201_nl <= MUX_s_1_2_2(mux_2200_nl, mux_2199_nl, fsm_output(0));
  mux_2195_nl <= MUX_s_1_2_2((fsm_output(7)), mux_tmp_2112, fsm_output(9));
  mux_2196_nl <= MUX_s_1_2_2(mux_2195_nl, or_tmp_2324, fsm_output(4));
  mux_2197_nl <= MUX_s_1_2_2(mux_2196_nl, mux_tmp_2135, fsm_output(0));
  mux_2202_nl <= MUX_s_1_2_2(mux_2201_nl, mux_2197_nl, fsm_output(1));
  mux_2203_nl <= MUX_s_1_2_2((NOT mux_2202_nl), mux_tmp_2139, fsm_output(5));
  mux_2191_nl <= MUX_s_1_2_2(mux_tmp_2139, mux_tmp_2132, fsm_output(0));
  mux_2189_nl <= MUX_s_1_2_2(mux_tmp_2130, mux_tmp_2127, fsm_output(0));
  mux_2192_nl <= MUX_s_1_2_2(mux_2191_nl, mux_2189_nl, fsm_output(1));
  mux_2194_nl <= MUX_s_1_2_2(mux_tmp_2142, mux_2192_nl, fsm_output(5));
  mux_2204_nl <= MUX_s_1_2_2(mux_2203_nl, mux_2194_nl, fsm_output(6));
  mux_2184_nl <= MUX_s_1_2_2(mux_tmp_2132, mux_tmp_2130, fsm_output(0));
  mux_2179_nl <= MUX_s_1_2_2(mux_tmp_2127, mux_tmp_2124, fsm_output(0));
  mux_2185_nl <= MUX_s_1_2_2(mux_2184_nl, mux_2179_nl, fsm_output(1));
  mux_2187_nl <= MUX_s_1_2_2((NOT mux_tmp_2135), mux_2185_nl, fsm_output(5));
  mux_2170_nl <= MUX_s_1_2_2(mux_tmp_2118, mux_tmp_2113, fsm_output(4));
  mux_2167_nl <= MUX_s_1_2_2((NOT or_tmp_2324), or_tmp_2322, fsm_output(9));
  mux_2168_nl <= MUX_s_1_2_2(mux_2167_nl, mux_tmp_2113, fsm_output(4));
  mux_2171_nl <= MUX_s_1_2_2(mux_2170_nl, mux_2168_nl, fsm_output(0));
  mux_2166_nl <= MUX_s_1_2_2(mux_tmp_2114, mux_tmp_2113, fsm_output(4));
  mux_2172_nl <= MUX_s_1_2_2(mux_2171_nl, mux_2166_nl, fsm_output(1));
  mux_2173_nl <= MUX_s_1_2_2(mux_2172_nl, mux_tmp_2111, fsm_output(5));
  mux_2188_nl <= MUX_s_1_2_2(mux_2187_nl, mux_2173_nl, fsm_output(6));
  mux_2205_nl <= MUX_s_1_2_2(mux_2204_nl, mux_2188_nl, fsm_output(3));
  mux_2240_itm <= MUX_s_1_2_2(mux_2239_nl, mux_2205_nl, fsm_output(2));
  nor_558_cse <= NOT((fsm_output(4)) OR (fsm_output(9)) OR (NOT (fsm_output(1)))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(2))) OR (fsm_output(8)) OR (NOT
      (fsm_output(5))));
  nor_368_cse <= NOT((fsm_output(7)) OR (NOT (fsm_output(4))));
  and_516_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"));
  and_515_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  or_602_cse <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"));
  or_2500_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"));
  mux_1016_nl <= MUX_s_1_2_2((fsm_output(6)), or_307_cse, fsm_output(5));
  mux_1031_cse <= MUX_s_1_2_2(mux_1016_nl, or_420_cse, fsm_output(4));
  nand_169_cse <= NOT((fsm_output(2)) AND (fsm_output(5)) AND (fsm_output(8)));
  or_2573_cse <= (fsm_output(4)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(2)))
      OR (fsm_output(5)) OR (fsm_output(8));
  or_598_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"));
  nor_813_cse <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 7)/=STD_LOGIC_VECTOR'("000")));
  and_330_rgt <= and_dcpl_294 AND and_dcpl_93;
  mux_79_cse <= MUX_s_1_2_2(and_711_cse, or_165_cse, fsm_output(2));
  nand_490_cse <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)=STD_LOGIC_VECTOR'("11")));
  nor_1039_cse <= NOT((fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)));
  or_111_cse <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  or_2700_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"));
  and_711_cse <= (fsm_output(3)) AND (fsm_output(6));
  or_165_cse <= (fsm_output(3)) OR (fsm_output(6));
  and_475_cse <= (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(8));
  nor_510_cse <= NOT((fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(8)));
  and_697_cse <= (fsm_output(0)) AND (fsm_output(2));
  nand_445_cse <= NOT((fsm_output(5)) AND (fsm_output(8)));
  and_679_cse <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11"));
  and_756_cse <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111"));
  nor_936_cse <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  or_307_cse <= (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6));
  or_2733_cse <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  and_459_cse <= (fsm_output(7)) AND (fsm_output(9));
  or_420_cse <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00"));
  and_623_cse <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"));
  and_613_cse <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("11"));
  nor_497_cse <= NOT((fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(9)));
  and_581_cse <= (fsm_output(4)) AND (fsm_output(0));
  nor_832_cse <= NOT((fsm_output(4)) OR (fsm_output(0)));
  nor_1040_cse <= NOT((fsm_output(0)) OR (NOT (fsm_output(9))));
  or_3018_cse <= (NOT (fsm_output(0))) OR (fsm_output(9));
  nor_569_cse <= NOT((fsm_output(9)) OR (fsm_output(7)));
  COMP_LOOP_1_operator_64_false_acc_tmp <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "0000")), 9), 10) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 1)), 9), 10), 10));
  COMP_LOOP_acc_8_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0(9
      DOWNTO 2)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 &
      STD_LOGIC_VECTOR'( "01")), 7), 8), 8));
  COMP_LOOP_acc_cse_4_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "0011")), 9), 10), 10));
  COMP_LOOP_acc_cse_2_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "0001")), 9), 10), 10));
  operator_64_false_acc_cse_2_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "0001")), 9), 10) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 1)), 9), 10), 10));
  operator_64_false_acc_cse_3_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "0010")), 9), 10) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 1)), 9), 10), 10));
  operator_64_false_acc_cse_4_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "0011")), 9), 10) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 1)), 9), 10), 10));
  operator_64_false_acc_cse_5_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "0100")), 9), 10) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 1)), 9), 10), 10));
  operator_64_false_acc_cse_6_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "0101")), 9), 10) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 1)), 9), 10), 10));
  operator_64_false_acc_cse_7_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "0110")), 9), 10) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 1)), 9), 10), 10));
  operator_64_false_acc_cse_8_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "0111")), 9), 10) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 1)), 9), 10), 10));
  operator_64_false_acc_cse_9_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "1000")), 9), 10) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 1)), 9), 10), 10));
  operator_64_false_acc_cse_10_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "1001")), 9), 10) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 1)), 9), 10), 10));
  operator_64_false_acc_cse_11_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "1010")), 9), 10) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 1)), 9), 10), 10));
  operator_64_false_acc_cse_12_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "1011")), 9), 10) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 1)), 9), 10), 10));
  operator_64_false_acc_cse_13_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "1100")), 9), 10) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 1)), 9), 10), 10));
  operator_64_false_acc_cse_14_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "1101")), 9), 10) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 1)), 9), 10), 10));
  operator_64_false_acc_cse_15_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "1110")), 9), 10) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 1)), 9), 10), 10));
  operator_64_false_acc_cse_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "1111")), 9), 10) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 1)), 9), 10), 10));
  or_tmp <= CONV_SL_1_1(fsm_output(6 DOWNTO 2)/=STD_LOGIC_VECTOR'("00000"));
  nor_tmp_1 <= (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(6));
  nor_tmp_3 <= (fsm_output(9)) AND (fsm_output(6));
  and_dcpl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_5 <= and_711_cse AND (NOT (fsm_output(2)));
  or_tmp_33 <= (fsm_output(3)) OR (NOT (fsm_output(6)));
  or_424_nl <= (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_tmp_79 <= MUX_s_1_2_2(or_420_cse, or_424_nl, fsm_output(4));
  nand_442_cse <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11")));
  mux_156_cse <= MUX_s_1_2_2((NOT (fsm_output(6))), (fsm_output(6)), fsm_output(5));
  or_204_cse <= (fsm_output(2)) OR (fsm_output(6));
  nor_tmp_87 <= CONV_SL_1_1(fsm_output(8 DOWNTO 5)=STD_LOGIC_VECTOR'("1111"));
  mux_tmp_302 <= MUX_s_1_2_2(nor_936_cse, and_756_cse, fsm_output(5));
  or_tmp_235 <= CONV_SL_1_1(fsm_output(8 DOWNTO 5)/=STD_LOGIC_VECTOR'("0000"));
  mux_494_cse <= MUX_s_1_2_2((NOT (fsm_output(9))), (fsm_output(9)), fsm_output(7));
  nor_tmp_130 <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)=STD_LOGIC_VECTOR'("11"));
  and_tmp_11 <= (fsm_output(9)) AND or_2733_cse;
  or_444_nl <= (fsm_output(0)) OR (fsm_output(6));
  or_533_nl <= (NOT (fsm_output(0))) OR (fsm_output(6));
  mux_792_cse <= MUX_s_1_2_2(or_444_nl, or_533_nl, fsm_output(9));
  and_dcpl_44 <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_70 <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)=STD_LOGIC_VECTOR'("10"));
  or_2836_nl <= (fsm_output(2)) OR (fsm_output(5)) OR (fsm_output(7)) OR (fsm_output(8))
      OR (fsm_output(9));
  nand_389_nl <= NOT((fsm_output(2)) AND (fsm_output(5)) AND (fsm_output(7)) AND
      (fsm_output(8)) AND (fsm_output(9)));
  mux_1048_nl <= MUX_s_1_2_2(or_2836_nl, nand_389_nl, or_2500_cse);
  nand_390_nl <= NOT((fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(8)) AND
      (fsm_output(9)));
  mux_1049_nl <= MUX_s_1_2_2(mux_1048_nl, nand_390_nl, or_602_cse);
  nand_391_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 7)=STD_LOGIC_VECTOR'("111")));
  not_tmp_266 <= MUX_s_1_2_2(mux_1049_nl, nand_391_nl, fsm_output(6));
  and_dcpl_91 <= (fsm_output(4)) AND (NOT (fsm_output(0)));
  and_dcpl_92 <= and_dcpl_91 AND (NOT (fsm_output(7)));
  and_dcpl_93 <= and_dcpl_92 AND and_dcpl;
  and_dcpl_94 <= (fsm_output(1)) AND (NOT (fsm_output(5)));
  and_dcpl_95 <= NOT((fsm_output(3)) OR (fsm_output(6)));
  and_dcpl_96 <= and_dcpl_95 AND (NOT (fsm_output(2)));
  and_dcpl_97 <= and_dcpl_96 AND and_dcpl_94;
  and_dcpl_98 <= and_dcpl_97 AND and_dcpl_93;
  or_tmp_546 <= (fsm_output(5)) OR (NOT (fsm_output(1)));
  and_dcpl_105 <= nor_832_cse AND (NOT (fsm_output(7)));
  and_dcpl_106 <= and_dcpl_105 AND and_dcpl;
  and_dcpl_109 <= and_dcpl_5 AND and_dcpl_94;
  xor_dcpl <= (fsm_output(4)) XOR (fsm_output(0));
  and_dcpl_113 <= and_dcpl_5 AND xor_dcpl;
  nor_809_nl <= NOT((fsm_output(4)) OR (fsm_output(1)) OR (NOT (fsm_output(2))));
  nor_810_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(1))) OR (fsm_output(2)));
  not_tmp_280 <= MUX_s_1_2_2(nor_809_nl, nor_810_nl, fsm_output(0));
  and_dcpl_125 <= (fsm_output(2)) AND (NOT (fsm_output(1))) AND (fsm_output(7)) AND
      and_dcpl;
  and_dcpl_131 <= and_623_cse AND (fsm_output(7));
  and_dcpl_135 <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_143 <= (fsm_output(1)) AND (fsm_output(5));
  and_dcpl_146 <= (fsm_output(3)) AND (NOT (fsm_output(6)));
  and_dcpl_147 <= and_dcpl_146 AND (fsm_output(2));
  and_dcpl_158 <= (NOT (fsm_output(1))) AND (fsm_output(5));
  and_dcpl_159 <= and_dcpl_158 AND (NOT (fsm_output(4)));
  and_741_nl <= (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6));
  nor_797_nl <= NOT((fsm_output(0)) OR (fsm_output(6)) OR (fsm_output(3)));
  not_tmp_292 <= MUX_s_1_2_2(and_741_nl, nor_797_nl, fsm_output(7));
  and_dcpl_176 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_192 <= NOT((fsm_output(1)) OR (fsm_output(5)));
  and_dcpl_199 <= and_dcpl_95 AND (fsm_output(2));
  or_tmp_591 <= (fsm_output(6)) OR (NOT (fsm_output(3)));
  and_dcpl_225 <= and_dcpl_158 AND (NOT (fsm_output(7))) AND nor_tmp_130;
  not_tmp_311 <= NOT((fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(5)));
  not_tmp_312 <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("11")));
  nor_775_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_312);
  nor_776_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_312);
  mux_1085_nl <= MUX_s_1_2_2(nor_775_nl, nor_776_nl, fsm_output(4));
  nand_tmp_16 <= NOT((fsm_output(8)) AND mux_1085_nl);
  or_694_cse <= (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("000")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  or_tmp_669 <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_735_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"));
  mux_1111_nl <= MUX_s_1_2_2(nand_442_cse, or_735_nl, fsm_output(6));
  nand_tmp_19 <= NOT((fsm_output(5)) AND (NOT mux_1111_nl));
  not_tmp_322 <= NOT((fsm_output(6)) AND (fsm_output(3)) AND (fsm_output(2)));
  nor_763_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_312);
  nor_764_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_312);
  mux_1153_nl <= MUX_s_1_2_2(nor_763_nl, nor_764_nl, fsm_output(4));
  nand_tmp_22 <= NOT((fsm_output(8)) AND mux_1153_nl);
  or_803_cse <= (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("001")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  nor_751_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_312);
  nor_752_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_312);
  mux_1221_nl <= MUX_s_1_2_2(nor_751_nl, nor_752_nl, fsm_output(4));
  nand_tmp_28 <= NOT((fsm_output(8)) AND mux_1221_nl);
  or_909_cse <= (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("010")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  nor_739_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_312);
  nor_740_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_312);
  mux_1289_nl <= MUX_s_1_2_2(nor_739_nl, nor_740_nl, fsm_output(4));
  nand_tmp_34 <= NOT((fsm_output(8)) AND mux_1289_nl);
  or_1018_cse <= (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("011")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  nor_727_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_312);
  nor_728_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_312);
  mux_1357_nl <= MUX_s_1_2_2(nor_727_nl, nor_728_nl, fsm_output(4));
  nand_tmp_40 <= NOT((fsm_output(8)) AND mux_1357_nl);
  or_1124_cse <= (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("100")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  nor_715_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_312);
  nor_716_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_312);
  mux_1425_nl <= MUX_s_1_2_2(nor_715_nl, nor_716_nl, fsm_output(4));
  nand_tmp_46 <= NOT((fsm_output(8)) AND mux_1425_nl);
  or_1233_cse <= (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("101")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  nor_703_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_312);
  nor_704_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_312);
  mux_1493_nl <= MUX_s_1_2_2(nor_703_nl, nor_704_nl, fsm_output(4));
  nand_tmp_52 <= NOT((fsm_output(8)) AND mux_1493_nl);
  or_1339_cse <= (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("110")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  nor_691_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_312);
  nor_692_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_312);
  mux_1561_nl <= MUX_s_1_2_2(nor_691_nl, nor_692_nl, fsm_output(4));
  nand_tmp_58 <= NOT((fsm_output(8)) AND mux_1561_nl);
  or_1448_cse <= (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("111")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  nor_679_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_312);
  nor_680_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_312);
  mux_1629_nl <= MUX_s_1_2_2(nor_679_nl, nor_680_nl, fsm_output(4));
  nand_tmp_64 <= NOT((fsm_output(8)) AND mux_1629_nl);
  nor_667_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_312);
  nor_668_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_312);
  mux_1697_nl <= MUX_s_1_2_2(nor_667_nl, nor_668_nl, fsm_output(4));
  nand_tmp_70 <= NOT((fsm_output(8)) AND mux_1697_nl);
  nor_655_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_312);
  nor_656_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_312);
  mux_1765_nl <= MUX_s_1_2_2(nor_655_nl, nor_656_nl, fsm_output(4));
  nand_tmp_76 <= NOT((fsm_output(8)) AND mux_1765_nl);
  nor_643_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_312);
  nor_644_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_312);
  mux_1833_nl <= MUX_s_1_2_2(nor_643_nl, nor_644_nl, fsm_output(4));
  nand_tmp_82 <= NOT((fsm_output(8)) AND mux_1833_nl);
  nor_631_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_312);
  nor_632_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_312);
  mux_1901_nl <= MUX_s_1_2_2(nor_631_nl, nor_632_nl, fsm_output(4));
  nand_tmp_88 <= NOT((fsm_output(8)) AND mux_1901_nl);
  nor_619_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_312);
  nor_620_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_312);
  mux_1969_nl <= MUX_s_1_2_2(nor_619_nl, nor_620_nl, fsm_output(4));
  nand_tmp_94 <= NOT((fsm_output(8)) AND mux_1969_nl);
  nor_607_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_312);
  nor_608_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_312);
  mux_2037_nl <= MUX_s_1_2_2(nor_607_nl, nor_608_nl, fsm_output(4));
  nand_tmp_100 <= NOT((fsm_output(8)) AND mux_2037_nl);
  nor_595_nl <= NOT((NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("01")))) OR not_tmp_312);
  nor_596_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (STAGE_VEC_LOOP_j_sva_9_0(0)) AND CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("01"))))
      OR not_tmp_312);
  mux_2105_nl <= MUX_s_1_2_2(nor_595_nl, nor_596_nl, fsm_output(4));
  nand_tmp_106 <= NOT((fsm_output(8)) AND mux_2105_nl);
  or_tmp_2322 <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"));
  mux_tmp_2110 <= MUX_s_1_2_2((NOT or_tmp_2322), (fsm_output(8)), fsm_output(9));
  mux_tmp_2111 <= MUX_s_1_2_2(and_679_cse, mux_tmp_2110, fsm_output(4));
  mux_tmp_2112 <= MUX_s_1_2_2((NOT (fsm_output(8))), (fsm_output(8)), fsm_output(7));
  mux_tmp_2113 <= MUX_s_1_2_2((NOT or_2733_cse), mux_tmp_2112, fsm_output(9));
  or_tmp_2324 <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"));
  mux_tmp_2114 <= MUX_s_1_2_2((NOT or_tmp_2324), (fsm_output(7)), fsm_output(9));
  mux_tmp_2118 <= MUX_s_1_2_2((NOT (fsm_output(8))), or_tmp_2324, fsm_output(9));
  or_2390_nl <= (fsm_output(9)) OR (NOT or_tmp_2322);
  mux_2174_nl <= MUX_s_1_2_2((NOT or_tmp_2322), or_2733_cse, fsm_output(9));
  mux_tmp_2124 <= MUX_s_1_2_2(or_2390_nl, mux_2174_nl, fsm_output(4));
  mux_2177_nl <= MUX_s_1_2_2((NOT and_679_cse), mux_tmp_2112, fsm_output(9));
  mux_2176_nl <= MUX_s_1_2_2((NOT mux_tmp_2112), (fsm_output(7)), fsm_output(9));
  mux_tmp_2127 <= MUX_s_1_2_2(mux_2177_nl, mux_2176_nl, fsm_output(4));
  mux_tmp_2129 <= MUX_s_1_2_2((fsm_output(7)), or_tmp_2322, fsm_output(9));
  mux_tmp_2130 <= MUX_s_1_2_2(mux_tmp_2113, mux_tmp_2129, fsm_output(4));
  mux_tmp_2131 <= MUX_s_1_2_2(or_tmp_2322, and_679_cse, fsm_output(9));
  mux_tmp_2132 <= MUX_s_1_2_2(mux_tmp_2113, mux_tmp_2131, fsm_output(4));
  mux_tmp_2135 <= MUX_s_1_2_2(mux_tmp_2129, or_tmp_2324, fsm_output(4));
  mux_tmp_2139 <= MUX_s_1_2_2(mux_tmp_2113, and_679_cse, fsm_output(4));
  mux_tmp_2142 <= MUX_s_1_2_2(mux_tmp_2110, mux_tmp_2114, fsm_output(4));
  nor_tmp_357 <= ((fsm_output(9)) OR (fsm_output(7))) AND (fsm_output(8));
  mux_tmp_2161 <= MUX_s_1_2_2(mux_tmp_2112, or_2733_cse, fsm_output(9));
  mux_2232_itm <= MUX_s_1_2_2(mux_tmp_2112, and_679_cse, fsm_output(9));
  and_dcpl_239 <= and_dcpl_199 AND and_dcpl_192;
  and_dcpl_240 <= and_dcpl_239 AND and_dcpl_93;
  or_2412_nl <= (fsm_output(8)) OR (NOT (fsm_output(5)));
  or_2411_nl <= (NOT (fsm_output(8))) OR (fsm_output(5));
  mux_2252_cse <= MUX_s_1_2_2(or_2412_nl, or_2411_nl, fsm_output(2));
  or_tmp_2348 <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      mux_2252_cse;
  or_tmp_2352 <= (NOT (fsm_output(1))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR (NOT (fsm_output(8))) OR (fsm_output(5));
  or_tmp_2355 <= (NOT (fsm_output(1))) OR (fsm_output(0)) OR (NOT (fsm_output(2)))
      OR (fsm_output(8)) OR (NOT (fsm_output(5)));
  and_dcpl_241 <= (NOT (fsm_output(4))) AND (fsm_output(0));
  and_dcpl_242 <= and_dcpl_241 AND (NOT (fsm_output(7)));
  and_dcpl_243 <= and_dcpl_242 AND and_dcpl;
  and_dcpl_244 <= nor_tmp_1 AND and_dcpl_192;
  and_dcpl_245 <= and_dcpl_244 AND and_dcpl_243;
  and_dcpl_246 <= nor_832_cse AND (fsm_output(7));
  and_dcpl_248 <= and_dcpl_199 AND and_dcpl_94;
  and_dcpl_249 <= and_dcpl_248 AND and_dcpl_246 AND and_dcpl;
  and_dcpl_251 <= and_581_cse AND (fsm_output(7));
  and_dcpl_252 <= and_dcpl_251 AND and_dcpl;
  and_dcpl_253 <= and_dcpl_147 AND and_dcpl_143;
  and_dcpl_254 <= and_dcpl_253 AND and_dcpl_252;
  and_dcpl_255 <= and_dcpl_91 AND (fsm_output(7));
  and_dcpl_256 <= and_dcpl_255 AND and_dcpl;
  and_dcpl_257 <= and_dcpl_5 AND and_dcpl_158;
  and_dcpl_258 <= and_dcpl_257 AND and_dcpl_256;
  and_dcpl_259 <= and_581_cse AND (NOT (fsm_output(7)));
  and_dcpl_260 <= and_dcpl_259 AND and_dcpl_44;
  and_dcpl_261 <= and_dcpl_96 AND and_dcpl_158;
  and_dcpl_262 <= and_dcpl_261 AND and_dcpl_260;
  and_dcpl_263 <= and_dcpl_105 AND and_dcpl_44;
  and_dcpl_264 <= and_dcpl_5 AND and_dcpl_143;
  and_dcpl_265 <= and_dcpl_264 AND and_dcpl_263;
  and_dcpl_266 <= and_dcpl_241 AND (fsm_output(7));
  and_dcpl_267 <= and_dcpl_266 AND and_dcpl_44;
  and_dcpl_268 <= and_dcpl_96 AND and_dcpl_143;
  and_dcpl_269 <= and_dcpl_268 AND and_dcpl_267;
  and_dcpl_270 <= and_dcpl_255 AND and_dcpl_44;
  and_dcpl_271 <= and_dcpl_244 AND and_dcpl_270;
  and_dcpl_273 <= and_dcpl_239 AND and_dcpl_259 AND and_dcpl_70;
  and_dcpl_275 <= nor_tmp_1 AND and_dcpl_94;
  and_dcpl_276 <= and_dcpl_275 AND and_dcpl_105 AND and_dcpl_70;
  and_dcpl_278 <= and_dcpl_248 AND and_dcpl_266 AND and_dcpl_70;
  and_dcpl_279 <= and_dcpl_246 AND and_dcpl_70;
  and_dcpl_280 <= (NOT (fsm_output(3))) AND (fsm_output(6));
  and_dcpl_282 <= and_dcpl_280 AND (NOT (fsm_output(2))) AND and_dcpl_192;
  and_dcpl_283 <= and_dcpl_282 AND and_dcpl_279;
  and_dcpl_284 <= and_dcpl_251 AND and_dcpl_70;
  and_dcpl_285 <= and_dcpl_257 AND and_dcpl_284;
  and_dcpl_286 <= and_dcpl_92 AND nor_tmp_130;
  and_dcpl_287 <= and_dcpl_268 AND and_dcpl_286;
  and_dcpl_288 <= and_dcpl_242 AND nor_tmp_130;
  and_dcpl_289 <= and_dcpl_264 AND and_dcpl_288;
  or_tmp_2368 <= (fsm_output(2)) OR nand_445_cse;
  or_2634_nl <= (NOT (fsm_output(8))) OR (fsm_output(2)) OR (fsm_output(5));
  mux_tmp_2215 <= MUX_s_1_2_2(or_tmp_2368, or_2634_nl, fsm_output(4));
  or_2431_nl <= (NOT (fsm_output(4))) OR (fsm_output(2)) OR (fsm_output(8)) OR (fsm_output(5));
  mux_tmp_2216 <= MUX_s_1_2_2(mux_tmp_2215, or_2431_nl, fsm_output(7));
  or_tmp_2373 <= (fsm_output(4)) OR mux_2252_cse;
  or_tmp_2381 <= (NOT (fsm_output(1))) OR (fsm_output(7)) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(2))) OR (fsm_output(8)) OR (NOT (fsm_output(5)));
  nand_180_nl <= NOT((fsm_output(1)) AND (fsm_output(7)) AND (fsm_output(4)) AND
      (fsm_output(2)) AND (fsm_output(8)) AND (fsm_output(5)));
  mux_tmp_2223 <= MUX_s_1_2_2(nand_180_nl, or_tmp_2381, fsm_output(9));
  mux_tmp_2226 <= MUX_s_1_2_2(or_tmp_2368, or_tmp_2373, fsm_output(7));
  and_dcpl_290 <= and_dcpl_239 AND and_dcpl_243;
  or_tmp_2391 <= (NOT (fsm_output(2))) OR (fsm_output(8)) OR (fsm_output(7));
  or_tmp_2393 <= (fsm_output(2)) OR (fsm_output(8)) OR (NOT (fsm_output(7)));
  or_tmp_2395 <= (fsm_output(5)) OR (fsm_output(8)) OR (NOT (fsm_output(7)));
  or_2464_nl <= (NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"));
  or_2462_nl <= (CONV_SL_1_1(fsm_output(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))) OR
      CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_2244 <= MUX_s_1_2_2(or_2464_nl, or_2462_nl, fsm_output(5));
  or_tmp_2401 <= (NOT (fsm_output(2))) OR (fsm_output(8)) OR (NOT (fsm_output(7)));
  or_tmp_2402 <= (fsm_output(2)) OR (NOT (fsm_output(8))) OR (fsm_output(7));
  mux_tmp_2247 <= MUX_s_1_2_2(or_tmp_2402, or_tmp_2401, and_515_cse);
  nor_554_cse <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  or_tmp_2406 <= nor_554_cse OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"));
  mux_tmp_2250 <= MUX_s_1_2_2(or_tmp_2393, or_tmp_2391, or_2500_cse);
  not_tmp_572 <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11")));
  or_tmp_2409 <= (or_2500_cse AND (fsm_output(2))) OR not_tmp_572;
  nor_552_nl <= NOT((fsm_output(0)) OR (NOT (fsm_output(2))));
  mux_2326_cse <= MUX_s_1_2_2(nor_552_nl, and_697_cse, fsm_output(9));
  nand_176_cse <= NOT((fsm_output(3)) AND (fsm_output(6)) AND mux_2326_cse);
  or_2486_nl <= (fsm_output(5)) OR nand_176_cse;
  or_2484_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (NOT (fsm_output(0))) OR (fsm_output(2));
  mux_tmp_2276 <= MUX_s_1_2_2(or_2486_nl, or_2484_nl, fsm_output(8));
  nor_550_nl <= NOT((fsm_output(0)) OR (fsm_output(2)));
  nor_551_nl <= NOT((NOT (fsm_output(0))) OR (fsm_output(2)));
  mux_2332_cse <= MUX_s_1_2_2(nor_550_nl, nor_551_nl, fsm_output(9));
  or_2497_nl <= (NOT (fsm_output(5))) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT
      (fsm_output(9))) OR (fsm_output(0)) OR (NOT (fsm_output(2)));
  nand_120_nl <= NOT((fsm_output(6)) AND mux_2332_cse);
  or_2492_nl <= (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(0)) OR (fsm_output(2));
  mux_2333_nl <= MUX_s_1_2_2(nand_120_nl, or_2492_nl, fsm_output(3));
  or_2495_nl <= (fsm_output(5)) OR mux_2333_nl;
  mux_2334_nl <= MUX_s_1_2_2(or_2497_nl, or_2495_nl, fsm_output(8));
  or_2498_nl <= (fsm_output(7)) OR mux_2334_nl;
  or_2491_nl <= (fsm_output(8)) OR (fsm_output(5)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (NOT and_697_cse);
  mux_2331_nl <= MUX_s_1_2_2(mux_tmp_2276, or_2491_nl, fsm_output(7));
  mux_2335_nl <= MUX_s_1_2_2(or_2498_nl, mux_2331_nl, fsm_output(4));
  or_2489_nl <= (NOT (fsm_output(5))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9))
      OR (NOT (fsm_output(0))) OR (fsm_output(2));
  or_2488_nl <= (fsm_output(5)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9))
      OR (NOT and_697_cse);
  mux_2328_nl <= MUX_s_1_2_2(or_2489_nl, or_2488_nl, fsm_output(8));
  mux_2329_nl <= MUX_s_1_2_2(mux_2328_nl, mux_tmp_2276, fsm_output(7));
  nand_175_nl <= NOT((fsm_output(8)) AND (fsm_output(5)) AND (fsm_output(3)) AND
      (fsm_output(6)) AND (fsm_output(9)) AND (NOT (fsm_output(0))) AND (NOT (fsm_output(2))));
  or_2482_nl <= (fsm_output(5)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9)))
      OR (fsm_output(0)) OR (NOT (fsm_output(2)));
  or_2480_nl <= (NOT (fsm_output(5))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_2324_nl <= MUX_s_1_2_2(or_2482_nl, or_2480_nl, fsm_output(8));
  mux_2325_nl <= MUX_s_1_2_2(nand_175_nl, mux_2324_nl, fsm_output(7));
  mux_2330_nl <= MUX_s_1_2_2(mux_2329_nl, mux_2325_nl, fsm_output(4));
  mux_2336_itm <= MUX_s_1_2_2(mux_2335_nl, mux_2330_nl, fsm_output(1));
  and_dcpl_293 <= and_dcpl_97 AND (NOT (fsm_output(4))) AND (NOT (fsm_output(7)))
      AND and_dcpl;
  and_dcpl_294 <= and_dcpl_96 AND and_dcpl_192;
  and_dcpl_295 <= and_dcpl_294 AND and_dcpl_243;
  or_tmp_2439 <= and_516_cse OR (fsm_output(6)) OR (fsm_output(3));
  and_tmp_24 <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11")) AND mux_1031_cse;
  nor_tmp_388 <= (fsm_output(0)) AND (fsm_output(6));
  or_tmp_2447 <= (NOT (fsm_output(2))) OR (fsm_output(5)) OR (NOT (fsm_output(9)))
      OR (fsm_output(0)) OR (NOT (fsm_output(6)));
  or_tmp_2451 <= (NOT (fsm_output(2))) OR (fsm_output(5)) OR mux_792_cse;
  nor_541_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(8))) OR (fsm_output(2)) OR
      (fsm_output(5)) OR (NOT (fsm_output(9))) OR (fsm_output(0)) OR (NOT (fsm_output(6))));
  nor_542_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(8)) OR (NOT (fsm_output(2)))
      OR (fsm_output(5)) OR (fsm_output(9)) OR (NOT nor_tmp_388));
  mux_2357_nl <= MUX_s_1_2_2(nor_541_nl, nor_542_nl, fsm_output(7));
  nor_825_nl <= NOT((fsm_output(0)) OR (NOT (fsm_output(6))));
  mux_2354_nl <= MUX_s_1_2_2(nor_825_nl, nor_tmp_388, fsm_output(9));
  or_2521_nl <= (fsm_output(2)) OR (NOT((fsm_output(5)) AND mux_2354_nl));
  mux_2355_nl <= MUX_s_1_2_2(or_tmp_2447, or_2521_nl, fsm_output(8));
  and_506_nl <= (fsm_output(3)) AND (NOT mux_2355_nl);
  or_2518_nl <= (fsm_output(2)) OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR (NOT
      (fsm_output(0))) OR (fsm_output(6));
  mux_2353_nl <= MUX_s_1_2_2(or_tmp_2451, or_2518_nl, fsm_output(8));
  nor_544_nl <= NOT((fsm_output(3)) OR mux_2353_nl);
  mux_2356_nl <= MUX_s_1_2_2(and_506_nl, nor_544_nl, fsm_output(7));
  mux_2358_nl <= MUX_s_1_2_2(mux_2357_nl, mux_2356_nl, fsm_output(4));
  or_2831_nl <= (fsm_output(2)) OR (NOT (fsm_output(5))) OR mux_792_cse;
  mux_2350_nl <= MUX_s_1_2_2(or_2831_nl, or_tmp_2451, fsm_output(8));
  nor_545_nl <= NOT((fsm_output(3)) OR mux_2350_nl);
  or_2510_nl <= (fsm_output(2)) OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR (fsm_output(0))
      OR (NOT (fsm_output(6)));
  mux_2348_nl <= MUX_s_1_2_2(or_tmp_2447, or_2510_nl, fsm_output(8));
  and_507_nl <= (fsm_output(3)) AND (NOT mux_2348_nl);
  mux_2351_nl <= MUX_s_1_2_2(nor_545_nl, and_507_nl, fsm_output(7));
  nor_546_nl <= NOT((fsm_output(2)) OR (fsm_output(5)) OR (fsm_output(9)) OR (NOT
      nor_tmp_388));
  nor_547_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(5))) OR (fsm_output(9))
      OR (NOT (fsm_output(0))) OR (fsm_output(6)));
  mux_2347_nl <= MUX_s_1_2_2(nor_546_nl, nor_547_nl, fsm_output(8));
  and_508_nl <= (NOT((fsm_output(7)) OR (NOT (fsm_output(3))))) AND mux_2347_nl;
  mux_2352_nl <= MUX_s_1_2_2(mux_2351_nl, and_508_nl, fsm_output(4));
  not_tmp_597 <= MUX_s_1_2_2(mux_2358_nl, mux_2352_nl, fsm_output(1));
  or_2549_cse <= (NOT (fsm_output(0))) OR (fsm_output(9)) OR (fsm_output(5)) OR (NOT
      (fsm_output(8))) OR (fsm_output(2));
  or_2555_nl <= (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(8)) OR (NOT
      (fsm_output(2)));
  nand_420_nl <= NOT((fsm_output(9)) AND (fsm_output(5)) AND (NOT (fsm_output(8)))
      AND (fsm_output(2)));
  mux_2374_cse <= MUX_s_1_2_2(or_2555_nl, nand_420_nl, fsm_output(0));
  or_2612_nl <= (fsm_output(5)) OR (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(6))
      OR (fsm_output(3));
  mux_tmp_2377 <= MUX_s_1_2_2(or_420_cse, or_2612_nl, fsm_output(4));
  or_tmp_2548 <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")) OR
      or_tmp_2439;
  or_tmp_2549 <= (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(3));
  mux_tmp_2380 <= MUX_s_1_2_2(and_dcpl_96, or_tmp_2549, fsm_output(5));
  nor_tmp_399 <= or_2700_cse AND (fsm_output(6)) AND (fsm_output(3));
  mux_tmp_2381 <= MUX_s_1_2_2((NOT nor_tmp_1), nor_tmp_399, fsm_output(5));
  mux_tmp_2382 <= MUX_s_1_2_2(mux_tmp_2381, mux_tmp_2380, fsm_output(4));
  not_tmp_617 <= NOT((fsm_output(1)) AND (fsm_output(2)) AND (fsm_output(6)) AND
      (fsm_output(3)));
  mux_2439_nl <= MUX_s_1_2_2(or_tmp_2439, (NOT or_tmp_2549), fsm_output(5));
  mux_2438_nl <= MUX_s_1_2_2((NOT nor_tmp_399), and_711_cse, fsm_output(5));
  mux_tmp_2389 <= MUX_s_1_2_2(mux_2439_nl, mux_2438_nl, fsm_output(4));
  or_tmp_2551 <= (fsm_output(5)) OR and_dcpl_96;
  or_tmp_2552 <= (fsm_output(5)) OR (NOT or_tmp_2439);
  mux_tmp_2400 <= MUX_s_1_2_2(and_711_cse, or_165_cse, and_516_cse);
  nor_tmp_403 <= (and_516_cse OR (fsm_output(6))) AND (fsm_output(3));
  and_dcpl_307 <= and_dcpl_266 AND and_dcpl;
  and_dcpl_311 <= and_dcpl_280 AND (fsm_output(2)) AND and_dcpl_143;
  and_dcpl_313 <= and_dcpl_92 AND and_dcpl_44;
  and_dcpl_317 <= and_dcpl_246 AND and_dcpl_44;
  and_dcpl_319 <= and_dcpl_251 AND and_dcpl_44;
  and_dcpl_321 <= and_dcpl_92 AND and_dcpl_70;
  and_dcpl_323 <= and_dcpl_242 AND and_dcpl_70;
  and_dcpl_329 <= and_dcpl_259 AND nor_tmp_130;
  and_dcpl_331 <= and_dcpl_105 AND nor_tmp_130;
  and_dcpl_345 <= and_dcpl_248 AND and_dcpl_246 AND nor_tmp_130;
  and_dcpl_346 <= and_dcpl_259 AND and_dcpl;
  mux_tmp_2449 <= MUX_s_1_2_2((fsm_output(6)), or_tmp_2549, fsm_output(5));
  mux_tmp_2450 <= MUX_s_1_2_2(mux_tmp_2449, or_420_cse, fsm_output(4));
  or_dcpl_72 <= or_307_cse OR or_tmp_546 OR (NOT (fsm_output(4))) OR (fsm_output(0))
      OR (fsm_output(7)) OR (fsm_output(8)) OR (fsm_output(9));
  mux_tmp_2457 <= MUX_s_1_2_2(and_dcpl_95, and_711_cse, fsm_output(2));
  mux_tmp_2458 <= MUX_s_1_2_2((NOT (fsm_output(3))), (fsm_output(3)), fsm_output(6));
  mux_tmp_2459 <= MUX_s_1_2_2(and_dcpl_95, mux_tmp_2458, fsm_output(2));
  mux_2511_nl <= MUX_s_1_2_2(mux_tmp_2459, mux_tmp_2457, fsm_output(1));
  or_tmp_2585 <= (fsm_output(5)) OR mux_2511_nl;
  mux_2507_nl <= MUX_s_1_2_2(and_dcpl_96, and_711_cse, fsm_output(5));
  mux_tmp_2461 <= MUX_s_1_2_2((NOT or_tmp_2585), mux_2507_nl, fsm_output(4));
  mux_tmp_2462 <= MUX_s_1_2_2(and_dcpl_96, nor_tmp_399, fsm_output(5));
  mux_tmp_2467 <= MUX_s_1_2_2(mux_tmp_2458, and_711_cse, fsm_output(2));
  mux_tmp_2468 <= MUX_s_1_2_2(mux_tmp_2457, mux_tmp_2467, fsm_output(1));
  or_tmp_2587 <= (fsm_output(5)) OR mux_tmp_2468;
  mux_tmp_2469 <= MUX_s_1_2_2(not_tmp_617, or_tmp_2549, fsm_output(5));
  mux_tmp_2470 <= MUX_s_1_2_2(mux_tmp_2469, or_tmp_2587, fsm_output(4));
  or_tmp_2588 <= (fsm_output(5)) OR (NOT nor_tmp_1);
  mux_2524_nl <= MUX_s_1_2_2(mux_tmp_2458, and_711_cse, or_2700_cse);
  nand_137_nl <= NOT((fsm_output(5)) AND (NOT mux_2524_nl));
  mux_tmp_2474 <= MUX_s_1_2_2(nand_137_nl, or_tmp_2588, fsm_output(4));
  and_494_nl <= or_204_cse AND (fsm_output(3));
  mux_2531_nl <= MUX_s_1_2_2(mux_tmp_2467, and_494_nl, fsm_output(1));
  nand_tmp_140 <= NOT((fsm_output(5)) AND (NOT mux_2531_nl));
  nor_tmp_417 <= (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(8)) AND (fsm_output(9));
  nor_516_nl <= NOT((fsm_output(6)) OR (fsm_output(8)) OR (fsm_output(9)));
  and_489_nl <= (fsm_output(6)) AND (fsm_output(8)) AND (fsm_output(9));
  mux_tmp_2529 <= MUX_s_1_2_2(nor_516_nl, and_489_nl, fsm_output(5));
  not_tmp_662 <= NOT((fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(8)) OR (fsm_output(9)));
  mux_2583_nl <= MUX_s_1_2_2(not_tmp_662, mux_tmp_2529, or_2700_cse);
  mux_2584_nl <= MUX_s_1_2_2(not_tmp_662, mux_2583_nl, fsm_output(3));
  mux_2581_nl <= MUX_s_1_2_2(mux_tmp_2529, nor_tmp_417, and_515_cse);
  mux_2582_nl <= MUX_s_1_2_2(mux_2581_nl, nor_tmp_417, or_598_cse);
  mux_2585_nl <= MUX_s_1_2_2(mux_2584_nl, mux_2582_nl, fsm_output(4));
  mux_2586_itm <= MUX_s_1_2_2(mux_2585_nl, nor_tmp_130, fsm_output(7));
  mux_tmp_2538 <= MUX_s_1_2_2(mux_tmp_79, mux_tmp_2377, fsm_output(0));
  not_tmp_664 <= NOT((fsm_output(7)) OR mux_tmp_2538);
  mux_2607_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), or_tmp_33, and_516_cse);
  mux_2608_nl <= MUX_s_1_2_2(mux_2607_nl, (fsm_output(6)), fsm_output(5));
  or_2877_nl <= (fsm_output(2)) OR (fsm_output(5));
  mux_2606_nl <= MUX_s_1_2_2(or_tmp_591, (fsm_output(6)), or_2877_nl);
  mux_2609_nl <= MUX_s_1_2_2(mux_2608_nl, mux_2606_nl, fsm_output(4));
  mux_2603_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), or_tmp_33, fsm_output(2));
  mux_2604_nl <= MUX_s_1_2_2(mux_2603_nl, (fsm_output(6)), fsm_output(5));
  or_2604_nl <= (fsm_output(5)) OR (fsm_output(1)) OR (fsm_output(2));
  mux_2602_nl <= MUX_s_1_2_2(or_tmp_591, (fsm_output(6)), or_2604_nl);
  mux_2605_nl <= MUX_s_1_2_2(mux_2604_nl, mux_2602_nl, fsm_output(4));
  mux_2610_nl <= MUX_s_1_2_2(mux_2609_nl, mux_2605_nl, fsm_output(0));
  and_dcpl_354 <= (NOT mux_2610_nl) AND nor_813_cse;
  mux_2613_nl <= MUX_s_1_2_2(mux_tmp_2538, (NOT or_tmp_2548), fsm_output(7));
  and_dcpl_357 <= mux_2613_nl AND and_dcpl;
  and_483_nl <= (fsm_output(0)) AND (fsm_output(4)) AND (fsm_output(5)) AND (fsm_output(1))
      AND (fsm_output(2));
  mux_2617_nl <= MUX_s_1_2_2((fsm_output(6)), or_165_cse, and_483_nl);
  mux_2618_nl <= MUX_s_1_2_2(mux_tmp_2538, (NOT mux_2617_nl), fsm_output(7));
  and_dcpl_359 <= mux_2618_nl AND and_dcpl;
  nor_tmp_427 <= CONV_SL_1_1(fsm_output(6 DOWNTO 3)=STD_LOGIC_VECTOR'("1111"));
  mux_2622_nl <= MUX_s_1_2_2(mux_tmp_2538, (NOT nor_tmp_427), fsm_output(7));
  and_dcpl_361 <= mux_2622_nl AND and_dcpl;
  nor_871_nl <= NOT((fsm_output(8)) OR (fsm_output(6)));
  and_684_nl <= (fsm_output(8)) AND (fsm_output(6));
  mux_tmp_2574 <= MUX_s_1_2_2(nor_871_nl, and_684_nl, fsm_output(5));
  or_tmp_2638 <= and_623_cse OR (fsm_output(6));
  mux_tmp_2583 <= MUX_s_1_2_2((fsm_output(6)), or_tmp_2549, and_623_cse);
  mux_2635_nl <= MUX_s_1_2_2(mux_tmp_2583, or_tmp_2638, fsm_output(0));
  or_2712_nl <= (fsm_output(7)) OR mux_2635_nl;
  mux_2636_nl <= MUX_s_1_2_2(not_tmp_664, or_2712_nl, fsm_output(8));
  and_dcpl_364 <= NOT(mux_2636_nl OR (fsm_output(9)));
  or_2719_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")) OR and_515_cse
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00"));
  mux_2643_nl <= MUX_s_1_2_2(or_420_cse, or_2719_nl, fsm_output(4));
  nor_940_nl <= NOT((fsm_output(7)) OR mux_2643_nl);
  and_395_nl <= (fsm_output(3)) AND or_2700_cse AND CONV_SL_1_1(fsm_output(6 DOWNTO
      5)=STD_LOGIC_VECTOR'("11"));
  mux_2642_nl <= MUX_s_1_2_2(and_395_nl, and_613_cse, fsm_output(4));
  or_2900_nl <= (fsm_output(7)) OR mux_2642_nl;
  mux_2644_nl <= MUX_s_1_2_2(nor_940_nl, or_2900_nl, fsm_output(8));
  and_dcpl_367 <= NOT(mux_2644_nl OR (fsm_output(9)));
  mux_2650_nl <= MUX_s_1_2_2(mux_1031_cse, mux_tmp_2450, fsm_output(0));
  and_400_nl <= (fsm_output(7)) AND mux_2650_nl;
  mux_2651_nl <= MUX_s_1_2_2(not_tmp_664, and_400_nl, fsm_output(8));
  and_dcpl_370 <= NOT(mux_2651_nl OR (fsm_output(9)));
  not_tmp_696 <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 5)/=STD_LOGIC_VECTOR'("0000")));
  not_tmp_698 <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_2538);
  mux_2659_nl <= MUX_s_1_2_2(nor_tmp_1, (fsm_output(6)), fsm_output(5));
  mux_2660_nl <= MUX_s_1_2_2(and_613_cse, mux_2659_nl, fsm_output(4));
  and_403_nl <= (fsm_output(7)) AND mux_2660_nl;
  mux_2661_nl <= MUX_s_1_2_2(not_tmp_664, and_403_nl, fsm_output(8));
  and_dcpl_372 <= NOT(mux_2661_nl OR (fsm_output(9)));
  mux_tmp_2612 <= MUX_s_1_2_2((NOT (fsm_output(9))), (fsm_output(9)), fsm_output(6));
  not_tmp_703 <= NOT((fsm_output(6)) OR (fsm_output(9)));
  mux_2664_nl <= MUX_s_1_2_2(not_tmp_703, mux_tmp_2612, fsm_output(3));
  mux_tmp_2614 <= MUX_s_1_2_2(mux_2664_nl, nor_tmp_3, fsm_output(4));
  or_2740_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")) OR and_515_cse
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 5)/=STD_LOGIC_VECTOR'("0000"));
  mux_2674_nl <= MUX_s_1_2_2(or_tmp_235, or_2740_nl, fsm_output(4));
  or_2735_nl <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(7)) OR (fsm_output(8));
  mux_2672_nl <= MUX_s_1_2_2(or_tmp_235, or_2735_nl, fsm_output(2));
  or_2737_nl <= (fsm_output(3)) OR mux_2672_nl;
  mux_2673_nl <= MUX_s_1_2_2(or_tmp_235, or_2737_nl, fsm_output(4));
  not_tmp_706 <= MUX_s_1_2_2(mux_2674_nl, (NOT mux_2673_nl), fsm_output(9));
  or_tmp_2668 <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000"));
  and_tmp_32 <= (fsm_output(9)) AND or_tmp_2668;
  mux_tmp_2625 <= MUX_s_1_2_2(and_tmp_11, and_tmp_32, fsm_output(3));
  mux_tmp_2626 <= MUX_s_1_2_2((NOT or_tmp_2668), or_2733_cse, fsm_output(9));
  or_2747_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")) OR and_515_cse
      OR (fsm_output(9));
  mux_2685_nl <= MUX_s_1_2_2((fsm_output(9)), or_2747_nl, fsm_output(4));
  and_461_nl <= (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(1)) AND (fsm_output(9));
  mux_2684_nl <= MUX_s_1_2_2(and_461_nl, (fsm_output(9)), fsm_output(4));
  mux_2686_nl <= MUX_s_1_2_2((NOT mux_2685_nl), mux_2684_nl, fsm_output(6));
  mux_2687_nl <= MUX_s_1_2_2(mux_2686_nl, nor_tmp_3, fsm_output(5));
  mux_2688_itm <= MUX_s_1_2_2(mux_2687_nl, (fsm_output(9)), or_2733_cse);
  mux_2698_nl <= MUX_s_1_2_2(mux_494_cse, and_459_cse, fsm_output(2));
  mux_2699_nl <= MUX_s_1_2_2(nor_569_cse, mux_2698_nl, fsm_output(4));
  mux_2696_nl <= MUX_s_1_2_2(nor_569_cse, mux_494_cse, fsm_output(2));
  mux_2697_nl <= MUX_s_1_2_2(mux_2696_nl, and_459_cse, fsm_output(4));
  mux_2700_nl <= MUX_s_1_2_2(mux_2699_nl, mux_2697_nl, and_515_cse);
  mux_2695_nl <= MUX_s_1_2_2(mux_494_cse, and_459_cse, fsm_output(4));
  mux_2701_nl <= MUX_s_1_2_2(mux_2700_nl, mux_2695_nl, fsm_output(3));
  mux_2702_nl <= MUX_s_1_2_2(mux_2701_nl, and_459_cse, or_420_cse);
  mux_2703_itm <= MUX_s_1_2_2(mux_2702_nl, (fsm_output(9)), fsm_output(8));
  nor_tmp_459 <= (fsm_output(6)) AND (fsm_output(7)) AND (fsm_output(9));
  mux_tmp_2653 <= MUX_s_1_2_2(nor_569_cse, and_459_cse, fsm_output(6));
  nor_tmp_463 <= (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(7)) AND (fsm_output(9));
  or_2762_nl <= (fsm_output(8)) OR (CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11")));
  mux_2715_itm <= MUX_s_1_2_2(not_tmp_698, or_2762_nl, fsm_output(9));
  nor_tmp_467 <= (fsm_output(5)) AND (fsm_output(8)) AND (fsm_output(9));
  mux_tmp_2666 <= MUX_s_1_2_2(and_dcpl, nor_tmp_130, fsm_output(5));
  not_tmp_729 <= NOT((fsm_output(5)) OR (fsm_output(8)) OR (fsm_output(9)));
  nor_494_nl <= NOT(and_515_cse OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(7))
      OR (fsm_output(9)));
  and_444_nl <= or_2500_cse AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(7))
      AND (fsm_output(9));
  mux_2724_nl <= MUX_s_1_2_2(nor_494_nl, and_444_nl, fsm_output(3));
  and_445_nl <= (fsm_output(3)) AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(7))
      AND (fsm_output(9));
  mux_2725_nl <= MUX_s_1_2_2(mux_2724_nl, and_445_nl, fsm_output(2));
  mux_2726_nl <= MUX_s_1_2_2(nor_497_cse, mux_2725_nl, fsm_output(4));
  mux_2727_itm <= MUX_s_1_2_2(mux_2726_nl, (fsm_output(9)), fsm_output(8));
  and_412_nl <= (fsm_output(8)) AND ((fsm_output(7)) OR mux_tmp_2583);
  mux_2734_itm <= MUX_s_1_2_2(not_tmp_698, and_412_nl, fsm_output(9));
  mux_2739_nl <= MUX_s_1_2_2(not_tmp_662, mux_tmp_2529, fsm_output(3));
  mux_tmp_2689 <= MUX_s_1_2_2(mux_2739_nl, nor_tmp_417, fsm_output(4));
  mux_2741_nl <= MUX_s_1_2_2(mux_tmp_2529, nor_tmp_417, fsm_output(3));
  mux_2742_nl <= MUX_s_1_2_2(not_tmp_662, mux_2741_nl, fsm_output(4));
  mux_2743_nl <= MUX_s_1_2_2(mux_2742_nl, mux_tmp_2689, and_515_cse);
  mux_2744_nl <= MUX_s_1_2_2(mux_2743_nl, mux_tmp_2689, fsm_output(2));
  mux_2745_itm <= MUX_s_1_2_2(mux_2744_nl, nor_tmp_130, fsm_output(7));
  and_694_cse <= (fsm_output(2)) AND (fsm_output(6));
  mux_2762_nl <= MUX_s_1_2_2((NOT (fsm_output(3))), (fsm_output(3)), and_694_cse);
  mux_2763_nl <= MUX_s_1_2_2(mux_2762_nl, mux_tmp_2459, fsm_output(1));
  nor_490_nl <= NOT((fsm_output(5)) OR mux_2763_nl);
  mux_tmp_2713 <= MUX_s_1_2_2(nor_490_nl, mux_tmp_2462, fsm_output(4));
  mux_tmp_2714 <= MUX_s_1_2_2(and_dcpl_96, nor_tmp_1, fsm_output(5));
  mux_tmp_2720 <= MUX_s_1_2_2(mux_tmp_2459, mux_tmp_2467, fsm_output(1));
  or_tmp_2733 <= (fsm_output(5)) OR mux_tmp_2720;
  or_tmp_2734 <= (NOT (fsm_output(5))) OR (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(6))
      OR (fsm_output(3));
  mux_tmp_2721 <= MUX_s_1_2_2(or_tmp_2734, or_tmp_2733, fsm_output(4));
  or_tmp_2735 <= (fsm_output(5)) OR mux_tmp_2459;
  or_tmp_2736 <= (fsm_output(5)) OR not_tmp_617;
  nand_145_nl <= NOT((fsm_output(5)) AND (NOT mux_tmp_2467));
  mux_tmp_2724 <= MUX_s_1_2_2(nand_145_nl, or_tmp_2736, fsm_output(4));
  mux_2782_nl <= MUX_s_1_2_2((NOT (fsm_output(3))), (fsm_output(3)), or_204_cse);
  mux_2783_nl <= MUX_s_1_2_2(mux_tmp_2467, mux_2782_nl, fsm_output(1));
  nand_tmp_148 <= NOT((fsm_output(5)) AND (NOT mux_2783_nl));
  mux_2793_nl <= MUX_s_1_2_2(nand_tmp_148, or_tmp_2588, fsm_output(4));
  mux_2794_nl <= MUX_s_1_2_2(mux_tmp_2724, mux_2793_nl, fsm_output(0));
  mux_2791_nl <= MUX_s_1_2_2(or_tmp_2736, or_tmp_2733, fsm_output(4));
  mux_2792_nl <= MUX_s_1_2_2(mux_tmp_2721, mux_2791_nl, fsm_output(0));
  mux_2795_nl <= MUX_s_1_2_2(mux_2794_nl, mux_2792_nl, fsm_output(7));
  mux_2787_nl <= MUX_s_1_2_2((NOT or_tmp_2549), nor_tmp_399, fsm_output(5));
  mux_2788_nl <= MUX_s_1_2_2((NOT or_tmp_2735), mux_2787_nl, fsm_output(4));
  mux_2789_nl <= MUX_s_1_2_2(mux_tmp_2713, mux_2788_nl, fsm_output(0));
  mux_2784_nl <= MUX_s_1_2_2(or_tmp_2439, (NOT nor_tmp_1), fsm_output(5));
  mux_2785_nl <= MUX_s_1_2_2(mux_2784_nl, nand_tmp_148, fsm_output(4));
  mux_2780_nl <= MUX_s_1_2_2(mux_tmp_2467, mux_79_cse, fsm_output(1));
  nand_147_nl <= NOT((fsm_output(5)) AND (NOT mux_2780_nl));
  mux_2781_nl <= MUX_s_1_2_2((NOT mux_tmp_2714), nand_147_nl, fsm_output(4));
  mux_2786_nl <= MUX_s_1_2_2(mux_2785_nl, mux_2781_nl, fsm_output(0));
  mux_2790_nl <= MUX_s_1_2_2((NOT mux_2789_nl), mux_2786_nl, fsm_output(7));
  mux_2796_nl <= MUX_s_1_2_2(mux_2795_nl, mux_2790_nl, fsm_output(8));
  nand_146_nl <= NOT((fsm_output(5)) AND (NOT mux_tmp_2720));
  mux_2776_nl <= MUX_s_1_2_2(nand_146_nl, or_tmp_2736, fsm_output(4));
  mux_2777_nl <= MUX_s_1_2_2(mux_2776_nl, mux_tmp_2724, fsm_output(0));
  mux_2773_nl <= MUX_s_1_2_2(or_tmp_2734, or_tmp_2735, fsm_output(4));
  mux_2774_nl <= MUX_s_1_2_2(mux_2773_nl, mux_tmp_2721, fsm_output(0));
  mux_2778_nl <= MUX_s_1_2_2(mux_2777_nl, mux_2774_nl, fsm_output(7));
  mux_2767_nl <= MUX_s_1_2_2((NOT mux_79_cse), mux_tmp_2459, fsm_output(1));
  nor_489_nl <= NOT((fsm_output(5)) OR mux_2767_nl);
  mux_2768_nl <= MUX_s_1_2_2(nor_489_nl, mux_tmp_2714, fsm_output(4));
  mux_2769_nl <= MUX_s_1_2_2(mux_2768_nl, mux_tmp_2713, fsm_output(0));
  mux_2770_nl <= MUX_s_1_2_2((NOT mux_2769_nl), or_tmp_2548, fsm_output(7));
  mux_2779_nl <= MUX_s_1_2_2(mux_2778_nl, mux_2770_nl, fsm_output(8));
  mux_2797_itm <= MUX_s_1_2_2(mux_2796_nl, mux_2779_nl, fsm_output(9));
  and_504_nl <= (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(0))) AND
      (fsm_output(9)) AND (NOT mux_2252_cse);
  or_2547_nl <= (fsm_output(9)) OR mux_2252_cse;
  nand_126_nl <= NOT((fsm_output(9)) AND (NOT mux_2252_cse));
  mux_2369_nl <= MUX_s_1_2_2(or_2547_nl, nand_126_nl, fsm_output(0));
  nor_534_nl <= NOT((fsm_output(3)) OR (fsm_output(6)) OR mux_2369_nl);
  mux_2370_nl <= MUX_s_1_2_2(and_504_nl, nor_534_nl, fsm_output(7));
  nor_535_nl <= NOT((NOT (fsm_output(0))) OR (fsm_output(9)) OR nand_169_cse);
  nor_536_nl <= NOT((NOT (fsm_output(0))) OR (fsm_output(9)) OR (fsm_output(2)) OR
      (fsm_output(8)) OR (fsm_output(5)));
  mux_2367_nl <= MUX_s_1_2_2(nor_535_nl, nor_536_nl, fsm_output(6));
  and_505_nl <= (fsm_output(7)) AND (fsm_output(3)) AND mux_2367_nl;
  mux_2371_nl <= MUX_s_1_2_2(mux_2370_nl, and_505_nl, fsm_output(4));
  or_2539_nl <= (NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(8)) OR (NOT (fsm_output(5)));
  mux_2364_nl <= MUX_s_1_2_2(mux_2374_cse, or_2549_cse, fsm_output(6));
  mux_2365_nl <= MUX_s_1_2_2(or_2539_nl, mux_2364_nl, fsm_output(3));
  nor_537_nl <= NOT((fsm_output(7)) OR mux_2365_nl);
  or_2531_nl <= (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(8))) OR (fsm_output(5));
  or_2530_nl <= (NOT (fsm_output(9))) OR (fsm_output(2)) OR (NOT (fsm_output(8)))
      OR (fsm_output(5));
  mux_2361_nl <= MUX_s_1_2_2(or_2531_nl, or_2530_nl, fsm_output(0));
  nor_538_nl <= NOT((fsm_output(3)) OR (fsm_output(6)) OR mux_2361_nl);
  nor_539_nl <= NOT((NOT (fsm_output(6))) OR (fsm_output(0)) OR (fsm_output(9)) OR
      nand_169_cse);
  nor_540_nl <= NOT((NOT (fsm_output(6))) OR (fsm_output(0)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(8)) OR (fsm_output(5)));
  mux_2360_nl <= MUX_s_1_2_2(nor_539_nl, nor_540_nl, fsm_output(3));
  mux_2362_nl <= MUX_s_1_2_2(nor_538_nl, mux_2360_nl, fsm_output(7));
  mux_2366_nl <= MUX_s_1_2_2(nor_537_nl, mux_2362_nl, fsm_output(4));
  COMP_LOOP_10_modExp_dev_1_while_mul_mut_mx0c4 <= MUX_s_1_2_2(mux_2371_nl, mux_2366_nl,
      fsm_output(1));
  or_2571_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(8))) OR (fsm_output(2));
  or_2625_nl <= (fsm_output(8)) OR (NOT (fsm_output(2))) OR (fsm_output(5));
  mux_2382_nl <= MUX_s_1_2_2(or_2571_nl, or_2625_nl, fsm_output(9));
  nand_172_nl <= NOT((fsm_output(9)) AND (fsm_output(5)) AND (fsm_output(8)) AND
      (NOT (fsm_output(2))));
  mux_2383_nl <= MUX_s_1_2_2(mux_2382_nl, nand_172_nl, fsm_output(0));
  nor_525_nl <= NOT((fsm_output(4)) OR (fsm_output(1)) OR mux_2383_nl);
  nor_526_nl <= NOT((NOT (fsm_output(0))) OR (fsm_output(9)) OR (NOT (fsm_output(5)))
      OR (fsm_output(8)) OR (NOT (fsm_output(2))));
  nor_527_nl <= NOT((fsm_output(0)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR (fsm_output(8)) OR (NOT (fsm_output(2))));
  mux_2381_nl <= MUX_s_1_2_2(nor_526_nl, nor_527_nl, fsm_output(1));
  and_501_nl <= (fsm_output(4)) AND mux_2381_nl;
  mux_2384_nl <= MUX_s_1_2_2(nor_525_nl, and_501_nl, fsm_output(6));
  nor_528_nl <= NOT((NOT (fsm_output(4))) OR (fsm_output(1)) OR mux_2374_cse);
  or_2560_nl <= (fsm_output(0)) OR (NOT (fsm_output(9))) OR (fsm_output(5)) OR (NOT
      (fsm_output(8))) OR (fsm_output(2));
  mux_2379_nl <= MUX_s_1_2_2(or_2549_cse, or_2560_nl, fsm_output(1));
  and_502_nl <= (fsm_output(4)) AND (NOT mux_2379_nl);
  mux_2380_nl <= MUX_s_1_2_2(nor_528_nl, and_502_nl, fsm_output(6));
  mux_2385_nl <= MUX_s_1_2_2(mux_2384_nl, mux_2380_nl, fsm_output(3));
  nor_529_nl <= NOT((fsm_output(9)) OR (fsm_output(5)) OR (NOT (fsm_output(8))) OR
      (fsm_output(2)));
  nor_530_nl <= NOT((NOT (fsm_output(9))) OR (fsm_output(5)) OR (NOT (fsm_output(8)))
      OR (fsm_output(2)));
  mux_2376_nl <= MUX_s_1_2_2(nor_529_nl, nor_530_nl, fsm_output(0));
  and_503_nl <= (fsm_output(4)) AND (fsm_output(1)) AND mux_2376_nl;
  mux_2377_nl <= MUX_s_1_2_2(and_503_nl, nor_558_cse, fsm_output(6));
  nor_532_nl <= NOT((fsm_output(4)) OR (NOT (fsm_output(1))) OR mux_2374_cse);
  or_2550_nl <= (fsm_output(0)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5)))
      OR (fsm_output(8)) OR (fsm_output(2));
  mux_2373_nl <= MUX_s_1_2_2(or_2550_nl, or_2549_cse, fsm_output(1));
  nor_533_nl <= NOT((fsm_output(4)) OR mux_2373_nl);
  mux_2375_nl <= MUX_s_1_2_2(nor_532_nl, nor_533_nl, fsm_output(6));
  mux_2378_nl <= MUX_s_1_2_2(mux_2377_nl, mux_2375_nl, fsm_output(3));
  COMP_LOOP_10_modExp_dev_1_while_mul_mut_mx0c5 <= MUX_s_1_2_2(mux_2385_nl, mux_2378_nl,
      fsm_output(7));
  STAGE_VEC_LOOP_j_sva_9_0_mx0c1 <= and_dcpl_268 AND and_dcpl_266 AND nor_tmp_130;
  COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c3 <= and_dcpl_253
      AND and_dcpl_243;
  COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c4 <= and_dcpl_257
      AND and_dcpl_106;
  COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c5 <= and_dcpl_109
      AND and_dcpl_256;
  COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c6 <= and_dcpl_97
      AND and_dcpl_260;
  COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c7 <= and_dcpl_244
      AND and_dcpl_263;
  COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c8 <= and_dcpl_253
      AND and_dcpl_270;
  COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c9 <= and_dcpl_311
      AND and_dcpl_319;
  COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c10 <= and_dcpl_261
      AND and_dcpl_321;
  COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c11 <= and_dcpl_268
      AND and_dcpl_279;
  COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c12 <= and_dcpl_109
      AND and_dcpl_284;
  COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c13 <= and_dcpl_239
      AND and_dcpl_286;
  or_2664_nl <= (fsm_output(5)) OR (NOT nor_tmp_399);
  mux_2541_nl <= MUX_s_1_2_2(nand_tmp_140, or_2664_nl, fsm_output(4));
  mux_2542_nl <= MUX_s_1_2_2(mux_tmp_2474, mux_2541_nl, fsm_output(0));
  mux_2539_nl <= MUX_s_1_2_2(or_tmp_2588, or_tmp_2587, fsm_output(4));
  mux_2540_nl <= MUX_s_1_2_2(mux_tmp_2470, mux_2539_nl, fsm_output(0));
  mux_2543_nl <= MUX_s_1_2_2(mux_2542_nl, mux_2540_nl, fsm_output(7));
  mux_2535_nl <= MUX_s_1_2_2((NOT or_tmp_2549), nor_tmp_403, fsm_output(5));
  mux_2536_nl <= MUX_s_1_2_2((NOT or_tmp_2585), mux_2535_nl, fsm_output(4));
  mux_2537_nl <= MUX_s_1_2_2(mux_tmp_2461, mux_2536_nl, fsm_output(0));
  mux_2532_nl <= MUX_s_1_2_2(or_tmp_2439, (NOT nor_tmp_399), fsm_output(5));
  mux_2533_nl <= MUX_s_1_2_2(mux_2532_nl, nand_tmp_140, fsm_output(4));
  nand_139_nl <= NOT((fsm_output(5)) AND (NOT mux_tmp_2400));
  mux_2530_nl <= MUX_s_1_2_2((NOT mux_tmp_2462), nand_139_nl, fsm_output(4));
  mux_2534_nl <= MUX_s_1_2_2(mux_2533_nl, mux_2530_nl, fsm_output(0));
  mux_2538_nl <= MUX_s_1_2_2((NOT mux_2537_nl), mux_2534_nl, fsm_output(7));
  mux_2544_nl <= MUX_s_1_2_2(mux_2543_nl, mux_2538_nl, fsm_output(8));
  nand_138_nl <= NOT((fsm_output(5)) AND (NOT mux_tmp_2468));
  mux_2526_nl <= MUX_s_1_2_2(nand_138_nl, or_tmp_2588, fsm_output(4));
  mux_2527_nl <= MUX_s_1_2_2(mux_2526_nl, mux_tmp_2474, fsm_output(0));
  mux_2522_nl <= MUX_s_1_2_2(mux_tmp_2469, or_tmp_2585, fsm_output(4));
  mux_2523_nl <= MUX_s_1_2_2(mux_2522_nl, mux_tmp_2470, fsm_output(0));
  mux_2528_nl <= MUX_s_1_2_2(mux_2527_nl, mux_2523_nl, fsm_output(7));
  mux_2514_nl <= MUX_s_1_2_2(and_dcpl_95, mux_tmp_2458, and_516_cse);
  nor_520_nl <= NOT((fsm_output(5)) OR mux_2514_nl);
  mux_2515_nl <= MUX_s_1_2_2(nor_520_nl, mux_tmp_2462, fsm_output(4));
  mux_2516_nl <= MUX_s_1_2_2(mux_2515_nl, mux_tmp_2461, fsm_output(0));
  mux_2517_nl <= MUX_s_1_2_2((NOT mux_2516_nl), or_tmp_2548, fsm_output(7));
  mux_2529_nl <= MUX_s_1_2_2(mux_2528_nl, mux_2517_nl, fsm_output(8));
  mux_2545_itm <= MUX_s_1_2_2(mux_2544_nl, mux_2529_nl, fsm_output(9));
  operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c1 <= and_dcpl_261 AND
      and_dcpl_307;
  operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c2 <= and_dcpl_239 AND
      and_dcpl_267;
  operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c3 <= and_dcpl_257 AND
      and_dcpl_323;
  operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c4 <= and_dcpl_244 AND
      and_dcpl_288;
  tmp_1_lpi_4_dfm_mx0c0 <= and_dcpl_97 AND and_dcpl_346;
  and_332_m1c <= and_dcpl_244 AND and_dcpl_106;
  and_334_m1c <= and_dcpl_239 AND and_dcpl_307;
  and_335_m1c <= and_dcpl_253 AND and_dcpl_256;
  and_338_m1c <= and_dcpl_311 AND and_dcpl_252;
  and_340_m1c <= and_dcpl_261 AND and_dcpl_313;
  and_342_m1c <= and_dcpl_257 AND and_dcpl_242 AND and_dcpl_44;
  and_344_m1c <= and_dcpl_268 AND and_dcpl_317;
  and_346_m1c <= and_dcpl_109 AND and_dcpl_319;
  and_348_m1c <= and_dcpl_239 AND and_dcpl_321;
  and_350_m1c <= and_dcpl_244 AND and_dcpl_323;
  and_351_m1c <= and_dcpl_248 AND and_dcpl_279;
  and_352_m1c <= and_dcpl_253 AND and_dcpl_284;
  and_354_m1c <= and_dcpl_257 AND and_dcpl_255 AND and_dcpl_70;
  and_356_m1c <= and_dcpl_261 AND and_dcpl_329;
  and_358_m1c <= and_dcpl_264 AND and_dcpl_331;
  or_508_nl <= (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1051_nl <= MUX_s_1_2_2(or_508_nl, or_tmp_546, fsm_output(4));
  and_125_nl <= (NOT mux_1051_nl) AND and_dcpl_95 AND (NOT (fsm_output(2))) AND (fsm_output(0))
      AND (NOT (fsm_output(7))) AND and_dcpl;
  and_132_nl <= and_dcpl_109 AND and_dcpl_106;
  and_136_nl <= and_dcpl_113 AND and_dcpl_94 AND (NOT (fsm_output(7))) AND and_dcpl;
  nor_811_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT nor_tmp_1));
  nor_812_nl <= NOT((NOT (fsm_output(0))) OR (NOT (fsm_output(1))) OR (fsm_output(2))
      OR (fsm_output(6)) OR (fsm_output(3)));
  mux_1052_nl <= MUX_s_1_2_2(nor_811_nl, nor_812_nl, fsm_output(7));
  and_139_nl <= mux_1052_nl AND CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("00"))
      AND and_dcpl;
  and_144_nl <= not_tmp_280 AND (NOT (fsm_output(3))) AND (NOT (fsm_output(6))) AND
      (NOT (fsm_output(5))) AND (fsm_output(7)) AND and_dcpl;
  and_556_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 3)=STD_LOGIC_VECTOR'("111"));
  nor_808_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 3)/=STD_LOGIC_VECTOR'("000")));
  mux_1054_nl <= MUX_s_1_2_2(and_556_nl, nor_808_nl, fsm_output(0));
  and_149_nl <= mux_1054_nl AND (NOT (fsm_output(6))) AND and_dcpl_125;
  nor_806_nl <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 4)/=STD_LOGIC_VECTOR'("100")));
  nor_807_nl <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 4)/=STD_LOGIC_VECTOR'("011")));
  mux_1055_nl <= MUX_s_1_2_2(nor_806_nl, nor_807_nl, fsm_output(0));
  and_151_nl <= mux_1055_nl AND (fsm_output(3)) AND and_dcpl_125;
  nor_804_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(6)) OR (NOT (fsm_output(3))));
  nor_805_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(6))) OR (fsm_output(3)));
  mux_1056_nl <= MUX_s_1_2_2(nor_804_nl, nor_805_nl, fsm_output(0));
  and_156_nl <= mux_1056_nl AND (fsm_output(2)) AND and_dcpl_131 AND and_dcpl;
  nor_802_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(0)) OR (NOT((fsm_output(4))
      AND (fsm_output(5)) AND (fsm_output(1)) AND (fsm_output(6)))));
  nor_803_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(0))) OR (fsm_output(4)) OR
      (fsm_output(5)) OR (fsm_output(1)) OR (fsm_output(6)));
  mux_1057_nl <= MUX_s_1_2_2(nor_802_nl, nor_803_nl, fsm_output(8));
  and_159_nl <= mux_1057_nl AND and_dcpl_135 AND (NOT (fsm_output(9)));
  and_555_nl <= (fsm_output(7)) AND (fsm_output(0)) AND (fsm_output(4)) AND (fsm_output(6))
      AND (NOT (fsm_output(3)));
  nor_801_nl <= NOT((fsm_output(7)) OR (fsm_output(0)) OR (fsm_output(4)) OR (fsm_output(6))
      OR (NOT (fsm_output(3))));
  mux_1058_nl <= MUX_s_1_2_2(and_555_nl, nor_801_nl, fsm_output(8));
  and_163_nl <= mux_1058_nl AND and_516_cse AND (fsm_output(5)) AND (NOT (fsm_output(9)));
  and_171_nl <= and_dcpl_147 AND xor_dcpl AND and_dcpl_143 AND (NOT (fsm_output(7)))
      AND and_dcpl_44;
  nor_799_nl <= NOT((NOT (fsm_output(4))) OR (fsm_output(1)) OR (fsm_output(2)) OR
      (fsm_output(6)));
  nor_800_nl <= NOT((fsm_output(4)) OR (NOT((fsm_output(1)) AND (fsm_output(2)) AND
      (fsm_output(6)))));
  mux_1059_nl <= MUX_s_1_2_2(nor_799_nl, nor_800_nl, fsm_output(0));
  and_175_nl <= mux_1059_nl AND (NOT (fsm_output(3))) AND (fsm_output(5)) AND (NOT
      (fsm_output(7))) AND and_dcpl_44;
  nor_798_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100")));
  and_554_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1011"));
  mux_1060_nl <= MUX_s_1_2_2(nor_798_nl, and_554_nl, fsm_output(0));
  and_179_nl <= mux_1060_nl AND and_613_cse AND (NOT (fsm_output(7))) AND and_dcpl_44;
  and_184_nl <= not_tmp_292 AND (NOT (fsm_output(2))) AND and_dcpl_159 AND and_dcpl_44;
  and_188_nl <= and_dcpl_96 AND xor_dcpl AND and_dcpl_158 AND (fsm_output(7)) AND
      and_dcpl_44;
  nor_795_nl <= NOT((fsm_output(4)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(1)))
      OR (fsm_output(6)) OR (fsm_output(3)));
  nor_796_nl <= NOT((NOT (fsm_output(4))) OR (fsm_output(5)) OR (fsm_output(1)) OR
      (NOT and_711_cse));
  mux_1062_nl <= MUX_s_1_2_2(nor_795_nl, nor_796_nl, fsm_output(0));
  and_191_nl <= mux_1062_nl AND (NOT (fsm_output(2))) AND (fsm_output(7)) AND and_dcpl_44;
  nor_793_nl <= NOT((NOT (fsm_output(4))) OR (fsm_output(5)) OR (NOT (fsm_output(1))));
  nor_794_nl <= NOT((fsm_output(4)) OR (NOT (fsm_output(5))) OR (fsm_output(1)));
  mux_1063_nl <= MUX_s_1_2_2(nor_793_nl, nor_794_nl, fsm_output(0));
  and_196_nl <= mux_1063_nl AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(2)))
      AND (fsm_output(7)) AND and_dcpl_44;
  and_552_nl <= (fsm_output(8)) AND (fsm_output(7)) AND (fsm_output(0)) AND (fsm_output(6))
      AND (fsm_output(3));
  nor_792_nl <= NOT((fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(0)) OR (fsm_output(6))
      OR (fsm_output(3)));
  mux_1064_nl <= MUX_s_1_2_2(and_552_nl, nor_792_nl, fsm_output(9));
  and_200_nl <= mux_1064_nl AND and_dcpl_176 AND CONV_SL_1_1(fsm_output(5 DOWNTO
      4)=STD_LOGIC_VECTOR'("01"));
  nor_790_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")));
  nor_791_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("01")));
  mux_1065_nl <= MUX_s_1_2_2(nor_790_nl, nor_791_nl, fsm_output(0));
  and_205_nl <= mux_1065_nl AND and_dcpl_95 AND and_dcpl_176 AND (NOT (fsm_output(7)))
      AND and_dcpl_70;
  nor_788_nl <= NOT((NOT (fsm_output(4))) OR (fsm_output(1)) OR (NOT (fsm_output(2)))
      OR (fsm_output(6)) OR (fsm_output(3)));
  nor_789_nl <= NOT((fsm_output(4)) OR (NOT (fsm_output(1))) OR (fsm_output(2)) OR
      (NOT and_711_cse));
  mux_1066_nl <= MUX_s_1_2_2(nor_788_nl, nor_789_nl, fsm_output(0));
  and_208_nl <= mux_1066_nl AND (NOT (fsm_output(5))) AND (NOT (fsm_output(7))) AND
      and_dcpl_70;
  and_213_nl <= not_tmp_280 AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(5)))
      AND (NOT (fsm_output(7))) AND and_dcpl_70;
  and_218_nl <= not_tmp_292 AND (fsm_output(2)) AND and_dcpl_192 AND (NOT (fsm_output(4)))
      AND and_dcpl_70;
  and_223_nl <= and_dcpl_199 AND xor_dcpl AND and_dcpl_192 AND (fsm_output(7)) AND
      and_dcpl_70;
  nor_786_nl <= NOT((fsm_output(4)) OR (fsm_output(5)) OR (NOT (fsm_output(1))) OR
      (fsm_output(3)));
  and_762_nl <= (fsm_output(4)) AND (fsm_output(5)) AND (NOT (fsm_output(1))) AND
      (fsm_output(3));
  mux_1067_nl <= MUX_s_1_2_2(nor_786_nl, and_762_nl, fsm_output(0));
  and_227_nl <= mux_1067_nl AND (NOT (fsm_output(6))) AND (fsm_output(2)) AND (fsm_output(7))
      AND and_dcpl_70;
  and_551_nl <= (fsm_output(4)) AND (fsm_output(5)) AND (fsm_output(1)) AND (NOT
      (fsm_output(6)));
  nor_785_nl <= NOT((fsm_output(4)) OR (fsm_output(5)) OR (fsm_output(1)) OR (NOT
      (fsm_output(6))));
  mux_1068_nl <= MUX_s_1_2_2(and_551_nl, nor_785_nl, fsm_output(0));
  and_231_nl <= mux_1068_nl AND (fsm_output(3)) AND (fsm_output(2)) AND (fsm_output(7))
      AND and_dcpl_70;
  mux_1069_nl <= MUX_s_1_2_2(or_tmp_33, or_tmp_591, fsm_output(0));
  and_234_nl <= (NOT mux_1069_nl) AND and_516_cse AND and_dcpl_131 AND and_dcpl_70;
  and_550_nl <= (fsm_output(7)) AND (fsm_output(0)) AND (fsm_output(4)) AND (fsm_output(5))
      AND (fsm_output(6));
  nor_784_nl <= NOT((fsm_output(7)) OR (fsm_output(0)) OR (fsm_output(4)) OR (fsm_output(5))
      OR (fsm_output(6)));
  mux_1070_nl <= MUX_s_1_2_2(and_550_nl, nor_784_nl, fsm_output(8));
  and_237_nl <= mux_1070_nl AND and_dcpl_135 AND (fsm_output(1)) AND (fsm_output(9));
  nor_782_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(0)) OR (NOT (fsm_output(4)))
      OR (fsm_output(1)) OR (fsm_output(2)) OR (NOT (fsm_output(6))));
  nor_783_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(0))) OR (fsm_output(4)) OR
      (NOT (fsm_output(1))) OR (NOT (fsm_output(2))) OR (fsm_output(6)));
  mux_1071_nl <= MUX_s_1_2_2(nor_782_nl, nor_783_nl, fsm_output(8));
  and_240_nl <= mux_1071_nl AND (fsm_output(3)) AND (fsm_output(5)) AND (fsm_output(9));
  nor_781_nl <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
  and_549_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111"));
  mux_1072_nl <= MUX_s_1_2_2(nor_781_nl, and_549_nl, fsm_output(0));
  and_245_nl <= mux_1072_nl AND (NOT (fsm_output(6))) AND and_623_cse AND (NOT (fsm_output(7)))
      AND nor_tmp_130;
  nor_779_nl <= NOT((fsm_output(4)) OR (NOT and_711_cse));
  nor_780_nl <= NOT((NOT (fsm_output(4))) OR (fsm_output(6)) OR (fsm_output(3)));
  mux_1073_nl <= MUX_s_1_2_2(nor_779_nl, nor_780_nl, fsm_output(0));
  and_249_nl <= mux_1073_nl AND (NOT (fsm_output(2))) AND and_dcpl_225;
  and_250_nl <= and_dcpl_113 AND and_dcpl_225;
  nor_777_nl <= NOT((fsm_output(0)) OR (NOT((fsm_output(1)) AND (fsm_output(6)) AND
      (fsm_output(3)))));
  nor_778_nl <= NOT((NOT (fsm_output(0))) OR (fsm_output(1)) OR (fsm_output(6)) OR
      (fsm_output(3)));
  mux_1074_nl <= MUX_s_1_2_2(nor_777_nl, nor_778_nl, fsm_output(7));
  and_254_nl <= mux_1074_nl AND (NOT (fsm_output(2))) AND (fsm_output(5)) AND (NOT
      (fsm_output(4))) AND nor_tmp_130;
  vec_rsc_0_0_i_adra_d_pff <= MUX1HOT_v_6_33_2((COMP_LOOP_1_operator_64_false_acc_tmp(9
      DOWNTO 4)), COMP_LOOP_acc_psp_sva, (operator_64_false_acc_cse_1_sva(9 DOWNTO
      4)), (COMP_LOOP_acc_cse_2_sva(9 DOWNTO 4)), (operator_64_false_acc_cse_2_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_7_psp_sva(8 DOWNTO 3)), (operator_64_false_acc_cse_3_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_cse_4_sva(9 DOWNTO 4)), (operator_64_false_acc_cse_4_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_8_psp_sva(7 DOWNTO 2)), (operator_64_false_acc_cse_5_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_cse_6_sva(9 DOWNTO 4)), (operator_64_false_acc_cse_6_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_9_psp_sva(8 DOWNTO 3)), (operator_64_false_acc_cse_7_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_cse_8_sva(9 DOWNTO 4)), (operator_64_false_acc_cse_8_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_10_psp_sva(6 DOWNTO 1)), (operator_64_false_acc_cse_9_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_cse_10_sva(9 DOWNTO 4)), (operator_64_false_acc_cse_10_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_11_psp_sva(8 DOWNTO 3)), (operator_64_false_acc_cse_11_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_cse_12_sva(9 DOWNTO 4)), (operator_64_false_acc_cse_12_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_12_psp_sva(7 DOWNTO 2)), (operator_64_false_acc_cse_13_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_cse_14_sva(9 DOWNTO 4)), (operator_64_false_acc_cse_14_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_13_psp_sva(8 DOWNTO 3)), (operator_64_false_acc_cse_15_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_cse_sva(9 DOWNTO 4)), (operator_64_false_acc_cse_sva(9
      DOWNTO 4)), STD_LOGIC_VECTOR'( and_dcpl_98 & and_125_nl & and_132_nl & and_136_nl
      & and_139_nl & and_144_nl & and_149_nl & and_151_nl & and_156_nl & and_159_nl
      & and_163_nl & and_171_nl & and_175_nl & and_179_nl & and_184_nl & and_188_nl
      & and_191_nl & and_196_nl & and_200_nl & and_205_nl & and_208_nl & and_213_nl
      & and_218_nl & and_223_nl & and_227_nl & and_231_nl & and_234_nl & and_237_nl
      & and_240_nl & and_245_nl & and_249_nl & and_250_nl & and_254_nl));
  vec_rsc_0_0_i_da_d_pff <= COMP_LOOP_1_modulo_dev_cmp_return_rsc_z;
  nor_765_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_766_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1103_nl <= MUX_s_1_2_2(nor_765_nl, nor_766_nl, fsm_output(4));
  nor_767_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_768_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  mux_1102_nl <= MUX_s_1_2_2(nor_767_nl, nor_768_nl, fsm_output(4));
  mux_1104_nl <= MUX_s_1_2_2(mux_1103_nl, mux_1102_nl, fsm_output(8));
  nand_18_nl <= NOT((fsm_output(1)) AND mux_1104_nl);
  nor_769_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(2)) OR not_tmp_311);
  nor_770_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(2)) OR not_tmp_311);
  mux_1100_nl <= MUX_s_1_2_2(nor_769_nl, nor_770_nl, fsm_output(4));
  nand_17_nl <= NOT((fsm_output(8)) AND mux_1100_nl);
  or_711_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_709_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1098_nl <= MUX_s_1_2_2(or_711_nl, or_709_nl, fsm_output(4));
  or_708_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1099_nl <= MUX_s_1_2_2(mux_1098_nl, or_708_nl, fsm_output(8));
  mux_1101_nl <= MUX_s_1_2_2(nand_17_nl, mux_1099_nl, fsm_output(1));
  mux_1105_nl <= MUX_s_1_2_2(nand_18_nl, mux_1101_nl, fsm_output(9));
  or_706_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_705_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1095_nl <= MUX_s_1_2_2(or_706_nl, or_705_nl, fsm_output(4));
  or_703_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_701_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_1094_nl <= MUX_s_1_2_2(or_703_nl, or_701_nl, fsm_output(4));
  mux_1096_nl <= MUX_s_1_2_2(mux_1095_nl, mux_1094_nl, fsm_output(8));
  or_707_nl <= (fsm_output(1)) OR mux_1096_nl;
  or_698_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_697_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1092_nl <= MUX_s_1_2_2(or_698_nl, or_697_nl, fsm_output(4));
  or_699_nl <= (fsm_output(8)) OR mux_1092_nl;
  or_696_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR not_tmp_312;
  mux_1093_nl <= MUX_s_1_2_2(or_699_nl, or_696_nl, fsm_output(1));
  mux_1097_nl <= MUX_s_1_2_2(or_707_nl, mux_1093_nl, fsm_output(9));
  mux_1106_nl <= MUX_s_1_2_2(mux_1105_nl, mux_1097_nl, fsm_output(7));
  or_692_nl <= CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1087_nl <= MUX_s_1_2_2(or_694_cse, or_692_nl, fsm_output(8));
  mux_1088_nl <= MUX_s_1_2_2(mux_1087_nl, nand_tmp_16, fsm_output(1));
  or_691_nl <= (NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1086_nl <= MUX_s_1_2_2(or_691_nl, nand_tmp_16, fsm_output(1));
  mux_1089_nl <= MUX_s_1_2_2(mux_1088_nl, mux_1086_nl, STAGE_VEC_LOOP_j_sva_9_0(3));
  nor_771_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_772_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1083_nl <= MUX_s_1_2_2(nor_771_nl, nor_772_nl, fsm_output(4));
  nor_773_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_774_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(5))));
  mux_1082_nl <= MUX_s_1_2_2(nor_773_nl, nor_774_nl, fsm_output(4));
  mux_1084_nl <= MUX_s_1_2_2(mux_1083_nl, mux_1082_nl, fsm_output(8));
  nand_15_nl <= NOT((fsm_output(1)) AND mux_1084_nl);
  mux_1090_nl <= MUX_s_1_2_2(mux_1089_nl, nand_15_nl, fsm_output(9));
  or_680_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("101")) OR not_tmp_312;
  or_678_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (COMP_LOOP_acc_10_psp_sva(0)) OR (fsm_output(2)) OR not_tmp_311;
  or_676_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5));
  mux_1078_nl <= MUX_s_1_2_2(or_678_nl, or_676_nl, fsm_output(4));
  mux_1079_nl <= MUX_s_1_2_2(or_680_nl, mux_1078_nl, fsm_output(8));
  or_674_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_673_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(5));
  mux_1077_nl <= MUX_s_1_2_2(or_674_nl, or_673_nl, fsm_output(4));
  or_675_nl <= (fsm_output(8)) OR mux_1077_nl;
  mux_1080_nl <= MUX_s_1_2_2(mux_1079_nl, or_675_nl, fsm_output(1));
  or_671_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_670_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1075_nl <= MUX_s_1_2_2(or_671_nl, or_670_nl, fsm_output(4));
  or_668_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  mux_1076_nl <= MUX_s_1_2_2(mux_1075_nl, or_668_nl, fsm_output(8));
  or_672_nl <= (fsm_output(1)) OR mux_1076_nl;
  mux_1081_nl <= MUX_s_1_2_2(mux_1080_nl, or_672_nl, fsm_output(9));
  mux_1091_nl <= MUX_s_1_2_2(mux_1090_nl, mux_1081_nl, fsm_output(7));
  mux_1107_nl <= MUX_s_1_2_2(mux_1106_nl, mux_1091_nl, fsm_output(0));
  vec_rsc_0_0_i_wea_d_pff <= NOT mux_1107_nl;
  or_775_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(5)) OR not_tmp_322;
  or_773_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_772_nl <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_771_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1137_nl <= MUX_s_1_2_2(or_772_nl, or_771_nl, fsm_output(0));
  mux_1138_nl <= MUX_s_1_2_2(or_773_nl, mux_1137_nl, fsm_output(4));
  mux_1139_nl <= MUX_s_1_2_2(or_775_nl, mux_1138_nl, fsm_output(1));
  or_770_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR not_tmp_322;
  or_768_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR not_tmp_322;
  mux_1134_nl <= MUX_s_1_2_2(or_770_nl, or_768_nl, fsm_output(0));
  or_766_nl <= (fsm_output(0)) OR CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1135_nl <= MUX_s_1_2_2(mux_1134_nl, or_766_nl, fsm_output(4));
  or_764_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1136_nl <= MUX_s_1_2_2(mux_1135_nl, or_764_nl, fsm_output(1));
  mux_1140_nl <= MUX_s_1_2_2(mux_1139_nl, mux_1136_nl, fsm_output(9));
  or_763_nl <= CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  or_762_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  mux_1130_nl <= MUX_s_1_2_2(or_763_nl, or_762_nl, fsm_output(0));
  or_761_nl <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  mux_1131_nl <= MUX_s_1_2_2(mux_1130_nl, or_761_nl, fsm_output(4));
  or_760_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(4)) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  mux_1132_nl <= MUX_s_1_2_2(mux_1131_nl, or_760_nl, fsm_output(1));
  or_758_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT (fsm_output(0)))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  or_757_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_756_nl <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1127_nl <= MUX_s_1_2_2(or_757_nl, or_756_nl, fsm_output(0));
  mux_1128_nl <= MUX_s_1_2_2(or_758_nl, mux_1127_nl, fsm_output(4));
  or_755_nl <= CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1129_nl <= MUX_s_1_2_2(mux_1128_nl, or_755_nl, fsm_output(1));
  mux_1133_nl <= MUX_s_1_2_2(mux_1132_nl, mux_1129_nl, fsm_output(9));
  mux_1141_nl <= MUX_s_1_2_2(mux_1140_nl, mux_1133_nl, fsm_output(8));
  or_754_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_752_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1122_nl <= MUX_s_1_2_2(or_754_nl, or_752_nl, fsm_output(0));
  or_750_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR nand_442_cse;
  mux_1123_nl <= MUX_s_1_2_2(mux_1122_nl, or_750_nl, fsm_output(4));
  or_748_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_1119_nl <= MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_748_nl);
  or_747_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_745_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"));
  mux_1120_nl <= MUX_s_1_2_2(mux_1119_nl, or_747_nl, or_745_nl);
  or_744_nl <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT
      (fsm_output(2)));
  mux_1121_nl <= MUX_s_1_2_2(mux_1120_nl, or_744_nl, fsm_output(0));
  nand_20_nl <= NOT((fsm_output(4)) AND (NOT mux_1121_nl));
  mux_1124_nl <= MUX_s_1_2_2(mux_1123_nl, nand_20_nl, fsm_output(1));
  or_742_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT (fsm_output(0)))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_740_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT
      (fsm_output(3))) OR (fsm_output(2));
  mux_1117_nl <= MUX_s_1_2_2(or_742_nl, or_740_nl, fsm_output(4));
  or_739_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3))
      OR (NOT (fsm_output(2)));
  or_737_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_730_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"));
  mux_1113_nl <= MUX_s_1_2_2(mux_1112_cse, nand_437_cse, or_730_nl);
  or_729_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_727_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"));
  mux_1114_nl <= MUX_s_1_2_2(mux_1113_nl, or_729_nl, or_727_nl);
  mux_1115_nl <= MUX_s_1_2_2(or_737_nl, mux_1114_nl, fsm_output(0));
  mux_1116_nl <= MUX_s_1_2_2(or_739_nl, mux_1115_nl, fsm_output(4));
  mux_1118_nl <= MUX_s_1_2_2(mux_1117_nl, mux_1116_nl, fsm_output(1));
  mux_1125_nl <= MUX_s_1_2_2(mux_1124_nl, mux_1118_nl, fsm_output(9));
  or_725_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(4)) OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm)
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_724_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_723_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (COMP_LOOP_acc_10_psp_sva(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_722_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1108_nl <= MUX_s_1_2_2(or_723_nl, or_722_nl, fsm_output(0));
  mux_1109_nl <= MUX_s_1_2_2(or_724_nl, mux_1108_nl, fsm_output(4));
  mux_1110_nl <= MUX_s_1_2_2(or_725_nl, mux_1109_nl, fsm_output(1));
  or_726_nl <= (fsm_output(9)) OR mux_1110_nl;
  mux_1126_nl <= MUX_s_1_2_2(mux_1125_nl, or_726_nl, fsm_output(8));
  mux_1142_nl <= MUX_s_1_2_2(mux_1141_nl, mux_1126_nl, fsm_output(7));
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= NOT mux_1142_nl;
  nor_753_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_754_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1171_nl <= MUX_s_1_2_2(nor_753_nl, nor_754_nl, fsm_output(4));
  nor_755_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_756_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  mux_1170_nl <= MUX_s_1_2_2(nor_755_nl, nor_756_nl, fsm_output(4));
  mux_1172_nl <= MUX_s_1_2_2(mux_1171_nl, mux_1170_nl, fsm_output(8));
  nand_24_nl <= NOT((fsm_output(1)) AND mux_1172_nl);
  nor_757_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(2)) OR not_tmp_311);
  nor_758_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(2)) OR not_tmp_311);
  mux_1168_nl <= MUX_s_1_2_2(nor_757_nl, nor_758_nl, fsm_output(4));
  nand_23_nl <= NOT((fsm_output(8)) AND mux_1168_nl);
  or_820_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_818_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1166_nl <= MUX_s_1_2_2(or_820_nl, or_818_nl, fsm_output(4));
  or_817_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1167_nl <= MUX_s_1_2_2(mux_1166_nl, or_817_nl, fsm_output(8));
  mux_1169_nl <= MUX_s_1_2_2(nand_23_nl, mux_1167_nl, fsm_output(1));
  mux_1173_nl <= MUX_s_1_2_2(nand_24_nl, mux_1169_nl, fsm_output(9));
  or_815_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_814_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1163_nl <= MUX_s_1_2_2(or_815_nl, or_814_nl, fsm_output(4));
  or_812_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_810_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_1162_nl <= MUX_s_1_2_2(or_812_nl, or_810_nl, fsm_output(4));
  mux_1164_nl <= MUX_s_1_2_2(mux_1163_nl, mux_1162_nl, fsm_output(8));
  or_816_nl <= (fsm_output(1)) OR mux_1164_nl;
  or_807_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_806_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1160_nl <= MUX_s_1_2_2(or_807_nl, or_806_nl, fsm_output(4));
  or_808_nl <= (fsm_output(8)) OR mux_1160_nl;
  or_805_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR not_tmp_312;
  mux_1161_nl <= MUX_s_1_2_2(or_808_nl, or_805_nl, fsm_output(1));
  mux_1165_nl <= MUX_s_1_2_2(or_816_nl, mux_1161_nl, fsm_output(9));
  mux_1174_nl <= MUX_s_1_2_2(mux_1173_nl, mux_1165_nl, fsm_output(7));
  or_801_nl <= CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1155_nl <= MUX_s_1_2_2(or_803_cse, or_801_nl, fsm_output(8));
  mux_1156_nl <= MUX_s_1_2_2(mux_1155_nl, nand_tmp_22, fsm_output(1));
  or_800_nl <= (NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1154_nl <= MUX_s_1_2_2(or_800_nl, nand_tmp_22, fsm_output(1));
  mux_1157_nl <= MUX_s_1_2_2(mux_1156_nl, mux_1154_nl, STAGE_VEC_LOOP_j_sva_9_0(3));
  nor_759_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_760_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1151_nl <= MUX_s_1_2_2(nor_759_nl, nor_760_nl, fsm_output(4));
  nor_761_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_762_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(5))));
  mux_1150_nl <= MUX_s_1_2_2(nor_761_nl, nor_762_nl, fsm_output(4));
  mux_1152_nl <= MUX_s_1_2_2(mux_1151_nl, mux_1150_nl, fsm_output(8));
  nand_21_nl <= NOT((fsm_output(1)) AND mux_1152_nl);
  mux_1158_nl <= MUX_s_1_2_2(mux_1157_nl, nand_21_nl, fsm_output(9));
  or_789_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("101")) OR not_tmp_312;
  or_787_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (COMP_LOOP_acc_10_psp_sva(0)) OR (fsm_output(2)) OR not_tmp_311;
  or_785_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5));
  mux_1146_nl <= MUX_s_1_2_2(or_787_nl, or_785_nl, fsm_output(4));
  mux_1147_nl <= MUX_s_1_2_2(or_789_nl, mux_1146_nl, fsm_output(8));
  or_783_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_782_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(2)) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1145_nl <= MUX_s_1_2_2(or_783_nl, or_782_nl, fsm_output(4));
  or_784_nl <= (fsm_output(8)) OR mux_1145_nl;
  mux_1148_nl <= MUX_s_1_2_2(mux_1147_nl, or_784_nl, fsm_output(1));
  or_780_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_779_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1143_nl <= MUX_s_1_2_2(or_780_nl, or_779_nl, fsm_output(4));
  or_777_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  mux_1144_nl <= MUX_s_1_2_2(mux_1143_nl, or_777_nl, fsm_output(8));
  or_781_nl <= (fsm_output(1)) OR mux_1144_nl;
  mux_1149_nl <= MUX_s_1_2_2(mux_1148_nl, or_781_nl, fsm_output(9));
  mux_1159_nl <= MUX_s_1_2_2(mux_1158_nl, mux_1149_nl, fsm_output(7));
  mux_1175_nl <= MUX_s_1_2_2(mux_1174_nl, mux_1159_nl, fsm_output(0));
  vec_rsc_0_1_i_wea_d_pff <= NOT mux_1175_nl;
  or_881_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(5)) OR not_tmp_322;
  or_879_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_878_nl <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_877_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1205_nl <= MUX_s_1_2_2(or_878_nl, or_877_nl, fsm_output(0));
  mux_1206_nl <= MUX_s_1_2_2(or_879_nl, mux_1205_nl, fsm_output(4));
  mux_1207_nl <= MUX_s_1_2_2(or_881_nl, mux_1206_nl, fsm_output(1));
  or_876_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR not_tmp_322;
  or_874_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(5)) OR not_tmp_322;
  mux_1202_nl <= MUX_s_1_2_2(or_876_nl, or_874_nl, fsm_output(0));
  or_872_nl <= (fsm_output(0)) OR CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1203_nl <= MUX_s_1_2_2(mux_1202_nl, or_872_nl, fsm_output(4));
  or_870_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1204_nl <= MUX_s_1_2_2(mux_1203_nl, or_870_nl, fsm_output(1));
  mux_1208_nl <= MUX_s_1_2_2(mux_1207_nl, mux_1204_nl, fsm_output(9));
  or_869_nl <= CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  or_868_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  mux_1198_nl <= MUX_s_1_2_2(or_869_nl, or_868_nl, fsm_output(0));
  or_867_nl <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  mux_1199_nl <= MUX_s_1_2_2(mux_1198_nl, or_867_nl, fsm_output(4));
  or_866_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(4)) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  mux_1200_nl <= MUX_s_1_2_2(mux_1199_nl, or_866_nl, fsm_output(1));
  or_864_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT (fsm_output(0)))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  or_863_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_862_nl <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1195_nl <= MUX_s_1_2_2(or_863_nl, or_862_nl, fsm_output(0));
  mux_1196_nl <= MUX_s_1_2_2(or_864_nl, mux_1195_nl, fsm_output(4));
  or_861_nl <= CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1197_nl <= MUX_s_1_2_2(mux_1196_nl, or_861_nl, fsm_output(1));
  mux_1201_nl <= MUX_s_1_2_2(mux_1200_nl, mux_1197_nl, fsm_output(9));
  mux_1209_nl <= MUX_s_1_2_2(mux_1208_nl, mux_1201_nl, fsm_output(8));
  or_860_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_858_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1190_nl <= MUX_s_1_2_2(or_860_nl, or_858_nl, fsm_output(0));
  or_856_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR nand_442_cse;
  mux_1191_nl <= MUX_s_1_2_2(mux_1190_nl, or_856_nl, fsm_output(4));
  or_854_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_852_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_1187_nl <= MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_852_nl);
  nor_277_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")));
  mux_1188_nl <= MUX_s_1_2_2(or_854_nl, mux_1187_nl, nor_277_nl);
  or_851_nl <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT
      (fsm_output(2)));
  mux_1189_nl <= MUX_s_1_2_2(mux_1188_nl, or_851_nl, fsm_output(0));
  nand_26_nl <= NOT((fsm_output(4)) AND (NOT mux_1189_nl));
  mux_1192_nl <= MUX_s_1_2_2(mux_1191_nl, nand_26_nl, fsm_output(1));
  or_849_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT (fsm_output(0)))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_847_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT
      (fsm_output(3))) OR (fsm_output(2));
  mux_1185_nl <= MUX_s_1_2_2(or_849_nl, or_847_nl, fsm_output(4));
  or_846_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3))
      OR (NOT (fsm_output(2)));
  or_844_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_842_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  nor_275_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")));
  mux_1181_nl <= MUX_s_1_2_2(nand_437_cse, mux_1112_cse, nor_275_nl);
  nor_274_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")));
  mux_1182_nl <= MUX_s_1_2_2(or_842_nl, mux_1181_nl, nor_274_nl);
  mux_1183_nl <= MUX_s_1_2_2(or_844_nl, mux_1182_nl, fsm_output(0));
  mux_1184_nl <= MUX_s_1_2_2(or_846_nl, mux_1183_nl, fsm_output(4));
  mux_1186_nl <= MUX_s_1_2_2(mux_1185_nl, mux_1184_nl, fsm_output(1));
  mux_1193_nl <= MUX_s_1_2_2(mux_1192_nl, mux_1186_nl, fsm_output(9));
  or_834_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(4)) OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm)
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_833_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_832_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (COMP_LOOP_acc_10_psp_sva(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_831_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1176_nl <= MUX_s_1_2_2(or_832_nl, or_831_nl, fsm_output(0));
  mux_1177_nl <= MUX_s_1_2_2(or_833_nl, mux_1176_nl, fsm_output(4));
  mux_1178_nl <= MUX_s_1_2_2(or_834_nl, mux_1177_nl, fsm_output(1));
  or_835_nl <= (fsm_output(9)) OR mux_1178_nl;
  mux_1194_nl <= MUX_s_1_2_2(mux_1193_nl, or_835_nl, fsm_output(8));
  mux_1210_nl <= MUX_s_1_2_2(mux_1209_nl, mux_1194_nl, fsm_output(7));
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= NOT mux_1210_nl;
  nor_741_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_742_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1239_nl <= MUX_s_1_2_2(nor_741_nl, nor_742_nl, fsm_output(4));
  nor_743_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_744_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  mux_1238_nl <= MUX_s_1_2_2(nor_743_nl, nor_744_nl, fsm_output(4));
  mux_1240_nl <= MUX_s_1_2_2(mux_1239_nl, mux_1238_nl, fsm_output(8));
  nand_30_nl <= NOT((fsm_output(1)) AND mux_1240_nl);
  nor_745_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(2)) OR not_tmp_311);
  nor_746_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(2)) OR not_tmp_311);
  mux_1236_nl <= MUX_s_1_2_2(nor_745_nl, nor_746_nl, fsm_output(4));
  nand_29_nl <= NOT((fsm_output(8)) AND mux_1236_nl);
  or_926_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_924_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1234_nl <= MUX_s_1_2_2(or_926_nl, or_924_nl, fsm_output(4));
  or_923_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1235_nl <= MUX_s_1_2_2(mux_1234_nl, or_923_nl, fsm_output(8));
  mux_1237_nl <= MUX_s_1_2_2(nand_29_nl, mux_1235_nl, fsm_output(1));
  mux_1241_nl <= MUX_s_1_2_2(nand_30_nl, mux_1237_nl, fsm_output(9));
  or_921_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_920_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1231_nl <= MUX_s_1_2_2(or_921_nl, or_920_nl, fsm_output(4));
  or_918_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_916_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_1230_nl <= MUX_s_1_2_2(or_918_nl, or_916_nl, fsm_output(4));
  mux_1232_nl <= MUX_s_1_2_2(mux_1231_nl, mux_1230_nl, fsm_output(8));
  or_922_nl <= (fsm_output(1)) OR mux_1232_nl;
  or_913_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_912_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1228_nl <= MUX_s_1_2_2(or_913_nl, or_912_nl, fsm_output(4));
  or_914_nl <= (fsm_output(8)) OR mux_1228_nl;
  or_911_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR not_tmp_312;
  mux_1229_nl <= MUX_s_1_2_2(or_914_nl, or_911_nl, fsm_output(1));
  mux_1233_nl <= MUX_s_1_2_2(or_922_nl, mux_1229_nl, fsm_output(9));
  mux_1242_nl <= MUX_s_1_2_2(mux_1241_nl, mux_1233_nl, fsm_output(7));
  or_907_nl <= CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1223_nl <= MUX_s_1_2_2(or_909_cse, or_907_nl, fsm_output(8));
  mux_1224_nl <= MUX_s_1_2_2(mux_1223_nl, nand_tmp_28, fsm_output(1));
  or_906_nl <= (NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1222_nl <= MUX_s_1_2_2(or_906_nl, nand_tmp_28, fsm_output(1));
  mux_1225_nl <= MUX_s_1_2_2(mux_1224_nl, mux_1222_nl, STAGE_VEC_LOOP_j_sva_9_0(3));
  nor_747_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_748_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1219_nl <= MUX_s_1_2_2(nor_747_nl, nor_748_nl, fsm_output(4));
  nor_749_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_750_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(5))));
  mux_1218_nl <= MUX_s_1_2_2(nor_749_nl, nor_750_nl, fsm_output(4));
  mux_1220_nl <= MUX_s_1_2_2(mux_1219_nl, mux_1218_nl, fsm_output(8));
  nand_27_nl <= NOT((fsm_output(1)) AND mux_1220_nl);
  mux_1226_nl <= MUX_s_1_2_2(mux_1225_nl, nand_27_nl, fsm_output(9));
  or_895_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("101")) OR not_tmp_312;
  or_893_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (COMP_LOOP_acc_10_psp_sva(0)) OR (fsm_output(2)) OR not_tmp_311;
  or_891_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5));
  mux_1214_nl <= MUX_s_1_2_2(or_893_nl, or_891_nl, fsm_output(4));
  mux_1215_nl <= MUX_s_1_2_2(or_895_nl, mux_1214_nl, fsm_output(8));
  or_889_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_888_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(5));
  mux_1213_nl <= MUX_s_1_2_2(or_889_nl, or_888_nl, fsm_output(4));
  or_890_nl <= (fsm_output(8)) OR mux_1213_nl;
  mux_1216_nl <= MUX_s_1_2_2(mux_1215_nl, or_890_nl, fsm_output(1));
  or_886_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_885_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1211_nl <= MUX_s_1_2_2(or_886_nl, or_885_nl, fsm_output(4));
  or_883_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  mux_1212_nl <= MUX_s_1_2_2(mux_1211_nl, or_883_nl, fsm_output(8));
  or_887_nl <= (fsm_output(1)) OR mux_1212_nl;
  mux_1217_nl <= MUX_s_1_2_2(mux_1216_nl, or_887_nl, fsm_output(9));
  mux_1227_nl <= MUX_s_1_2_2(mux_1226_nl, mux_1217_nl, fsm_output(7));
  mux_1243_nl <= MUX_s_1_2_2(mux_1242_nl, mux_1227_nl, fsm_output(0));
  vec_rsc_0_2_i_wea_d_pff <= NOT mux_1243_nl;
  or_990_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(5)) OR not_tmp_322;
  or_988_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_987_nl <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_986_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1273_nl <= MUX_s_1_2_2(or_987_nl, or_986_nl, fsm_output(0));
  mux_1274_nl <= MUX_s_1_2_2(or_988_nl, mux_1273_nl, fsm_output(4));
  mux_1275_nl <= MUX_s_1_2_2(or_990_nl, mux_1274_nl, fsm_output(1));
  or_985_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR not_tmp_322;
  or_983_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR not_tmp_322;
  mux_1270_nl <= MUX_s_1_2_2(or_985_nl, or_983_nl, fsm_output(0));
  or_981_nl <= (fsm_output(0)) OR CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1271_nl <= MUX_s_1_2_2(mux_1270_nl, or_981_nl, fsm_output(4));
  or_979_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1272_nl <= MUX_s_1_2_2(mux_1271_nl, or_979_nl, fsm_output(1));
  mux_1276_nl <= MUX_s_1_2_2(mux_1275_nl, mux_1272_nl, fsm_output(9));
  or_978_nl <= CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  or_977_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  mux_1266_nl <= MUX_s_1_2_2(or_978_nl, or_977_nl, fsm_output(0));
  or_976_nl <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  mux_1267_nl <= MUX_s_1_2_2(mux_1266_nl, or_976_nl, fsm_output(4));
  or_975_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(4)) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  mux_1268_nl <= MUX_s_1_2_2(mux_1267_nl, or_975_nl, fsm_output(1));
  or_973_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT
      (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  or_972_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_971_nl <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1263_nl <= MUX_s_1_2_2(or_972_nl, or_971_nl, fsm_output(0));
  mux_1264_nl <= MUX_s_1_2_2(or_973_nl, mux_1263_nl, fsm_output(4));
  or_970_nl <= CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1265_nl <= MUX_s_1_2_2(mux_1264_nl, or_970_nl, fsm_output(1));
  mux_1269_nl <= MUX_s_1_2_2(mux_1268_nl, mux_1265_nl, fsm_output(9));
  mux_1277_nl <= MUX_s_1_2_2(mux_1276_nl, mux_1269_nl, fsm_output(8));
  or_969_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_967_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1258_nl <= MUX_s_1_2_2(or_969_nl, or_967_nl, fsm_output(0));
  or_965_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR nand_442_cse;
  mux_1259_nl <= MUX_s_1_2_2(mux_1258_nl, or_965_nl, fsm_output(4));
  or_963_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_1255_nl <= MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_963_nl);
  or_962_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_960_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"));
  mux_1256_nl <= MUX_s_1_2_2(mux_1255_nl, or_962_nl, or_960_nl);
  or_959_nl <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT
      (fsm_output(2)));
  mux_1257_nl <= MUX_s_1_2_2(mux_1256_nl, or_959_nl, fsm_output(0));
  nand_32_nl <= NOT((fsm_output(4)) AND (NOT mux_1257_nl));
  mux_1260_nl <= MUX_s_1_2_2(mux_1259_nl, nand_32_nl, fsm_output(1));
  or_957_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT
      (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_955_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT
      (fsm_output(3))) OR (fsm_output(2));
  mux_1253_nl <= MUX_s_1_2_2(or_957_nl, or_955_nl, fsm_output(4));
  or_954_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3))
      OR (NOT (fsm_output(2)));
  or_952_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_945_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"));
  mux_1249_nl <= MUX_s_1_2_2(mux_1112_cse, nand_437_cse, or_945_nl);
  or_944_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_942_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"));
  mux_1250_nl <= MUX_s_1_2_2(mux_1249_nl, or_944_nl, or_942_nl);
  mux_1251_nl <= MUX_s_1_2_2(or_952_nl, mux_1250_nl, fsm_output(0));
  mux_1252_nl <= MUX_s_1_2_2(or_954_nl, mux_1251_nl, fsm_output(4));
  mux_1254_nl <= MUX_s_1_2_2(mux_1253_nl, mux_1252_nl, fsm_output(1));
  mux_1261_nl <= MUX_s_1_2_2(mux_1260_nl, mux_1254_nl, fsm_output(9));
  or_940_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(4)) OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm)
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_939_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_938_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (COMP_LOOP_acc_10_psp_sva(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_937_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1244_nl <= MUX_s_1_2_2(or_938_nl, or_937_nl, fsm_output(0));
  mux_1245_nl <= MUX_s_1_2_2(or_939_nl, mux_1244_nl, fsm_output(4));
  mux_1246_nl <= MUX_s_1_2_2(or_940_nl, mux_1245_nl, fsm_output(1));
  or_941_nl <= (fsm_output(9)) OR mux_1246_nl;
  mux_1262_nl <= MUX_s_1_2_2(mux_1261_nl, or_941_nl, fsm_output(8));
  mux_1278_nl <= MUX_s_1_2_2(mux_1277_nl, mux_1262_nl, fsm_output(7));
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= NOT mux_1278_nl;
  nor_729_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_730_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1307_nl <= MUX_s_1_2_2(nor_729_nl, nor_730_nl, fsm_output(4));
  nor_731_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_732_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  mux_1306_nl <= MUX_s_1_2_2(nor_731_nl, nor_732_nl, fsm_output(4));
  mux_1308_nl <= MUX_s_1_2_2(mux_1307_nl, mux_1306_nl, fsm_output(8));
  nand_36_nl <= NOT((fsm_output(1)) AND mux_1308_nl);
  nor_733_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(2)) OR not_tmp_311);
  nor_734_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(2)) OR not_tmp_311);
  mux_1304_nl <= MUX_s_1_2_2(nor_733_nl, nor_734_nl, fsm_output(4));
  nand_35_nl <= NOT((fsm_output(8)) AND mux_1304_nl);
  or_1035_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1033_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1302_nl <= MUX_s_1_2_2(or_1035_nl, or_1033_nl, fsm_output(4));
  or_1032_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0011")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1303_nl <= MUX_s_1_2_2(mux_1302_nl, or_1032_nl, fsm_output(8));
  mux_1305_nl <= MUX_s_1_2_2(nand_35_nl, mux_1303_nl, fsm_output(1));
  mux_1309_nl <= MUX_s_1_2_2(nand_36_nl, mux_1305_nl, fsm_output(9));
  or_1030_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_1029_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1299_nl <= MUX_s_1_2_2(or_1030_nl, or_1029_nl, fsm_output(4));
  or_1027_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1025_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_1298_nl <= MUX_s_1_2_2(or_1027_nl, or_1025_nl, fsm_output(4));
  mux_1300_nl <= MUX_s_1_2_2(mux_1299_nl, mux_1298_nl, fsm_output(8));
  or_1031_nl <= (fsm_output(1)) OR mux_1300_nl;
  or_1022_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1021_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1296_nl <= MUX_s_1_2_2(or_1022_nl, or_1021_nl, fsm_output(4));
  or_1023_nl <= (fsm_output(8)) OR mux_1296_nl;
  or_1020_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR not_tmp_312;
  mux_1297_nl <= MUX_s_1_2_2(or_1023_nl, or_1020_nl, fsm_output(1));
  mux_1301_nl <= MUX_s_1_2_2(or_1031_nl, mux_1297_nl, fsm_output(9));
  mux_1310_nl <= MUX_s_1_2_2(mux_1309_nl, mux_1301_nl, fsm_output(7));
  or_1016_nl <= CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1291_nl <= MUX_s_1_2_2(or_1018_cse, or_1016_nl, fsm_output(8));
  mux_1292_nl <= MUX_s_1_2_2(mux_1291_nl, nand_tmp_34, fsm_output(1));
  or_1015_nl <= (NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1290_nl <= MUX_s_1_2_2(or_1015_nl, nand_tmp_34, fsm_output(1));
  mux_1293_nl <= MUX_s_1_2_2(mux_1292_nl, mux_1290_nl, STAGE_VEC_LOOP_j_sva_9_0(3));
  nor_735_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_736_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1287_nl <= MUX_s_1_2_2(nor_735_nl, nor_736_nl, fsm_output(4));
  nor_737_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_738_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(5))));
  mux_1286_nl <= MUX_s_1_2_2(nor_737_nl, nor_738_nl, fsm_output(4));
  mux_1288_nl <= MUX_s_1_2_2(mux_1287_nl, mux_1286_nl, fsm_output(8));
  nand_33_nl <= NOT((fsm_output(1)) AND mux_1288_nl);
  mux_1294_nl <= MUX_s_1_2_2(mux_1293_nl, nand_33_nl, fsm_output(9));
  or_1004_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("101")) OR not_tmp_312;
  or_1002_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (COMP_LOOP_acc_10_psp_sva(0)) OR (fsm_output(2)) OR not_tmp_311;
  or_1000_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5));
  mux_1282_nl <= MUX_s_1_2_2(or_1002_nl, or_1000_nl, fsm_output(4));
  mux_1283_nl <= MUX_s_1_2_2(or_1004_nl, mux_1282_nl, fsm_output(8));
  or_998_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_997_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(2)) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1281_nl <= MUX_s_1_2_2(or_998_nl, or_997_nl, fsm_output(4));
  or_999_nl <= (fsm_output(8)) OR mux_1281_nl;
  mux_1284_nl <= MUX_s_1_2_2(mux_1283_nl, or_999_nl, fsm_output(1));
  or_995_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_994_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1279_nl <= MUX_s_1_2_2(or_995_nl, or_994_nl, fsm_output(4));
  or_992_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  mux_1280_nl <= MUX_s_1_2_2(mux_1279_nl, or_992_nl, fsm_output(8));
  or_996_nl <= (fsm_output(1)) OR mux_1280_nl;
  mux_1285_nl <= MUX_s_1_2_2(mux_1284_nl, or_996_nl, fsm_output(9));
  mux_1295_nl <= MUX_s_1_2_2(mux_1294_nl, mux_1285_nl, fsm_output(7));
  mux_1311_nl <= MUX_s_1_2_2(mux_1310_nl, mux_1295_nl, fsm_output(0));
  vec_rsc_0_3_i_wea_d_pff <= NOT mux_1311_nl;
  or_1096_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(5)) OR not_tmp_322;
  or_1094_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_1093_nl <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1092_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1341_nl <= MUX_s_1_2_2(or_1093_nl, or_1092_nl, fsm_output(0));
  mux_1342_nl <= MUX_s_1_2_2(or_1094_nl, mux_1341_nl, fsm_output(4));
  mux_1343_nl <= MUX_s_1_2_2(or_1096_nl, mux_1342_nl, fsm_output(1));
  or_1091_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR not_tmp_322;
  or_1089_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR not_tmp_322;
  mux_1338_nl <= MUX_s_1_2_2(or_1091_nl, or_1089_nl, fsm_output(0));
  or_1087_nl <= (fsm_output(0)) OR CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1339_nl <= MUX_s_1_2_2(mux_1338_nl, or_1087_nl, fsm_output(4));
  or_1085_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1340_nl <= MUX_s_1_2_2(mux_1339_nl, or_1085_nl, fsm_output(1));
  mux_1344_nl <= MUX_s_1_2_2(mux_1343_nl, mux_1340_nl, fsm_output(9));
  or_1084_nl <= CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  or_1083_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  mux_1334_nl <= MUX_s_1_2_2(or_1084_nl, or_1083_nl, fsm_output(0));
  or_1082_nl <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  mux_1335_nl <= MUX_s_1_2_2(mux_1334_nl, or_1082_nl, fsm_output(4));
  or_1081_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(4)) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  mux_1336_nl <= MUX_s_1_2_2(mux_1335_nl, or_1081_nl, fsm_output(1));
  nand_357_nl <= NOT(operator_64_false_slc_operator_64_false_acc_1_60_itm AND (fsm_output(0))
      AND CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0011"))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  or_1078_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1077_nl <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1331_nl <= MUX_s_1_2_2(or_1078_nl, or_1077_nl, fsm_output(0));
  mux_1332_nl <= MUX_s_1_2_2(nand_357_nl, mux_1331_nl, fsm_output(4));
  or_1076_nl <= CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1333_nl <= MUX_s_1_2_2(mux_1332_nl, or_1076_nl, fsm_output(1));
  mux_1337_nl <= MUX_s_1_2_2(mux_1336_nl, mux_1333_nl, fsm_output(9));
  mux_1345_nl <= MUX_s_1_2_2(mux_1344_nl, mux_1337_nl, fsm_output(8));
  or_1075_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1073_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1326_nl <= MUX_s_1_2_2(or_1075_nl, or_1073_nl, fsm_output(0));
  or_1071_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR nand_442_cse;
  mux_1327_nl <= MUX_s_1_2_2(mux_1326_nl, or_1071_nl, fsm_output(4));
  or_1069_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1067_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_1323_nl <= MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_1067_nl);
  nor_288_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")));
  mux_1324_nl <= MUX_s_1_2_2(or_1069_nl, mux_1323_nl, nor_288_nl);
  or_1066_nl <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT
      (fsm_output(2)));
  mux_1325_nl <= MUX_s_1_2_2(mux_1324_nl, or_1066_nl, fsm_output(0));
  nand_38_nl <= NOT((fsm_output(4)) AND (NOT mux_1325_nl));
  mux_1328_nl <= MUX_s_1_2_2(mux_1327_nl, nand_38_nl, fsm_output(1));
  or_1064_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT
      (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1062_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT
      (fsm_output(3))) OR (fsm_output(2));
  mux_1321_nl <= MUX_s_1_2_2(or_1064_nl, or_1062_nl, fsm_output(4));
  or_1061_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3))
      OR (NOT (fsm_output(2)));
  or_1059_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_1057_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  nor_286_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")));
  mux_1317_nl <= MUX_s_1_2_2(nand_437_cse, mux_1112_cse, nor_286_nl);
  nor_285_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")));
  mux_1318_nl <= MUX_s_1_2_2(or_1057_nl, mux_1317_nl, nor_285_nl);
  mux_1319_nl <= MUX_s_1_2_2(or_1059_nl, mux_1318_nl, fsm_output(0));
  mux_1320_nl <= MUX_s_1_2_2(or_1061_nl, mux_1319_nl, fsm_output(4));
  mux_1322_nl <= MUX_s_1_2_2(mux_1321_nl, mux_1320_nl, fsm_output(1));
  mux_1329_nl <= MUX_s_1_2_2(mux_1328_nl, mux_1322_nl, fsm_output(9));
  or_1049_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(4)) OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm)
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1048_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1047_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (COMP_LOOP_acc_10_psp_sva(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_1046_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1312_nl <= MUX_s_1_2_2(or_1047_nl, or_1046_nl, fsm_output(0));
  mux_1313_nl <= MUX_s_1_2_2(or_1048_nl, mux_1312_nl, fsm_output(4));
  mux_1314_nl <= MUX_s_1_2_2(or_1049_nl, mux_1313_nl, fsm_output(1));
  or_1050_nl <= (fsm_output(9)) OR mux_1314_nl;
  mux_1330_nl <= MUX_s_1_2_2(mux_1329_nl, or_1050_nl, fsm_output(8));
  mux_1346_nl <= MUX_s_1_2_2(mux_1345_nl, mux_1330_nl, fsm_output(7));
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= NOT mux_1346_nl;
  nor_717_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_718_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1375_nl <= MUX_s_1_2_2(nor_717_nl, nor_718_nl, fsm_output(4));
  nor_719_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_720_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  mux_1374_nl <= MUX_s_1_2_2(nor_719_nl, nor_720_nl, fsm_output(4));
  mux_1376_nl <= MUX_s_1_2_2(mux_1375_nl, mux_1374_nl, fsm_output(8));
  nand_42_nl <= NOT((fsm_output(1)) AND mux_1376_nl);
  nor_721_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(2)) OR not_tmp_311);
  nor_722_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(2)) OR not_tmp_311);
  mux_1372_nl <= MUX_s_1_2_2(nor_721_nl, nor_722_nl, fsm_output(4));
  nand_41_nl <= NOT((fsm_output(8)) AND mux_1372_nl);
  or_1141_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1139_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1370_nl <= MUX_s_1_2_2(or_1141_nl, or_1139_nl, fsm_output(4));
  or_1138_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1371_nl <= MUX_s_1_2_2(mux_1370_nl, or_1138_nl, fsm_output(8));
  mux_1373_nl <= MUX_s_1_2_2(nand_41_nl, mux_1371_nl, fsm_output(1));
  mux_1377_nl <= MUX_s_1_2_2(nand_42_nl, mux_1373_nl, fsm_output(9));
  or_1136_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_1135_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1367_nl <= MUX_s_1_2_2(or_1136_nl, or_1135_nl, fsm_output(4));
  or_1133_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1131_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_1366_nl <= MUX_s_1_2_2(or_1133_nl, or_1131_nl, fsm_output(4));
  mux_1368_nl <= MUX_s_1_2_2(mux_1367_nl, mux_1366_nl, fsm_output(8));
  or_1137_nl <= (fsm_output(1)) OR mux_1368_nl;
  or_1128_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1127_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1364_nl <= MUX_s_1_2_2(or_1128_nl, or_1127_nl, fsm_output(4));
  or_1129_nl <= (fsm_output(8)) OR mux_1364_nl;
  or_1126_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR not_tmp_312;
  mux_1365_nl <= MUX_s_1_2_2(or_1129_nl, or_1126_nl, fsm_output(1));
  mux_1369_nl <= MUX_s_1_2_2(or_1137_nl, mux_1365_nl, fsm_output(9));
  mux_1378_nl <= MUX_s_1_2_2(mux_1377_nl, mux_1369_nl, fsm_output(7));
  or_1122_nl <= CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1359_nl <= MUX_s_1_2_2(or_1124_cse, or_1122_nl, fsm_output(8));
  mux_1360_nl <= MUX_s_1_2_2(mux_1359_nl, nand_tmp_40, fsm_output(1));
  or_1121_nl <= (NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1358_nl <= MUX_s_1_2_2(or_1121_nl, nand_tmp_40, fsm_output(1));
  mux_1361_nl <= MUX_s_1_2_2(mux_1360_nl, mux_1358_nl, STAGE_VEC_LOOP_j_sva_9_0(3));
  nor_723_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_724_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1355_nl <= MUX_s_1_2_2(nor_723_nl, nor_724_nl, fsm_output(4));
  nor_725_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_726_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(5))));
  mux_1354_nl <= MUX_s_1_2_2(nor_725_nl, nor_726_nl, fsm_output(4));
  mux_1356_nl <= MUX_s_1_2_2(mux_1355_nl, mux_1354_nl, fsm_output(8));
  nand_39_nl <= NOT((fsm_output(1)) AND mux_1356_nl);
  mux_1362_nl <= MUX_s_1_2_2(mux_1361_nl, nand_39_nl, fsm_output(9));
  or_1110_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("101")) OR not_tmp_312;
  or_1108_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (COMP_LOOP_acc_10_psp_sva(0)) OR (fsm_output(2)) OR not_tmp_311;
  or_1106_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5));
  mux_1350_nl <= MUX_s_1_2_2(or_1108_nl, or_1106_nl, fsm_output(4));
  mux_1351_nl <= MUX_s_1_2_2(or_1110_nl, mux_1350_nl, fsm_output(8));
  or_1104_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1103_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(5));
  mux_1349_nl <= MUX_s_1_2_2(or_1104_nl, or_1103_nl, fsm_output(4));
  or_1105_nl <= (fsm_output(8)) OR mux_1349_nl;
  mux_1352_nl <= MUX_s_1_2_2(mux_1351_nl, or_1105_nl, fsm_output(1));
  or_1101_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_1100_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1347_nl <= MUX_s_1_2_2(or_1101_nl, or_1100_nl, fsm_output(4));
  or_1098_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  mux_1348_nl <= MUX_s_1_2_2(mux_1347_nl, or_1098_nl, fsm_output(8));
  or_1102_nl <= (fsm_output(1)) OR mux_1348_nl;
  mux_1353_nl <= MUX_s_1_2_2(mux_1352_nl, or_1102_nl, fsm_output(9));
  mux_1363_nl <= MUX_s_1_2_2(mux_1362_nl, mux_1353_nl, fsm_output(7));
  mux_1379_nl <= MUX_s_1_2_2(mux_1378_nl, mux_1363_nl, fsm_output(0));
  vec_rsc_0_4_i_wea_d_pff <= NOT mux_1379_nl;
  or_1205_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(5)) OR not_tmp_322;
  or_1203_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_1202_nl <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1201_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1409_nl <= MUX_s_1_2_2(or_1202_nl, or_1201_nl, fsm_output(0));
  mux_1410_nl <= MUX_s_1_2_2(or_1203_nl, mux_1409_nl, fsm_output(4));
  mux_1411_nl <= MUX_s_1_2_2(or_1205_nl, mux_1410_nl, fsm_output(1));
  or_1200_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR not_tmp_322;
  or_1198_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR not_tmp_322;
  mux_1406_nl <= MUX_s_1_2_2(or_1200_nl, or_1198_nl, fsm_output(0));
  or_1196_nl <= (fsm_output(0)) OR CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1407_nl <= MUX_s_1_2_2(mux_1406_nl, or_1196_nl, fsm_output(4));
  or_1194_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1408_nl <= MUX_s_1_2_2(mux_1407_nl, or_1194_nl, fsm_output(1));
  mux_1412_nl <= MUX_s_1_2_2(mux_1411_nl, mux_1408_nl, fsm_output(9));
  or_1193_nl <= CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  or_1192_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  mux_1402_nl <= MUX_s_1_2_2(or_1193_nl, or_1192_nl, fsm_output(0));
  or_1191_nl <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  mux_1403_nl <= MUX_s_1_2_2(mux_1402_nl, or_1191_nl, fsm_output(4));
  or_1190_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(4)) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  mux_1404_nl <= MUX_s_1_2_2(mux_1403_nl, or_1190_nl, fsm_output(1));
  or_1188_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT (fsm_output(0)))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  or_1187_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1186_nl <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1399_nl <= MUX_s_1_2_2(or_1187_nl, or_1186_nl, fsm_output(0));
  mux_1400_nl <= MUX_s_1_2_2(or_1188_nl, mux_1399_nl, fsm_output(4));
  or_1185_nl <= CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1401_nl <= MUX_s_1_2_2(mux_1400_nl, or_1185_nl, fsm_output(1));
  mux_1405_nl <= MUX_s_1_2_2(mux_1404_nl, mux_1401_nl, fsm_output(9));
  mux_1413_nl <= MUX_s_1_2_2(mux_1412_nl, mux_1405_nl, fsm_output(8));
  or_1184_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1182_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1394_nl <= MUX_s_1_2_2(or_1184_nl, or_1182_nl, fsm_output(0));
  or_1180_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR nand_442_cse;
  mux_1395_nl <= MUX_s_1_2_2(mux_1394_nl, or_1180_nl, fsm_output(4));
  or_1178_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_1391_nl <= MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_1178_nl);
  or_1177_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1175_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"));
  mux_1392_nl <= MUX_s_1_2_2(mux_1391_nl, or_1177_nl, or_1175_nl);
  or_1174_nl <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT
      (fsm_output(2)));
  mux_1393_nl <= MUX_s_1_2_2(mux_1392_nl, or_1174_nl, fsm_output(0));
  nand_44_nl <= NOT((fsm_output(4)) AND (NOT mux_1393_nl));
  mux_1396_nl <= MUX_s_1_2_2(mux_1395_nl, nand_44_nl, fsm_output(1));
  or_1172_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT (fsm_output(0)))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1170_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT
      (fsm_output(3))) OR (fsm_output(2));
  mux_1389_nl <= MUX_s_1_2_2(or_1172_nl, or_1170_nl, fsm_output(4));
  or_1169_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3))
      OR (NOT (fsm_output(2)));
  or_1167_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_1160_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"));
  mux_1385_nl <= MUX_s_1_2_2(mux_1112_cse, nand_437_cse, or_1160_nl);
  or_1159_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_1157_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"));
  mux_1386_nl <= MUX_s_1_2_2(mux_1385_nl, or_1159_nl, or_1157_nl);
  mux_1387_nl <= MUX_s_1_2_2(or_1167_nl, mux_1386_nl, fsm_output(0));
  mux_1388_nl <= MUX_s_1_2_2(or_1169_nl, mux_1387_nl, fsm_output(4));
  mux_1390_nl <= MUX_s_1_2_2(mux_1389_nl, mux_1388_nl, fsm_output(1));
  mux_1397_nl <= MUX_s_1_2_2(mux_1396_nl, mux_1390_nl, fsm_output(9));
  or_1155_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(4)) OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm)
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1154_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1153_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (COMP_LOOP_acc_10_psp_sva(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_1152_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1380_nl <= MUX_s_1_2_2(or_1153_nl, or_1152_nl, fsm_output(0));
  mux_1381_nl <= MUX_s_1_2_2(or_1154_nl, mux_1380_nl, fsm_output(4));
  mux_1382_nl <= MUX_s_1_2_2(or_1155_nl, mux_1381_nl, fsm_output(1));
  or_1156_nl <= (fsm_output(9)) OR mux_1382_nl;
  mux_1398_nl <= MUX_s_1_2_2(mux_1397_nl, or_1156_nl, fsm_output(8));
  mux_1414_nl <= MUX_s_1_2_2(mux_1413_nl, mux_1398_nl, fsm_output(7));
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= NOT mux_1414_nl;
  nor_705_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_706_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1443_nl <= MUX_s_1_2_2(nor_705_nl, nor_706_nl, fsm_output(4));
  nor_707_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_708_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  mux_1442_nl <= MUX_s_1_2_2(nor_707_nl, nor_708_nl, fsm_output(4));
  mux_1444_nl <= MUX_s_1_2_2(mux_1443_nl, mux_1442_nl, fsm_output(8));
  nand_48_nl <= NOT((fsm_output(1)) AND mux_1444_nl);
  nor_709_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(2)) OR not_tmp_311);
  nor_710_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(2)) OR not_tmp_311);
  mux_1440_nl <= MUX_s_1_2_2(nor_709_nl, nor_710_nl, fsm_output(4));
  nand_47_nl <= NOT((fsm_output(8)) AND mux_1440_nl);
  or_1250_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1248_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1438_nl <= MUX_s_1_2_2(or_1250_nl, or_1248_nl, fsm_output(4));
  or_1247_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0101")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1439_nl <= MUX_s_1_2_2(mux_1438_nl, or_1247_nl, fsm_output(8));
  mux_1441_nl <= MUX_s_1_2_2(nand_47_nl, mux_1439_nl, fsm_output(1));
  mux_1445_nl <= MUX_s_1_2_2(nand_48_nl, mux_1441_nl, fsm_output(9));
  or_1245_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_1244_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1435_nl <= MUX_s_1_2_2(or_1245_nl, or_1244_nl, fsm_output(4));
  or_1242_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1240_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_1434_nl <= MUX_s_1_2_2(or_1242_nl, or_1240_nl, fsm_output(4));
  mux_1436_nl <= MUX_s_1_2_2(mux_1435_nl, mux_1434_nl, fsm_output(8));
  or_1246_nl <= (fsm_output(1)) OR mux_1436_nl;
  or_1237_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1236_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1432_nl <= MUX_s_1_2_2(or_1237_nl, or_1236_nl, fsm_output(4));
  or_1238_nl <= (fsm_output(8)) OR mux_1432_nl;
  or_1235_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR not_tmp_312;
  mux_1433_nl <= MUX_s_1_2_2(or_1238_nl, or_1235_nl, fsm_output(1));
  mux_1437_nl <= MUX_s_1_2_2(or_1246_nl, mux_1433_nl, fsm_output(9));
  mux_1446_nl <= MUX_s_1_2_2(mux_1445_nl, mux_1437_nl, fsm_output(7));
  or_1231_nl <= CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1427_nl <= MUX_s_1_2_2(or_1233_cse, or_1231_nl, fsm_output(8));
  mux_1428_nl <= MUX_s_1_2_2(mux_1427_nl, nand_tmp_46, fsm_output(1));
  or_1230_nl <= (NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1426_nl <= MUX_s_1_2_2(or_1230_nl, nand_tmp_46, fsm_output(1));
  mux_1429_nl <= MUX_s_1_2_2(mux_1428_nl, mux_1426_nl, STAGE_VEC_LOOP_j_sva_9_0(3));
  nor_711_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_712_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1423_nl <= MUX_s_1_2_2(nor_711_nl, nor_712_nl, fsm_output(4));
  nor_713_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_714_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(5))));
  mux_1422_nl <= MUX_s_1_2_2(nor_713_nl, nor_714_nl, fsm_output(4));
  mux_1424_nl <= MUX_s_1_2_2(mux_1423_nl, mux_1422_nl, fsm_output(8));
  nand_45_nl <= NOT((fsm_output(1)) AND mux_1424_nl);
  mux_1430_nl <= MUX_s_1_2_2(mux_1429_nl, nand_45_nl, fsm_output(9));
  or_1219_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("101")) OR not_tmp_312;
  or_1217_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (COMP_LOOP_acc_10_psp_sva(0)) OR (fsm_output(2)) OR not_tmp_311;
  or_1215_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5));
  mux_1418_nl <= MUX_s_1_2_2(or_1217_nl, or_1215_nl, fsm_output(4));
  mux_1419_nl <= MUX_s_1_2_2(or_1219_nl, mux_1418_nl, fsm_output(8));
  or_1213_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1212_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(2)) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1417_nl <= MUX_s_1_2_2(or_1213_nl, or_1212_nl, fsm_output(4));
  or_1214_nl <= (fsm_output(8)) OR mux_1417_nl;
  mux_1420_nl <= MUX_s_1_2_2(mux_1419_nl, or_1214_nl, fsm_output(1));
  or_1210_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_1209_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1415_nl <= MUX_s_1_2_2(or_1210_nl, or_1209_nl, fsm_output(4));
  or_1207_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  mux_1416_nl <= MUX_s_1_2_2(mux_1415_nl, or_1207_nl, fsm_output(8));
  or_1211_nl <= (fsm_output(1)) OR mux_1416_nl;
  mux_1421_nl <= MUX_s_1_2_2(mux_1420_nl, or_1211_nl, fsm_output(9));
  mux_1431_nl <= MUX_s_1_2_2(mux_1430_nl, mux_1421_nl, fsm_output(7));
  mux_1447_nl <= MUX_s_1_2_2(mux_1446_nl, mux_1431_nl, fsm_output(0));
  vec_rsc_0_5_i_wea_d_pff <= NOT mux_1447_nl;
  or_1311_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(5)) OR not_tmp_322;
  or_1309_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_1308_nl <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1307_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1477_nl <= MUX_s_1_2_2(or_1308_nl, or_1307_nl, fsm_output(0));
  mux_1478_nl <= MUX_s_1_2_2(or_1309_nl, mux_1477_nl, fsm_output(4));
  mux_1479_nl <= MUX_s_1_2_2(or_1311_nl, mux_1478_nl, fsm_output(1));
  or_1306_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR not_tmp_322;
  or_1304_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(5)) OR not_tmp_322;
  mux_1474_nl <= MUX_s_1_2_2(or_1306_nl, or_1304_nl, fsm_output(0));
  or_1302_nl <= (fsm_output(0)) OR CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1475_nl <= MUX_s_1_2_2(mux_1474_nl, or_1302_nl, fsm_output(4));
  or_1300_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1476_nl <= MUX_s_1_2_2(mux_1475_nl, or_1300_nl, fsm_output(1));
  mux_1480_nl <= MUX_s_1_2_2(mux_1479_nl, mux_1476_nl, fsm_output(9));
  or_1299_nl <= CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  or_1298_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  mux_1470_nl <= MUX_s_1_2_2(or_1299_nl, or_1298_nl, fsm_output(0));
  or_1297_nl <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  mux_1471_nl <= MUX_s_1_2_2(mux_1470_nl, or_1297_nl, fsm_output(4));
  or_1296_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(4)) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  mux_1472_nl <= MUX_s_1_2_2(mux_1471_nl, or_1296_nl, fsm_output(1));
  nand_346_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0101"))
      AND operator_64_false_slc_operator_64_false_acc_1_60_itm AND (fsm_output(0))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  or_1293_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1292_nl <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1467_nl <= MUX_s_1_2_2(or_1293_nl, or_1292_nl, fsm_output(0));
  mux_1468_nl <= MUX_s_1_2_2(nand_346_nl, mux_1467_nl, fsm_output(4));
  or_1291_nl <= CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1469_nl <= MUX_s_1_2_2(mux_1468_nl, or_1291_nl, fsm_output(1));
  mux_1473_nl <= MUX_s_1_2_2(mux_1472_nl, mux_1469_nl, fsm_output(9));
  mux_1481_nl <= MUX_s_1_2_2(mux_1480_nl, mux_1473_nl, fsm_output(8));
  or_1290_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1288_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1462_nl <= MUX_s_1_2_2(or_1290_nl, or_1288_nl, fsm_output(0));
  or_1286_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR nand_442_cse;
  mux_1463_nl <= MUX_s_1_2_2(mux_1462_nl, or_1286_nl, fsm_output(4));
  or_1284_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1282_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_1459_nl <= MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_1282_nl);
  nor_299_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")));
  mux_1460_nl <= MUX_s_1_2_2(or_1284_nl, mux_1459_nl, nor_299_nl);
  or_1281_nl <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT
      (fsm_output(2)));
  mux_1461_nl <= MUX_s_1_2_2(mux_1460_nl, or_1281_nl, fsm_output(0));
  nand_50_nl <= NOT((fsm_output(4)) AND (NOT mux_1461_nl));
  mux_1464_nl <= MUX_s_1_2_2(mux_1463_nl, nand_50_nl, fsm_output(1));
  or_1279_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT (fsm_output(0)))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1277_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT
      (fsm_output(3))) OR (fsm_output(2));
  mux_1457_nl <= MUX_s_1_2_2(or_1279_nl, or_1277_nl, fsm_output(4));
  or_1276_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3))
      OR (NOT (fsm_output(2)));
  or_1274_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_1272_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  nor_297_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")));
  mux_1453_nl <= MUX_s_1_2_2(nand_437_cse, mux_1112_cse, nor_297_nl);
  nor_296_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")));
  mux_1454_nl <= MUX_s_1_2_2(or_1272_nl, mux_1453_nl, nor_296_nl);
  mux_1455_nl <= MUX_s_1_2_2(or_1274_nl, mux_1454_nl, fsm_output(0));
  mux_1456_nl <= MUX_s_1_2_2(or_1276_nl, mux_1455_nl, fsm_output(4));
  mux_1458_nl <= MUX_s_1_2_2(mux_1457_nl, mux_1456_nl, fsm_output(1));
  mux_1465_nl <= MUX_s_1_2_2(mux_1464_nl, mux_1458_nl, fsm_output(9));
  or_1264_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(4)) OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm)
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1263_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1262_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (COMP_LOOP_acc_10_psp_sva(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_1261_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1448_nl <= MUX_s_1_2_2(or_1262_nl, or_1261_nl, fsm_output(0));
  mux_1449_nl <= MUX_s_1_2_2(or_1263_nl, mux_1448_nl, fsm_output(4));
  mux_1450_nl <= MUX_s_1_2_2(or_1264_nl, mux_1449_nl, fsm_output(1));
  or_1265_nl <= (fsm_output(9)) OR mux_1450_nl;
  mux_1466_nl <= MUX_s_1_2_2(mux_1465_nl, or_1265_nl, fsm_output(8));
  mux_1482_nl <= MUX_s_1_2_2(mux_1481_nl, mux_1466_nl, fsm_output(7));
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= NOT mux_1482_nl;
  nor_693_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_694_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1511_nl <= MUX_s_1_2_2(nor_693_nl, nor_694_nl, fsm_output(4));
  nor_695_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_696_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  mux_1510_nl <= MUX_s_1_2_2(nor_695_nl, nor_696_nl, fsm_output(4));
  mux_1512_nl <= MUX_s_1_2_2(mux_1511_nl, mux_1510_nl, fsm_output(8));
  nand_54_nl <= NOT((fsm_output(1)) AND mux_1512_nl);
  nor_697_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(2)) OR not_tmp_311);
  nor_698_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(2)) OR not_tmp_311);
  mux_1508_nl <= MUX_s_1_2_2(nor_697_nl, nor_698_nl, fsm_output(4));
  nand_53_nl <= NOT((fsm_output(8)) AND mux_1508_nl);
  or_1356_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1354_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1506_nl <= MUX_s_1_2_2(or_1356_nl, or_1354_nl, fsm_output(4));
  or_1353_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0110")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1507_nl <= MUX_s_1_2_2(mux_1506_nl, or_1353_nl, fsm_output(8));
  mux_1509_nl <= MUX_s_1_2_2(nand_53_nl, mux_1507_nl, fsm_output(1));
  mux_1513_nl <= MUX_s_1_2_2(nand_54_nl, mux_1509_nl, fsm_output(9));
  or_1351_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_1350_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1503_nl <= MUX_s_1_2_2(or_1351_nl, or_1350_nl, fsm_output(4));
  or_1348_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1346_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_1502_nl <= MUX_s_1_2_2(or_1348_nl, or_1346_nl, fsm_output(4));
  mux_1504_nl <= MUX_s_1_2_2(mux_1503_nl, mux_1502_nl, fsm_output(8));
  or_1352_nl <= (fsm_output(1)) OR mux_1504_nl;
  or_1343_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1342_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1500_nl <= MUX_s_1_2_2(or_1343_nl, or_1342_nl, fsm_output(4));
  or_1344_nl <= (fsm_output(8)) OR mux_1500_nl;
  or_1341_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR not_tmp_312;
  mux_1501_nl <= MUX_s_1_2_2(or_1344_nl, or_1341_nl, fsm_output(1));
  mux_1505_nl <= MUX_s_1_2_2(or_1352_nl, mux_1501_nl, fsm_output(9));
  mux_1514_nl <= MUX_s_1_2_2(mux_1513_nl, mux_1505_nl, fsm_output(7));
  or_1337_nl <= CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1495_nl <= MUX_s_1_2_2(or_1339_cse, or_1337_nl, fsm_output(8));
  mux_1496_nl <= MUX_s_1_2_2(mux_1495_nl, nand_tmp_52, fsm_output(1));
  or_1336_nl <= (NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1494_nl <= MUX_s_1_2_2(or_1336_nl, nand_tmp_52, fsm_output(1));
  mux_1497_nl <= MUX_s_1_2_2(mux_1496_nl, mux_1494_nl, STAGE_VEC_LOOP_j_sva_9_0(3));
  nor_699_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_700_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1491_nl <= MUX_s_1_2_2(nor_699_nl, nor_700_nl, fsm_output(4));
  nor_701_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_702_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(5))));
  mux_1490_nl <= MUX_s_1_2_2(nor_701_nl, nor_702_nl, fsm_output(4));
  mux_1492_nl <= MUX_s_1_2_2(mux_1491_nl, mux_1490_nl, fsm_output(8));
  nand_51_nl <= NOT((fsm_output(1)) AND mux_1492_nl);
  mux_1498_nl <= MUX_s_1_2_2(mux_1497_nl, nand_51_nl, fsm_output(9));
  or_1325_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("101")) OR not_tmp_312;
  or_1323_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (COMP_LOOP_acc_10_psp_sva(0)) OR (fsm_output(2)) OR not_tmp_311;
  or_1321_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5));
  mux_1486_nl <= MUX_s_1_2_2(or_1323_nl, or_1321_nl, fsm_output(4));
  mux_1487_nl <= MUX_s_1_2_2(or_1325_nl, mux_1486_nl, fsm_output(8));
  or_1319_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1318_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(5));
  mux_1485_nl <= MUX_s_1_2_2(or_1319_nl, or_1318_nl, fsm_output(4));
  or_1320_nl <= (fsm_output(8)) OR mux_1485_nl;
  mux_1488_nl <= MUX_s_1_2_2(mux_1487_nl, or_1320_nl, fsm_output(1));
  or_1316_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_1315_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1483_nl <= MUX_s_1_2_2(or_1316_nl, or_1315_nl, fsm_output(4));
  or_1313_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  mux_1484_nl <= MUX_s_1_2_2(mux_1483_nl, or_1313_nl, fsm_output(8));
  or_1317_nl <= (fsm_output(1)) OR mux_1484_nl;
  mux_1489_nl <= MUX_s_1_2_2(mux_1488_nl, or_1317_nl, fsm_output(9));
  mux_1499_nl <= MUX_s_1_2_2(mux_1498_nl, mux_1489_nl, fsm_output(7));
  mux_1515_nl <= MUX_s_1_2_2(mux_1514_nl, mux_1499_nl, fsm_output(0));
  vec_rsc_0_6_i_wea_d_pff <= NOT mux_1515_nl;
  or_1420_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(5)) OR not_tmp_322;
  or_1418_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_1417_nl <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1416_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1545_nl <= MUX_s_1_2_2(or_1417_nl, or_1416_nl, fsm_output(0));
  mux_1546_nl <= MUX_s_1_2_2(or_1418_nl, mux_1545_nl, fsm_output(4));
  mux_1547_nl <= MUX_s_1_2_2(or_1420_nl, mux_1546_nl, fsm_output(1));
  or_1415_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR not_tmp_322;
  or_1413_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR not_tmp_322;
  mux_1542_nl <= MUX_s_1_2_2(or_1415_nl, or_1413_nl, fsm_output(0));
  or_1411_nl <= (fsm_output(0)) OR CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1543_nl <= MUX_s_1_2_2(mux_1542_nl, or_1411_nl, fsm_output(4));
  or_1409_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1544_nl <= MUX_s_1_2_2(mux_1543_nl, or_1409_nl, fsm_output(1));
  mux_1548_nl <= MUX_s_1_2_2(mux_1547_nl, mux_1544_nl, fsm_output(9));
  or_1408_nl <= CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  or_1407_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  mux_1538_nl <= MUX_s_1_2_2(or_1408_nl, or_1407_nl, fsm_output(0));
  or_1406_nl <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  mux_1539_nl <= MUX_s_1_2_2(mux_1538_nl, or_1406_nl, fsm_output(4));
  or_1405_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(4)) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  mux_1540_nl <= MUX_s_1_2_2(mux_1539_nl, or_1405_nl, fsm_output(1));
  nand_340_nl <= NOT(operator_64_false_slc_operator_64_false_acc_1_60_itm AND (fsm_output(0))
      AND CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0110"))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  or_1402_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1401_nl <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1535_nl <= MUX_s_1_2_2(or_1402_nl, or_1401_nl, fsm_output(0));
  mux_1536_nl <= MUX_s_1_2_2(nand_340_nl, mux_1535_nl, fsm_output(4));
  or_1400_nl <= CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1537_nl <= MUX_s_1_2_2(mux_1536_nl, or_1400_nl, fsm_output(1));
  mux_1541_nl <= MUX_s_1_2_2(mux_1540_nl, mux_1537_nl, fsm_output(9));
  mux_1549_nl <= MUX_s_1_2_2(mux_1548_nl, mux_1541_nl, fsm_output(8));
  or_1399_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1397_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1530_nl <= MUX_s_1_2_2(or_1399_nl, or_1397_nl, fsm_output(0));
  or_1395_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR nand_442_cse;
  mux_1531_nl <= MUX_s_1_2_2(mux_1530_nl, or_1395_nl, fsm_output(4));
  or_1393_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_1527_nl <= MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_1393_nl);
  or_1392_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1390_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"));
  mux_1528_nl <= MUX_s_1_2_2(mux_1527_nl, or_1392_nl, or_1390_nl);
  or_1389_nl <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT
      (fsm_output(2)));
  mux_1529_nl <= MUX_s_1_2_2(mux_1528_nl, or_1389_nl, fsm_output(0));
  nand_56_nl <= NOT((fsm_output(4)) AND (NOT mux_1529_nl));
  mux_1532_nl <= MUX_s_1_2_2(mux_1531_nl, nand_56_nl, fsm_output(1));
  or_1387_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT
      (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1385_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT
      (fsm_output(3))) OR (fsm_output(2));
  mux_1525_nl <= MUX_s_1_2_2(or_1387_nl, or_1385_nl, fsm_output(4));
  or_1384_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3))
      OR (NOT (fsm_output(2)));
  or_1382_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_1375_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"));
  mux_1521_nl <= MUX_s_1_2_2(mux_1112_cse, nand_437_cse, or_1375_nl);
  or_1374_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_1372_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"));
  mux_1522_nl <= MUX_s_1_2_2(mux_1521_nl, or_1374_nl, or_1372_nl);
  mux_1523_nl <= MUX_s_1_2_2(or_1382_nl, mux_1522_nl, fsm_output(0));
  mux_1524_nl <= MUX_s_1_2_2(or_1384_nl, mux_1523_nl, fsm_output(4));
  mux_1526_nl <= MUX_s_1_2_2(mux_1525_nl, mux_1524_nl, fsm_output(1));
  mux_1533_nl <= MUX_s_1_2_2(mux_1532_nl, mux_1526_nl, fsm_output(9));
  or_1370_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(4)) OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm)
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1369_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1368_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (COMP_LOOP_acc_10_psp_sva(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_1367_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1516_nl <= MUX_s_1_2_2(or_1368_nl, or_1367_nl, fsm_output(0));
  mux_1517_nl <= MUX_s_1_2_2(or_1369_nl, mux_1516_nl, fsm_output(4));
  mux_1518_nl <= MUX_s_1_2_2(or_1370_nl, mux_1517_nl, fsm_output(1));
  or_1371_nl <= (fsm_output(9)) OR mux_1518_nl;
  mux_1534_nl <= MUX_s_1_2_2(mux_1533_nl, or_1371_nl, fsm_output(8));
  mux_1550_nl <= MUX_s_1_2_2(mux_1549_nl, mux_1534_nl, fsm_output(7));
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= NOT mux_1550_nl;
  nor_681_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_682_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1579_nl <= MUX_s_1_2_2(nor_681_nl, nor_682_nl, fsm_output(4));
  and_773_nl <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  and_779_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  mux_1578_nl <= MUX_s_1_2_2(and_773_nl, and_779_nl, fsm_output(4));
  mux_1580_nl <= MUX_s_1_2_2(mux_1579_nl, mux_1578_nl, fsm_output(8));
  nand_60_nl <= NOT((fsm_output(1)) AND mux_1580_nl);
  nor_685_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(2)) OR not_tmp_311);
  nor_686_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(2)) OR not_tmp_311);
  mux_1576_nl <= MUX_s_1_2_2(nor_685_nl, nor_686_nl, fsm_output(4));
  nand_59_nl <= NOT((fsm_output(8)) AND mux_1576_nl);
  or_1465_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1463_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1574_nl <= MUX_s_1_2_2(or_1465_nl, or_1463_nl, fsm_output(4));
  or_1462_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0111")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1575_nl <= MUX_s_1_2_2(mux_1574_nl, or_1462_nl, fsm_output(8));
  mux_1577_nl <= MUX_s_1_2_2(nand_59_nl, mux_1575_nl, fsm_output(1));
  mux_1581_nl <= MUX_s_1_2_2(nand_60_nl, mux_1577_nl, fsm_output(9));
  nand_331_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(5))));
  nand_472_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5)));
  mux_1571_nl <= MUX_s_1_2_2(nand_331_nl, nand_472_nl, fsm_output(4));
  or_1457_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1455_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_1570_nl <= MUX_s_1_2_2(or_1457_nl, or_1455_nl, fsm_output(4));
  mux_1572_nl <= MUX_s_1_2_2(mux_1571_nl, mux_1570_nl, fsm_output(8));
  or_1461_nl <= (fsm_output(1)) OR mux_1572_nl;
  or_1452_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1451_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1568_nl <= MUX_s_1_2_2(or_1452_nl, or_1451_nl, fsm_output(4));
  or_1453_nl <= (fsm_output(8)) OR mux_1568_nl;
  or_1450_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR not_tmp_312;
  mux_1569_nl <= MUX_s_1_2_2(or_1453_nl, or_1450_nl, fsm_output(1));
  mux_1573_nl <= MUX_s_1_2_2(or_1461_nl, mux_1569_nl, fsm_output(9));
  mux_1582_nl <= MUX_s_1_2_2(mux_1581_nl, mux_1573_nl, fsm_output(7));
  or_1446_nl <= CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1563_nl <= MUX_s_1_2_2(or_1448_cse, or_1446_nl, fsm_output(8));
  mux_1564_nl <= MUX_s_1_2_2(mux_1563_nl, nand_tmp_58, fsm_output(1));
  or_1445_nl <= (NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1562_nl <= MUX_s_1_2_2(or_1445_nl, nand_tmp_58, fsm_output(1));
  mux_1565_nl <= MUX_s_1_2_2(mux_1564_nl, mux_1562_nl, STAGE_VEC_LOOP_j_sva_9_0(3));
  nor_687_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_688_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1559_nl <= MUX_s_1_2_2(nor_687_nl, nor_688_nl, fsm_output(4));
  and_789_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  and_790_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))
      AND (STAGE_VEC_LOOP_j_sva_9_0(0)) AND (fsm_output(2)) AND (fsm_output(3)) AND
      (NOT (fsm_output(6))) AND (fsm_output(5));
  mux_1558_nl <= MUX_s_1_2_2(and_789_nl, and_790_nl, fsm_output(4));
  mux_1560_nl <= MUX_s_1_2_2(mux_1559_nl, mux_1558_nl, fsm_output(8));
  nand_57_nl <= NOT((fsm_output(1)) AND mux_1560_nl);
  mux_1566_nl <= MUX_s_1_2_2(mux_1565_nl, nand_57_nl, fsm_output(9));
  or_1434_nl <= (NOT(CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("101")))) OR not_tmp_312;
  or_1432_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (COMP_LOOP_acc_10_psp_sva(0)) OR (fsm_output(2)) OR not_tmp_311;
  or_1430_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5));
  mux_1554_nl <= MUX_s_1_2_2(or_1432_nl, or_1430_nl, fsm_output(4));
  mux_1555_nl <= MUX_s_1_2_2(or_1434_nl, mux_1554_nl, fsm_output(8));
  or_1428_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1427_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(2)) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1553_nl <= MUX_s_1_2_2(or_1428_nl, or_1427_nl, fsm_output(4));
  or_1429_nl <= (fsm_output(8)) OR mux_1553_nl;
  mux_1556_nl <= MUX_s_1_2_2(mux_1555_nl, or_1429_nl, fsm_output(1));
  nand_336_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(5))));
  nand_453_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5)));
  mux_1551_nl <= MUX_s_1_2_2(nand_336_nl, nand_453_nl, fsm_output(4));
  or_1422_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0111")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  mux_1552_nl <= MUX_s_1_2_2(mux_1551_nl, or_1422_nl, fsm_output(8));
  or_1426_nl <= (fsm_output(1)) OR mux_1552_nl;
  mux_1557_nl <= MUX_s_1_2_2(mux_1556_nl, or_1426_nl, fsm_output(9));
  mux_1567_nl <= MUX_s_1_2_2(mux_1566_nl, mux_1557_nl, fsm_output(7));
  mux_1583_nl <= MUX_s_1_2_2(mux_1582_nl, mux_1567_nl, fsm_output(0));
  vec_rsc_0_7_i_wea_d_pff <= NOT mux_1583_nl;
  or_1526_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(5)) OR not_tmp_322;
  nand_317_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(0)) AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      AND (NOT (fsm_output(5))) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT
      (fsm_output(2))));
  or_1523_nl <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1522_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1613_nl <= MUX_s_1_2_2(or_1523_nl, or_1522_nl, fsm_output(0));
  mux_1614_nl <= MUX_s_1_2_2(nand_317_nl, mux_1613_nl, fsm_output(4));
  mux_1615_nl <= MUX_s_1_2_2(or_1526_nl, mux_1614_nl, fsm_output(1));
  or_1521_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR not_tmp_322;
  or_1519_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR not_tmp_322;
  mux_1610_nl <= MUX_s_1_2_2(or_1521_nl, or_1519_nl, fsm_output(0));
  or_1517_nl <= (fsm_output(0)) OR CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1611_nl <= MUX_s_1_2_2(mux_1610_nl, or_1517_nl, fsm_output(4));
  or_1515_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1612_nl <= MUX_s_1_2_2(mux_1611_nl, or_1515_nl, fsm_output(1));
  mux_1616_nl <= MUX_s_1_2_2(mux_1615_nl, mux_1612_nl, fsm_output(9));
  nand_318_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))
      AND (STAGE_VEC_LOOP_j_sva_9_0(0)) AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  nand_319_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  mux_1606_nl <= MUX_s_1_2_2(nand_318_nl, nand_319_nl, fsm_output(0));
  or_1512_nl <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  mux_1607_nl <= MUX_s_1_2_2(mux_1606_nl, or_1512_nl, fsm_output(4));
  or_1511_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(4)) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  mux_1608_nl <= MUX_s_1_2_2(mux_1607_nl, or_1511_nl, fsm_output(1));
  nand_320_nl <= NOT(operator_64_false_slc_operator_64_false_acc_1_60_itm AND (fsm_output(0))
      AND CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  or_1508_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1507_nl <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1603_nl <= MUX_s_1_2_2(or_1508_nl, or_1507_nl, fsm_output(0));
  mux_1604_nl <= MUX_s_1_2_2(nand_320_nl, mux_1603_nl, fsm_output(4));
  or_1506_nl <= CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1605_nl <= MUX_s_1_2_2(mux_1604_nl, or_1506_nl, fsm_output(1));
  mux_1609_nl <= MUX_s_1_2_2(mux_1608_nl, mux_1605_nl, fsm_output(9));
  mux_1617_nl <= MUX_s_1_2_2(mux_1616_nl, mux_1609_nl, fsm_output(8));
  or_1505_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1503_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1598_nl <= MUX_s_1_2_2(or_1505_nl, or_1503_nl, fsm_output(0));
  or_1501_nl <= (NOT(operator_64_false_slc_operator_64_false_acc_1_60_itm AND CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("0111")) AND (fsm_output(0)) AND (fsm_output(5))
      AND (NOT (fsm_output(6))))) OR nand_442_cse;
  mux_1599_nl <= MUX_s_1_2_2(mux_1598_nl, or_1501_nl, fsm_output(4));
  nand_467_nl <= NOT(CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm AND (fsm_output(5))
      AND (fsm_output(6)) AND (NOT (fsm_output(3))) AND (fsm_output(2)));
  nand_323_nl <= NOT(CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_1595_nl <= MUX_s_1_2_2(nand_tmp_19, or_tmp_669, nand_323_nl);
  and_546_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
  mux_1596_nl <= MUX_s_1_2_2(nand_467_nl, mux_1595_nl, and_546_nl);
  nand_463_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (NOT (fsm_output(3))) AND (fsm_output(2)));
  mux_1597_nl <= MUX_s_1_2_2(mux_1596_nl, nand_463_nl, fsm_output(0));
  nand_62_nl <= NOT((fsm_output(4)) AND (NOT mux_1597_nl));
  mux_1600_nl <= MUX_s_1_2_2(mux_1599_nl, nand_62_nl, fsm_output(1));
  or_1494_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT
      (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1492_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT
      (fsm_output(3))) OR (fsm_output(2));
  mux_1593_nl <= MUX_s_1_2_2(or_1494_nl, or_1492_nl, fsm_output(4));
  or_1491_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3))
      OR (NOT (fsm_output(2)));
  or_1489_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm AND CONV_SL_1_1(fsm_output(6
      DOWNTO 5)=STD_LOGIC_VECTOR'("01")))) OR nand_442_cse;
  or_1487_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  and_547_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
  mux_1589_nl <= MUX_s_1_2_2(nand_437_cse, mux_1112_cse, and_547_nl);
  and_548_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
  mux_1590_nl <= MUX_s_1_2_2(or_1487_nl, mux_1589_nl, and_548_nl);
  mux_1591_nl <= MUX_s_1_2_2(or_1489_nl, mux_1590_nl, fsm_output(0));
  mux_1592_nl <= MUX_s_1_2_2(or_1491_nl, mux_1591_nl, fsm_output(4));
  mux_1594_nl <= MUX_s_1_2_2(mux_1593_nl, mux_1592_nl, fsm_output(1));
  mux_1601_nl <= MUX_s_1_2_2(mux_1600_nl, mux_1594_nl, fsm_output(9));
  or_1479_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(4)) OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm)
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1478_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1477_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (COMP_LOOP_acc_10_psp_sva(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_1476_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1584_nl <= MUX_s_1_2_2(or_1477_nl, or_1476_nl, fsm_output(0));
  mux_1585_nl <= MUX_s_1_2_2(or_1478_nl, mux_1584_nl, fsm_output(4));
  mux_1586_nl <= MUX_s_1_2_2(or_1479_nl, mux_1585_nl, fsm_output(1));
  or_1480_nl <= (fsm_output(9)) OR mux_1586_nl;
  mux_1602_nl <= MUX_s_1_2_2(mux_1601_nl, or_1480_nl, fsm_output(8));
  mux_1618_nl <= MUX_s_1_2_2(mux_1617_nl, mux_1602_nl, fsm_output(7));
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= NOT mux_1618_nl;
  nor_669_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_670_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1647_nl <= MUX_s_1_2_2(nor_669_nl, nor_670_nl, fsm_output(4));
  nor_671_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_672_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  mux_1646_nl <= MUX_s_1_2_2(nor_671_nl, nor_672_nl, fsm_output(4));
  mux_1648_nl <= MUX_s_1_2_2(mux_1647_nl, mux_1646_nl, fsm_output(8));
  nand_66_nl <= NOT((fsm_output(1)) AND mux_1648_nl);
  nor_673_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(2)) OR not_tmp_311);
  nor_674_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(2)) OR not_tmp_311);
  mux_1644_nl <= MUX_s_1_2_2(nor_673_nl, nor_674_nl, fsm_output(4));
  nand_65_nl <= NOT((fsm_output(8)) AND mux_1644_nl);
  or_1571_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1569_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1642_nl <= MUX_s_1_2_2(or_1571_nl, or_1569_nl, fsm_output(4));
  or_1568_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1000")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1643_nl <= MUX_s_1_2_2(mux_1642_nl, or_1568_nl, fsm_output(8));
  mux_1645_nl <= MUX_s_1_2_2(nand_65_nl, mux_1643_nl, fsm_output(1));
  mux_1649_nl <= MUX_s_1_2_2(nand_66_nl, mux_1645_nl, fsm_output(9));
  or_1566_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_1565_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1639_nl <= MUX_s_1_2_2(or_1566_nl, or_1565_nl, fsm_output(4));
  or_1563_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1561_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_1638_nl <= MUX_s_1_2_2(or_1563_nl, or_1561_nl, fsm_output(4));
  mux_1640_nl <= MUX_s_1_2_2(mux_1639_nl, mux_1638_nl, fsm_output(8));
  or_1567_nl <= (fsm_output(1)) OR mux_1640_nl;
  or_1558_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1557_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1636_nl <= MUX_s_1_2_2(or_1558_nl, or_1557_nl, fsm_output(4));
  or_1559_nl <= (fsm_output(8)) OR mux_1636_nl;
  or_1556_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR not_tmp_312;
  mux_1637_nl <= MUX_s_1_2_2(or_1559_nl, or_1556_nl, fsm_output(1));
  mux_1641_nl <= MUX_s_1_2_2(or_1567_nl, mux_1637_nl, fsm_output(9));
  mux_1650_nl <= MUX_s_1_2_2(mux_1649_nl, mux_1641_nl, fsm_output(7));
  or_1554_nl <= (NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1632_nl <= MUX_s_1_2_2(or_1554_nl, nand_tmp_64, fsm_output(1));
  or_1551_nl <= CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1630_nl <= MUX_s_1_2_2(or_694_cse, or_1551_nl, fsm_output(8));
  mux_1631_nl <= MUX_s_1_2_2(mux_1630_nl, nand_tmp_64, fsm_output(1));
  mux_1633_nl <= MUX_s_1_2_2(mux_1632_nl, mux_1631_nl, STAGE_VEC_LOOP_j_sva_9_0(3));
  nor_675_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_676_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1627_nl <= MUX_s_1_2_2(nor_675_nl, nor_676_nl, fsm_output(4));
  nor_677_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_678_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(5))));
  mux_1626_nl <= MUX_s_1_2_2(nor_677_nl, nor_678_nl, fsm_output(4));
  mux_1628_nl <= MUX_s_1_2_2(mux_1627_nl, mux_1626_nl, fsm_output(8));
  nand_63_nl <= NOT((fsm_output(1)) AND mux_1628_nl);
  mux_1634_nl <= MUX_s_1_2_2(mux_1633_nl, nand_63_nl, fsm_output(9));
  or_1540_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("101")) OR not_tmp_312;
  or_1538_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (COMP_LOOP_acc_10_psp_sva(0))) OR (fsm_output(2)) OR not_tmp_311;
  or_1536_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5));
  mux_1622_nl <= MUX_s_1_2_2(or_1538_nl, or_1536_nl, fsm_output(4));
  mux_1623_nl <= MUX_s_1_2_2(or_1540_nl, mux_1622_nl, fsm_output(8));
  or_1534_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1533_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(5));
  mux_1621_nl <= MUX_s_1_2_2(or_1534_nl, or_1533_nl, fsm_output(4));
  or_1535_nl <= (fsm_output(8)) OR mux_1621_nl;
  mux_1624_nl <= MUX_s_1_2_2(mux_1623_nl, or_1535_nl, fsm_output(1));
  or_1531_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_1530_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1619_nl <= MUX_s_1_2_2(or_1531_nl, or_1530_nl, fsm_output(4));
  or_1528_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  mux_1620_nl <= MUX_s_1_2_2(mux_1619_nl, or_1528_nl, fsm_output(8));
  or_1532_nl <= (fsm_output(1)) OR mux_1620_nl;
  mux_1625_nl <= MUX_s_1_2_2(mux_1624_nl, or_1532_nl, fsm_output(9));
  mux_1635_nl <= MUX_s_1_2_2(mux_1634_nl, mux_1625_nl, fsm_output(7));
  mux_1651_nl <= MUX_s_1_2_2(mux_1650_nl, mux_1635_nl, fsm_output(0));
  vec_rsc_0_8_i_wea_d_pff <= NOT mux_1651_nl;
  or_1635_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(5)) OR not_tmp_322;
  or_1633_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_1632_nl <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1631_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1681_nl <= MUX_s_1_2_2(or_1632_nl, or_1631_nl, fsm_output(0));
  mux_1682_nl <= MUX_s_1_2_2(or_1633_nl, mux_1681_nl, fsm_output(4));
  mux_1683_nl <= MUX_s_1_2_2(or_1635_nl, mux_1682_nl, fsm_output(1));
  or_1630_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR not_tmp_322;
  or_1628_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR not_tmp_322;
  mux_1678_nl <= MUX_s_1_2_2(or_1630_nl, or_1628_nl, fsm_output(0));
  or_1626_nl <= (fsm_output(0)) OR CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1679_nl <= MUX_s_1_2_2(mux_1678_nl, or_1626_nl, fsm_output(4));
  or_1624_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1680_nl <= MUX_s_1_2_2(mux_1679_nl, or_1624_nl, fsm_output(1));
  mux_1684_nl <= MUX_s_1_2_2(mux_1683_nl, mux_1680_nl, fsm_output(9));
  or_1623_nl <= CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  or_1622_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  mux_1674_nl <= MUX_s_1_2_2(or_1623_nl, or_1622_nl, fsm_output(0));
  or_1621_nl <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  mux_1675_nl <= MUX_s_1_2_2(mux_1674_nl, or_1621_nl, fsm_output(4));
  or_1620_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(4)) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  mux_1676_nl <= MUX_s_1_2_2(mux_1675_nl, or_1620_nl, fsm_output(1));
  or_1618_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT (fsm_output(0)))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  or_1617_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1616_nl <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1671_nl <= MUX_s_1_2_2(or_1617_nl, or_1616_nl, fsm_output(0));
  mux_1672_nl <= MUX_s_1_2_2(or_1618_nl, mux_1671_nl, fsm_output(4));
  or_1615_nl <= CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1673_nl <= MUX_s_1_2_2(mux_1672_nl, or_1615_nl, fsm_output(1));
  mux_1677_nl <= MUX_s_1_2_2(mux_1676_nl, mux_1673_nl, fsm_output(9));
  mux_1685_nl <= MUX_s_1_2_2(mux_1684_nl, mux_1677_nl, fsm_output(8));
  or_1614_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1612_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1666_nl <= MUX_s_1_2_2(or_1614_nl, or_1612_nl, fsm_output(0));
  or_1610_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR nand_442_cse;
  mux_1667_nl <= MUX_s_1_2_2(mux_1666_nl, or_1610_nl, fsm_output(4));
  or_1608_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_1663_nl <= MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_1608_nl);
  or_1607_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1605_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"));
  mux_1664_nl <= MUX_s_1_2_2(mux_1663_nl, or_1607_nl, or_1605_nl);
  or_1604_nl <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT
      (fsm_output(2)));
  mux_1665_nl <= MUX_s_1_2_2(mux_1664_nl, or_1604_nl, fsm_output(0));
  nand_68_nl <= NOT((fsm_output(4)) AND (NOT mux_1665_nl));
  mux_1668_nl <= MUX_s_1_2_2(mux_1667_nl, nand_68_nl, fsm_output(1));
  or_1602_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT (fsm_output(0)))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1600_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT
      (fsm_output(3))) OR (fsm_output(2));
  mux_1661_nl <= MUX_s_1_2_2(or_1602_nl, or_1600_nl, fsm_output(4));
  or_1599_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3))
      OR (NOT (fsm_output(2)));
  or_1597_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_1590_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"));
  mux_1657_nl <= MUX_s_1_2_2(mux_1112_cse, nand_437_cse, or_1590_nl);
  or_1589_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_1587_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"));
  mux_1658_nl <= MUX_s_1_2_2(mux_1657_nl, or_1589_nl, or_1587_nl);
  mux_1659_nl <= MUX_s_1_2_2(or_1597_nl, mux_1658_nl, fsm_output(0));
  mux_1660_nl <= MUX_s_1_2_2(or_1599_nl, mux_1659_nl, fsm_output(4));
  mux_1662_nl <= MUX_s_1_2_2(mux_1661_nl, mux_1660_nl, fsm_output(1));
  mux_1669_nl <= MUX_s_1_2_2(mux_1668_nl, mux_1662_nl, fsm_output(9));
  or_1585_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(4)) OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm)
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1584_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1583_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (COMP_LOOP_acc_10_psp_sva(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_1582_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1652_nl <= MUX_s_1_2_2(or_1583_nl, or_1582_nl, fsm_output(0));
  mux_1653_nl <= MUX_s_1_2_2(or_1584_nl, mux_1652_nl, fsm_output(4));
  mux_1654_nl <= MUX_s_1_2_2(or_1585_nl, mux_1653_nl, fsm_output(1));
  or_1586_nl <= (fsm_output(9)) OR mux_1654_nl;
  mux_1670_nl <= MUX_s_1_2_2(mux_1669_nl, or_1586_nl, fsm_output(8));
  mux_1686_nl <= MUX_s_1_2_2(mux_1685_nl, mux_1670_nl, fsm_output(7));
  vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= NOT mux_1686_nl;
  nor_657_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_658_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1715_nl <= MUX_s_1_2_2(nor_657_nl, nor_658_nl, fsm_output(4));
  nor_659_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_660_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  mux_1714_nl <= MUX_s_1_2_2(nor_659_nl, nor_660_nl, fsm_output(4));
  mux_1716_nl <= MUX_s_1_2_2(mux_1715_nl, mux_1714_nl, fsm_output(8));
  nand_72_nl <= NOT((fsm_output(1)) AND mux_1716_nl);
  nor_661_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(2)) OR not_tmp_311);
  nor_662_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(2)) OR not_tmp_311);
  mux_1712_nl <= MUX_s_1_2_2(nor_661_nl, nor_662_nl, fsm_output(4));
  nand_71_nl <= NOT((fsm_output(8)) AND mux_1712_nl);
  or_1680_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1678_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1710_nl <= MUX_s_1_2_2(or_1680_nl, or_1678_nl, fsm_output(4));
  or_1677_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1001")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1711_nl <= MUX_s_1_2_2(mux_1710_nl, or_1677_nl, fsm_output(8));
  mux_1713_nl <= MUX_s_1_2_2(nand_71_nl, mux_1711_nl, fsm_output(1));
  mux_1717_nl <= MUX_s_1_2_2(nand_72_nl, mux_1713_nl, fsm_output(9));
  or_1675_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_1674_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1707_nl <= MUX_s_1_2_2(or_1675_nl, or_1674_nl, fsm_output(4));
  or_1672_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1670_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_1706_nl <= MUX_s_1_2_2(or_1672_nl, or_1670_nl, fsm_output(4));
  mux_1708_nl <= MUX_s_1_2_2(mux_1707_nl, mux_1706_nl, fsm_output(8));
  or_1676_nl <= (fsm_output(1)) OR mux_1708_nl;
  or_1667_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1666_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1704_nl <= MUX_s_1_2_2(or_1667_nl, or_1666_nl, fsm_output(4));
  or_1668_nl <= (fsm_output(8)) OR mux_1704_nl;
  or_1665_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR not_tmp_312;
  mux_1705_nl <= MUX_s_1_2_2(or_1668_nl, or_1665_nl, fsm_output(1));
  mux_1709_nl <= MUX_s_1_2_2(or_1676_nl, mux_1705_nl, fsm_output(9));
  mux_1718_nl <= MUX_s_1_2_2(mux_1717_nl, mux_1709_nl, fsm_output(7));
  or_1663_nl <= (NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1700_nl <= MUX_s_1_2_2(or_1663_nl, nand_tmp_70, fsm_output(1));
  or_1660_nl <= CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1698_nl <= MUX_s_1_2_2(or_803_cse, or_1660_nl, fsm_output(8));
  mux_1699_nl <= MUX_s_1_2_2(mux_1698_nl, nand_tmp_70, fsm_output(1));
  mux_1701_nl <= MUX_s_1_2_2(mux_1700_nl, mux_1699_nl, STAGE_VEC_LOOP_j_sva_9_0(3));
  nor_663_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_664_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1695_nl <= MUX_s_1_2_2(nor_663_nl, nor_664_nl, fsm_output(4));
  nor_665_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_666_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(5))));
  mux_1694_nl <= MUX_s_1_2_2(nor_665_nl, nor_666_nl, fsm_output(4));
  mux_1696_nl <= MUX_s_1_2_2(mux_1695_nl, mux_1694_nl, fsm_output(8));
  nand_69_nl <= NOT((fsm_output(1)) AND mux_1696_nl);
  mux_1702_nl <= MUX_s_1_2_2(mux_1701_nl, nand_69_nl, fsm_output(9));
  or_1649_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("101")) OR not_tmp_312;
  or_1647_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (COMP_LOOP_acc_10_psp_sva(0))) OR (fsm_output(2)) OR not_tmp_311;
  or_1645_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5));
  mux_1690_nl <= MUX_s_1_2_2(or_1647_nl, or_1645_nl, fsm_output(4));
  mux_1691_nl <= MUX_s_1_2_2(or_1649_nl, mux_1690_nl, fsm_output(8));
  or_1643_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1642_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(2)) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1689_nl <= MUX_s_1_2_2(or_1643_nl, or_1642_nl, fsm_output(4));
  or_1644_nl <= (fsm_output(8)) OR mux_1689_nl;
  mux_1692_nl <= MUX_s_1_2_2(mux_1691_nl, or_1644_nl, fsm_output(1));
  or_1640_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_1639_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1687_nl <= MUX_s_1_2_2(or_1640_nl, or_1639_nl, fsm_output(4));
  or_1637_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  mux_1688_nl <= MUX_s_1_2_2(mux_1687_nl, or_1637_nl, fsm_output(8));
  or_1641_nl <= (fsm_output(1)) OR mux_1688_nl;
  mux_1693_nl <= MUX_s_1_2_2(mux_1692_nl, or_1641_nl, fsm_output(9));
  mux_1703_nl <= MUX_s_1_2_2(mux_1702_nl, mux_1693_nl, fsm_output(7));
  mux_1719_nl <= MUX_s_1_2_2(mux_1718_nl, mux_1703_nl, fsm_output(0));
  vec_rsc_0_9_i_wea_d_pff <= NOT mux_1719_nl;
  or_1741_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(5)) OR not_tmp_322;
  or_1739_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_1738_nl <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1737_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1749_nl <= MUX_s_1_2_2(or_1738_nl, or_1737_nl, fsm_output(0));
  mux_1750_nl <= MUX_s_1_2_2(or_1739_nl, mux_1749_nl, fsm_output(4));
  mux_1751_nl <= MUX_s_1_2_2(or_1741_nl, mux_1750_nl, fsm_output(1));
  or_1736_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR not_tmp_322;
  or_1734_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(5)) OR not_tmp_322;
  mux_1746_nl <= MUX_s_1_2_2(or_1736_nl, or_1734_nl, fsm_output(0));
  or_1732_nl <= (fsm_output(0)) OR CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1747_nl <= MUX_s_1_2_2(mux_1746_nl, or_1732_nl, fsm_output(4));
  or_1730_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1748_nl <= MUX_s_1_2_2(mux_1747_nl, or_1730_nl, fsm_output(1));
  mux_1752_nl <= MUX_s_1_2_2(mux_1751_nl, mux_1748_nl, fsm_output(9));
  or_1729_nl <= CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  or_1728_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  mux_1742_nl <= MUX_s_1_2_2(or_1729_nl, or_1728_nl, fsm_output(0));
  or_1727_nl <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  mux_1743_nl <= MUX_s_1_2_2(mux_1742_nl, or_1727_nl, fsm_output(4));
  or_1726_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(4)) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  mux_1744_nl <= MUX_s_1_2_2(mux_1743_nl, or_1726_nl, fsm_output(1));
  nand_306_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1001"))
      AND operator_64_false_slc_operator_64_false_acc_1_60_itm AND (fsm_output(0))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  or_1723_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1722_nl <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1739_nl <= MUX_s_1_2_2(or_1723_nl, or_1722_nl, fsm_output(0));
  mux_1740_nl <= MUX_s_1_2_2(nand_306_nl, mux_1739_nl, fsm_output(4));
  or_1721_nl <= CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1741_nl <= MUX_s_1_2_2(mux_1740_nl, or_1721_nl, fsm_output(1));
  mux_1745_nl <= MUX_s_1_2_2(mux_1744_nl, mux_1741_nl, fsm_output(9));
  mux_1753_nl <= MUX_s_1_2_2(mux_1752_nl, mux_1745_nl, fsm_output(8));
  or_1720_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1718_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1734_nl <= MUX_s_1_2_2(or_1720_nl, or_1718_nl, fsm_output(0));
  or_1716_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR nand_442_cse;
  mux_1735_nl <= MUX_s_1_2_2(mux_1734_nl, or_1716_nl, fsm_output(4));
  or_1714_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1712_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_1731_nl <= MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_1712_nl);
  nor_321_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")));
  mux_1732_nl <= MUX_s_1_2_2(or_1714_nl, mux_1731_nl, nor_321_nl);
  or_1711_nl <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT
      (fsm_output(2)));
  mux_1733_nl <= MUX_s_1_2_2(mux_1732_nl, or_1711_nl, fsm_output(0));
  nand_74_nl <= NOT((fsm_output(4)) AND (NOT mux_1733_nl));
  mux_1736_nl <= MUX_s_1_2_2(mux_1735_nl, nand_74_nl, fsm_output(1));
  or_1709_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT (fsm_output(0)))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1707_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT
      (fsm_output(3))) OR (fsm_output(2));
  mux_1729_nl <= MUX_s_1_2_2(or_1709_nl, or_1707_nl, fsm_output(4));
  or_1706_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3))
      OR (NOT (fsm_output(2)));
  or_1704_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_1702_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  nor_319_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")));
  mux_1725_nl <= MUX_s_1_2_2(nand_437_cse, mux_1112_cse, nor_319_nl);
  nor_318_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")));
  mux_1726_nl <= MUX_s_1_2_2(or_1702_nl, mux_1725_nl, nor_318_nl);
  mux_1727_nl <= MUX_s_1_2_2(or_1704_nl, mux_1726_nl, fsm_output(0));
  mux_1728_nl <= MUX_s_1_2_2(or_1706_nl, mux_1727_nl, fsm_output(4));
  mux_1730_nl <= MUX_s_1_2_2(mux_1729_nl, mux_1728_nl, fsm_output(1));
  mux_1737_nl <= MUX_s_1_2_2(mux_1736_nl, mux_1730_nl, fsm_output(9));
  or_1694_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(4)) OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm)
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1693_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1692_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (COMP_LOOP_acc_10_psp_sva(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_1691_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1720_nl <= MUX_s_1_2_2(or_1692_nl, or_1691_nl, fsm_output(0));
  mux_1721_nl <= MUX_s_1_2_2(or_1693_nl, mux_1720_nl, fsm_output(4));
  mux_1722_nl <= MUX_s_1_2_2(or_1694_nl, mux_1721_nl, fsm_output(1));
  or_1695_nl <= (fsm_output(9)) OR mux_1722_nl;
  mux_1738_nl <= MUX_s_1_2_2(mux_1737_nl, or_1695_nl, fsm_output(8));
  mux_1754_nl <= MUX_s_1_2_2(mux_1753_nl, mux_1738_nl, fsm_output(7));
  vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= NOT mux_1754_nl;
  nor_645_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_646_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1783_nl <= MUX_s_1_2_2(nor_645_nl, nor_646_nl, fsm_output(4));
  nor_647_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_648_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  mux_1782_nl <= MUX_s_1_2_2(nor_647_nl, nor_648_nl, fsm_output(4));
  mux_1784_nl <= MUX_s_1_2_2(mux_1783_nl, mux_1782_nl, fsm_output(8));
  nand_78_nl <= NOT((fsm_output(1)) AND mux_1784_nl);
  nor_649_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(2)) OR not_tmp_311);
  nor_650_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(2)) OR not_tmp_311);
  mux_1780_nl <= MUX_s_1_2_2(nor_649_nl, nor_650_nl, fsm_output(4));
  nand_77_nl <= NOT((fsm_output(8)) AND mux_1780_nl);
  or_1786_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1784_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1778_nl <= MUX_s_1_2_2(or_1786_nl, or_1784_nl, fsm_output(4));
  or_1783_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1010")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1779_nl <= MUX_s_1_2_2(mux_1778_nl, or_1783_nl, fsm_output(8));
  mux_1781_nl <= MUX_s_1_2_2(nand_77_nl, mux_1779_nl, fsm_output(1));
  mux_1785_nl <= MUX_s_1_2_2(nand_78_nl, mux_1781_nl, fsm_output(9));
  or_1781_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_1780_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1775_nl <= MUX_s_1_2_2(or_1781_nl, or_1780_nl, fsm_output(4));
  or_1778_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1776_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_1774_nl <= MUX_s_1_2_2(or_1778_nl, or_1776_nl, fsm_output(4));
  mux_1776_nl <= MUX_s_1_2_2(mux_1775_nl, mux_1774_nl, fsm_output(8));
  or_1782_nl <= (fsm_output(1)) OR mux_1776_nl;
  or_1773_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1772_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1772_nl <= MUX_s_1_2_2(or_1773_nl, or_1772_nl, fsm_output(4));
  or_1774_nl <= (fsm_output(8)) OR mux_1772_nl;
  or_1771_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR not_tmp_312;
  mux_1773_nl <= MUX_s_1_2_2(or_1774_nl, or_1771_nl, fsm_output(1));
  mux_1777_nl <= MUX_s_1_2_2(or_1782_nl, mux_1773_nl, fsm_output(9));
  mux_1786_nl <= MUX_s_1_2_2(mux_1785_nl, mux_1777_nl, fsm_output(7));
  or_1769_nl <= (NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1768_nl <= MUX_s_1_2_2(or_1769_nl, nand_tmp_76, fsm_output(1));
  or_1766_nl <= CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1766_nl <= MUX_s_1_2_2(or_909_cse, or_1766_nl, fsm_output(8));
  mux_1767_nl <= MUX_s_1_2_2(mux_1766_nl, nand_tmp_76, fsm_output(1));
  mux_1769_nl <= MUX_s_1_2_2(mux_1768_nl, mux_1767_nl, STAGE_VEC_LOOP_j_sva_9_0(3));
  nor_651_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_652_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1763_nl <= MUX_s_1_2_2(nor_651_nl, nor_652_nl, fsm_output(4));
  nor_653_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_654_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(5))));
  mux_1762_nl <= MUX_s_1_2_2(nor_653_nl, nor_654_nl, fsm_output(4));
  mux_1764_nl <= MUX_s_1_2_2(mux_1763_nl, mux_1762_nl, fsm_output(8));
  nand_75_nl <= NOT((fsm_output(1)) AND mux_1764_nl);
  mux_1770_nl <= MUX_s_1_2_2(mux_1769_nl, nand_75_nl, fsm_output(9));
  or_1755_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("101")) OR not_tmp_312;
  or_1753_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (COMP_LOOP_acc_10_psp_sva(0))) OR (fsm_output(2)) OR not_tmp_311;
  or_1751_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5));
  mux_1758_nl <= MUX_s_1_2_2(or_1753_nl, or_1751_nl, fsm_output(4));
  mux_1759_nl <= MUX_s_1_2_2(or_1755_nl, mux_1758_nl, fsm_output(8));
  or_1749_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1748_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(5));
  mux_1757_nl <= MUX_s_1_2_2(or_1749_nl, or_1748_nl, fsm_output(4));
  or_1750_nl <= (fsm_output(8)) OR mux_1757_nl;
  mux_1760_nl <= MUX_s_1_2_2(mux_1759_nl, or_1750_nl, fsm_output(1));
  or_1746_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_1745_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1755_nl <= MUX_s_1_2_2(or_1746_nl, or_1745_nl, fsm_output(4));
  or_1743_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  mux_1756_nl <= MUX_s_1_2_2(mux_1755_nl, or_1743_nl, fsm_output(8));
  or_1747_nl <= (fsm_output(1)) OR mux_1756_nl;
  mux_1761_nl <= MUX_s_1_2_2(mux_1760_nl, or_1747_nl, fsm_output(9));
  mux_1771_nl <= MUX_s_1_2_2(mux_1770_nl, mux_1761_nl, fsm_output(7));
  mux_1787_nl <= MUX_s_1_2_2(mux_1786_nl, mux_1771_nl, fsm_output(0));
  vec_rsc_0_10_i_wea_d_pff <= NOT mux_1787_nl;
  or_1850_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(5)) OR not_tmp_322;
  or_1848_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_1847_nl <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1846_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1817_nl <= MUX_s_1_2_2(or_1847_nl, or_1846_nl, fsm_output(0));
  mux_1818_nl <= MUX_s_1_2_2(or_1848_nl, mux_1817_nl, fsm_output(4));
  mux_1819_nl <= MUX_s_1_2_2(or_1850_nl, mux_1818_nl, fsm_output(1));
  or_1845_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR not_tmp_322;
  or_1843_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR not_tmp_322;
  mux_1814_nl <= MUX_s_1_2_2(or_1845_nl, or_1843_nl, fsm_output(0));
  or_1841_nl <= (fsm_output(0)) OR CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1815_nl <= MUX_s_1_2_2(mux_1814_nl, or_1841_nl, fsm_output(4));
  or_1839_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1816_nl <= MUX_s_1_2_2(mux_1815_nl, or_1839_nl, fsm_output(1));
  mux_1820_nl <= MUX_s_1_2_2(mux_1819_nl, mux_1816_nl, fsm_output(9));
  or_1838_nl <= CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  or_1837_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  mux_1810_nl <= MUX_s_1_2_2(or_1838_nl, or_1837_nl, fsm_output(0));
  or_1836_nl <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  mux_1811_nl <= MUX_s_1_2_2(mux_1810_nl, or_1836_nl, fsm_output(4));
  or_1835_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(4)) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  mux_1812_nl <= MUX_s_1_2_2(mux_1811_nl, or_1835_nl, fsm_output(1));
  nand_300_nl <= NOT(operator_64_false_slc_operator_64_false_acc_1_60_itm AND (fsm_output(0))
      AND CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1010"))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  or_1832_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1831_nl <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1807_nl <= MUX_s_1_2_2(or_1832_nl, or_1831_nl, fsm_output(0));
  mux_1808_nl <= MUX_s_1_2_2(nand_300_nl, mux_1807_nl, fsm_output(4));
  or_1830_nl <= CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1809_nl <= MUX_s_1_2_2(mux_1808_nl, or_1830_nl, fsm_output(1));
  mux_1813_nl <= MUX_s_1_2_2(mux_1812_nl, mux_1809_nl, fsm_output(9));
  mux_1821_nl <= MUX_s_1_2_2(mux_1820_nl, mux_1813_nl, fsm_output(8));
  or_1829_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1827_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1802_nl <= MUX_s_1_2_2(or_1829_nl, or_1827_nl, fsm_output(0));
  or_1825_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR nand_442_cse;
  mux_1803_nl <= MUX_s_1_2_2(mux_1802_nl, or_1825_nl, fsm_output(4));
  or_1823_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_1799_nl <= MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_1823_nl);
  or_1822_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1820_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"));
  mux_1800_nl <= MUX_s_1_2_2(mux_1799_nl, or_1822_nl, or_1820_nl);
  or_1819_nl <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT
      (fsm_output(2)));
  mux_1801_nl <= MUX_s_1_2_2(mux_1800_nl, or_1819_nl, fsm_output(0));
  nand_80_nl <= NOT((fsm_output(4)) AND (NOT mux_1801_nl));
  mux_1804_nl <= MUX_s_1_2_2(mux_1803_nl, nand_80_nl, fsm_output(1));
  or_1817_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT
      (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1815_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT
      (fsm_output(3))) OR (fsm_output(2));
  mux_1797_nl <= MUX_s_1_2_2(or_1817_nl, or_1815_nl, fsm_output(4));
  or_1814_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3))
      OR (NOT (fsm_output(2)));
  or_1812_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_1805_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"));
  mux_1793_nl <= MUX_s_1_2_2(mux_1112_cse, nand_437_cse, or_1805_nl);
  or_1804_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_1802_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"));
  mux_1794_nl <= MUX_s_1_2_2(mux_1793_nl, or_1804_nl, or_1802_nl);
  mux_1795_nl <= MUX_s_1_2_2(or_1812_nl, mux_1794_nl, fsm_output(0));
  mux_1796_nl <= MUX_s_1_2_2(or_1814_nl, mux_1795_nl, fsm_output(4));
  mux_1798_nl <= MUX_s_1_2_2(mux_1797_nl, mux_1796_nl, fsm_output(1));
  mux_1805_nl <= MUX_s_1_2_2(mux_1804_nl, mux_1798_nl, fsm_output(9));
  or_1800_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(4)) OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm)
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1799_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1798_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (COMP_LOOP_acc_10_psp_sva(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_1797_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1788_nl <= MUX_s_1_2_2(or_1798_nl, or_1797_nl, fsm_output(0));
  mux_1789_nl <= MUX_s_1_2_2(or_1799_nl, mux_1788_nl, fsm_output(4));
  mux_1790_nl <= MUX_s_1_2_2(or_1800_nl, mux_1789_nl, fsm_output(1));
  or_1801_nl <= (fsm_output(9)) OR mux_1790_nl;
  mux_1806_nl <= MUX_s_1_2_2(mux_1805_nl, or_1801_nl, fsm_output(8));
  mux_1822_nl <= MUX_s_1_2_2(mux_1821_nl, mux_1806_nl, fsm_output(7));
  vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= NOT mux_1822_nl;
  nor_633_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_634_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1851_nl <= MUX_s_1_2_2(nor_633_nl, nor_634_nl, fsm_output(4));
  and_772_nl <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  and_778_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  mux_1850_nl <= MUX_s_1_2_2(and_772_nl, and_778_nl, fsm_output(4));
  mux_1852_nl <= MUX_s_1_2_2(mux_1851_nl, mux_1850_nl, fsm_output(8));
  nand_84_nl <= NOT((fsm_output(1)) AND mux_1852_nl);
  nor_637_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(2)) OR not_tmp_311);
  nor_638_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(2)) OR not_tmp_311);
  mux_1848_nl <= MUX_s_1_2_2(nor_637_nl, nor_638_nl, fsm_output(4));
  nand_83_nl <= NOT((fsm_output(8)) AND mux_1848_nl);
  or_1895_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1893_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1846_nl <= MUX_s_1_2_2(or_1895_nl, or_1893_nl, fsm_output(4));
  or_1892_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1011")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1847_nl <= MUX_s_1_2_2(mux_1846_nl, or_1892_nl, fsm_output(8));
  mux_1849_nl <= MUX_s_1_2_2(nand_83_nl, mux_1847_nl, fsm_output(1));
  mux_1853_nl <= MUX_s_1_2_2(nand_84_nl, mux_1849_nl, fsm_output(9));
  nand_291_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(5))));
  nand_471_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5)));
  mux_1843_nl <= MUX_s_1_2_2(nand_291_nl, nand_471_nl, fsm_output(4));
  or_1887_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1885_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_1842_nl <= MUX_s_1_2_2(or_1887_nl, or_1885_nl, fsm_output(4));
  mux_1844_nl <= MUX_s_1_2_2(mux_1843_nl, mux_1842_nl, fsm_output(8));
  or_1891_nl <= (fsm_output(1)) OR mux_1844_nl;
  or_1882_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1881_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1840_nl <= MUX_s_1_2_2(or_1882_nl, or_1881_nl, fsm_output(4));
  or_1883_nl <= (fsm_output(8)) OR mux_1840_nl;
  or_1880_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR not_tmp_312;
  mux_1841_nl <= MUX_s_1_2_2(or_1883_nl, or_1880_nl, fsm_output(1));
  mux_1845_nl <= MUX_s_1_2_2(or_1891_nl, mux_1841_nl, fsm_output(9));
  mux_1854_nl <= MUX_s_1_2_2(mux_1853_nl, mux_1845_nl, fsm_output(7));
  or_1878_nl <= (NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1836_nl <= MUX_s_1_2_2(or_1878_nl, nand_tmp_82, fsm_output(1));
  or_1875_nl <= CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1834_nl <= MUX_s_1_2_2(or_1018_cse, or_1875_nl, fsm_output(8));
  mux_1835_nl <= MUX_s_1_2_2(mux_1834_nl, nand_tmp_82, fsm_output(1));
  mux_1837_nl <= MUX_s_1_2_2(mux_1836_nl, mux_1835_nl, STAGE_VEC_LOOP_j_sva_9_0(3));
  nor_639_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_640_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1831_nl <= MUX_s_1_2_2(nor_639_nl, nor_640_nl, fsm_output(4));
  and_787_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  and_788_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("101"))
      AND (STAGE_VEC_LOOP_j_sva_9_0(0)) AND (fsm_output(2)) AND (fsm_output(3)) AND
      (NOT (fsm_output(6))) AND (fsm_output(5));
  mux_1830_nl <= MUX_s_1_2_2(and_787_nl, and_788_nl, fsm_output(4));
  mux_1832_nl <= MUX_s_1_2_2(mux_1831_nl, mux_1830_nl, fsm_output(8));
  nand_81_nl <= NOT((fsm_output(1)) AND mux_1832_nl);
  mux_1838_nl <= MUX_s_1_2_2(mux_1837_nl, nand_81_nl, fsm_output(9));
  or_1864_nl <= (NOT(CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("101")))) OR not_tmp_312;
  or_1862_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (COMP_LOOP_acc_10_psp_sva(0))) OR (fsm_output(2)) OR not_tmp_311;
  or_1860_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5));
  mux_1826_nl <= MUX_s_1_2_2(or_1862_nl, or_1860_nl, fsm_output(4));
  mux_1827_nl <= MUX_s_1_2_2(or_1864_nl, mux_1826_nl, fsm_output(8));
  or_1858_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1857_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(2)) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1825_nl <= MUX_s_1_2_2(or_1858_nl, or_1857_nl, fsm_output(4));
  or_1859_nl <= (fsm_output(8)) OR mux_1825_nl;
  mux_1828_nl <= MUX_s_1_2_2(mux_1827_nl, or_1859_nl, fsm_output(1));
  nand_296_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(5))));
  nand_452_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5)));
  mux_1823_nl <= MUX_s_1_2_2(nand_296_nl, nand_452_nl, fsm_output(4));
  or_1852_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  mux_1824_nl <= MUX_s_1_2_2(mux_1823_nl, or_1852_nl, fsm_output(8));
  or_1856_nl <= (fsm_output(1)) OR mux_1824_nl;
  mux_1829_nl <= MUX_s_1_2_2(mux_1828_nl, or_1856_nl, fsm_output(9));
  mux_1839_nl <= MUX_s_1_2_2(mux_1838_nl, mux_1829_nl, fsm_output(7));
  mux_1855_nl <= MUX_s_1_2_2(mux_1854_nl, mux_1839_nl, fsm_output(0));
  vec_rsc_0_11_i_wea_d_pff <= NOT mux_1855_nl;
  or_1956_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(5)) OR not_tmp_322;
  nand_277_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(0)) AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      AND (NOT (fsm_output(5))) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT
      (fsm_output(2))));
  or_1953_nl <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1952_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1885_nl <= MUX_s_1_2_2(or_1953_nl, or_1952_nl, fsm_output(0));
  mux_1886_nl <= MUX_s_1_2_2(nand_277_nl, mux_1885_nl, fsm_output(4));
  mux_1887_nl <= MUX_s_1_2_2(or_1956_nl, mux_1886_nl, fsm_output(1));
  or_1951_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR not_tmp_322;
  or_1949_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR not_tmp_322;
  mux_1882_nl <= MUX_s_1_2_2(or_1951_nl, or_1949_nl, fsm_output(0));
  or_1947_nl <= (fsm_output(0)) OR CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1883_nl <= MUX_s_1_2_2(mux_1882_nl, or_1947_nl, fsm_output(4));
  or_1945_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1884_nl <= MUX_s_1_2_2(mux_1883_nl, or_1945_nl, fsm_output(1));
  mux_1888_nl <= MUX_s_1_2_2(mux_1887_nl, mux_1884_nl, fsm_output(9));
  nand_278_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("101"))
      AND (STAGE_VEC_LOOP_j_sva_9_0(0)) AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  nand_279_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  mux_1878_nl <= MUX_s_1_2_2(nand_278_nl, nand_279_nl, fsm_output(0));
  or_1942_nl <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  mux_1879_nl <= MUX_s_1_2_2(mux_1878_nl, or_1942_nl, fsm_output(4));
  or_1941_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(4)) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  mux_1880_nl <= MUX_s_1_2_2(mux_1879_nl, or_1941_nl, fsm_output(1));
  nand_280_nl <= NOT(operator_64_false_slc_operator_64_false_acc_1_60_itm AND (fsm_output(0))
      AND CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  or_1938_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_1937_nl <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1875_nl <= MUX_s_1_2_2(or_1938_nl, or_1937_nl, fsm_output(0));
  mux_1876_nl <= MUX_s_1_2_2(nand_280_nl, mux_1875_nl, fsm_output(4));
  or_1936_nl <= CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1877_nl <= MUX_s_1_2_2(mux_1876_nl, or_1936_nl, fsm_output(1));
  mux_1881_nl <= MUX_s_1_2_2(mux_1880_nl, mux_1877_nl, fsm_output(9));
  mux_1889_nl <= MUX_s_1_2_2(mux_1888_nl, mux_1881_nl, fsm_output(8));
  or_1935_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1933_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1870_nl <= MUX_s_1_2_2(or_1935_nl, or_1933_nl, fsm_output(0));
  or_1931_nl <= (NOT(operator_64_false_slc_operator_64_false_acc_1_60_itm AND CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1011")) AND (fsm_output(0)) AND (fsm_output(5))
      AND (NOT (fsm_output(6))))) OR nand_442_cse;
  mux_1871_nl <= MUX_s_1_2_2(mux_1870_nl, or_1931_nl, fsm_output(4));
  nand_466_nl <= NOT(CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm AND (fsm_output(5))
      AND (fsm_output(6)) AND (NOT (fsm_output(3))) AND (fsm_output(2)));
  nand_283_nl <= NOT(CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_1867_nl <= MUX_s_1_2_2(nand_tmp_19, or_tmp_669, nand_283_nl);
  and_543_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
  mux_1868_nl <= MUX_s_1_2_2(nand_466_nl, mux_1867_nl, and_543_nl);
  nand_462_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (NOT (fsm_output(3))) AND (fsm_output(2)));
  mux_1869_nl <= MUX_s_1_2_2(mux_1868_nl, nand_462_nl, fsm_output(0));
  nand_86_nl <= NOT((fsm_output(4)) AND (NOT mux_1869_nl));
  mux_1872_nl <= MUX_s_1_2_2(mux_1871_nl, nand_86_nl, fsm_output(1));
  or_1924_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT
      (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_1922_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT
      (fsm_output(3))) OR (fsm_output(2));
  mux_1865_nl <= MUX_s_1_2_2(or_1924_nl, or_1922_nl, fsm_output(4));
  or_1921_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3))
      OR (NOT (fsm_output(2)));
  or_1919_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm AND CONV_SL_1_1(fsm_output(6
      DOWNTO 5)=STD_LOGIC_VECTOR'("01")))) OR nand_442_cse;
  or_1917_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  and_544_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
  mux_1861_nl <= MUX_s_1_2_2(nand_437_cse, mux_1112_cse, and_544_nl);
  and_545_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
  mux_1862_nl <= MUX_s_1_2_2(or_1917_nl, mux_1861_nl, and_545_nl);
  mux_1863_nl <= MUX_s_1_2_2(or_1919_nl, mux_1862_nl, fsm_output(0));
  mux_1864_nl <= MUX_s_1_2_2(or_1921_nl, mux_1863_nl, fsm_output(4));
  mux_1866_nl <= MUX_s_1_2_2(mux_1865_nl, mux_1864_nl, fsm_output(1));
  mux_1873_nl <= MUX_s_1_2_2(mux_1872_nl, mux_1866_nl, fsm_output(9));
  or_1909_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(4)) OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm)
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1908_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_1907_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (COMP_LOOP_acc_10_psp_sva(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_1906_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1856_nl <= MUX_s_1_2_2(or_1907_nl, or_1906_nl, fsm_output(0));
  mux_1857_nl <= MUX_s_1_2_2(or_1908_nl, mux_1856_nl, fsm_output(4));
  mux_1858_nl <= MUX_s_1_2_2(or_1909_nl, mux_1857_nl, fsm_output(1));
  or_1910_nl <= (fsm_output(9)) OR mux_1858_nl;
  mux_1874_nl <= MUX_s_1_2_2(mux_1873_nl, or_1910_nl, fsm_output(8));
  mux_1890_nl <= MUX_s_1_2_2(mux_1889_nl, mux_1874_nl, fsm_output(7));
  vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= NOT mux_1890_nl;
  nor_621_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_622_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1919_nl <= MUX_s_1_2_2(nor_621_nl, nor_622_nl, fsm_output(4));
  nor_623_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_624_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  mux_1918_nl <= MUX_s_1_2_2(nor_623_nl, nor_624_nl, fsm_output(4));
  mux_1920_nl <= MUX_s_1_2_2(mux_1919_nl, mux_1918_nl, fsm_output(8));
  nand_90_nl <= NOT((fsm_output(1)) AND mux_1920_nl);
  nor_625_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(2)) OR not_tmp_311);
  nor_626_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(2)) OR not_tmp_311);
  mux_1916_nl <= MUX_s_1_2_2(nor_625_nl, nor_626_nl, fsm_output(4));
  nand_89_nl <= NOT((fsm_output(8)) AND mux_1916_nl);
  or_2001_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1999_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1914_nl <= MUX_s_1_2_2(or_2001_nl, or_1999_nl, fsm_output(4));
  or_1998_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1100")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1915_nl <= MUX_s_1_2_2(mux_1914_nl, or_1998_nl, fsm_output(8));
  mux_1917_nl <= MUX_s_1_2_2(nand_89_nl, mux_1915_nl, fsm_output(1));
  mux_1921_nl <= MUX_s_1_2_2(nand_90_nl, mux_1917_nl, fsm_output(9));
  or_1996_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_1995_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1911_nl <= MUX_s_1_2_2(or_1996_nl, or_1995_nl, fsm_output(4));
  or_1993_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_1991_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_1910_nl <= MUX_s_1_2_2(or_1993_nl, or_1991_nl, fsm_output(4));
  mux_1912_nl <= MUX_s_1_2_2(mux_1911_nl, mux_1910_nl, fsm_output(8));
  or_1997_nl <= (fsm_output(1)) OR mux_1912_nl;
  or_1988_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1987_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1908_nl <= MUX_s_1_2_2(or_1988_nl, or_1987_nl, fsm_output(4));
  or_1989_nl <= (fsm_output(8)) OR mux_1908_nl;
  or_1986_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR not_tmp_312;
  mux_1909_nl <= MUX_s_1_2_2(or_1989_nl, or_1986_nl, fsm_output(1));
  mux_1913_nl <= MUX_s_1_2_2(or_1997_nl, mux_1909_nl, fsm_output(9));
  mux_1922_nl <= MUX_s_1_2_2(mux_1921_nl, mux_1913_nl, fsm_output(7));
  or_1984_nl <= (NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1904_nl <= MUX_s_1_2_2(or_1984_nl, nand_tmp_88, fsm_output(1));
  or_1981_nl <= CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1902_nl <= MUX_s_1_2_2(or_1124_cse, or_1981_nl, fsm_output(8));
  mux_1903_nl <= MUX_s_1_2_2(mux_1902_nl, nand_tmp_88, fsm_output(1));
  mux_1905_nl <= MUX_s_1_2_2(mux_1904_nl, mux_1903_nl, STAGE_VEC_LOOP_j_sva_9_0(3));
  nor_627_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_628_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1899_nl <= MUX_s_1_2_2(nor_627_nl, nor_628_nl, fsm_output(4));
  nor_629_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))));
  nor_630_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(5))));
  mux_1898_nl <= MUX_s_1_2_2(nor_629_nl, nor_630_nl, fsm_output(4));
  mux_1900_nl <= MUX_s_1_2_2(mux_1899_nl, mux_1898_nl, fsm_output(8));
  nand_87_nl <= NOT((fsm_output(1)) AND mux_1900_nl);
  mux_1906_nl <= MUX_s_1_2_2(mux_1905_nl, nand_87_nl, fsm_output(9));
  or_1970_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("101")) OR not_tmp_312;
  or_1968_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (COMP_LOOP_acc_10_psp_sva(0))) OR (fsm_output(2)) OR not_tmp_311;
  or_1966_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5));
  mux_1894_nl <= MUX_s_1_2_2(or_1968_nl, or_1966_nl, fsm_output(4));
  mux_1895_nl <= MUX_s_1_2_2(or_1970_nl, mux_1894_nl, fsm_output(8));
  or_1964_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_1963_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(5));
  mux_1893_nl <= MUX_s_1_2_2(or_1964_nl, or_1963_nl, fsm_output(4));
  or_1965_nl <= (fsm_output(8)) OR mux_1893_nl;
  mux_1896_nl <= MUX_s_1_2_2(mux_1895_nl, or_1965_nl, fsm_output(1));
  or_1961_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5));
  or_1960_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT
      (fsm_output(5)));
  mux_1891_nl <= MUX_s_1_2_2(or_1961_nl, or_1960_nl, fsm_output(4));
  or_1958_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  mux_1892_nl <= MUX_s_1_2_2(mux_1891_nl, or_1958_nl, fsm_output(8));
  or_1962_nl <= (fsm_output(1)) OR mux_1892_nl;
  mux_1897_nl <= MUX_s_1_2_2(mux_1896_nl, or_1962_nl, fsm_output(9));
  mux_1907_nl <= MUX_s_1_2_2(mux_1906_nl, mux_1897_nl, fsm_output(7));
  mux_1923_nl <= MUX_s_1_2_2(mux_1922_nl, mux_1907_nl, fsm_output(0));
  vec_rsc_0_12_i_wea_d_pff <= NOT mux_1923_nl;
  or_2065_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(5)) OR not_tmp_322;
  or_2063_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_2062_nl <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_2061_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1953_nl <= MUX_s_1_2_2(or_2062_nl, or_2061_nl, fsm_output(0));
  mux_1954_nl <= MUX_s_1_2_2(or_2063_nl, mux_1953_nl, fsm_output(4));
  mux_1955_nl <= MUX_s_1_2_2(or_2065_nl, mux_1954_nl, fsm_output(1));
  or_2060_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR not_tmp_322;
  or_2058_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR not_tmp_322;
  mux_1950_nl <= MUX_s_1_2_2(or_2060_nl, or_2058_nl, fsm_output(0));
  or_2056_nl <= (fsm_output(0)) OR CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1951_nl <= MUX_s_1_2_2(mux_1950_nl, or_2056_nl, fsm_output(4));
  or_2054_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1952_nl <= MUX_s_1_2_2(mux_1951_nl, or_2054_nl, fsm_output(1));
  mux_1956_nl <= MUX_s_1_2_2(mux_1955_nl, mux_1952_nl, fsm_output(9));
  or_2053_nl <= CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  or_2052_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2));
  mux_1946_nl <= MUX_s_1_2_2(or_2053_nl, or_2052_nl, fsm_output(0));
  or_2051_nl <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  mux_1947_nl <= MUX_s_1_2_2(mux_1946_nl, or_2051_nl, fsm_output(4));
  or_2050_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(4)) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  mux_1948_nl <= MUX_s_1_2_2(mux_1947_nl, or_2050_nl, fsm_output(1));
  nand_271_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1100"))
      AND operator_64_false_slc_operator_64_false_acc_1_60_itm AND (fsm_output(0))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  or_2047_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_2046_nl <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_1943_nl <= MUX_s_1_2_2(or_2047_nl, or_2046_nl, fsm_output(0));
  mux_1944_nl <= MUX_s_1_2_2(nand_271_nl, mux_1943_nl, fsm_output(4));
  or_2045_nl <= CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1945_nl <= MUX_s_1_2_2(mux_1944_nl, or_2045_nl, fsm_output(1));
  mux_1949_nl <= MUX_s_1_2_2(mux_1948_nl, mux_1945_nl, fsm_output(9));
  mux_1957_nl <= MUX_s_1_2_2(mux_1956_nl, mux_1949_nl, fsm_output(8));
  or_2044_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_2042_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_1938_nl <= MUX_s_1_2_2(or_2044_nl, or_2042_nl, fsm_output(0));
  or_2040_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5)))
      OR (fsm_output(6)) OR nand_442_cse;
  mux_1939_nl <= MUX_s_1_2_2(mux_1938_nl, or_2040_nl, fsm_output(4));
  or_2038_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_1935_nl <= MUX_s_1_2_2(nand_tmp_19, or_tmp_669, or_2038_nl);
  or_2037_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_2035_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"));
  mux_1936_nl <= MUX_s_1_2_2(mux_1935_nl, or_2037_nl, or_2035_nl);
  or_2034_nl <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT
      (fsm_output(2)));
  mux_1937_nl <= MUX_s_1_2_2(mux_1936_nl, or_2034_nl, fsm_output(0));
  nand_92_nl <= NOT((fsm_output(4)) AND (NOT mux_1937_nl));
  mux_1940_nl <= MUX_s_1_2_2(mux_1939_nl, nand_92_nl, fsm_output(1));
  or_2032_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT (fsm_output(0)))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_2030_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT
      (fsm_output(3))) OR (fsm_output(2));
  mux_1933_nl <= MUX_s_1_2_2(or_2032_nl, or_2030_nl, fsm_output(4));
  or_2029_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3))
      OR (NOT (fsm_output(2)));
  or_2027_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm) OR
      CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_2020_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"));
  mux_1929_nl <= MUX_s_1_2_2(mux_1112_cse, nand_437_cse, or_2020_nl);
  or_2019_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  or_2017_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"));
  mux_1930_nl <= MUX_s_1_2_2(mux_1929_nl, or_2019_nl, or_2017_nl);
  mux_1931_nl <= MUX_s_1_2_2(or_2027_nl, mux_1930_nl, fsm_output(0));
  mux_1932_nl <= MUX_s_1_2_2(or_2029_nl, mux_1931_nl, fsm_output(4));
  mux_1934_nl <= MUX_s_1_2_2(mux_1933_nl, mux_1932_nl, fsm_output(1));
  mux_1941_nl <= MUX_s_1_2_2(mux_1940_nl, mux_1934_nl, fsm_output(9));
  or_2015_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(4)) OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm)
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_2014_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_2013_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (COMP_LOOP_acc_10_psp_sva(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_2012_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1924_nl <= MUX_s_1_2_2(or_2013_nl, or_2012_nl, fsm_output(0));
  mux_1925_nl <= MUX_s_1_2_2(or_2014_nl, mux_1924_nl, fsm_output(4));
  mux_1926_nl <= MUX_s_1_2_2(or_2015_nl, mux_1925_nl, fsm_output(1));
  or_2016_nl <= (fsm_output(9)) OR mux_1926_nl;
  mux_1942_nl <= MUX_s_1_2_2(mux_1941_nl, or_2016_nl, fsm_output(8));
  mux_1958_nl <= MUX_s_1_2_2(mux_1957_nl, mux_1942_nl, fsm_output(7));
  vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= NOT mux_1958_nl;
  nor_609_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_610_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1987_nl <= MUX_s_1_2_2(nor_609_nl, nor_610_nl, fsm_output(4));
  and_771_nl <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  and_777_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  mux_1986_nl <= MUX_s_1_2_2(and_771_nl, and_777_nl, fsm_output(4));
  mux_1988_nl <= MUX_s_1_2_2(mux_1987_nl, mux_1986_nl, fsm_output(8));
  nand_96_nl <= NOT((fsm_output(1)) AND mux_1988_nl);
  nor_613_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(2)) OR not_tmp_311);
  nor_614_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(2)) OR not_tmp_311);
  mux_1984_nl <= MUX_s_1_2_2(nor_613_nl, nor_614_nl, fsm_output(4));
  nand_95_nl <= NOT((fsm_output(8)) AND mux_1984_nl);
  or_2110_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_2108_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1982_nl <= MUX_s_1_2_2(or_2110_nl, or_2108_nl, fsm_output(4));
  or_2107_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1101")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1983_nl <= MUX_s_1_2_2(mux_1982_nl, or_2107_nl, fsm_output(8));
  mux_1985_nl <= MUX_s_1_2_2(nand_95_nl, mux_1983_nl, fsm_output(1));
  mux_1989_nl <= MUX_s_1_2_2(nand_96_nl, mux_1985_nl, fsm_output(9));
  nand_262_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(5))));
  nand_470_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5)));
  mux_1979_nl <= MUX_s_1_2_2(nand_262_nl, nand_470_nl, fsm_output(4));
  or_2102_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_2100_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_1978_nl <= MUX_s_1_2_2(or_2102_nl, or_2100_nl, fsm_output(4));
  mux_1980_nl <= MUX_s_1_2_2(mux_1979_nl, mux_1978_nl, fsm_output(8));
  or_2106_nl <= (fsm_output(1)) OR mux_1980_nl;
  or_2097_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_2096_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1976_nl <= MUX_s_1_2_2(or_2097_nl, or_2096_nl, fsm_output(4));
  or_2098_nl <= (fsm_output(8)) OR mux_1976_nl;
  or_2095_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR not_tmp_312;
  mux_1977_nl <= MUX_s_1_2_2(or_2098_nl, or_2095_nl, fsm_output(1));
  mux_1981_nl <= MUX_s_1_2_2(or_2106_nl, mux_1977_nl, fsm_output(9));
  mux_1990_nl <= MUX_s_1_2_2(mux_1989_nl, mux_1981_nl, fsm_output(7));
  or_2093_nl <= (NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1972_nl <= MUX_s_1_2_2(or_2093_nl, nand_tmp_94, fsm_output(1));
  or_2090_nl <= CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_1970_nl <= MUX_s_1_2_2(or_1233_cse, or_2090_nl, fsm_output(8));
  mux_1971_nl <= MUX_s_1_2_2(mux_1970_nl, nand_tmp_94, fsm_output(1));
  mux_1973_nl <= MUX_s_1_2_2(mux_1972_nl, mux_1971_nl, STAGE_VEC_LOOP_j_sva_9_0(3));
  nor_615_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_616_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_1967_nl <= MUX_s_1_2_2(nor_615_nl, nor_616_nl, fsm_output(4));
  and_785_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  and_786_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("110"))
      AND (STAGE_VEC_LOOP_j_sva_9_0(0)) AND (fsm_output(2)) AND (fsm_output(3)) AND
      (NOT (fsm_output(6))) AND (fsm_output(5));
  mux_1966_nl <= MUX_s_1_2_2(and_785_nl, and_786_nl, fsm_output(4));
  mux_1968_nl <= MUX_s_1_2_2(mux_1967_nl, mux_1966_nl, fsm_output(8));
  nand_93_nl <= NOT((fsm_output(1)) AND mux_1968_nl);
  mux_1974_nl <= MUX_s_1_2_2(mux_1973_nl, nand_93_nl, fsm_output(9));
  or_2079_nl <= (NOT(CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("101")))) OR not_tmp_312;
  or_2077_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (COMP_LOOP_acc_10_psp_sva(0))) OR (fsm_output(2)) OR not_tmp_311;
  or_2075_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5));
  mux_1962_nl <= MUX_s_1_2_2(or_2077_nl, or_2075_nl, fsm_output(4));
  mux_1963_nl <= MUX_s_1_2_2(or_2079_nl, mux_1962_nl, fsm_output(8));
  or_2073_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_2072_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(2)) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_1961_nl <= MUX_s_1_2_2(or_2073_nl, or_2072_nl, fsm_output(4));
  or_2074_nl <= (fsm_output(8)) OR mux_1961_nl;
  mux_1964_nl <= MUX_s_1_2_2(mux_1963_nl, or_2074_nl, fsm_output(1));
  nand_267_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(5))));
  nand_451_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5)));
  mux_1959_nl <= MUX_s_1_2_2(nand_267_nl, nand_451_nl, fsm_output(4));
  or_2067_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  mux_1960_nl <= MUX_s_1_2_2(mux_1959_nl, or_2067_nl, fsm_output(8));
  or_2071_nl <= (fsm_output(1)) OR mux_1960_nl;
  mux_1965_nl <= MUX_s_1_2_2(mux_1964_nl, or_2071_nl, fsm_output(9));
  mux_1975_nl <= MUX_s_1_2_2(mux_1974_nl, mux_1965_nl, fsm_output(7));
  mux_1991_nl <= MUX_s_1_2_2(mux_1990_nl, mux_1975_nl, fsm_output(0));
  vec_rsc_0_13_i_wea_d_pff <= NOT mux_1991_nl;
  or_2171_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(5)) OR not_tmp_322;
  nand_248_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(0)) AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      AND (NOT (fsm_output(5))) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT
      (fsm_output(2))));
  or_2168_nl <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_2167_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_2021_nl <= MUX_s_1_2_2(or_2168_nl, or_2167_nl, fsm_output(0));
  mux_2022_nl <= MUX_s_1_2_2(nand_248_nl, mux_2021_nl, fsm_output(4));
  mux_2023_nl <= MUX_s_1_2_2(or_2171_nl, mux_2022_nl, fsm_output(1));
  or_2166_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR not_tmp_322;
  or_2164_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(5)) OR not_tmp_322;
  mux_2018_nl <= MUX_s_1_2_2(or_2166_nl, or_2164_nl, fsm_output(0));
  or_2162_nl <= (fsm_output(0)) OR CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_2019_nl <= MUX_s_1_2_2(mux_2018_nl, or_2162_nl, fsm_output(4));
  or_2160_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_2020_nl <= MUX_s_1_2_2(mux_2019_nl, or_2160_nl, fsm_output(1));
  mux_2024_nl <= MUX_s_1_2_2(mux_2023_nl, mux_2020_nl, fsm_output(9));
  nand_249_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("110"))
      AND (STAGE_VEC_LOOP_j_sva_9_0(0)) AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  nand_250_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  mux_2014_nl <= MUX_s_1_2_2(nand_249_nl, nand_250_nl, fsm_output(0));
  or_2157_nl <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  mux_2015_nl <= MUX_s_1_2_2(mux_2014_nl, or_2157_nl, fsm_output(4));
  or_2156_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(4)) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  mux_2016_nl <= MUX_s_1_2_2(mux_2015_nl, or_2156_nl, fsm_output(1));
  nand_251_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND operator_64_false_slc_operator_64_false_acc_1_60_itm AND (fsm_output(0))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  or_2153_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_2152_nl <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_2011_nl <= MUX_s_1_2_2(or_2153_nl, or_2152_nl, fsm_output(0));
  mux_2012_nl <= MUX_s_1_2_2(nand_251_nl, mux_2011_nl, fsm_output(4));
  or_2151_nl <= CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_2013_nl <= MUX_s_1_2_2(mux_2012_nl, or_2151_nl, fsm_output(1));
  mux_2017_nl <= MUX_s_1_2_2(mux_2016_nl, mux_2013_nl, fsm_output(9));
  mux_2025_nl <= MUX_s_1_2_2(mux_2024_nl, mux_2017_nl, fsm_output(8));
  or_2150_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_2148_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_2006_nl <= MUX_s_1_2_2(or_2150_nl, or_2148_nl, fsm_output(0));
  or_2146_nl <= (NOT(operator_64_false_slc_operator_64_false_acc_1_60_itm AND CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1101")) AND (fsm_output(0)) AND (fsm_output(5))
      AND (NOT (fsm_output(6))))) OR nand_442_cse;
  mux_2007_nl <= MUX_s_1_2_2(mux_2006_nl, or_2146_nl, fsm_output(4));
  nand_465_nl <= NOT(CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm AND (fsm_output(5))
      AND (fsm_output(6)) AND (NOT (fsm_output(3))) AND (fsm_output(2)));
  nand_254_nl <= NOT(CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_2003_nl <= MUX_s_1_2_2(nand_tmp_19, or_tmp_669, nand_254_nl);
  and_540_nl <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
  mux_2004_nl <= MUX_s_1_2_2(nand_465_nl, mux_2003_nl, and_540_nl);
  nand_461_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (NOT (fsm_output(3))) AND (fsm_output(2)));
  mux_2005_nl <= MUX_s_1_2_2(mux_2004_nl, nand_461_nl, fsm_output(0));
  nand_98_nl <= NOT((fsm_output(4)) AND (NOT mux_2005_nl));
  mux_2008_nl <= MUX_s_1_2_2(mux_2007_nl, nand_98_nl, fsm_output(1));
  or_2139_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT (fsm_output(0)))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_2137_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT
      (fsm_output(3))) OR (fsm_output(2));
  mux_2001_nl <= MUX_s_1_2_2(or_2139_nl, or_2137_nl, fsm_output(4));
  or_2136_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3))
      OR (NOT (fsm_output(2)));
  or_2134_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm AND CONV_SL_1_1(fsm_output(6
      DOWNTO 5)=STD_LOGIC_VECTOR'("01")))) OR nand_442_cse;
  or_2132_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  and_541_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
  mux_1997_nl <= MUX_s_1_2_2(nand_437_cse, mux_1112_cse, and_541_nl);
  and_542_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
  mux_1998_nl <= MUX_s_1_2_2(or_2132_nl, mux_1997_nl, and_542_nl);
  mux_1999_nl <= MUX_s_1_2_2(or_2134_nl, mux_1998_nl, fsm_output(0));
  mux_2000_nl <= MUX_s_1_2_2(or_2136_nl, mux_1999_nl, fsm_output(4));
  mux_2002_nl <= MUX_s_1_2_2(mux_2001_nl, mux_2000_nl, fsm_output(1));
  mux_2009_nl <= MUX_s_1_2_2(mux_2008_nl, mux_2002_nl, fsm_output(9));
  or_2124_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(4)) OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm)
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_2123_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_2122_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (COMP_LOOP_acc_10_psp_sva(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_2121_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_1992_nl <= MUX_s_1_2_2(or_2122_nl, or_2121_nl, fsm_output(0));
  mux_1993_nl <= MUX_s_1_2_2(or_2123_nl, mux_1992_nl, fsm_output(4));
  mux_1994_nl <= MUX_s_1_2_2(or_2124_nl, mux_1993_nl, fsm_output(1));
  or_2125_nl <= (fsm_output(9)) OR mux_1994_nl;
  mux_2010_nl <= MUX_s_1_2_2(mux_2009_nl, or_2125_nl, fsm_output(8));
  mux_2026_nl <= MUX_s_1_2_2(mux_2025_nl, mux_2010_nl, fsm_output(7));
  vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= NOT mux_2026_nl;
  nor_597_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_598_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_2055_nl <= MUX_s_1_2_2(nor_597_nl, nor_598_nl, fsm_output(4));
  and_770_nl <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  and_776_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  mux_2054_nl <= MUX_s_1_2_2(and_770_nl, and_776_nl, fsm_output(4));
  mux_2056_nl <= MUX_s_1_2_2(mux_2055_nl, mux_2054_nl, fsm_output(8));
  nand_102_nl <= NOT((fsm_output(1)) AND mux_2056_nl);
  nor_601_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(2)) OR not_tmp_311);
  nor_602_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(2)) OR not_tmp_311);
  mux_2052_nl <= MUX_s_1_2_2(nor_601_nl, nor_602_nl, fsm_output(4));
  nand_101_nl <= NOT((fsm_output(8)) AND mux_2052_nl);
  or_2216_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_2214_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_2050_nl <= MUX_s_1_2_2(or_2216_nl, or_2214_nl, fsm_output(4));
  or_2213_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1110")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_2051_nl <= MUX_s_1_2_2(mux_2050_nl, or_2213_nl, fsm_output(8));
  mux_2053_nl <= MUX_s_1_2_2(nand_101_nl, mux_2051_nl, fsm_output(1));
  mux_2057_nl <= MUX_s_1_2_2(nand_102_nl, mux_2053_nl, fsm_output(9));
  nand_239_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(5))));
  nand_469_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5)));
  mux_2047_nl <= MUX_s_1_2_2(nand_239_nl, nand_469_nl, fsm_output(4));
  or_2208_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_2206_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_2046_nl <= MUX_s_1_2_2(or_2208_nl, or_2206_nl, fsm_output(4));
  mux_2048_nl <= MUX_s_1_2_2(mux_2047_nl, mux_2046_nl, fsm_output(8));
  or_2212_nl <= (fsm_output(1)) OR mux_2048_nl;
  or_2203_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_2202_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_2044_nl <= MUX_s_1_2_2(or_2203_nl, or_2202_nl, fsm_output(4));
  or_2204_nl <= (fsm_output(8)) OR mux_2044_nl;
  or_2201_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR not_tmp_312;
  mux_2045_nl <= MUX_s_1_2_2(or_2204_nl, or_2201_nl, fsm_output(1));
  mux_2049_nl <= MUX_s_1_2_2(or_2212_nl, mux_2045_nl, fsm_output(9));
  mux_2058_nl <= MUX_s_1_2_2(mux_2057_nl, mux_2049_nl, fsm_output(7));
  or_2199_nl <= (NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_2040_nl <= MUX_s_1_2_2(or_2199_nl, nand_tmp_100, fsm_output(1));
  or_2196_nl <= CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_2038_nl <= MUX_s_1_2_2(or_1339_cse, or_2196_nl, fsm_output(8));
  mux_2039_nl <= MUX_s_1_2_2(mux_2038_nl, nand_tmp_100, fsm_output(1));
  mux_2041_nl <= MUX_s_1_2_2(mux_2040_nl, mux_2039_nl, STAGE_VEC_LOOP_j_sva_9_0(3));
  nor_603_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nor_604_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  mux_2035_nl <= MUX_s_1_2_2(nor_603_nl, nor_604_nl, fsm_output(4));
  and_783_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  and_784_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) AND (fsm_output(2)) AND (fsm_output(3))
      AND (NOT (fsm_output(6))) AND (fsm_output(5));
  mux_2034_nl <= MUX_s_1_2_2(and_783_nl, and_784_nl, fsm_output(4));
  mux_2036_nl <= MUX_s_1_2_2(mux_2035_nl, mux_2034_nl, fsm_output(8));
  nand_99_nl <= NOT((fsm_output(1)) AND mux_2036_nl);
  mux_2042_nl <= MUX_s_1_2_2(mux_2041_nl, nand_99_nl, fsm_output(9));
  or_2185_nl <= (NOT(CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("101")))) OR not_tmp_312;
  or_2183_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (COMP_LOOP_acc_10_psp_sva(0))) OR (fsm_output(2)) OR not_tmp_311;
  or_2181_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(5));
  mux_2030_nl <= MUX_s_1_2_2(or_2183_nl, or_2181_nl, fsm_output(4));
  mux_2031_nl <= MUX_s_1_2_2(or_2185_nl, mux_2030_nl, fsm_output(8));
  or_2179_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_2178_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(5));
  mux_2029_nl <= MUX_s_1_2_2(or_2179_nl, or_2178_nl, fsm_output(4));
  or_2180_nl <= (fsm_output(8)) OR mux_2029_nl;
  mux_2032_nl <= MUX_s_1_2_2(mux_2031_nl, or_2180_nl, fsm_output(1));
  nand_244_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(5))));
  nand_450_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5)));
  mux_2027_nl <= MUX_s_1_2_2(nand_244_nl, nand_450_nl, fsm_output(4));
  or_2173_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  mux_2028_nl <= MUX_s_1_2_2(mux_2027_nl, or_2173_nl, fsm_output(8));
  or_2177_nl <= (fsm_output(1)) OR mux_2028_nl;
  mux_2033_nl <= MUX_s_1_2_2(mux_2032_nl, or_2177_nl, fsm_output(9));
  mux_2043_nl <= MUX_s_1_2_2(mux_2042_nl, mux_2033_nl, fsm_output(7));
  mux_2059_nl <= MUX_s_1_2_2(mux_2058_nl, mux_2043_nl, fsm_output(0));
  vec_rsc_0_14_i_wea_d_pff <= NOT mux_2059_nl;
  or_2280_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(5)) OR not_tmp_322;
  nand_222_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(0)) AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      AND (NOT (fsm_output(5))) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT
      (fsm_output(2))));
  or_2277_nl <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_2276_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_2089_nl <= MUX_s_1_2_2(or_2277_nl, or_2276_nl, fsm_output(0));
  mux_2090_nl <= MUX_s_1_2_2(nand_222_nl, mux_2089_nl, fsm_output(4));
  mux_2091_nl <= MUX_s_1_2_2(or_2280_nl, mux_2090_nl, fsm_output(1));
  or_2275_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR not_tmp_322;
  or_2273_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR not_tmp_322;
  mux_2086_nl <= MUX_s_1_2_2(or_2275_nl, or_2273_nl, fsm_output(0));
  or_2271_nl <= (fsm_output(0)) OR CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_2087_nl <= MUX_s_1_2_2(mux_2086_nl, or_2271_nl, fsm_output(4));
  or_2269_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_2088_nl <= MUX_s_1_2_2(mux_2087_nl, or_2269_nl, fsm_output(1));
  mux_2092_nl <= MUX_s_1_2_2(mux_2091_nl, mux_2088_nl, fsm_output(9));
  nand_223_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  nand_224_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  mux_2082_nl <= MUX_s_1_2_2(nand_223_nl, nand_224_nl, fsm_output(0));
  or_2266_nl <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  mux_2083_nl <= MUX_s_1_2_2(mux_2082_nl, or_2266_nl, fsm_output(4));
  or_2265_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(4)) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  mux_2084_nl <= MUX_s_1_2_2(mux_2083_nl, or_2265_nl, fsm_output(1));
  nand_225_nl <= NOT(operator_64_false_slc_operator_64_false_acc_1_60_itm AND (fsm_output(0))
      AND CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(3)) AND (NOT (fsm_output(2))));
  or_2262_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  or_2261_nl <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(2));
  mux_2079_nl <= MUX_s_1_2_2(or_2262_nl, or_2261_nl, fsm_output(0));
  mux_2080_nl <= MUX_s_1_2_2(nand_225_nl, mux_2079_nl, fsm_output(4));
  or_2260_nl <= CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_2081_nl <= MUX_s_1_2_2(mux_2080_nl, or_2260_nl, fsm_output(1));
  mux_2085_nl <= MUX_s_1_2_2(mux_2084_nl, mux_2081_nl, fsm_output(9));
  mux_2093_nl <= MUX_s_1_2_2(mux_2092_nl, mux_2085_nl, fsm_output(8));
  or_2259_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (STAGE_VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_2257_nl <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  mux_2074_nl <= MUX_s_1_2_2(or_2259_nl, or_2257_nl, fsm_output(0));
  or_2255_nl <= (NOT(operator_64_false_slc_operator_64_false_acc_1_60_itm AND CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1110")) AND (fsm_output(0)) AND (fsm_output(5))
      AND (NOT (fsm_output(6))))) OR nand_442_cse;
  mux_2075_nl <= MUX_s_1_2_2(mux_2074_nl, or_2255_nl, fsm_output(4));
  nand_227_nl <= NOT(CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_2071_nl <= MUX_s_1_2_2(nand_tmp_19, or_tmp_669, nand_227_nl);
  nand_464_nl <= NOT(CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm AND (fsm_output(5))
      AND (fsm_output(6)) AND (NOT (fsm_output(3))) AND (fsm_output(2)));
  nand_229_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110")));
  mux_2072_nl <= MUX_s_1_2_2(mux_2071_nl, nand_464_nl, nand_229_nl);
  nand_460_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(5)) AND (fsm_output(6)) AND (NOT (fsm_output(3))) AND (fsm_output(2)));
  mux_2073_nl <= MUX_s_1_2_2(mux_2072_nl, nand_460_nl, fsm_output(0));
  nand_104_nl <= NOT((fsm_output(4)) AND (NOT mux_2073_nl));
  mux_2076_nl <= MUX_s_1_2_2(mux_2075_nl, nand_104_nl, fsm_output(1));
  or_2247_nl <= (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm) OR (NOT
      (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(2)));
  or_2245_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (NOT
      (fsm_output(3))) OR (fsm_output(2));
  mux_2069_nl <= MUX_s_1_2_2(or_2247_nl, or_2245_nl, fsm_output(4));
  or_2244_nl <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3))
      OR (NOT (fsm_output(2)));
  or_2242_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm AND CONV_SL_1_1(fsm_output(6
      DOWNTO 5)=STD_LOGIC_VECTOR'("01")))) OR nand_442_cse;
  nand_233_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110")));
  mux_2065_nl <= MUX_s_1_2_2(mux_1112_cse, nand_437_cse, nand_233_nl);
  or_2234_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01")) OR nand_442_cse;
  nand_234_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110")));
  mux_2066_nl <= MUX_s_1_2_2(mux_2065_nl, or_2234_nl, nand_234_nl);
  mux_2067_nl <= MUX_s_1_2_2(or_2242_nl, mux_2066_nl, fsm_output(0));
  mux_2068_nl <= MUX_s_1_2_2(or_2244_nl, mux_2067_nl, fsm_output(4));
  mux_2070_nl <= MUX_s_1_2_2(mux_2069_nl, mux_2068_nl, fsm_output(1));
  mux_2077_nl <= MUX_s_1_2_2(mux_2076_nl, mux_2070_nl, fsm_output(9));
  or_2230_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(4)) OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm)
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_2229_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(2));
  or_2228_nl <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (COMP_LOOP_acc_10_psp_sva(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  or_2227_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(2));
  mux_2060_nl <= MUX_s_1_2_2(or_2228_nl, or_2227_nl, fsm_output(0));
  mux_2061_nl <= MUX_s_1_2_2(or_2229_nl, mux_2060_nl, fsm_output(4));
  mux_2062_nl <= MUX_s_1_2_2(or_2230_nl, mux_2061_nl, fsm_output(1));
  or_2231_nl <= (fsm_output(9)) OR mux_2062_nl;
  mux_2078_nl <= MUX_s_1_2_2(mux_2077_nl, or_2231_nl, fsm_output(8));
  mux_2094_nl <= MUX_s_1_2_2(mux_2093_nl, mux_2078_nl, fsm_output(7));
  vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= NOT mux_2094_nl;
  and_536_nl <= CONV_SL_1_1(operator_64_false_acc_cse_1_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(2))) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT
      (fsm_output(5)));
  and_537_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(2))) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT
      (fsm_output(5)));
  mux_2123_nl <= MUX_s_1_2_2(and_536_nl, and_537_nl, fsm_output(4));
  and_769_nl <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  and_775_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  mux_2122_nl <= MUX_s_1_2_2(and_769_nl, and_775_nl, fsm_output(4));
  mux_2124_nl <= MUX_s_1_2_2(mux_2123_nl, mux_2122_nl, fsm_output(8));
  nand_108_nl <= NOT((fsm_output(1)) AND mux_2124_nl);
  nor_591_nl <= NOT((NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(2))))) OR not_tmp_311);
  nor_592_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(2))))) OR not_tmp_311);
  mux_2120_nl <= MUX_s_1_2_2(nor_591_nl, nor_592_nl, fsm_output(4));
  nand_107_nl <= NOT((fsm_output(8)) AND mux_2120_nl);
  or_2325_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_2323_nl <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_2118_nl <= MUX_s_1_2_2(or_2325_nl, or_2323_nl, fsm_output(4));
  or_2322_nl <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1111")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_2119_nl <= MUX_s_1_2_2(mux_2118_nl, or_2322_nl, fsm_output(8));
  mux_2121_nl <= MUX_s_1_2_2(nand_107_nl, mux_2119_nl, fsm_output(1));
  mux_2125_nl <= MUX_s_1_2_2(nand_108_nl, mux_2121_nl, fsm_output(9));
  nand_208_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(5))));
  nand_468_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5)));
  mux_2115_nl <= MUX_s_1_2_2(nand_208_nl, nand_468_nl, fsm_output(4));
  or_2317_nl <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  or_2315_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_2114_nl <= MUX_s_1_2_2(or_2317_nl, or_2315_nl, fsm_output(4));
  mux_2116_nl <= MUX_s_1_2_2(mux_2115_nl, mux_2114_nl, fsm_output(8));
  or_2321_nl <= (fsm_output(1)) OR mux_2116_nl;
  or_2312_nl <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_2311_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_2112_nl <= MUX_s_1_2_2(or_2312_nl, or_2311_nl, fsm_output(4));
  or_2313_nl <= (fsm_output(8)) OR mux_2112_nl;
  or_2310_nl <= (NOT(CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(8))) AND (fsm_output(4)) AND (fsm_output(2)) AND (NOT
      (fsm_output(3))))) OR not_tmp_312;
  mux_2113_nl <= MUX_s_1_2_2(or_2313_nl, or_2310_nl, fsm_output(1));
  mux_2117_nl <= MUX_s_1_2_2(or_2321_nl, mux_2113_nl, fsm_output(9));
  mux_2126_nl <= MUX_s_1_2_2(mux_2125_nl, mux_2117_nl, fsm_output(7));
  or_2308_nl <= (NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (NOT (fsm_output(2))) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_2108_nl <= MUX_s_1_2_2(or_2308_nl, nand_tmp_106, fsm_output(1));
  or_2305_nl <= CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(4)) OR CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  mux_2106_nl <= MUX_s_1_2_2(or_1448_cse, or_2305_nl, fsm_output(8));
  mux_2107_nl <= MUX_s_1_2_2(mux_2106_nl, nand_tmp_106, fsm_output(1));
  mux_2109_nl <= MUX_s_1_2_2(mux_2108_nl, mux_2107_nl, STAGE_VEC_LOOP_j_sva_9_0(3));
  and_538_nl <= CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(2))) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT
      (fsm_output(5)));
  and_539_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (STAGE_VEC_LOOP_j_sva_9_0(0)) AND (NOT (fsm_output(2))) AND (fsm_output(3))
      AND (fsm_output(6)) AND (NOT (fsm_output(5)));
  mux_2103_nl <= MUX_s_1_2_2(and_538_nl, and_539_nl, fsm_output(4));
  and_781_nl <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  and_782_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (STAGE_VEC_LOOP_j_sva_9_0(0)) AND (fsm_output(2)) AND (fsm_output(3)) AND
      (NOT (fsm_output(6))) AND (fsm_output(5));
  mux_2102_nl <= MUX_s_1_2_2(and_781_nl, and_782_nl, fsm_output(4));
  mux_2104_nl <= MUX_s_1_2_2(mux_2103_nl, mux_2102_nl, fsm_output(8));
  nand_105_nl <= NOT((fsm_output(1)) AND mux_2104_nl);
  mux_2110_nl <= MUX_s_1_2_2(mux_2109_nl, nand_105_nl, fsm_output(9));
  or_2294_nl <= (NOT(CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("101")))) OR not_tmp_312;
  or_2292_nl <= (NOT(CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (COMP_LOOP_acc_10_psp_sva(0)) AND (NOT (fsm_output(2))))) OR not_tmp_311;
  nand_215_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(2))) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT
      (fsm_output(5))));
  mux_2098_nl <= MUX_s_1_2_2(or_2292_nl, nand_215_nl, fsm_output(4));
  mux_2099_nl <= MUX_s_1_2_2(or_2294_nl, mux_2098_nl, fsm_output(8));
  or_2288_nl <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5));
  or_2287_nl <= CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(2)) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(5));
  mux_2097_nl <= MUX_s_1_2_2(or_2288_nl, or_2287_nl, fsm_output(4));
  or_2289_nl <= (fsm_output(8)) OR mux_2097_nl;
  mux_2100_nl <= MUX_s_1_2_2(mux_2099_nl, or_2289_nl, fsm_output(1));
  nand_216_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(5))));
  nand_449_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5)));
  mux_2095_nl <= MUX_s_1_2_2(nand_216_nl, nand_449_nl, fsm_output(4));
  or_2282_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1111")) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(5)));
  mux_2096_nl <= MUX_s_1_2_2(mux_2095_nl, or_2282_nl, fsm_output(8));
  or_2286_nl <= (fsm_output(1)) OR mux_2096_nl;
  mux_2101_nl <= MUX_s_1_2_2(mux_2100_nl, or_2286_nl, fsm_output(9));
  mux_2111_nl <= MUX_s_1_2_2(mux_2110_nl, mux_2101_nl, fsm_output(7));
  mux_2127_nl <= MUX_s_1_2_2(mux_2126_nl, mux_2111_nl, fsm_output(0));
  vec_rsc_0_15_i_wea_d_pff <= NOT mux_2127_nl;
  and_531_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(0)) AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(5)));
  nor_570_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5)));
  nor_571_nl <= NOT(CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5)));
  mux_2155_nl <= MUX_s_1_2_2(nor_570_nl, nor_571_nl, fsm_output(0));
  mux_2156_nl <= MUX_s_1_2_2(and_531_nl, mux_2155_nl, fsm_output(4));
  and_530_nl <= (fsm_output(1)) AND mux_2156_nl;
  and_532_nl <= (fsm_output(1)) AND (fsm_output(4)) AND (fsm_output(0)) AND CONV_SL_1_1(COMP_LOOP_acc_cse_10_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      AND (NOT (fsm_output(3))) AND (NOT (fsm_output(6))) AND (NOT (fsm_output(5)));
  mux_2157_nl <= MUX_s_1_2_2(and_530_nl, and_532_nl, fsm_output(9));
  nor_572_nl <= NOT((NOT(CONV_SL_1_1(operator_64_false_acc_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(9)) AND (NOT (fsm_output(1))) AND (fsm_output(4)) AND (NOT
      (fsm_output(0))))) OR not_tmp_311);
  mux_2158_nl <= MUX_s_1_2_2(mux_2157_nl, nor_572_nl, fsm_output(7));
  or_2835_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_9_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (STAGE_VEC_LOOP_j_sva_9_0(0)) AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm))
      OR not_tmp_311;
  nand_188_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_7_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(5)));
  mux_2151_nl <= MUX_s_1_2_2(or_2835_nl, nand_188_nl, fsm_output(0));
  or_2377_nl <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  mux_2152_nl <= MUX_s_1_2_2(mux_2151_nl, or_2377_nl, fsm_output(4));
  nor_573_nl <= NOT((fsm_output(1)) OR mux_2152_nl);
  and_533_nl <= operator_64_false_slc_operator_64_false_acc_1_60_itm AND (fsm_output(0))
      AND CONV_SL_1_1(COMP_LOOP_acc_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(5));
  and_766_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (STAGE_VEC_LOOP_j_sva_9_0(0)) AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      AND (NOT (fsm_output(3))) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  and_767_nl <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(3))) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  mux_2148_nl <= MUX_s_1_2_2(and_766_nl, and_767_nl, fsm_output(0));
  mux_2149_nl <= MUX_s_1_2_2(and_533_nl, mux_2148_nl, fsm_output(4));
  nor_576_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(4)) OR (fsm_output(0)) OR not_tmp_311);
  mux_2150_nl <= MUX_s_1_2_2(mux_2149_nl, nor_576_nl, fsm_output(1));
  mux_2153_nl <= MUX_s_1_2_2(nor_573_nl, mux_2150_nl, fsm_output(9));
  nand_459_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(4))) AND operator_64_false_slc_operator_64_false_acc_1_60_itm
      AND (fsm_output(0)) AND (NOT (fsm_output(3))) AND (NOT (fsm_output(6))) AND
      (fsm_output(5)));
  or_2365_nl <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(5)));
  nand_190_nl <= NOT(CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"))
      AND (COMP_LOOP_acc_10_psp_sva(0)) AND (STAGE_VEC_LOOP_j_sva_9_0(0)) AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(5))));
  nand_191_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_9_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(5))));
  mux_2145_nl <= MUX_s_1_2_2(nand_190_nl, nand_191_nl, fsm_output(0));
  mux_2146_nl <= MUX_s_1_2_2(or_2365_nl, mux_2145_nl, fsm_output(4));
  mux_2147_nl <= MUX_s_1_2_2(nand_459_nl, mux_2146_nl, fsm_output(1));
  nor_577_nl <= NOT((fsm_output(9)) OR mux_2147_nl);
  mux_2154_nl <= MUX_s_1_2_2(mux_2153_nl, nor_577_nl, fsm_output(7));
  mux_2159_nl <= MUX_s_1_2_2(mux_2158_nl, mux_2154_nl, fsm_output(8));
  nor_578_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(1)) OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(5)));
  nand_192_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (STAGE_VEC_LOOP_j_sva_9_0(0)) AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(5))));
  nand_193_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_11_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(5))));
  mux_2140_nl <= MUX_s_1_2_2(nand_192_nl, nand_193_nl, fsm_output(0));
  or_2357_nl <= (fsm_output(0)) OR CONV_SL_1_1(operator_64_false_acc_cse_10_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1111")) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(5));
  mux_2141_nl <= MUX_s_1_2_2(mux_2140_nl, or_2357_nl, fsm_output(4));
  nor_579_nl <= NOT((fsm_output(1)) OR mux_2141_nl);
  mux_2142_nl <= MUX_s_1_2_2(nor_578_nl, nor_579_nl, fsm_output(9));
  nor_580_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_7_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (NOT (STAGE_VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm)
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5)));
  nor_581_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5)));
  mux_2136_nl <= MUX_s_1_2_2(nor_580_nl, nor_581_nl, fsm_output(0));
  and_768_nl <= operator_64_false_slc_operator_64_false_acc_1_60_itm AND CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(0)) AND (fsm_output(3))
      AND (NOT (fsm_output(6))) AND (fsm_output(5));
  mux_2137_nl <= MUX_s_1_2_2(mux_2136_nl, and_768_nl, fsm_output(4));
  nand_448_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("01")));
  mux_2133_nl <= MUX_s_1_2_2(not_tmp_312, nand_448_nl, fsm_output(3));
  nand_422_nl <= NOT((fsm_output(3)) AND CONV_SL_1_1(operator_64_false_acc_cse_4_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("01")));
  nand_197_nl <= NOT((STAGE_VEC_LOOP_j_sva_9_0(1)) AND CONV_SL_1_1(COMP_LOOP_acc_8_psp_sva(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (STAGE_VEC_LOOP_j_sva_9_0(0)) AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_2134_nl <= MUX_s_1_2_2(mux_2133_nl, nand_422_nl, nand_197_nl);
  or_2347_nl <= (NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(3))))) OR not_tmp_312;
  mux_2135_nl <= MUX_s_1_2_2(mux_2134_nl, or_2347_nl, fsm_output(0));
  and_534_nl <= (fsm_output(4)) AND (NOT mux_2135_nl);
  mux_2138_nl <= MUX_s_1_2_2(mux_2137_nl, and_534_nl, fsm_output(1));
  nor_583_nl <= NOT((fsm_output(4)) OR (NOT operator_64_false_slc_operator_64_false_acc_1_60_itm)
      OR (NOT (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5)));
  nor_584_nl <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5)));
  and_774_nl <= CONV_SL_1_1(COMP_LOOP_acc_12_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm AND (fsm_output(3))
      AND (NOT (fsm_output(6))) AND (fsm_output(5));
  and_780_nl <= (fsm_output(3)) AND CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("01"));
  and_535_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("11"));
  and_791_nl <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("01"));
  mux_2128_nl <= MUX_s_1_2_2(and_535_nl, and_791_nl, fsm_output(3));
  mux_2129_nl <= MUX_s_1_2_2(and_780_nl, mux_2128_nl, COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm);
  mux_2130_nl <= MUX_s_1_2_2(and_774_nl, mux_2129_nl, fsm_output(0));
  mux_2131_nl <= MUX_s_1_2_2(nor_584_nl, mux_2130_nl, fsm_output(4));
  mux_2132_nl <= MUX_s_1_2_2(nor_583_nl, mux_2131_nl, fsm_output(1));
  mux_2139_nl <= MUX_s_1_2_2(mux_2138_nl, mux_2132_nl, fsm_output(9));
  mux_2143_nl <= MUX_s_1_2_2(mux_2142_nl, mux_2139_nl, fsm_output(7));
  and_792_nl <= CONV_SL_1_1(COMP_LOOP_acc_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(7))) AND (NOT (fsm_output(9))) AND (fsm_output(1)) AND
      (NOT (fsm_output(4))) AND (fsm_output(0)) AND COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  mux_2144_nl <= MUX_s_1_2_2(mux_2143_nl, and_792_nl, fsm_output(8));
  vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_2159_nl, mux_2144_nl,
      fsm_output(2));
  or_tmp_2740 <= NOT((fsm_output(5)) AND (fsm_output(3)) AND (NOT (fsm_output(8)))
      AND (fsm_output(2)));
  or_2912_nl <= (NOT (fsm_output(5))) OR (fsm_output(3)) OR (NOT (fsm_output(8)))
      OR (fsm_output(2));
  mux_2799_nl <= MUX_s_1_2_2(or_2912_nl, or_tmp_2740, fsm_output(4));
  or_2913_nl <= (fsm_output(7)) OR mux_2799_nl;
  or_2999_nl <= (fsm_output(5)) OR (fsm_output(3)) OR (NOT (fsm_output(8))) OR (fsm_output(2));
  mux_nl <= MUX_s_1_2_2(or_tmp_2740, or_2999_nl, fsm_output(4));
  nand_481_nl <= NOT((fsm_output(7)) AND (NOT mux_nl));
  mux_2800_nl <= MUX_s_1_2_2(or_2913_nl, nand_481_nl, fsm_output(1));
  or_tmp_2743 <= (fsm_output(6)) OR mux_2800_nl;
  or_2918_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(8))) OR (fsm_output(2));
  or_2917_nl <= (fsm_output(3)) OR (fsm_output(8)) OR (NOT (fsm_output(2)));
  mux_tmp_2749 <= MUX_s_1_2_2(or_2918_nl, or_2917_nl, fsm_output(5));
  nand_tmp_150 <= (fsm_output(7)) OR (NOT (fsm_output(4))) OR mux_tmp_2749;
  and_dcpl_402 <= CONV_SL_1_1(fsm_output=STD_LOGIC_VECTOR'("0000000101"));
  or_2929_cse <= (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT and_697_cse);
  or_2938_cse <= (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(0))
      OR (NOT (fsm_output(2)));
  and_dcpl_418 <= (NOT (fsm_output(2))) AND (fsm_output(1)) AND (fsm_output(8)) AND
      (fsm_output(0)) AND (fsm_output(7)) AND and_dcpl_95 AND (fsm_output(5)) AND
      (fsm_output(9)) AND (NOT (fsm_output(4)));
  and_dcpl_419 <= NOT((fsm_output(9)) OR (fsm_output(4)));
  and_dcpl_421 <= (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  and_dcpl_423 <= (fsm_output(0)) AND (NOT (fsm_output(7)));
  and_dcpl_424 <= (NOT (fsm_output(8))) AND (fsm_output(2));
  and_dcpl_427 <= and_dcpl_424 AND (fsm_output(1)) AND and_dcpl_423 AND and_dcpl_421
      AND and_dcpl_419;
  and_dcpl_429 <= and_711_cse AND (fsm_output(5));
  and_dcpl_431 <= NOT((fsm_output(0)) OR (fsm_output(7)));
  and_dcpl_432 <= NOT((fsm_output(8)) OR (fsm_output(2)));
  and_dcpl_433 <= and_dcpl_432 AND (NOT (fsm_output(1)));
  and_dcpl_434 <= and_dcpl_433 AND and_dcpl_431;
  and_dcpl_435 <= and_dcpl_434 AND and_dcpl_429 AND and_dcpl_419;
  and_dcpl_436 <= (NOT (fsm_output(9))) AND (fsm_output(4));
  and_dcpl_437 <= and_711_cse AND (NOT (fsm_output(5)));
  and_dcpl_439 <= (NOT (fsm_output(0))) AND (fsm_output(7));
  and_dcpl_440 <= and_dcpl_432 AND (fsm_output(1));
  and_dcpl_441 <= and_dcpl_440 AND and_dcpl_439;
  and_dcpl_442 <= and_dcpl_441 AND and_dcpl_437 AND and_dcpl_436;
  and_dcpl_444 <= and_dcpl_95 AND (NOT (fsm_output(5)));
  and_dcpl_445 <= and_dcpl_444 AND and_dcpl_436;
  and_dcpl_449 <= (fsm_output(8)) AND (NOT (fsm_output(2))) AND (fsm_output(1)) AND
      and_dcpl_423 AND and_dcpl_445;
  and_dcpl_451 <= (fsm_output(8)) AND (fsm_output(2));
  and_dcpl_452 <= and_dcpl_451 AND (NOT (fsm_output(1)));
  and_dcpl_453 <= and_dcpl_452 AND and_dcpl_431;
  and_dcpl_454 <= and_dcpl_453 AND and_dcpl_437 AND and_dcpl_419;
  and_dcpl_456 <= and_dcpl_451 AND (fsm_output(1));
  and_dcpl_457 <= and_dcpl_456 AND and_dcpl_439;
  and_dcpl_458 <= and_dcpl_457 AND and_dcpl_421 AND and_dcpl_436;
  and_dcpl_462 <= (fsm_output(0)) AND (fsm_output(7));
  and_dcpl_464 <= and_dcpl_456 AND and_dcpl_462 AND (NOT (fsm_output(3))) AND (fsm_output(6))
      AND (fsm_output(5)) AND and_dcpl_436;
  and_dcpl_465 <= (fsm_output(9)) AND (fsm_output(4));
  and_dcpl_466 <= and_dcpl_95 AND (fsm_output(5));
  and_dcpl_468 <= and_dcpl_434 AND and_dcpl_466 AND and_dcpl_465;
  and_dcpl_469 <= (fsm_output(9)) AND (NOT (fsm_output(4)));
  and_dcpl_470 <= and_dcpl_466 AND and_dcpl_469;
  and_dcpl_471 <= and_dcpl_441 AND and_dcpl_470;
  and_dcpl_474 <= and_dcpl_440 AND and_dcpl_462 AND and_dcpl_437 AND and_dcpl_465;
  and_dcpl_476 <= and_dcpl_453 AND and_dcpl_444 AND and_dcpl_465;
  and_dcpl_478 <= and_dcpl_440 AND and_dcpl_431 AND and_dcpl_445;
  and_dcpl_481 <= and_dcpl_433 AND and_dcpl_462 AND and_dcpl_466 AND and_dcpl_419;
  and_dcpl_483 <= and_dcpl_433 AND and_dcpl_423;
  and_dcpl_484 <= and_dcpl_483 AND and_dcpl_429 AND and_dcpl_469;
  and_dcpl_487 <= and_dcpl_452 AND and_dcpl_423 AND and_dcpl_437 AND and_dcpl_469;
  or_2955_cse <= (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(0)))
      OR (fsm_output(2));
  mux_2829_cse <= MUX_s_1_2_2(or_2938_cse, or_2955_cse, fsm_output(1));
  mux_2830_cse <= MUX_s_1_2_2(or_2929_cse, or_2938_cse, fsm_output(1));
  or_2960_cse <= (fsm_output(1)) OR nand_176_cse;
  nand_484_nl <= NOT((fsm_output(7)) AND (fsm_output(1)) AND (fsm_output(6)) AND
      (fsm_output(3)) AND mux_2326_cse);
  mux_2832_nl <= MUX_s_1_2_2(or_2960_cse, mux_2830_cse, fsm_output(7));
  mux_2833_nl <= MUX_s_1_2_2(nand_484_nl, mux_2832_nl, fsm_output(4));
  or_2958_nl <= (fsm_output(4)) OR (fsm_output(7)) OR mux_2829_cse;
  mux_2834_nl <= MUX_s_1_2_2(mux_2833_nl, or_2958_nl, fsm_output(5));
  or_2952_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(0))
      OR (fsm_output(2));
  or_2950_nl <= (fsm_output(0)) OR (fsm_output(2));
  or_2949_nl <= (NOT (fsm_output(0))) OR (fsm_output(2));
  mux_2825_nl <= MUX_s_1_2_2(or_2950_nl, or_2949_nl, fsm_output(9));
  or_2951_nl <= (fsm_output(3)) OR mux_2825_nl;
  mux_2826_nl <= MUX_s_1_2_2(or_2952_nl, or_2951_nl, fsm_output(6));
  mux_2827_nl <= MUX_s_1_2_2(mux_2826_nl, or_2929_cse, fsm_output(1));
  or_2953_nl <= (fsm_output(4)) OR (fsm_output(7)) OR mux_2827_nl;
  nand_479_nl <= NOT((fsm_output(7)) AND (fsm_output(1)) AND (fsm_output(6)) AND
      (fsm_output(3)) AND (NOT (fsm_output(9))) AND (fsm_output(0)) AND (NOT (fsm_output(2))));
  or_2944_nl <= (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(0))) OR (fsm_output(2));
  or_2943_nl <= (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_2822_nl <= MUX_s_1_2_2(or_2944_nl, or_2943_nl, fsm_output(1));
  or_2942_nl <= (NOT (fsm_output(1))) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_2823_nl <= MUX_s_1_2_2(mux_2822_nl, or_2942_nl, fsm_output(7));
  mux_2824_nl <= MUX_s_1_2_2(nand_479_nl, mux_2823_nl, fsm_output(4));
  mux_2828_nl <= MUX_s_1_2_2(or_2953_nl, mux_2824_nl, fsm_output(5));
  mux_2835_cse <= MUX_s_1_2_2(mux_2834_nl, mux_2828_nl, fsm_output(8));
  and_dcpl_489 <= and_dcpl_452 AND and_dcpl_439 AND and_dcpl_470;
  and_dcpl_490 <= and_dcpl_444 AND and_dcpl_419;
  and_dcpl_491 <= and_dcpl_424 AND (NOT (fsm_output(1)));
  and_dcpl_493 <= and_dcpl_491 AND and_dcpl_431 AND and_dcpl_490;
  and_dcpl_495 <= and_dcpl_491 AND and_dcpl_423 AND and_dcpl_490;
  and_dcpl_496 <= and_dcpl_483 AND and_dcpl_445;
  and_dcpl_498 <= and_dcpl_457 AND and_dcpl_444 AND and_dcpl_469;
  and_dcpl_505 <= nor_554_cse AND (NOT (fsm_output(8)));
  and_dcpl_507 <= and_dcpl_505 AND and_dcpl_423 AND and_dcpl_490;
  and_dcpl_508 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_509 <= and_dcpl_508 AND (NOT (fsm_output(8)));
  and_dcpl_510 <= and_dcpl_509 AND and_dcpl_423;
  and_dcpl_511 <= and_dcpl_510 AND and_dcpl_490;
  and_920_cse <= and_dcpl_509 AND and_dcpl_431 AND and_dcpl_444 AND and_dcpl_436;
  nand_477_nl <= NOT((fsm_output(7)) AND (fsm_output(4)) AND (fsm_output(1)) AND
      (fsm_output(6)) AND (fsm_output(3)) AND mux_2332_cse);
  mux_2860_nl <= MUX_s_1_2_2(or_2960_cse, mux_2829_cse, fsm_output(4));
  or_2996_nl <= (fsm_output(4)) OR mux_2830_cse;
  mux_2861_nl <= MUX_s_1_2_2(mux_2860_nl, or_2996_nl, fsm_output(7));
  mux_2862_nl <= MUX_s_1_2_2(nand_477_nl, mux_2861_nl, fsm_output(8));
  nand_476_nl <= NOT((fsm_output(6)) AND (fsm_output(3)) AND mux_2332_cse);
  or_2989_nl <= (fsm_output(6)) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT
      and_697_cse);
  mux_2853_nl <= MUX_s_1_2_2(nand_476_nl, or_2989_nl, fsm_output(1));
  or_2987_nl <= (fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_2854_nl <= MUX_s_1_2_2(mux_2853_nl, or_2987_nl, fsm_output(4));
  or_2984_nl <= (fsm_output(6)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(0))
      OR (fsm_output(2));
  mux_2851_nl <= MUX_s_1_2_2(or_2955_cse, or_2984_nl, fsm_output(1));
  or_2986_nl <= (fsm_output(4)) OR mux_2851_nl;
  mux_2855_nl <= MUX_s_1_2_2(mux_2854_nl, or_2986_nl, fsm_output(7));
  nor_1007_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(0))
      OR (NOT (fsm_output(2))));
  nor_1008_nl <= NOT((fsm_output(3)) OR (fsm_output(9)) OR (NOT and_697_cse));
  mux_2850_nl <= MUX_s_1_2_2(nor_1007_nl, nor_1008_nl, fsm_output(6));
  nand_475_nl <= NOT((fsm_output(7)) AND (fsm_output(4)) AND (fsm_output(1)) AND
      mux_2850_nl);
  mux_2856_nl <= MUX_s_1_2_2(mux_2855_nl, nand_475_nl, fsm_output(8));
  mux_2863_itm <= MUX_s_1_2_2(mux_2862_nl, mux_2856_nl, fsm_output(5));
  and_925_cse <= and_dcpl_510 AND and_dcpl_437 AND and_dcpl_419;
  and_dcpl_523 <= (fsm_output(2)) AND (fsm_output(1)) AND (NOT (fsm_output(8)));
  and_dcpl_525 <= and_dcpl_523 AND and_dcpl_439 AND and_dcpl_490;
  and_dcpl_530 <= and_dcpl_523 AND and_dcpl_462;
  and_936_cse <= and_dcpl_530 AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(5))
      AND and_dcpl_436;
  and_dcpl_534 <= and_dcpl_505 AND and_dcpl_439;
  and_940_cse <= and_dcpl_534 AND and_dcpl_429 AND and_dcpl_436;
  and_945_cse <= nor_554_cse AND (fsm_output(8)) AND and_dcpl_423 AND and_dcpl_466
      AND and_dcpl_436;
  and_dcpl_543 <= (NOT (fsm_output(2))) AND (fsm_output(1)) AND (fsm_output(8));
  and_dcpl_544 <= and_dcpl_543 AND and_dcpl_431;
  and_950_cse <= and_dcpl_544 AND and_dcpl_429 AND and_dcpl_419;
  and_953_cse <= and_dcpl_543 AND and_dcpl_462 AND and_dcpl_466 AND and_dcpl_419;
  and_957_cse <= and_dcpl_508 AND (fsm_output(8)) AND and_dcpl_439 AND and_dcpl_437
      AND and_dcpl_436;
  and_960_cse <= and_dcpl_510 AND and_dcpl_444 AND and_dcpl_465;
  and_964_cse <= and_dcpl_523 AND and_dcpl_431 AND and_dcpl_437 AND and_dcpl_469;
  and_966_cse <= and_dcpl_530 AND and_dcpl_444 AND and_dcpl_469;
  and_970_cse <= and_dcpl_534 AND (NOT (fsm_output(3))) AND (fsm_output(6)) AND (NOT
      (fsm_output(5))) AND and_dcpl_469;
  and_973_cse <= and_dcpl_505 AND and_dcpl_462 AND and_dcpl_429 AND and_dcpl_465;
  and_975_cse <= and_dcpl_544 AND and_dcpl_466 AND and_dcpl_465;
  and_978_cse <= and_dcpl_543 AND and_dcpl_423 AND and_dcpl_429 AND and_dcpl_469;
  and_dcpl_582 <= and_dcpl_432 AND (fsm_output(1)) AND (NOT (fsm_output(0))) AND
      (NOT (fsm_output(7))) AND nor_1039_cse AND (NOT (fsm_output(9))) AND (fsm_output(4));
  and_dcpl_584 <= nor_1039_cse AND (NOT (fsm_output(9))) AND (NOT (fsm_output(4)));
  and_dcpl_589 <= and_dcpl_451 AND (NOT (fsm_output(1))) AND (fsm_output(0)) AND
      (fsm_output(7)) AND and_dcpl_584;
  and_dcpl_593 <= and_dcpl_432 AND (NOT (fsm_output(1))) AND (fsm_output(0)) AND
      (NOT (fsm_output(7))) AND and_dcpl_584;
  and_dcpl_599 <= and_dcpl_451 AND (fsm_output(1)) AND (NOT (fsm_output(0))) AND
      (fsm_output(7)) AND nor_1039_cse AND (fsm_output(9)) AND (NOT (fsm_output(4)));
  and_dcpl_621 <= and_dcpl_523 AND and_dcpl_439 AND and_dcpl_444 AND and_dcpl_419;
  mux_tmp_2812 <= MUX_s_1_2_2(and_694_cse, or_204_cse, fsm_output(3));
  mux_tmp_2813 <= MUX_s_1_2_2((NOT or_204_cse), or_204_cse, fsm_output(3));
  mux_tmp_2815 <= MUX_s_1_2_2((NOT or_204_cse), (fsm_output(6)), fsm_output(3));
  mux_tmp_2823 <= MUX_s_1_2_2((NOT (fsm_output(6))), and_694_cse, fsm_output(3));
  mux_tmp_2824 <= MUX_s_1_2_2((NOT and_694_cse), and_694_cse, fsm_output(3));
  operator_64_false_or_120_itm <= and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442 OR
      and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_or_121_cse <= (NOT mux_2835_cse) OR and_dcpl_495;
  operator_64_false_operator_64_false_or_1_cse <= (NOT(and_dcpl_427 OR and_dcpl_435
      OR and_dcpl_442 OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464
      OR and_dcpl_468 OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_478
      OR and_dcpl_481 OR and_dcpl_484 OR and_dcpl_487 OR (NOT mux_2835_cse) OR and_dcpl_493
      OR and_dcpl_495 OR and_dcpl_496 OR and_dcpl_498)) OR and_dcpl_489;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( not_tmp_266 = '0' ) THEN
        p_sva <= p_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( not_tmp_266 = '0' ) THEN
        r_sva <= r_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_vec_rsc_triosy_0_15_obj_ld_cse <= '0';
        reg_ensig_cgo_cse <= '0';
        COMP_LOOP_COMP_LOOP_nor_1_itm <= '0';
        COMP_LOOP_nor_12_itm <= '0';
        COMP_LOOP_nor_14_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_19_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_20_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_21_itm <= '0';
        COMP_LOOP_nor_17_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_23_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_24_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_25_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_26_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_27_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_28_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_29_itm <= '0';
      ELSE
        reg_vec_rsc_triosy_0_15_obj_ld_cse <= and_dcpl_199 AND and_dcpl_159 AND (NOT
            (fsm_output(0))) AND (fsm_output(7)) AND (fsm_output(8)) AND (fsm_output(9))
            AND (z_out_2(4));
        reg_ensig_cgo_cse <= NOT mux_2240_itm;
        COMP_LOOP_COMP_LOOP_nor_1_itm <= NOT(CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_12_itm <= NOT((COMP_LOOP_1_operator_64_false_acc_tmp(3)) OR
            (COMP_LOOP_1_operator_64_false_acc_tmp(2)) OR (COMP_LOOP_1_operator_64_false_acc_tmp(0)));
        COMP_LOOP_nor_14_itm <= NOT((COMP_LOOP_1_operator_64_false_acc_tmp(3)) OR
            (COMP_LOOP_1_operator_64_false_acc_tmp(1)) OR (COMP_LOOP_1_operator_64_false_acc_tmp(0)));
        COMP_LOOP_COMP_LOOP_and_19_itm <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_20_itm <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_21_itm <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_nor_17_itm <= NOT(CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_23_itm <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_24_itm <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_25_itm <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_26_itm <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_27_itm <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_28_itm <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_29_itm <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      reg_COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat_cse <= p_sva;
      modExp_dev_while_rem_cmp_a <= MUX_v_64_2_2(COMP_LOOP_10_modExp_dev_1_while_mul_mut,
          z_out, mux_2323_nl);
      STAGE_MAIN_LOOP_div_cmp_a <= MUX_v_64_2_2(z_out_3, COMP_LOOP_10_modExp_dev_1_while_mul_mut,
          and_dcpl_293);
      STAGE_MAIN_LOOP_div_cmp_b <= MUX_v_10_2_2(STAGE_MAIN_LOOP_lshift_psp_1_sva_mx0w0,
          STAGE_MAIN_LOOP_lshift_psp_1_sva, and_dcpl_293);
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_2339_nl OR and_dcpl_295) = '1' ) THEN
        STAGE_MAIN_LOOP_acc_1_psp_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'( "1010"),
            (COMP_LOOP_slc_acc_3_12_1_slc(3 DOWNTO 0)), and_dcpl_295);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(nor_548_nl, and_tmp_24, fsm_output(9))) = '1' ) THEN
        STAGE_MAIN_LOOP_lshift_psp_1_sva <= STAGE_MAIN_LOOP_lshift_psp_1_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (and_dcpl_295 OR and_dcpl_290 OR not_tmp_597 OR (NOT mux_2336_itm) OR
          COMP_LOOP_10_modExp_dev_1_while_mul_mut_mx0c4 OR COMP_LOOP_10_modExp_dev_1_while_mul_mut_mx0c5)
          = '1' ) THEN
        COMP_LOOP_10_modExp_dev_1_while_mul_mut <= MUX1HOT_v_64_4_2(z_out_3, z_out,
            STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000001"),
            modExp_dev_while_rem_cmp_z, STD_LOGIC_VECTOR'( and_dcpl_295 & operator_64_false_or_2_nl
            & not_tmp_597 & COMP_LOOP_10_modExp_dev_1_while_mul_mut_mx0c4));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        STAGE_VEC_LOOP_j_sva_9_0 <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( ((and_dcpl_95 AND (NOT (fsm_output(1))) AND ((fsm_output(2)) XOR (fsm_output(4)))
          AND (NOT (fsm_output(5))) AND (NOT (fsm_output(0))) AND (NOT (fsm_output(7)))
          AND and_dcpl) OR STAGE_VEC_LOOP_j_sva_9_0_mx0c1) = '1' ) THEN
        STAGE_VEC_LOOP_j_sva_9_0 <= MUX_v_10_2_2(STD_LOGIC_VECTOR'("0000000000"),
            (z_out_1(9 DOWNTO 0)), STAGE_VEC_LOOP_j_sva_9_0_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_2427_nl OR and_330_rgt) = '1' ) THEN
        modExp_dev_result_sva <= MUX_v_64_2_2(STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000001"),
            modExp_dev_while_rem_cmp_z, and_330_rgt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_2475_nl, mux_2450_nl, fsm_output(9))) = '1' ) THEN
        tmp_10_lpi_4_dfm <= MUX1HOT_v_64_18_2(STAGE_MAIN_LOOP_div_cmp_z, z_out_3,
            vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d,
            vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_6_i_qa_d, vec_rsc_0_7_i_qa_d,
            vec_rsc_0_8_i_qa_d, vec_rsc_0_9_i_qa_d, vec_rsc_0_10_i_qa_d, vec_rsc_0_11_i_qa_d,
            vec_rsc_0_12_i_qa_d, vec_rsc_0_13_i_qa_d, vec_rsc_0_14_i_qa_d, vec_rsc_0_15_i_qa_d,
            STD_LOGIC_VECTOR'( and_331_nl & and_dcpl_290 & COMP_LOOP_or_2_nl & COMP_LOOP_or_3_nl
            & COMP_LOOP_or_4_nl & COMP_LOOP_or_5_nl & COMP_LOOP_or_6_nl & COMP_LOOP_or_7_nl
            & COMP_LOOP_or_8_nl & COMP_LOOP_or_9_nl & COMP_LOOP_or_10_nl & COMP_LOOP_or_11_nl
            & COMP_LOOP_or_12_nl & COMP_LOOP_or_13_nl & COMP_LOOP_or_14_nl & COMP_LOOP_or_15_nl
            & COMP_LOOP_or_16_nl & COMP_LOOP_or_17_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm <= '0';
      ELSIF ( (and_dcpl_290 OR and_dcpl_98 OR (NOT mux_2336_itm) OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c3
          OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c4
          OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c5
          OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c6
          OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c7
          OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c8
          OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c9
          OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c10
          OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c11
          OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c12
          OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c13
          OR and_dcpl_345) = '1' ) THEN
        COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm <= MUX1HOT_s_1_4_2((NOT
            (z_out_2(64))), COMP_LOOP_COMP_LOOP_and_17_nl, (z_out_2(63)), (NOT (z_out_2(63))),
            STD_LOGIC_VECTOR'( modExp_dev_while_or_nl & and_dcpl_98 & modExp_dev_while_or_1_nl
            & and_dcpl_345));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_2864_nl AND nor_1039_cse) = '1' ) THEN
        COMP_LOOP_k_9_4_sva_4_0 <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), (COMP_LOOP_slc_acc_3_12_1_slc(4
            DOWNTO 0)), nand_486_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_acc_cse_1_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( or_dcpl_72 = '0' ) THEN
        operator_64_false_acc_cse_1_sva <= COMP_LOOP_1_operator_64_false_acc_tmp;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (and_dcpl_98 OR (NOT mux_2545_itm)) = '1' ) THEN
        COMP_LOOP_acc_psp_sva <= MUX_v_6_2_2((STD_LOGIC_VECTOR'( "00") & operator_64_false_or_2_nl_1),
            (z_out_1(5 DOWNTO 0)), mux_2545_itm);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_72 = '0' ) THEN
        operator_64_false_1_slc_operator_64_false_1_acc_5_itm <= operator_64_false_1_acc_nl(5);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_244_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_62_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_185_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_64_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_65_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_66_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_6_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_68_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_69_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_70_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_10_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_72_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_12_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_13_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_14_itm <= '0';
      ELSIF ( mux_2586_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_itm <= NOT(CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_COMP_LOOP_and_244_itm <= (COMP_LOOP_acc_8_psp_sva_1(0)) AND (STAGE_VEC_LOOP_j_sva_9_0(0))
            AND (NOT((COMP_LOOP_acc_8_psp_sva_1(1)) OR (STAGE_VEC_LOOP_j_sva_9_0(1))));
        COMP_LOOP_COMP_LOOP_and_62_itm <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_COMP_LOOP_and_185_itm <= CONV_SL_1_1(COMP_LOOP_acc_cse_4_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_64_itm <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_65_itm <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_66_itm <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_COMP_LOOP_and_6_itm <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_COMP_LOOP_and_68_itm <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_69_itm <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_70_itm <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_10_itm <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_72_itm <= CONV_SL_1_1(COMP_LOOP_acc_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_12_itm <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_13_itm <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_14_itm <= CONV_SL_1_1(STAGE_VEC_LOOP_j_sva_9_0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_8_psp_sva <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( (mux_2590_nl OR (fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_8_psp_sva <= COMP_LOOP_acc_8_psp_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_cse_4_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (NOT(mux_2592_nl AND and_dcpl)) = '1' ) THEN
        COMP_LOOP_acc_cse_4_sva <= COMP_LOOP_acc_cse_4_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_cse_2_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (NOT((NOT mux_2599_nl) AND nor_813_cse)) = '1' ) THEN
        COMP_LOOP_acc_cse_2_sva <= COMP_LOOP_acc_cse_2_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_acc_cse_2_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (NOT(mux_2601_nl AND and_dcpl)) = '1' ) THEN
        operator_64_false_acc_cse_2_sva <= operator_64_false_acc_cse_2_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_5_itm <= '0';
      ELSIF ( and_dcpl_354 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_5_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_2_sva_mx0w0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_51_itm <= '0';
      ELSIF ( and_dcpl_354 = '0' ) THEN
        COMP_LOOP_nor_51_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_2_sva_mx0w0(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_52_itm <= '0';
      ELSIF ( and_dcpl_354 = '0' ) THEN
        COMP_LOOP_nor_52_itm <= NOT((operator_64_false_acc_cse_2_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_2_sva_mx0w0(2)) OR (operator_64_false_acc_cse_2_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_77_itm <= '0';
      ELSIF ( and_dcpl_354 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_77_itm <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_54_itm <= '0';
      ELSIF ( and_dcpl_354 = '0' ) THEN
        COMP_LOOP_nor_54_itm <= NOT((operator_64_false_acc_cse_2_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_2_sva_mx0w0(1)) OR (operator_64_false_acc_cse_2_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_79_itm <= '0';
      ELSIF ( and_dcpl_354 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_79_itm <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_80_itm <= '0';
      ELSIF ( and_dcpl_354 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_80_itm <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_81_itm <= '0';
      ELSIF ( and_dcpl_354 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_81_itm <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_57_itm <= '0';
      ELSIF ( and_dcpl_354 = '0' ) THEN
        COMP_LOOP_nor_57_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_2_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_83_itm <= '0';
      ELSIF ( and_dcpl_354 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_83_itm <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_84_itm <= '0';
      ELSIF ( and_dcpl_354 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_84_itm <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_85_itm <= '0';
      ELSIF ( and_dcpl_354 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_85_itm <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_86_itm <= '0';
      ELSIF ( and_dcpl_354 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_86_itm <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_87_itm <= '0';
      ELSIF ( and_dcpl_354 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_87_itm <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_88_itm <= '0';
      ELSIF ( and_dcpl_354 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_88_itm <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_89_itm <= '0';
      ELSIF ( and_dcpl_354 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_89_itm <= CONV_SL_1_1(operator_64_false_acc_cse_2_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_7_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( (NOT((mux_tmp_2538 XOR (fsm_output(7))) AND and_dcpl)) = '1' ) THEN
        COMP_LOOP_acc_7_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0(9
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & STD_LOGIC_VECTOR'( "001")), 8), 9), 9));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_acc_cse_3_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (NOT(mux_2612_nl AND and_dcpl)) = '1' ) THEN
        operator_64_false_acc_cse_3_sva <= operator_64_false_acc_cse_3_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_9_itm <= '0';
      ELSIF ( and_dcpl_357 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_9_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_3_sva_mx0w0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_91_itm <= '0';
      ELSIF ( and_dcpl_357 = '0' ) THEN
        COMP_LOOP_nor_91_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_3_sva_mx0w0(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_92_itm <= '0';
      ELSIF ( and_dcpl_357 = '0' ) THEN
        COMP_LOOP_nor_92_itm <= NOT((operator_64_false_acc_cse_3_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_3_sva_mx0w0(2)) OR (operator_64_false_acc_cse_3_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_137_itm <= '0';
      ELSIF ( and_dcpl_357 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_137_itm <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_94_itm <= '0';
      ELSIF ( and_dcpl_357 = '0' ) THEN
        COMP_LOOP_nor_94_itm <= NOT((operator_64_false_acc_cse_3_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_3_sva_mx0w0(1)) OR (operator_64_false_acc_cse_3_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_139_itm <= '0';
      ELSIF ( and_dcpl_357 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_139_itm <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_140_itm <= '0';
      ELSIF ( and_dcpl_357 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_140_itm <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_141_itm <= '0';
      ELSIF ( and_dcpl_357 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_141_itm <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_97_itm <= '0';
      ELSIF ( and_dcpl_357 = '0' ) THEN
        COMP_LOOP_nor_97_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_3_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_143_itm <= '0';
      ELSIF ( and_dcpl_357 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_143_itm <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_144_itm <= '0';
      ELSIF ( and_dcpl_357 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_144_itm <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_145_itm <= '0';
      ELSIF ( and_dcpl_357 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_145_itm <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_146_itm <= '0';
      ELSIF ( and_dcpl_357 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_146_itm <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_147_itm <= '0';
      ELSIF ( and_dcpl_357 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_147_itm <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_148_itm <= '0';
      ELSIF ( and_dcpl_357 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_148_itm <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_149_itm <= '0';
      ELSIF ( and_dcpl_357 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_149_itm <= CONV_SL_1_1(operator_64_false_acc_cse_3_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_acc_cse_4_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (NOT(mux_2616_nl AND and_dcpl)) = '1' ) THEN
        operator_64_false_acc_cse_4_sva <= operator_64_false_acc_cse_4_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_13_itm <= '0';
      ELSIF ( and_dcpl_359 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_13_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_4_sva_mx0w0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_131_itm <= '0';
      ELSIF ( and_dcpl_359 = '0' ) THEN
        COMP_LOOP_nor_131_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_4_sva_mx0w0(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_132_itm <= '0';
      ELSIF ( and_dcpl_359 = '0' ) THEN
        COMP_LOOP_nor_132_itm <= NOT((operator_64_false_acc_cse_4_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_4_sva_mx0w0(2)) OR (operator_64_false_acc_cse_4_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_197_itm <= '0';
      ELSIF ( and_dcpl_359 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_197_itm <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_134_itm <= '0';
      ELSIF ( and_dcpl_359 = '0' ) THEN
        COMP_LOOP_nor_134_itm <= NOT((operator_64_false_acc_cse_4_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_4_sva_mx0w0(1)) OR (operator_64_false_acc_cse_4_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_199_itm <= '0';
      ELSIF ( and_dcpl_359 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_199_itm <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_200_itm <= '0';
      ELSIF ( and_dcpl_359 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_200_itm <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_201_itm <= '0';
      ELSIF ( and_dcpl_359 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_201_itm <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_137_itm <= '0';
      ELSIF ( and_dcpl_359 = '0' ) THEN
        COMP_LOOP_nor_137_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_4_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_203_itm <= '0';
      ELSIF ( and_dcpl_359 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_203_itm <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_204_itm <= '0';
      ELSIF ( and_dcpl_359 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_204_itm <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_205_itm <= '0';
      ELSIF ( and_dcpl_359 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_205_itm <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_206_itm <= '0';
      ELSIF ( and_dcpl_359 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_206_itm <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_207_itm <= '0';
      ELSIF ( and_dcpl_359 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_207_itm <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_208_itm <= '0';
      ELSIF ( and_dcpl_359 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_208_itm <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_209_itm <= '0';
      ELSIF ( and_dcpl_359 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_209_itm <= CONV_SL_1_1(operator_64_false_acc_cse_4_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_acc_cse_5_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_2621_nl OR (fsm_output(9))) = '1' ) THEN
        operator_64_false_acc_cse_5_sva <= operator_64_false_acc_cse_5_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_17_itm <= '0';
      ELSIF ( and_dcpl_361 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_17_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva_mx0w0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_171_itm <= '0';
      ELSIF ( and_dcpl_361 = '0' ) THEN
        COMP_LOOP_nor_171_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva_mx0w0(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_172_itm <= '0';
      ELSIF ( and_dcpl_361 = '0' ) THEN
        COMP_LOOP_nor_172_itm <= NOT((operator_64_false_acc_cse_5_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_5_sva_mx0w0(2)) OR (operator_64_false_acc_cse_5_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_257_itm <= '0';
      ELSIF ( and_dcpl_361 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_257_itm <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_174_itm <= '0';
      ELSIF ( and_dcpl_361 = '0' ) THEN
        COMP_LOOP_nor_174_itm <= NOT((operator_64_false_acc_cse_5_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_5_sva_mx0w0(1)) OR (operator_64_false_acc_cse_5_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_259_itm <= '0';
      ELSIF ( and_dcpl_361 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_259_itm <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_260_itm <= '0';
      ELSIF ( and_dcpl_361 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_260_itm <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_261_itm <= '0';
      ELSIF ( and_dcpl_361 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_261_itm <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_177_itm <= '0';
      ELSIF ( and_dcpl_361 = '0' ) THEN
        COMP_LOOP_nor_177_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_5_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_263_itm <= '0';
      ELSIF ( and_dcpl_361 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_263_itm <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_264_itm <= '0';
      ELSIF ( and_dcpl_361 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_264_itm <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_265_itm <= '0';
      ELSIF ( and_dcpl_361 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_265_itm <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_266_itm <= '0';
      ELSIF ( and_dcpl_361 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_266_itm <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_267_itm <= '0';
      ELSIF ( and_dcpl_361 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_267_itm <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_268_itm <= '0';
      ELSIF ( and_dcpl_361 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_268_itm <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_269_itm <= '0';
      ELSIF ( and_dcpl_361 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_269_itm <= CONV_SL_1_1(operator_64_false_acc_cse_5_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_cse_6_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_2624_nl OR (fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_cse_6_sva <= COMP_LOOP_slc_acc_3_12_1_slc(9 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_acc_cse_6_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_2633_nl OR (fsm_output(9))) = '1' ) THEN
        operator_64_false_acc_cse_6_sva <= operator_64_false_acc_cse_6_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_21_itm <= '0';
      ELSIF ( and_dcpl_364 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_21_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva_mx0w0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_211_itm <= '0';
      ELSIF ( and_dcpl_364 = '0' ) THEN
        COMP_LOOP_nor_211_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva_mx0w0(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_212_itm <= '0';
      ELSIF ( and_dcpl_364 = '0' ) THEN
        COMP_LOOP_nor_212_itm <= NOT((operator_64_false_acc_cse_6_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_6_sva_mx0w0(2)) OR (operator_64_false_acc_cse_6_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_317_itm <= '0';
      ELSIF ( and_dcpl_364 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_317_itm <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_214_itm <= '0';
      ELSIF ( and_dcpl_364 = '0' ) THEN
        COMP_LOOP_nor_214_itm <= NOT((operator_64_false_acc_cse_6_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_6_sva_mx0w0(1)) OR (operator_64_false_acc_cse_6_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_319_itm <= '0';
      ELSIF ( and_dcpl_364 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_319_itm <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_320_itm <= '0';
      ELSIF ( and_dcpl_364 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_320_itm <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_321_itm <= '0';
      ELSIF ( and_dcpl_364 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_321_itm <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_217_itm <= '0';
      ELSIF ( and_dcpl_364 = '0' ) THEN
        COMP_LOOP_nor_217_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_6_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_323_itm <= '0';
      ELSIF ( and_dcpl_364 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_323_itm <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_324_itm <= '0';
      ELSIF ( and_dcpl_364 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_324_itm <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_325_itm <= '0';
      ELSIF ( and_dcpl_364 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_325_itm <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_326_itm <= '0';
      ELSIF ( and_dcpl_364 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_326_itm <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_327_itm <= '0';
      ELSIF ( and_dcpl_364 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_327_itm <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_328_itm <= '0';
      ELSIF ( and_dcpl_364 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_328_itm <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_329_itm <= '0';
      ELSIF ( and_dcpl_364 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_329_itm <= CONV_SL_1_1(operator_64_false_acc_cse_6_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_9_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( (mux_2640_nl OR (fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_9_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0(9
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & STD_LOGIC_VECTOR'( "011")), 8), 9), 9));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_acc_cse_7_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_2641_nl OR (fsm_output(9))) = '1' ) THEN
        operator_64_false_acc_cse_7_sva <= operator_64_false_acc_cse_7_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_25_itm <= '0';
      ELSIF ( and_dcpl_367 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_25_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_7_sva_mx0w0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_251_itm <= '0';
      ELSIF ( and_dcpl_367 = '0' ) THEN
        COMP_LOOP_nor_251_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_7_sva_mx0w0(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_252_itm <= '0';
      ELSIF ( and_dcpl_367 = '0' ) THEN
        COMP_LOOP_nor_252_itm <= NOT((operator_64_false_acc_cse_7_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_7_sva_mx0w0(2)) OR (operator_64_false_acc_cse_7_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_377_itm <= '0';
      ELSIF ( and_dcpl_367 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_377_itm <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_254_itm <= '0';
      ELSIF ( and_dcpl_367 = '0' ) THEN
        COMP_LOOP_nor_254_itm <= NOT((operator_64_false_acc_cse_7_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_7_sva_mx0w0(1)) OR (operator_64_false_acc_cse_7_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_379_itm <= '0';
      ELSIF ( and_dcpl_367 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_379_itm <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_380_itm <= '0';
      ELSIF ( and_dcpl_367 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_380_itm <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_381_itm <= '0';
      ELSIF ( and_dcpl_367 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_381_itm <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_257_itm <= '0';
      ELSIF ( and_dcpl_367 = '0' ) THEN
        COMP_LOOP_nor_257_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_7_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_383_itm <= '0';
      ELSIF ( and_dcpl_367 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_383_itm <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_384_itm <= '0';
      ELSIF ( and_dcpl_367 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_384_itm <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_385_itm <= '0';
      ELSIF ( and_dcpl_367 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_385_itm <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_386_itm <= '0';
      ELSIF ( and_dcpl_367 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_386_itm <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_387_itm <= '0';
      ELSIF ( and_dcpl_367 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_387_itm <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_388_itm <= '0';
      ELSIF ( and_dcpl_367 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_388_itm <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_389_itm <= '0';
      ELSIF ( and_dcpl_367 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_389_itm <= CONV_SL_1_1(operator_64_false_acc_cse_7_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_cse_8_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_2645_nl OR (fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_cse_8_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "0111")), 9), 10), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_acc_cse_8_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_2649_nl OR (fsm_output(9))) = '1' ) THEN
        operator_64_false_acc_cse_8_sva <= operator_64_false_acc_cse_8_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_29_itm <= '0';
      ELSIF ( and_dcpl_370 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_29_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_8_sva_mx0w0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_291_itm <= '0';
      ELSIF ( and_dcpl_370 = '0' ) THEN
        COMP_LOOP_nor_291_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_8_sva_mx0w0(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_292_itm <= '0';
      ELSIF ( and_dcpl_370 = '0' ) THEN
        COMP_LOOP_nor_292_itm <= NOT((operator_64_false_acc_cse_8_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_8_sva_mx0w0(2)) OR (operator_64_false_acc_cse_8_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_437_itm <= '0';
      ELSIF ( and_dcpl_370 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_437_itm <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_294_itm <= '0';
      ELSIF ( and_dcpl_370 = '0' ) THEN
        COMP_LOOP_nor_294_itm <= NOT((operator_64_false_acc_cse_8_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_8_sva_mx0w0(1)) OR (operator_64_false_acc_cse_8_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_439_itm <= '0';
      ELSIF ( and_dcpl_370 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_439_itm <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_440_itm <= '0';
      ELSIF ( and_dcpl_370 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_440_itm <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_441_itm <= '0';
      ELSIF ( and_dcpl_370 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_441_itm <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_297_itm <= '0';
      ELSIF ( and_dcpl_370 = '0' ) THEN
        COMP_LOOP_nor_297_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_8_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_443_itm <= '0';
      ELSIF ( and_dcpl_370 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_443_itm <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_444_itm <= '0';
      ELSIF ( and_dcpl_370 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_444_itm <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_445_itm <= '0';
      ELSIF ( and_dcpl_370 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_445_itm <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_446_itm <= '0';
      ELSIF ( and_dcpl_370 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_446_itm <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_447_itm <= '0';
      ELSIF ( and_dcpl_370 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_447_itm <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_448_itm <= '0';
      ELSIF ( and_dcpl_370 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_448_itm <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_449_itm <= '0';
      ELSIF ( and_dcpl_370 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_449_itm <= CONV_SL_1_1(operator_64_false_acc_cse_8_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_psp_sva <= STD_LOGIC_VECTOR'( "0000000");
      ELSIF ( (mux_2657_nl OR (fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_10_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0(9
            DOWNTO 3)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & '1'), 6), 7), 7));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_acc_cse_9_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(not_tmp_698, or_2651_nl, fsm_output(9))) = '1' ) THEN
        operator_64_false_acc_cse_9_sva <= operator_64_false_acc_cse_9_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_33_itm <= '0';
      ELSIF ( and_dcpl_372 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_33_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_9_sva_mx0w0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_331_itm <= '0';
      ELSIF ( and_dcpl_372 = '0' ) THEN
        COMP_LOOP_nor_331_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_9_sva_mx0w0(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_332_itm <= '0';
      ELSIF ( and_dcpl_372 = '0' ) THEN
        COMP_LOOP_nor_332_itm <= NOT((operator_64_false_acc_cse_9_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_9_sva_mx0w0(2)) OR (operator_64_false_acc_cse_9_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_497_itm <= '0';
      ELSIF ( and_dcpl_372 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_497_itm <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_334_itm <= '0';
      ELSIF ( and_dcpl_372 = '0' ) THEN
        COMP_LOOP_nor_334_itm <= NOT((operator_64_false_acc_cse_9_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_9_sva_mx0w0(1)) OR (operator_64_false_acc_cse_9_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_499_itm <= '0';
      ELSIF ( and_dcpl_372 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_499_itm <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_500_itm <= '0';
      ELSIF ( and_dcpl_372 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_500_itm <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_501_itm <= '0';
      ELSIF ( and_dcpl_372 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_501_itm <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_337_itm <= '0';
      ELSIF ( and_dcpl_372 = '0' ) THEN
        COMP_LOOP_nor_337_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_9_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_503_itm <= '0';
      ELSIF ( and_dcpl_372 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_503_itm <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_504_itm <= '0';
      ELSIF ( and_dcpl_372 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_504_itm <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_505_itm <= '0';
      ELSIF ( and_dcpl_372 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_505_itm <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_506_itm <= '0';
      ELSIF ( and_dcpl_372 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_506_itm <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_507_itm <= '0';
      ELSIF ( and_dcpl_372 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_507_itm <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_508_itm <= '0';
      ELSIF ( and_dcpl_372 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_508_itm <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_509_itm <= '0';
      ELSIF ( and_dcpl_372 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_509_itm <= CONV_SL_1_1(operator_64_false_acc_cse_9_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_cse_10_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(not_tmp_698, or_2732_nl, fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_cse_10_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "1001")), 9), 10), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_acc_cse_10_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_2670_nl, (fsm_output(9)), or_2733_cse)) = '1' ) THEN
        operator_64_false_acc_cse_10_sva <= operator_64_false_acc_cse_10_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_37_itm <= '0';
      ELSIF ( not_tmp_706 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_37_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva_mx0w0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_371_itm <= '0';
      ELSIF ( not_tmp_706 = '0' ) THEN
        COMP_LOOP_nor_371_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva_mx0w0(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_372_itm <= '0';
      ELSIF ( not_tmp_706 = '0' ) THEN
        COMP_LOOP_nor_372_itm <= NOT((operator_64_false_acc_cse_10_sva_mx0w0(3))
            OR (operator_64_false_acc_cse_10_sva_mx0w0(2)) OR (operator_64_false_acc_cse_10_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_557_itm <= '0';
      ELSIF ( not_tmp_706 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_557_itm <= CONV_SL_1_1(operator_64_false_acc_cse_10_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_374_itm <= '0';
      ELSIF ( not_tmp_706 = '0' ) THEN
        COMP_LOOP_nor_374_itm <= NOT((operator_64_false_acc_cse_10_sva_mx0w0(3))
            OR (operator_64_false_acc_cse_10_sva_mx0w0(1)) OR (operator_64_false_acc_cse_10_sva_mx0w0(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_559_itm <= '0';
      ELSIF ( not_tmp_706 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_559_itm <= CONV_SL_1_1(operator_64_false_acc_cse_10_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_560_itm <= '0';
      ELSIF ( not_tmp_706 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_560_itm <= CONV_SL_1_1(operator_64_false_acc_cse_10_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_561_itm <= '0';
      ELSIF ( not_tmp_706 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_561_itm <= CONV_SL_1_1(operator_64_false_acc_cse_10_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_377_itm <= '0';
      ELSIF ( not_tmp_706 = '0' ) THEN
        COMP_LOOP_nor_377_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_10_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_563_itm <= '0';
      ELSIF ( not_tmp_706 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_563_itm <= CONV_SL_1_1(operator_64_false_acc_cse_10_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_564_itm <= '0';
      ELSIF ( not_tmp_706 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_564_itm <= CONV_SL_1_1(operator_64_false_acc_cse_10_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_565_itm <= '0';
      ELSIF ( not_tmp_706 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_565_itm <= CONV_SL_1_1(operator_64_false_acc_cse_10_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_566_itm <= '0';
      ELSIF ( not_tmp_706 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_566_itm <= CONV_SL_1_1(operator_64_false_acc_cse_10_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_567_itm <= '0';
      ELSIF ( not_tmp_706 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_567_itm <= CONV_SL_1_1(operator_64_false_acc_cse_10_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_568_itm <= '0';
      ELSIF ( not_tmp_706 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_568_itm <= CONV_SL_1_1(operator_64_false_acc_cse_10_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_569_itm <= '0';
      ELSIF ( not_tmp_706 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_569_itm <= CONV_SL_1_1(operator_64_false_acc_cse_10_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_11_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( (MUX_s_1_2_2(mux_2681_nl, and_tmp_32, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_11_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0(9
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & STD_LOGIC_VECTOR'( "101")), 8), 9), 9));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_acc_cse_11_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(not_tmp_698, or_2743_nl, fsm_output(9))) = '1' ) THEN
        operator_64_false_acc_cse_11_sva <= operator_64_false_acc_cse_11_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_41_itm <= '0';
        COMP_LOOP_nor_411_itm <= '0';
        COMP_LOOP_nor_412_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_617_itm <= '0';
        COMP_LOOP_nor_414_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_619_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_620_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_621_itm <= '0';
        COMP_LOOP_nor_417_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_623_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_624_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_625_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_626_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_627_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_628_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_629_itm <= '0';
      ELSIF ( mux_2688_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_41_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_11_sva_mx0w0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_411_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_11_sva_mx0w0(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_nor_412_itm <= NOT((operator_64_false_acc_cse_11_sva_mx0w0(3))
            OR (operator_64_false_acc_cse_11_sva_mx0w0(2)) OR (operator_64_false_acc_cse_11_sva_mx0w0(0)));
        COMP_LOOP_COMP_LOOP_and_617_itm <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_nor_414_itm <= NOT((operator_64_false_acc_cse_11_sva_mx0w0(3))
            OR (operator_64_false_acc_cse_11_sva_mx0w0(1)) OR (operator_64_false_acc_cse_11_sva_mx0w0(0)));
        COMP_LOOP_COMP_LOOP_and_619_itm <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_620_itm <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_621_itm <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_nor_417_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_11_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_623_itm <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_624_itm <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_625_itm <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_626_itm <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_627_itm <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_628_itm <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_629_itm <= CONV_SL_1_1(operator_64_false_acc_cse_11_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_cse_12_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(not_tmp_698, or_2748_nl, fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_cse_12_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "1011")), 9), 10), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_acc_cse_12_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_2692_nl, (fsm_output(9)), fsm_output(8))) = '1' )
          THEN
        operator_64_false_acc_cse_12_sva <= operator_64_false_acc_cse_12_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_45_itm <= '0';
        COMP_LOOP_nor_451_itm <= '0';
        COMP_LOOP_nor_452_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_677_itm <= '0';
        COMP_LOOP_nor_454_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_679_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_680_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_681_itm <= '0';
        COMP_LOOP_nor_457_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_683_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_684_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_685_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_686_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_687_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_688_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_689_itm <= '0';
      ELSIF ( mux_2703_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_45_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_12_sva_mx0w0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_451_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_12_sva_mx0w0(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_nor_452_itm <= NOT((operator_64_false_acc_cse_12_sva_mx0w0(3))
            OR (operator_64_false_acc_cse_12_sva_mx0w0(2)) OR (operator_64_false_acc_cse_12_sva_mx0w0(0)));
        COMP_LOOP_COMP_LOOP_and_677_itm <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_nor_454_itm <= NOT((operator_64_false_acc_cse_12_sva_mx0w0(3))
            OR (operator_64_false_acc_cse_12_sva_mx0w0(1)) OR (operator_64_false_acc_cse_12_sva_mx0w0(0)));
        COMP_LOOP_COMP_LOOP_and_679_itm <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_680_itm <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_681_itm <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_nor_457_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_12_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_683_itm <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_684_itm <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_685_itm <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_686_itm <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_687_itm <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_688_itm <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_689_itm <= CONV_SL_1_1(operator_64_false_acc_cse_12_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_12_psp_sva <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( (MUX_s_1_2_2(mux_2708_nl, (fsm_output(9)), fsm_output(8))) = '1' )
          THEN
        COMP_LOOP_acc_12_psp_sva <= z_out_2(7 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_acc_cse_13_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_2713_nl, (fsm_output(9)), fsm_output(8))) = '1' )
          THEN
        operator_64_false_acc_cse_13_sva <= operator_64_false_acc_cse_13_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_49_itm <= '0';
        COMP_LOOP_nor_491_itm <= '0';
        COMP_LOOP_nor_492_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_737_itm <= '0';
        COMP_LOOP_nor_494_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_739_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_740_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_741_itm <= '0';
        COMP_LOOP_nor_497_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_743_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_744_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_745_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_746_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_747_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_748_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_749_itm <= '0';
      ELSIF ( mux_2715_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_49_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_13_sva_mx0w0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_491_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_13_sva_mx0w0(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_nor_492_itm <= NOT((operator_64_false_acc_cse_13_sva_mx0w0(3))
            OR (operator_64_false_acc_cse_13_sva_mx0w0(2)) OR (operator_64_false_acc_cse_13_sva_mx0w0(0)));
        COMP_LOOP_COMP_LOOP_and_737_itm <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_nor_494_itm <= NOT((operator_64_false_acc_cse_13_sva_mx0w0(3))
            OR (operator_64_false_acc_cse_13_sva_mx0w0(1)) OR (operator_64_false_acc_cse_13_sva_mx0w0(0)));
        COMP_LOOP_COMP_LOOP_and_739_itm <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_740_itm <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_741_itm <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_nor_497_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_13_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_743_itm <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_744_itm <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_745_itm <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_746_itm <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_747_itm <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_748_itm <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_749_itm <= CONV_SL_1_1(operator_64_false_acc_cse_13_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_cse_14_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(not_tmp_698, and_410_nl, fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_cse_14_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "1101")), 9), 10), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_acc_cse_14_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_2722_nl, nor_tmp_130, or_111_cse)) = '1' ) THEN
        operator_64_false_acc_cse_14_sva <= operator_64_false_acc_cse_14_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_53_itm <= '0';
        COMP_LOOP_nor_531_itm <= '0';
        COMP_LOOP_nor_532_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_797_itm <= '0';
        COMP_LOOP_nor_534_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_799_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_800_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_801_itm <= '0';
        COMP_LOOP_nor_537_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_803_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_804_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_805_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_806_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_807_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_808_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_809_itm <= '0';
      ELSIF ( mux_2727_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_53_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_14_sva_mx0w0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_531_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_14_sva_mx0w0(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_nor_532_itm <= NOT((operator_64_false_acc_cse_14_sva_mx0w0(3))
            OR (operator_64_false_acc_cse_14_sva_mx0w0(2)) OR (operator_64_false_acc_cse_14_sva_mx0w0(0)));
        COMP_LOOP_COMP_LOOP_and_797_itm <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_nor_534_itm <= NOT((operator_64_false_acc_cse_14_sva_mx0w0(3))
            OR (operator_64_false_acc_cse_14_sva_mx0w0(1)) OR (operator_64_false_acc_cse_14_sva_mx0w0(0)));
        COMP_LOOP_COMP_LOOP_and_799_itm <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_800_itm <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_801_itm <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_nor_537_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_14_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_803_itm <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_804_itm <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_805_itm <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_806_itm <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_807_itm <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_808_itm <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_809_itm <= CONV_SL_1_1(operator_64_false_acc_cse_14_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_13_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( mux_2730_nl = '0' ) THEN
        COMP_LOOP_acc_13_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0(9
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & STD_LOGIC_VECTOR'( "111")), 8), 9), 9));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_acc_cse_15_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( mux_2733_nl = '0' ) THEN
        operator_64_false_acc_cse_15_sva <= operator_64_false_acc_cse_15_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_57_itm <= '0';
        COMP_LOOP_nor_571_itm <= '0';
        COMP_LOOP_nor_572_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_857_itm <= '0';
        COMP_LOOP_nor_574_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_859_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_860_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_861_itm <= '0';
        COMP_LOOP_nor_577_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_863_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_864_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_865_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_866_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_867_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_868_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_869_itm <= '0';
      ELSIF ( mux_2734_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_57_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva_mx0w0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_571_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva_mx0w0(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_nor_572_itm <= NOT((operator_64_false_acc_cse_15_sva_mx0w0(3))
            OR (operator_64_false_acc_cse_15_sva_mx0w0(2)) OR (operator_64_false_acc_cse_15_sva_mx0w0(0)));
        COMP_LOOP_COMP_LOOP_and_857_itm <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_nor_574_itm <= NOT((operator_64_false_acc_cse_15_sva_mx0w0(3))
            OR (operator_64_false_acc_cse_15_sva_mx0w0(1)) OR (operator_64_false_acc_cse_15_sva_mx0w0(0)));
        COMP_LOOP_COMP_LOOP_and_859_itm <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_860_itm <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_861_itm <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_nor_577_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_15_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_863_itm <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_864_itm <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_865_itm <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_866_itm <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_867_itm <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_868_itm <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_869_itm <= CONV_SL_1_1(operator_64_false_acc_cse_15_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_cse_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(not_tmp_698, and_413_nl, fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_cse_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_VEC_LOOP_j_sva_9_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "1111")), 9), 10), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_acc_cse_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(not_tmp_698, and_414_nl, fsm_output(9))) = '1' ) THEN
        operator_64_false_acc_cse_sva <= operator_64_false_acc_cse_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_61_itm <= '0';
        COMP_LOOP_nor_611_itm <= '0';
        COMP_LOOP_nor_612_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_917_itm <= '0';
        COMP_LOOP_nor_614_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_919_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_920_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_921_itm <= '0';
        COMP_LOOP_nor_617_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_923_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_924_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_925_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_926_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_927_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_928_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_929_itm <= '0';
      ELSIF ( mux_2745_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_61_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_sva_mx0w0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_611_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_sva_mx0w0(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_nor_612_itm <= NOT((operator_64_false_acc_cse_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_sva_mx0w0(2)) OR (operator_64_false_acc_cse_sva_mx0w0(0)));
        COMP_LOOP_COMP_LOOP_and_917_itm <= CONV_SL_1_1(operator_64_false_acc_cse_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_nor_614_itm <= NOT((operator_64_false_acc_cse_sva_mx0w0(3)) OR
            (operator_64_false_acc_cse_sva_mx0w0(1)) OR (operator_64_false_acc_cse_sva_mx0w0(0)));
        COMP_LOOP_COMP_LOOP_and_919_itm <= CONV_SL_1_1(operator_64_false_acc_cse_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_920_itm <= CONV_SL_1_1(operator_64_false_acc_cse_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_921_itm <= CONV_SL_1_1(operator_64_false_acc_cse_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_nor_617_itm <= NOT(CONV_SL_1_1(operator_64_false_acc_cse_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_923_itm <= CONV_SL_1_1(operator_64_false_acc_cse_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_924_itm <= CONV_SL_1_1(operator_64_false_acc_cse_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_925_itm <= CONV_SL_1_1(operator_64_false_acc_cse_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_926_itm <= CONV_SL_1_1(operator_64_false_acc_cse_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_927_itm <= CONV_SL_1_1(operator_64_false_acc_cse_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_928_itm <= CONV_SL_1_1(operator_64_false_acc_cse_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_929_itm <= CONV_SL_1_1(operator_64_false_acc_cse_sva_mx0w0(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_64_false_slc_operator_64_false_acc_1_60_itm <= '0';
      ELSIF ( (and_dcpl_98 OR operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c1
          OR operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c2 OR operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c3
          OR operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c4) = '1' )
          THEN
        operator_64_false_slc_operator_64_false_acc_1_60_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_11_nl,
            (z_out_2(61)), (COMP_LOOP_slc_acc_3_12_1_slc(11)), (z_out_2(59)), STD_LOGIC_VECTOR'(
            and_dcpl_98 & COMP_LOOP_or_35_nl & operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c2
            & operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c4));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (tmp_1_lpi_4_dfm_mx0c0 OR and_dcpl_245 OR and_dcpl_249 OR and_dcpl_254
          OR and_dcpl_258 OR and_dcpl_262 OR and_dcpl_265 OR and_dcpl_269 OR and_dcpl_271
          OR and_dcpl_273 OR and_dcpl_276 OR and_dcpl_278 OR and_dcpl_283 OR and_dcpl_285
          OR and_dcpl_287 OR and_dcpl_289) = '1' ) THEN
        tmp_1_lpi_4_dfm <= MUX1HOT_v_64_16_2(vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d,
            vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d, vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d,
            vec_rsc_0_6_i_qa_d, vec_rsc_0_7_i_qa_d, vec_rsc_0_8_i_qa_d, vec_rsc_0_9_i_qa_d,
            vec_rsc_0_10_i_qa_d, vec_rsc_0_11_i_qa_d, vec_rsc_0_12_i_qa_d, vec_rsc_0_13_i_qa_d,
            vec_rsc_0_14_i_qa_d, vec_rsc_0_15_i_qa_d, STD_LOGIC_VECTOR'( COMP_LOOP_or_18_nl
            & COMP_LOOP_or_19_nl & COMP_LOOP_or_20_nl & COMP_LOOP_or_21_nl & COMP_LOOP_or_22_nl
            & COMP_LOOP_or_23_nl & COMP_LOOP_or_24_nl & COMP_LOOP_or_25_nl & COMP_LOOP_or_26_nl
            & COMP_LOOP_or_27_nl & COMP_LOOP_or_28_nl & COMP_LOOP_or_29_nl & COMP_LOOP_or_30_nl
            & COMP_LOOP_or_31_nl & COMP_LOOP_or_32_nl & COMP_LOOP_or_33_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mux_2797_itm = '1' ) THEN
        modExp_dev_exp_1_sva_8_4 <= MUX_v_5_2_2((z_out_3(8 DOWNTO 4)), COMP_LOOP_k_9_4_sva_4_0,
            mux_2336_itm);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_2893_nl, mux_2884_nl, fsm_output(8))) = '1' ) THEN
        modExp_dev_exp_1_sva_63_9 <= MUX_v_55_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000000000000000000"),
            (z_out_3(63 DOWNTO 9)), not_7089_nl);
      END IF;
    END IF;
  END PROCESS;
  or_2479_nl <= (fsm_output(2)) OR not_tmp_572;
  mux_2317_nl <= MUX_s_1_2_2(not_tmp_572, or_2733_cse, fsm_output(2));
  mux_2318_nl <= MUX_s_1_2_2(or_2479_nl, mux_2317_nl, fsm_output(1));
  mux_2319_nl <= MUX_s_1_2_2(mux_2318_nl, or_tmp_2391, fsm_output(5));
  mux_2320_nl <= MUX_s_1_2_2(mux_2319_nl, mux_tmp_2244, fsm_output(6));
  mux_2314_nl <= MUX_s_1_2_2(or_tmp_2402, or_tmp_2401, fsm_output(1));
  nand_177_nl <= NOT((and_515_cse OR (fsm_output(2))) AND CONV_SL_1_1(fsm_output(8
      DOWNTO 7)=STD_LOGIC_VECTOR'("11")));
  mux_2315_nl <= MUX_s_1_2_2(mux_2314_nl, nand_177_nl, fsm_output(5));
  or_2477_nl <= and_516_cse OR not_tmp_572;
  mux_2313_nl <= MUX_s_1_2_2(or_tmp_2324, or_2477_nl, fsm_output(5));
  mux_2316_nl <= MUX_s_1_2_2(mux_2315_nl, mux_2313_nl, fsm_output(6));
  mux_2321_nl <= MUX_s_1_2_2(mux_2320_nl, mux_2316_nl, fsm_output(4));
  or_2476_nl <= and_516_cse OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_2310_nl <= MUX_s_1_2_2((fsm_output(7)), or_2476_nl, fsm_output(5));
  nand_178_nl <= NOT((fsm_output(2)) AND (fsm_output(8)) AND (fsm_output(7)));
  mux_2309_nl <= MUX_s_1_2_2(mux_tmp_2247, nand_178_nl, fsm_output(5));
  mux_2311_nl <= MUX_s_1_2_2(mux_2310_nl, mux_2309_nl, fsm_output(6));
  mux_2307_nl <= MUX_s_1_2_2(or_tmp_2324, or_tmp_2409, fsm_output(5));
  mux_2306_nl <= MUX_s_1_2_2(mux_tmp_2250, or_tmp_2406, fsm_output(5));
  mux_2308_nl <= MUX_s_1_2_2(mux_2307_nl, mux_2306_nl, fsm_output(6));
  mux_2312_nl <= MUX_s_1_2_2(mux_2311_nl, mux_2308_nl, fsm_output(4));
  mux_2322_nl <= MUX_s_1_2_2(mux_2321_nl, mux_2312_nl, fsm_output(3));
  mux_2302_nl <= MUX_s_1_2_2(or_tmp_2409, mux_tmp_2250, fsm_output(5));
  mux_2300_nl <= MUX_s_1_2_2(or_tmp_2406, or_2733_cse, fsm_output(5));
  mux_2303_nl <= MUX_s_1_2_2(mux_2302_nl, mux_2300_nl, fsm_output(6));
  or_2468_nl <= (fsm_output(5)) OR mux_tmp_2247;
  mux_2299_nl <= MUX_s_1_2_2(or_2468_nl, or_tmp_2395, fsm_output(6));
  mux_2304_nl <= MUX_s_1_2_2(mux_2303_nl, mux_2299_nl, fsm_output(4));
  or_2461_nl <= (fsm_output(5)) OR (fsm_output(2)) OR (NOT (fsm_output(8))) OR (fsm_output(7));
  mux_2296_nl <= MUX_s_1_2_2(mux_tmp_2244, or_2461_nl, fsm_output(6));
  mux_2292_nl <= MUX_s_1_2_2(or_tmp_2393, or_tmp_2391, fsm_output(1));
  or_2455_nl <= (NOT(and_515_cse OR (fsm_output(2)))) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 7)/=STD_LOGIC_VECTOR'("10"));
  mux_2293_nl <= MUX_s_1_2_2(mux_2292_nl, or_2455_nl, fsm_output(5));
  mux_2294_nl <= MUX_s_1_2_2(or_tmp_2395, mux_2293_nl, fsm_output(6));
  mux_2297_nl <= MUX_s_1_2_2(mux_2296_nl, mux_2294_nl, fsm_output(4));
  mux_2305_nl <= MUX_s_1_2_2(mux_2304_nl, mux_2297_nl, fsm_output(3));
  mux_2323_nl <= MUX_s_1_2_2(mux_2322_nl, mux_2305_nl, fsm_output(9));
  nor_549_nl <= NOT((fsm_output(2)) OR (fsm_output(5)) OR (fsm_output(7)) OR (fsm_output(8))
      OR (fsm_output(9)));
  and_511_nl <= (fsm_output(2)) AND (fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(8))
      AND (fsm_output(9));
  mux_2337_nl <= MUX_s_1_2_2(nor_549_nl, and_511_nl, or_2500_cse);
  and_512_nl <= (fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(8)) AND (fsm_output(9));
  mux_2338_nl <= MUX_s_1_2_2(mux_2337_nl, and_512_nl, or_602_cse);
  and_513_nl <= CONV_SL_1_1(fsm_output(9 DOWNTO 7)=STD_LOGIC_VECTOR'("111"));
  mux_2339_nl <= MUX_s_1_2_2(mux_2338_nl, and_513_nl, fsm_output(6));
  nor_548_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 1)/=STD_LOGIC_VECTOR'("00000000")));
  operator_64_false_or_2_nl <= and_dcpl_290 OR COMP_LOOP_10_modExp_dev_1_while_mul_mut_mx0c5
      OR (NOT mux_2336_itm);
  nor_524_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 4)/=STD_LOGIC_VECTOR'("00000")));
  mux_2427_nl <= MUX_s_1_2_2(nor_524_nl, and_tmp_24, fsm_output(9));
  and_331_nl <= and_dcpl_239 AND and_dcpl_106;
  COMP_LOOP_or_2_nl <= (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_240) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_332_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_335_m1c) OR (COMP_LOOP_COMP_LOOP_and_72_itm AND and_338_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_340_m1c) OR (COMP_LOOP_COMP_LOOP_and_70_itm AND and_342_m1c) OR (COMP_LOOP_COMP_LOOP_and_69_itm
      AND and_344_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_346_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_348_m1c) OR (COMP_LOOP_COMP_LOOP_and_66_itm AND and_350_m1c) OR (COMP_LOOP_COMP_LOOP_and_65_itm
      AND and_351_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_352_m1c) OR (COMP_LOOP_COMP_LOOP_and_185_itm
      AND and_354_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_356_m1c) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_358_m1c);
  COMP_LOOP_or_3_nl <= (COMP_LOOP_COMP_LOOP_and_244_itm AND and_dcpl_240) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_332_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_335_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_338_m1c) OR (COMP_LOOP_COMP_LOOP_and_72_itm
      AND and_340_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_342_m1c) OR (COMP_LOOP_COMP_LOOP_and_70_itm
      AND and_344_m1c) OR (COMP_LOOP_COMP_LOOP_and_69_itm AND and_346_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_348_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_350_m1c) OR (COMP_LOOP_COMP_LOOP_and_66_itm
      AND and_351_m1c) OR (COMP_LOOP_COMP_LOOP_and_65_itm AND and_352_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_354_m1c) OR (COMP_LOOP_COMP_LOOP_and_185_itm AND and_356_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_358_m1c);
  COMP_LOOP_or_4_nl <= (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_240) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_332_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_335_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_338_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_340_m1c) OR (COMP_LOOP_COMP_LOOP_and_72_itm AND and_342_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_344_m1c) OR (COMP_LOOP_COMP_LOOP_and_70_itm AND and_346_m1c) OR (COMP_LOOP_COMP_LOOP_and_69_itm
      AND and_348_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_350_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_351_m1c) OR (COMP_LOOP_COMP_LOOP_and_66_itm AND and_352_m1c) OR (COMP_LOOP_COMP_LOOP_and_65_itm
      AND and_354_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_356_m1c) OR (COMP_LOOP_COMP_LOOP_and_185_itm
      AND and_358_m1c);
  COMP_LOOP_or_5_nl <= (COMP_LOOP_COMP_LOOP_and_185_itm AND and_dcpl_240) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_332_m1c) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_335_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_338_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_340_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_342_m1c) OR (COMP_LOOP_COMP_LOOP_and_72_itm
      AND and_344_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_346_m1c) OR (COMP_LOOP_COMP_LOOP_and_70_itm
      AND and_348_m1c) OR (COMP_LOOP_COMP_LOOP_and_69_itm AND and_350_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_351_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_352_m1c) OR (COMP_LOOP_COMP_LOOP_and_66_itm
      AND and_354_m1c) OR (COMP_LOOP_COMP_LOOP_and_65_itm AND and_356_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_358_m1c);
  COMP_LOOP_or_6_nl <= (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_240) OR (COMP_LOOP_COMP_LOOP_and_185_itm
      AND and_332_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_335_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_338_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_340_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_342_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_344_m1c) OR (COMP_LOOP_COMP_LOOP_and_72_itm AND and_346_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_348_m1c) OR (COMP_LOOP_COMP_LOOP_and_70_itm AND and_350_m1c) OR (COMP_LOOP_COMP_LOOP_and_69_itm
      AND and_351_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_352_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_354_m1c) OR (COMP_LOOP_COMP_LOOP_and_66_itm AND and_356_m1c) OR (COMP_LOOP_COMP_LOOP_and_65_itm
      AND and_358_m1c);
  COMP_LOOP_or_7_nl <= (COMP_LOOP_COMP_LOOP_and_65_itm AND and_dcpl_240) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_332_m1c) OR (COMP_LOOP_COMP_LOOP_and_185_itm AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_335_m1c) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_338_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_340_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_342_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_344_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_346_m1c) OR (COMP_LOOP_COMP_LOOP_and_72_itm
      AND and_348_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_350_m1c) OR (COMP_LOOP_COMP_LOOP_and_70_itm
      AND and_351_m1c) OR (COMP_LOOP_COMP_LOOP_and_69_itm AND and_352_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_354_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_356_m1c) OR (COMP_LOOP_COMP_LOOP_and_66_itm
      AND and_358_m1c);
  COMP_LOOP_or_8_nl <= (COMP_LOOP_COMP_LOOP_and_66_itm AND and_dcpl_240) OR (COMP_LOOP_COMP_LOOP_and_65_itm
      AND and_332_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_185_itm
      AND and_335_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_338_m1c) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_340_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_342_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_344_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_346_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_348_m1c) OR (COMP_LOOP_COMP_LOOP_and_72_itm AND and_350_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_351_m1c) OR (COMP_LOOP_COMP_LOOP_and_70_itm AND and_352_m1c) OR (COMP_LOOP_COMP_LOOP_and_69_itm
      AND and_354_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_356_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_358_m1c);
  COMP_LOOP_or_9_nl <= (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_240) OR (COMP_LOOP_COMP_LOOP_and_66_itm
      AND and_332_m1c) OR (COMP_LOOP_COMP_LOOP_and_65_itm AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_335_m1c) OR (COMP_LOOP_COMP_LOOP_and_185_itm AND and_338_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_340_m1c) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_342_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_344_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_346_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_348_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_350_m1c) OR (COMP_LOOP_COMP_LOOP_and_72_itm
      AND and_351_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_352_m1c) OR (COMP_LOOP_COMP_LOOP_and_70_itm
      AND and_354_m1c) OR (COMP_LOOP_COMP_LOOP_and_69_itm AND and_356_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_358_m1c);
  COMP_LOOP_or_10_nl <= (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_240) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_332_m1c) OR (COMP_LOOP_COMP_LOOP_and_66_itm AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_65_itm
      AND and_335_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_338_m1c) OR (COMP_LOOP_COMP_LOOP_and_185_itm
      AND and_340_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_342_m1c) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_344_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_346_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_348_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_350_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_351_m1c) OR (COMP_LOOP_COMP_LOOP_and_72_itm AND and_352_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_354_m1c) OR (COMP_LOOP_COMP_LOOP_and_70_itm AND and_356_m1c) OR (COMP_LOOP_COMP_LOOP_and_69_itm
      AND and_358_m1c);
  COMP_LOOP_or_11_nl <= (COMP_LOOP_COMP_LOOP_and_69_itm AND and_dcpl_240) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_332_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_66_itm
      AND and_335_m1c) OR (COMP_LOOP_COMP_LOOP_and_65_itm AND and_338_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_340_m1c) OR (COMP_LOOP_COMP_LOOP_and_185_itm AND and_342_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_344_m1c) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_346_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_348_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_350_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_351_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_352_m1c) OR (COMP_LOOP_COMP_LOOP_and_72_itm
      AND and_354_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_356_m1c) OR (COMP_LOOP_COMP_LOOP_and_70_itm
      AND and_358_m1c);
  COMP_LOOP_or_12_nl <= (COMP_LOOP_COMP_LOOP_and_70_itm AND and_dcpl_240) OR (COMP_LOOP_COMP_LOOP_and_69_itm
      AND and_332_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_335_m1c) OR (COMP_LOOP_COMP_LOOP_and_66_itm AND and_338_m1c) OR (COMP_LOOP_COMP_LOOP_and_65_itm
      AND and_340_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_342_m1c) OR (COMP_LOOP_COMP_LOOP_and_185_itm
      AND and_344_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_346_m1c) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_348_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_350_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_351_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_352_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_354_m1c) OR (COMP_LOOP_COMP_LOOP_and_72_itm AND and_356_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_358_m1c);
  COMP_LOOP_or_13_nl <= (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_240) OR (COMP_LOOP_COMP_LOOP_and_70_itm
      AND and_332_m1c) OR (COMP_LOOP_COMP_LOOP_and_69_itm AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_335_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_338_m1c) OR (COMP_LOOP_COMP_LOOP_and_66_itm
      AND and_340_m1c) OR (COMP_LOOP_COMP_LOOP_and_65_itm AND and_342_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_344_m1c) OR (COMP_LOOP_COMP_LOOP_and_185_itm AND and_346_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_348_m1c) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_350_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_351_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_352_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_354_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_356_m1c) OR (COMP_LOOP_COMP_LOOP_and_72_itm
      AND and_358_m1c);
  COMP_LOOP_or_14_nl <= (COMP_LOOP_COMP_LOOP_and_72_itm AND and_dcpl_240) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_332_m1c) OR (COMP_LOOP_COMP_LOOP_and_70_itm AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_69_itm
      AND and_335_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_338_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_340_m1c) OR (COMP_LOOP_COMP_LOOP_and_66_itm AND and_342_m1c) OR (COMP_LOOP_COMP_LOOP_and_65_itm
      AND and_344_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_346_m1c) OR (COMP_LOOP_COMP_LOOP_and_185_itm
      AND and_348_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_350_m1c) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_351_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_352_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_354_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_356_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_358_m1c);
  COMP_LOOP_or_15_nl <= (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_240) OR (COMP_LOOP_COMP_LOOP_and_72_itm
      AND and_332_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_70_itm
      AND and_335_m1c) OR (COMP_LOOP_COMP_LOOP_and_69_itm AND and_338_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_340_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_342_m1c) OR (COMP_LOOP_COMP_LOOP_and_66_itm
      AND and_344_m1c) OR (COMP_LOOP_COMP_LOOP_and_65_itm AND and_346_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_348_m1c) OR (COMP_LOOP_COMP_LOOP_and_185_itm AND and_350_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_351_m1c) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_352_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_354_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_356_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_358_m1c);
  COMP_LOOP_or_16_nl <= (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_240) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_332_m1c) OR (COMP_LOOP_COMP_LOOP_and_72_itm AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_335_m1c) OR (COMP_LOOP_COMP_LOOP_and_70_itm AND and_338_m1c) OR (COMP_LOOP_COMP_LOOP_and_69_itm
      AND and_340_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_342_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_344_m1c) OR (COMP_LOOP_COMP_LOOP_and_66_itm AND and_346_m1c) OR (COMP_LOOP_COMP_LOOP_and_65_itm
      AND and_348_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_350_m1c) OR (COMP_LOOP_COMP_LOOP_and_185_itm
      AND and_351_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_352_m1c) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_354_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_356_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_358_m1c);
  COMP_LOOP_or_17_nl <= (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_240) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_332_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_72_itm
      AND and_335_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_338_m1c) OR (COMP_LOOP_COMP_LOOP_and_70_itm
      AND and_340_m1c) OR (COMP_LOOP_COMP_LOOP_and_69_itm AND and_342_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_344_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_346_m1c) OR (COMP_LOOP_COMP_LOOP_and_66_itm
      AND and_348_m1c) OR (COMP_LOOP_COMP_LOOP_and_65_itm AND and_350_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_351_m1c) OR (COMP_LOOP_COMP_LOOP_and_185_itm AND and_352_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_354_m1c) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_356_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_358_m1c);
  mux_2470_nl <= MUX_s_1_2_2(and_dcpl_146, or_tmp_33, and_516_cse);
  mux_2471_nl <= MUX_s_1_2_2((NOT mux_2470_nl), and_711_cse, fsm_output(5));
  or_2622_nl <= (NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(3));
  mux_2469_nl <= MUX_s_1_2_2(or_2622_nl, or_307_cse, fsm_output(1));
  or_2623_nl <= (fsm_output(5)) OR (NOT mux_2469_nl);
  mux_2472_nl <= MUX_s_1_2_2(mux_2471_nl, or_2623_nl, fsm_output(4));
  mux_2465_nl <= MUX_s_1_2_2(and_dcpl_146, (fsm_output(3)), fsm_output(2));
  mux_2464_nl <= MUX_s_1_2_2(and_dcpl_146, or_tmp_33, fsm_output(2));
  mux_2466_nl <= MUX_s_1_2_2(mux_2465_nl, mux_2464_nl, fsm_output(1));
  mux_2467_nl <= MUX_s_1_2_2((NOT mux_2466_nl), nor_tmp_403, fsm_output(5));
  mux_2468_nl <= MUX_s_1_2_2(mux_2467_nl, or_tmp_2551, fsm_output(4));
  mux_2473_nl <= MUX_s_1_2_2(mux_2472_nl, mux_2468_nl, fsm_output(0));
  mux_2461_nl <= MUX_s_1_2_2((NOT nor_tmp_399), nor_tmp_403, fsm_output(5));
  mux_2462_nl <= MUX_s_1_2_2((NOT or_tmp_2552), mux_2461_nl, fsm_output(4));
  mux_2463_nl <= MUX_s_1_2_2(mux_tmp_2389, mux_2462_nl, fsm_output(0));
  mux_2474_nl <= MUX_s_1_2_2(mux_2473_nl, (NOT mux_2463_nl), fsm_output(7));
  or_2621_nl <= (fsm_output(5)) OR (NOT or_tmp_2549);
  mux_2458_nl <= MUX_s_1_2_2(mux_tmp_2381, or_2621_nl, fsm_output(4));
  mux_2459_nl <= MUX_s_1_2_2(mux_tmp_2382, mux_2458_nl, fsm_output(0));
  mux_2455_nl <= MUX_s_1_2_2(or_tmp_2439, (NOT or_307_cse), fsm_output(5));
  mux_2454_nl <= MUX_s_1_2_2((NOT nor_tmp_1), nor_tmp_403, fsm_output(5));
  mux_2456_nl <= MUX_s_1_2_2(mux_2455_nl, mux_2454_nl, fsm_output(4));
  mux_2452_nl <= MUX_s_1_2_2((NOT nor_tmp_1), mux_tmp_2400, fsm_output(5));
  mux_2453_nl <= MUX_s_1_2_2((NOT mux_tmp_2380), mux_2452_nl, fsm_output(4));
  mux_2457_nl <= MUX_s_1_2_2(mux_2456_nl, mux_2453_nl, fsm_output(0));
  mux_2460_nl <= MUX_s_1_2_2((NOT mux_2459_nl), mux_2457_nl, fsm_output(7));
  mux_2475_nl <= MUX_s_1_2_2(mux_2474_nl, mux_2460_nl, fsm_output(8));
  mux_2446_nl <= MUX_s_1_2_2(not_tmp_617, nor_tmp_399, fsm_output(5));
  mux_2447_nl <= MUX_s_1_2_2(mux_2446_nl, or_tmp_2552, fsm_output(4));
  mux_2444_nl <= MUX_s_1_2_2(not_tmp_617, and_711_cse, fsm_output(5));
  mux_2445_nl <= MUX_s_1_2_2(mux_2444_nl, or_tmp_2551, fsm_output(4));
  mux_2448_nl <= MUX_s_1_2_2(mux_2447_nl, mux_2445_nl, fsm_output(0));
  mux_2441_nl <= MUX_s_1_2_2(and_dcpl_95, or_tmp_2549, fsm_output(5));
  mux_2442_nl <= MUX_s_1_2_2((NOT mux_2441_nl), mux_tmp_2381, fsm_output(4));
  mux_2443_nl <= MUX_s_1_2_2(mux_2442_nl, mux_tmp_2389, fsm_output(0));
  mux_2449_nl <= MUX_s_1_2_2(mux_2448_nl, (NOT mux_2443_nl), fsm_output(7));
  mux_2434_nl <= MUX_s_1_2_2(not_tmp_617, nor_tmp_1, fsm_output(5));
  mux_2435_nl <= MUX_s_1_2_2(mux_2434_nl, mux_tmp_2380, fsm_output(4));
  mux_2436_nl <= MUX_s_1_2_2(mux_2435_nl, mux_tmp_2382, fsm_output(0));
  mux_2437_nl <= MUX_s_1_2_2((NOT mux_2436_nl), or_tmp_2548, fsm_output(7));
  mux_2450_nl <= MUX_s_1_2_2(mux_2449_nl, mux_2437_nl, fsm_output(8));
  COMP_LOOP_COMP_LOOP_and_17_nl <= CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
  modExp_dev_while_or_nl <= and_dcpl_290 OR (NOT mux_2336_itm);
  modExp_dev_while_or_1_nl <= COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c3
      OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c4 OR
      COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c5 OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c6
      OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c7 OR
      COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c8 OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c9
      OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c10 OR
      COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c11 OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c12
      OR COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm_mx0c13;
  nand_486_nl <= NOT(and_dcpl_294 AND and_dcpl_346);
  nor_nl <= NOT((fsm_output(1)) OR (fsm_output(7)) OR (NOT (fsm_output(0))) OR (NOT
      (fsm_output(4))) OR (fsm_output(9)) OR (fsm_output(8)));
  nor_1038_nl <= NOT((NOT (fsm_output(1))) OR (NOT (fsm_output(7))) OR (fsm_output(0))
      OR (fsm_output(4)) OR nand_490_cse);
  mux_2864_nl <= MUX_s_1_2_2(nor_nl, nor_1038_nl, fsm_output(2));
  and_421_nl <= and_dcpl_109 AND and_dcpl_346;
  and_422_nl <= and_dcpl_239 AND and_dcpl_256;
  and_423_nl <= and_dcpl_244 AND and_dcpl_307;
  and_424_nl <= and_dcpl_248 AND and_dcpl_263;
  and_425_nl <= and_dcpl_253 AND and_dcpl_260;
  and_426_nl <= and_dcpl_257 AND and_dcpl_313;
  and_427_nl <= and_dcpl_261 AND and_dcpl_319;
  and_428_nl <= and_dcpl_264 AND and_dcpl_317;
  and_429_nl <= and_dcpl_268 AND and_dcpl_323;
  and_430_nl <= and_dcpl_244 AND and_dcpl_321;
  and_431_nl <= and_dcpl_239 AND and_dcpl_284;
  and_432_nl <= and_dcpl_275 AND and_dcpl_279;
  and_433_nl <= and_dcpl_248 AND and_dcpl_288;
  and_434_nl <= and_dcpl_282 AND and_dcpl_331;
  operator_64_false_mux1h_nl <= MUX1HOT_v_4_16_2((z_out_3(3 DOWNTO 0)), (COMP_LOOP_acc_psp_sva(3
      DOWNTO 0)), STD_LOGIC_VECTOR'( "0001"), STD_LOGIC_VECTOR'( "0010"), STD_LOGIC_VECTOR'(
      "0011"), STD_LOGIC_VECTOR'( "0100"), STD_LOGIC_VECTOR'( "0101"), STD_LOGIC_VECTOR'(
      "0110"), STD_LOGIC_VECTOR'( "0111"), STD_LOGIC_VECTOR'( "1000"), STD_LOGIC_VECTOR'(
      "1001"), STD_LOGIC_VECTOR'( "1010"), STD_LOGIC_VECTOR'( "1011"), STD_LOGIC_VECTOR'(
      "1100"), STD_LOGIC_VECTOR'( "1101"), STD_LOGIC_VECTOR'( "1110"), STD_LOGIC_VECTOR'(
      (NOT mux_2336_itm) & (NOT mux_2797_itm) & and_421_nl & and_422_nl & and_423_nl
      & and_424_nl & and_425_nl & and_426_nl & and_427_nl & and_428_nl & and_429_nl
      & and_430_nl & and_431_nl & and_432_nl & and_433_nl & and_434_nl));
  COMP_LOOP_nand_nl <= NOT(and_dcpl_268 AND and_dcpl_106);
  operator_64_false_and_nl <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), operator_64_false_mux1h_nl,
      COMP_LOOP_nand_nl);
  and_435_nl <= and_dcpl_257 AND and_dcpl_329;
  operator_64_false_or_2_nl_1 <= MUX_v_4_2_2(operator_64_false_and_nl, STD_LOGIC_VECTOR'("1111"),
      and_435_nl);
  operator_64_false_1_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & (NOT
      COMP_LOOP_k_9_4_sva_4_0)) + UNSIGNED'( "000001"), 6));
  mux_2587_nl <= MUX_s_1_2_2(or_tmp_2548, or_tmp, fsm_output(0));
  or_2696_nl <= (fsm_output(7)) OR mux_2587_nl;
  mux_2590_nl <= MUX_s_1_2_2(not_tmp_664, or_2696_nl, fsm_output(8));
  or_2699_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00"));
  mux_2591_nl <= MUX_s_1_2_2(nor_tmp_1, (fsm_output(6)), or_2699_nl);
  mux_2592_nl <= MUX_s_1_2_2(mux_tmp_2538, (NOT mux_2591_nl), fsm_output(7));
  mux_2597_nl <= MUX_s_1_2_2(mux_tmp_2468, (fsm_output(6)), fsm_output(5));
  mux_2598_nl <= MUX_s_1_2_2(mux_156_cse, mux_2597_nl, fsm_output(4));
  mux_2593_nl <= MUX_s_1_2_2(and_dcpl_95, and_711_cse, or_2700_cse);
  mux_2594_nl <= MUX_s_1_2_2(mux_2593_nl, (fsm_output(6)), fsm_output(5));
  mux_2596_nl <= MUX_s_1_2_2(mux_156_cse, mux_2594_nl, fsm_output(4));
  mux_2599_nl <= MUX_s_1_2_2(mux_2598_nl, mux_2596_nl, fsm_output(0));
  or_2701_nl <= CONV_SL_1_1(fsm_output(6 DOWNTO 1)/=STD_LOGIC_VECTOR'("000000"));
  mux_2600_nl <= MUX_s_1_2_2(or_tmp, or_2701_nl, fsm_output(0));
  mux_2601_nl <= MUX_s_1_2_2(mux_tmp_2538, (NOT mux_2600_nl), fsm_output(7));
  and_485_nl <= (fsm_output(4)) AND (fsm_output(5)) AND (fsm_output(2));
  mux_2611_nl <= MUX_s_1_2_2((fsm_output(6)), or_165_cse, and_485_nl);
  mux_2612_nl <= MUX_s_1_2_2(mux_tmp_2538, (NOT mux_2611_nl), fsm_output(7));
  or_2824_nl <= CONV_SL_1_1(fsm_output(7 DOWNTO 5)/=STD_LOGIC_VECTOR'("000"));
  or_2825_nl <= and_515_cse OR CONV_SL_1_1(fsm_output(7 DOWNTO 5)/=STD_LOGIC_VECTOR'("000"));
  nand_161_nl <= NOT(or_2500_cse AND CONV_SL_1_1(fsm_output(7 DOWNTO 5)=STD_LOGIC_VECTOR'("111")));
  mux_2614_nl <= MUX_s_1_2_2(or_2825_nl, nand_161_nl, fsm_output(2));
  nand_162_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 5)=STD_LOGIC_VECTOR'("111")));
  mux_2615_nl <= MUX_s_1_2_2(mux_2614_nl, nand_162_nl, fsm_output(3));
  mux_2616_nl <= MUX_s_1_2_2(or_2824_nl, mux_2615_nl, fsm_output(4));
  and_482_nl <= (fsm_output(5)) AND (fsm_output(1)) AND (fsm_output(2));
  mux_2619_nl <= MUX_s_1_2_2((fsm_output(6)), or_165_cse, and_482_nl);
  mux_2620_nl <= MUX_s_1_2_2(mux_2619_nl, or_420_cse, fsm_output(4));
  or_2707_nl <= (fsm_output(7)) OR mux_2620_nl;
  mux_2621_nl <= MUX_s_1_2_2(not_tmp_664, or_2707_nl, fsm_output(8));
  and_480_nl <= (fsm_output(4)) AND (fsm_output(5)) AND (fsm_output(1)) AND (fsm_output(2));
  mux_2623_nl <= MUX_s_1_2_2((fsm_output(6)), or_165_cse, and_480_nl);
  or_2708_nl <= (fsm_output(7)) OR mux_2623_nl;
  mux_2624_nl <= MUX_s_1_2_2(not_tmp_664, or_2708_nl, fsm_output(8));
  mux_2629_nl <= MUX_s_1_2_2(mux_tmp_2574, and_475_cse, fsm_output(2));
  mux_2630_nl <= MUX_s_1_2_2(nor_510_cse, mux_2629_nl, fsm_output(4));
  mux_2627_nl <= MUX_s_1_2_2(nor_510_cse, mux_tmp_2574, fsm_output(2));
  mux_2628_nl <= MUX_s_1_2_2(mux_2627_nl, and_475_cse, fsm_output(4));
  mux_2631_nl <= MUX_s_1_2_2(mux_2630_nl, mux_2628_nl, and_515_cse);
  mux_2626_nl <= MUX_s_1_2_2(mux_tmp_2574, and_475_cse, fsm_output(4));
  mux_2632_nl <= MUX_s_1_2_2(mux_2631_nl, mux_2626_nl, fsm_output(3));
  mux_2633_nl <= MUX_s_1_2_2(mux_2632_nl, (fsm_output(8)), fsm_output(7));
  nor_511_nl <= NOT((fsm_output(2)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(8)));
  and_473_nl <= (fsm_output(2)) AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(8));
  mux_2637_nl <= MUX_s_1_2_2(nor_511_nl, and_473_nl, and_515_cse);
  mux_2638_nl <= MUX_s_1_2_2(mux_2637_nl, and_475_cse, fsm_output(3));
  mux_2639_nl <= MUX_s_1_2_2(nor_510_cse, mux_2638_nl, fsm_output(4));
  mux_2640_nl <= MUX_s_1_2_2(mux_2639_nl, (fsm_output(8)), fsm_output(7));
  and_393_nl <= (fsm_output(7)) AND or_420_cse;
  mux_2641_nl <= MUX_s_1_2_2(not_tmp_664, and_393_nl, fsm_output(8));
  and_397_nl <= (fsm_output(7)) AND or_tmp_2638;
  mux_2645_nl <= MUX_s_1_2_2(not_tmp_664, and_397_nl, fsm_output(8));
  nor_937_nl <= NOT(and_515_cse OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  and_754_nl <= or_2500_cse AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111"));
  mux_2646_nl <= MUX_s_1_2_2(nor_937_nl, and_754_nl, fsm_output(3));
  and_755_nl <= (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(7)) AND (fsm_output(8));
  mux_2647_nl <= MUX_s_1_2_2(mux_2646_nl, and_755_nl, fsm_output(2));
  mux_2648_nl <= MUX_s_1_2_2(nor_936_cse, mux_2647_nl, fsm_output(4));
  mux_2649_nl <= MUX_s_1_2_2(mux_2648_nl, and_756_cse, fsm_output(5));
  or_196_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_2655_nl <= MUX_s_1_2_2(not_tmp_696, mux_tmp_302, or_196_nl);
  mux_2656_nl <= MUX_s_1_2_2(not_tmp_696, mux_2655_nl, fsm_output(3));
  mux_2653_nl <= MUX_s_1_2_2(mux_tmp_302, nor_tmp_87, and_515_cse);
  mux_2654_nl <= MUX_s_1_2_2(mux_2653_nl, nor_tmp_87, or_598_cse);
  mux_2657_nl <= MUX_s_1_2_2(mux_2656_nl, mux_2654_nl, fsm_output(4));
  or_2651_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00")) OR mux_tmp_2377;
  or_2732_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00")) OR mux_tmp_2450;
  mux_2666_nl <= MUX_s_1_2_2(mux_tmp_2612, nor_tmp_3, fsm_output(3));
  mux_2667_nl <= MUX_s_1_2_2(not_tmp_703, mux_2666_nl, fsm_output(4));
  mux_2668_nl <= MUX_s_1_2_2(mux_2667_nl, mux_tmp_2614, and_515_cse);
  mux_2669_nl <= MUX_s_1_2_2(mux_2668_nl, mux_tmp_2614, fsm_output(2));
  mux_2670_nl <= MUX_s_1_2_2(mux_2669_nl, nor_tmp_3, fsm_output(5));
  mux_2678_nl <= MUX_s_1_2_2(mux_tmp_2626, and_tmp_11, fsm_output(3));
  mux_2679_nl <= MUX_s_1_2_2(mux_2678_nl, mux_tmp_2625, and_515_cse);
  mux_2680_nl <= MUX_s_1_2_2(mux_2679_nl, mux_tmp_2625, fsm_output(2));
  mux_2681_nl <= MUX_s_1_2_2(mux_tmp_2626, mux_2680_nl, fsm_output(4));
  or_2743_nl <= (fsm_output(8)) OR ((fsm_output(7)) AND or_tmp);
  or_2748_nl <= (fsm_output(8)) OR ((fsm_output(7)) AND mux_tmp_79);
  nor_503_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (fsm_output(9)));
  nor_504_nl <= NOT((fsm_output(3)) OR and_515_cse OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(9)));
  and_409_nl <= (fsm_output(3)) AND or_2500_cse AND (fsm_output(5)) AND (fsm_output(7))
      AND (fsm_output(9));
  mux_2690_nl <= MUX_s_1_2_2(nor_504_nl, and_409_nl, fsm_output(2));
  mux_2691_nl <= MUX_s_1_2_2(nor_503_nl, mux_2690_nl, fsm_output(4));
  mux_2692_nl <= MUX_s_1_2_2(mux_2691_nl, and_459_cse, fsm_output(6));
  nor_500_nl <= NOT((fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(9)));
  and_452_nl <= or_2500_cse AND CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"));
  mux_2706_nl <= MUX_s_1_2_2(nor_500_nl, mux_tmp_2653, and_452_nl);
  or_2755_nl <= and_515_cse OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"));
  mux_2705_nl <= MUX_s_1_2_2(mux_tmp_2653, nor_tmp_459, or_2755_nl);
  mux_2707_nl <= MUX_s_1_2_2(mux_2706_nl, mux_2705_nl, fsm_output(4));
  mux_2708_nl <= MUX_s_1_2_2(mux_2707_nl, nor_tmp_459, fsm_output(5));
  nor_498_nl <= NOT((fsm_output(2)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(7))
      OR (fsm_output(9)));
  nor_499_nl <= NOT((fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(7))
      OR (fsm_output(9)));
  mux_2710_nl <= MUX_s_1_2_2(nor_499_nl, nor_tmp_463, fsm_output(2));
  mux_2711_nl <= MUX_s_1_2_2(nor_498_nl, mux_2710_nl, fsm_output(1));
  mux_2712_nl <= MUX_s_1_2_2(mux_2711_nl, nor_tmp_463, fsm_output(3));
  mux_2713_nl <= MUX_s_1_2_2(nor_497_cse, mux_2712_nl, fsm_output(4));
  and_410_nl <= (fsm_output(8)) AND ((fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(5))
      OR or_tmp_2439);
  mux_2720_nl <= MUX_s_1_2_2(mux_tmp_2666, nor_tmp_467, or_598_cse);
  mux_2721_nl <= MUX_s_1_2_2(not_tmp_729, mux_2720_nl, fsm_output(4));
  and_636_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"));
  mux_2718_nl <= MUX_s_1_2_2(not_tmp_729, mux_tmp_2666, and_636_nl);
  mux_2719_nl <= MUX_s_1_2_2(mux_2718_nl, nor_tmp_467, fsm_output(4));
  mux_2722_nl <= MUX_s_1_2_2(mux_2721_nl, mux_2719_nl, and_515_cse);
  or_2814_nl <= (fsm_output(5)) OR (fsm_output(8)) OR (fsm_output(9));
  or_2815_nl <= (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(5)) OR (fsm_output(8))
      OR (fsm_output(9));
  nand_156_nl <= NOT((fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(5)) AND
      (fsm_output(8)) AND (fsm_output(9)));
  mux_2728_nl <= MUX_s_1_2_2(or_2815_nl, nand_156_nl, and_515_cse);
  mux_2729_nl <= MUX_s_1_2_2(or_2814_nl, mux_2728_nl, fsm_output(4));
  mux_2730_nl <= MUX_s_1_2_2(mux_2729_nl, nand_490_cse, or_111_cse);
  or_411_nl <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("00"));
  or_2777_nl <= (fsm_output(2)) OR and_515_cse OR (fsm_output(3)) OR (fsm_output(8))
      OR (fsm_output(9));
  mux_2731_nl <= MUX_s_1_2_2(or_411_nl, or_2777_nl, fsm_output(4));
  or_2812_nl <= (fsm_output(6)) OR mux_2731_nl;
  nand_154_nl <= NOT((fsm_output(6)) AND or_602_cse AND CONV_SL_1_1(fsm_output(9
      DOWNTO 8)=STD_LOGIC_VECTOR'("11")));
  mux_2732_nl <= MUX_s_1_2_2(or_2812_nl, nand_154_nl, fsm_output(5));
  mux_2733_nl <= MUX_s_1_2_2(mux_2732_nl, nand_490_cse, fsm_output(7));
  and_413_nl <= (fsm_output(8)) AND ((fsm_output(7)) OR nor_tmp_427);
  or_2891_nl <= (fsm_output(0)) OR (fsm_output(4));
  mux_2736_nl <= MUX_s_1_2_2(mux_tmp_2449, or_420_cse, or_2891_nl);
  and_414_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11")) AND mux_2736_nl;
  COMP_LOOP_nor_11_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_operator_64_false_acc_tmp(3
      DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
  COMP_LOOP_or_35_nl <= operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c1
      OR operator_64_false_slc_operator_64_false_acc_1_60_itm_mx0c3;
  COMP_LOOP_or_18_nl <= (COMP_LOOP_COMP_LOOP_nor_1_itm AND tmp_1_lpi_4_dfm_mx0c0)
      OR (COMP_LOOP_COMP_LOOP_nor_5_itm AND and_dcpl_245) OR (COMP_LOOP_COMP_LOOP_nor_9_itm
      AND and_dcpl_249) OR (COMP_LOOP_COMP_LOOP_nor_13_itm AND and_dcpl_254) OR (COMP_LOOP_COMP_LOOP_nor_17_itm
      AND and_dcpl_258) OR (COMP_LOOP_COMP_LOOP_nor_21_itm AND and_dcpl_262) OR (COMP_LOOP_COMP_LOOP_nor_25_itm
      AND and_dcpl_265) OR (COMP_LOOP_COMP_LOOP_nor_29_itm AND and_dcpl_269) OR (COMP_LOOP_COMP_LOOP_nor_33_itm
      AND and_dcpl_271) OR (COMP_LOOP_COMP_LOOP_nor_37_itm AND and_dcpl_273) OR (COMP_LOOP_COMP_LOOP_nor_41_itm
      AND and_dcpl_276) OR (COMP_LOOP_COMP_LOOP_nor_45_itm AND and_dcpl_278) OR (COMP_LOOP_COMP_LOOP_nor_49_itm
      AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_nor_53_itm AND and_dcpl_285) OR (COMP_LOOP_COMP_LOOP_nor_57_itm
      AND and_dcpl_287) OR (COMP_LOOP_COMP_LOOP_nor_61_itm AND and_dcpl_289);
  COMP_LOOP_or_19_nl <= ((operator_64_false_acc_cse_1_sva(0)) AND operator_64_false_slc_operator_64_false_acc_1_60_itm
      AND tmp_1_lpi_4_dfm_mx0c0) OR ((operator_64_false_acc_cse_2_sva(0)) AND COMP_LOOP_nor_51_itm
      AND and_dcpl_245) OR ((operator_64_false_acc_cse_3_sva(0)) AND COMP_LOOP_nor_91_itm
      AND and_dcpl_249) OR ((operator_64_false_acc_cse_4_sva(0)) AND COMP_LOOP_nor_131_itm
      AND and_dcpl_254) OR ((operator_64_false_acc_cse_5_sva(0)) AND COMP_LOOP_nor_171_itm
      AND and_dcpl_258) OR ((operator_64_false_acc_cse_6_sva(0)) AND COMP_LOOP_nor_211_itm
      AND and_dcpl_262) OR ((operator_64_false_acc_cse_7_sva(0)) AND COMP_LOOP_nor_251_itm
      AND and_dcpl_265) OR ((operator_64_false_acc_cse_8_sva(0)) AND COMP_LOOP_nor_291_itm
      AND and_dcpl_269) OR ((operator_64_false_acc_cse_9_sva(0)) AND COMP_LOOP_nor_331_itm
      AND and_dcpl_271) OR ((operator_64_false_acc_cse_10_sva(0)) AND COMP_LOOP_nor_371_itm
      AND and_dcpl_273) OR ((operator_64_false_acc_cse_11_sva(0)) AND COMP_LOOP_nor_411_itm
      AND and_dcpl_276) OR ((operator_64_false_acc_cse_12_sva(0)) AND COMP_LOOP_nor_451_itm
      AND and_dcpl_278) OR ((operator_64_false_acc_cse_13_sva(0)) AND COMP_LOOP_nor_491_itm
      AND and_dcpl_283) OR ((operator_64_false_acc_cse_14_sva(0)) AND COMP_LOOP_nor_531_itm
      AND and_dcpl_285) OR ((operator_64_false_acc_cse_15_sva(0)) AND COMP_LOOP_nor_571_itm
      AND and_dcpl_287) OR ((operator_64_false_acc_cse_sva(0)) AND COMP_LOOP_nor_611_itm
      AND and_dcpl_289);
  COMP_LOOP_or_20_nl <= ((operator_64_false_acc_cse_1_sva(1)) AND COMP_LOOP_nor_12_itm
      AND tmp_1_lpi_4_dfm_mx0c0) OR ((operator_64_false_acc_cse_2_sva(1)) AND COMP_LOOP_nor_52_itm
      AND and_dcpl_245) OR ((operator_64_false_acc_cse_3_sva(1)) AND COMP_LOOP_nor_92_itm
      AND and_dcpl_249) OR ((operator_64_false_acc_cse_4_sva(1)) AND COMP_LOOP_nor_132_itm
      AND and_dcpl_254) OR ((operator_64_false_acc_cse_5_sva(1)) AND COMP_LOOP_nor_172_itm
      AND and_dcpl_258) OR ((operator_64_false_acc_cse_6_sva(1)) AND COMP_LOOP_nor_212_itm
      AND and_dcpl_262) OR ((operator_64_false_acc_cse_7_sva(1)) AND COMP_LOOP_nor_252_itm
      AND and_dcpl_265) OR ((operator_64_false_acc_cse_8_sva(1)) AND COMP_LOOP_nor_292_itm
      AND and_dcpl_269) OR ((operator_64_false_acc_cse_9_sva(1)) AND COMP_LOOP_nor_332_itm
      AND and_dcpl_271) OR ((operator_64_false_acc_cse_10_sva(1)) AND COMP_LOOP_nor_372_itm
      AND and_dcpl_273) OR ((operator_64_false_acc_cse_11_sva(1)) AND COMP_LOOP_nor_412_itm
      AND and_dcpl_276) OR ((operator_64_false_acc_cse_12_sva(1)) AND COMP_LOOP_nor_452_itm
      AND and_dcpl_278) OR ((operator_64_false_acc_cse_13_sva(1)) AND COMP_LOOP_nor_492_itm
      AND and_dcpl_283) OR ((operator_64_false_acc_cse_14_sva(1)) AND COMP_LOOP_nor_532_itm
      AND and_dcpl_285) OR ((operator_64_false_acc_cse_15_sva(1)) AND COMP_LOOP_nor_572_itm
      AND and_dcpl_287) OR ((operator_64_false_acc_cse_sva(1)) AND COMP_LOOP_nor_612_itm
      AND and_dcpl_289);
  COMP_LOOP_or_21_nl <= (COMP_LOOP_10_operator_64_false_slc_operator_64_false_acc_63_itm
      AND tmp_1_lpi_4_dfm_mx0c0) OR (COMP_LOOP_COMP_LOOP_and_77_itm AND and_dcpl_245)
      OR (COMP_LOOP_COMP_LOOP_and_137_itm AND and_dcpl_249) OR (COMP_LOOP_COMP_LOOP_and_197_itm
      AND and_dcpl_254) OR (COMP_LOOP_COMP_LOOP_and_257_itm AND and_dcpl_258) OR
      (COMP_LOOP_COMP_LOOP_and_317_itm AND and_dcpl_262) OR (COMP_LOOP_COMP_LOOP_and_377_itm
      AND and_dcpl_265) OR (COMP_LOOP_COMP_LOOP_and_437_itm AND and_dcpl_269) OR
      (COMP_LOOP_COMP_LOOP_and_497_itm AND and_dcpl_271) OR (COMP_LOOP_COMP_LOOP_and_557_itm
      AND and_dcpl_273) OR (COMP_LOOP_COMP_LOOP_and_617_itm AND and_dcpl_276) OR
      (COMP_LOOP_COMP_LOOP_and_677_itm AND and_dcpl_278) OR (COMP_LOOP_COMP_LOOP_and_737_itm
      AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_and_797_itm AND and_dcpl_285) OR
      (COMP_LOOP_COMP_LOOP_and_857_itm AND and_dcpl_287) OR (COMP_LOOP_COMP_LOOP_and_917_itm
      AND and_dcpl_289);
  COMP_LOOP_or_22_nl <= ((operator_64_false_acc_cse_1_sva(2)) AND COMP_LOOP_nor_14_itm
      AND tmp_1_lpi_4_dfm_mx0c0) OR ((operator_64_false_acc_cse_2_sva(2)) AND COMP_LOOP_nor_54_itm
      AND and_dcpl_245) OR ((operator_64_false_acc_cse_3_sva(2)) AND COMP_LOOP_nor_94_itm
      AND and_dcpl_249) OR ((operator_64_false_acc_cse_4_sva(2)) AND COMP_LOOP_nor_134_itm
      AND and_dcpl_254) OR ((operator_64_false_acc_cse_5_sva(2)) AND COMP_LOOP_nor_174_itm
      AND and_dcpl_258) OR ((operator_64_false_acc_cse_6_sva(2)) AND COMP_LOOP_nor_214_itm
      AND and_dcpl_262) OR ((operator_64_false_acc_cse_7_sva(2)) AND COMP_LOOP_nor_254_itm
      AND and_dcpl_265) OR ((operator_64_false_acc_cse_8_sva(2)) AND COMP_LOOP_nor_294_itm
      AND and_dcpl_269) OR ((operator_64_false_acc_cse_9_sva(2)) AND COMP_LOOP_nor_334_itm
      AND and_dcpl_271) OR ((operator_64_false_acc_cse_10_sva(2)) AND COMP_LOOP_nor_374_itm
      AND and_dcpl_273) OR ((operator_64_false_acc_cse_11_sva(2)) AND COMP_LOOP_nor_414_itm
      AND and_dcpl_276) OR ((operator_64_false_acc_cse_12_sva(2)) AND COMP_LOOP_nor_454_itm
      AND and_dcpl_278) OR ((operator_64_false_acc_cse_13_sva(2)) AND COMP_LOOP_nor_494_itm
      AND and_dcpl_283) OR ((operator_64_false_acc_cse_14_sva(2)) AND COMP_LOOP_nor_534_itm
      AND and_dcpl_285) OR ((operator_64_false_acc_cse_15_sva(2)) AND COMP_LOOP_nor_574_itm
      AND and_dcpl_287) OR ((operator_64_false_acc_cse_sva(2)) AND COMP_LOOP_nor_614_itm
      AND and_dcpl_289);
  COMP_LOOP_or_23_nl <= (COMP_LOOP_COMP_LOOP_and_19_itm AND tmp_1_lpi_4_dfm_mx0c0)
      OR (COMP_LOOP_COMP_LOOP_and_79_itm AND and_dcpl_245) OR (COMP_LOOP_COMP_LOOP_and_139_itm
      AND and_dcpl_249) OR (COMP_LOOP_COMP_LOOP_and_199_itm AND and_dcpl_254) OR
      (COMP_LOOP_COMP_LOOP_and_259_itm AND and_dcpl_258) OR (COMP_LOOP_COMP_LOOP_and_319_itm
      AND and_dcpl_262) OR (COMP_LOOP_COMP_LOOP_and_379_itm AND and_dcpl_265) OR
      (COMP_LOOP_COMP_LOOP_and_439_itm AND and_dcpl_269) OR (COMP_LOOP_COMP_LOOP_and_499_itm
      AND and_dcpl_271) OR (COMP_LOOP_COMP_LOOP_and_559_itm AND and_dcpl_273) OR
      (COMP_LOOP_COMP_LOOP_and_619_itm AND and_dcpl_276) OR (COMP_LOOP_COMP_LOOP_and_679_itm
      AND and_dcpl_278) OR (COMP_LOOP_COMP_LOOP_and_739_itm AND and_dcpl_283) OR
      (COMP_LOOP_COMP_LOOP_and_799_itm AND and_dcpl_285) OR (COMP_LOOP_COMP_LOOP_and_859_itm
      AND and_dcpl_287) OR (COMP_LOOP_COMP_LOOP_and_919_itm AND and_dcpl_289);
  COMP_LOOP_or_24_nl <= (COMP_LOOP_COMP_LOOP_and_20_itm AND tmp_1_lpi_4_dfm_mx0c0)
      OR (COMP_LOOP_COMP_LOOP_and_80_itm AND and_dcpl_245) OR (COMP_LOOP_COMP_LOOP_and_140_itm
      AND and_dcpl_249) OR (COMP_LOOP_COMP_LOOP_and_200_itm AND and_dcpl_254) OR
      (COMP_LOOP_COMP_LOOP_and_260_itm AND and_dcpl_258) OR (COMP_LOOP_COMP_LOOP_and_320_itm
      AND and_dcpl_262) OR (COMP_LOOP_COMP_LOOP_and_380_itm AND and_dcpl_265) OR
      (COMP_LOOP_COMP_LOOP_and_440_itm AND and_dcpl_269) OR (COMP_LOOP_COMP_LOOP_and_500_itm
      AND and_dcpl_271) OR (COMP_LOOP_COMP_LOOP_and_560_itm AND and_dcpl_273) OR
      (COMP_LOOP_COMP_LOOP_and_620_itm AND and_dcpl_276) OR (COMP_LOOP_COMP_LOOP_and_680_itm
      AND and_dcpl_278) OR (COMP_LOOP_COMP_LOOP_and_740_itm AND and_dcpl_283) OR
      (COMP_LOOP_COMP_LOOP_and_800_itm AND and_dcpl_285) OR (COMP_LOOP_COMP_LOOP_and_860_itm
      AND and_dcpl_287) OR (COMP_LOOP_COMP_LOOP_and_920_itm AND and_dcpl_289);
  COMP_LOOP_or_25_nl <= (COMP_LOOP_COMP_LOOP_and_21_itm AND tmp_1_lpi_4_dfm_mx0c0)
      OR (COMP_LOOP_COMP_LOOP_and_81_itm AND and_dcpl_245) OR (COMP_LOOP_COMP_LOOP_and_141_itm
      AND and_dcpl_249) OR (COMP_LOOP_COMP_LOOP_and_201_itm AND and_dcpl_254) OR
      (COMP_LOOP_COMP_LOOP_and_261_itm AND and_dcpl_258) OR (COMP_LOOP_COMP_LOOP_and_321_itm
      AND and_dcpl_262) OR (COMP_LOOP_COMP_LOOP_and_381_itm AND and_dcpl_265) OR
      (COMP_LOOP_COMP_LOOP_and_441_itm AND and_dcpl_269) OR (COMP_LOOP_COMP_LOOP_and_501_itm
      AND and_dcpl_271) OR (COMP_LOOP_COMP_LOOP_and_561_itm AND and_dcpl_273) OR
      (COMP_LOOP_COMP_LOOP_and_621_itm AND and_dcpl_276) OR (COMP_LOOP_COMP_LOOP_and_681_itm
      AND and_dcpl_278) OR (COMP_LOOP_COMP_LOOP_and_741_itm AND and_dcpl_283) OR
      (COMP_LOOP_COMP_LOOP_and_801_itm AND and_dcpl_285) OR (COMP_LOOP_COMP_LOOP_and_861_itm
      AND and_dcpl_287) OR (COMP_LOOP_COMP_LOOP_and_921_itm AND and_dcpl_289);
  COMP_LOOP_or_26_nl <= ((operator_64_false_acc_cse_1_sva(3)) AND COMP_LOOP_nor_17_itm
      AND tmp_1_lpi_4_dfm_mx0c0) OR ((operator_64_false_acc_cse_2_sva(3)) AND COMP_LOOP_nor_57_itm
      AND and_dcpl_245) OR ((operator_64_false_acc_cse_3_sva(3)) AND COMP_LOOP_nor_97_itm
      AND and_dcpl_249) OR ((operator_64_false_acc_cse_4_sva(3)) AND COMP_LOOP_nor_137_itm
      AND and_dcpl_254) OR ((operator_64_false_acc_cse_5_sva(3)) AND COMP_LOOP_nor_177_itm
      AND and_dcpl_258) OR ((operator_64_false_acc_cse_6_sva(3)) AND COMP_LOOP_nor_217_itm
      AND and_dcpl_262) OR ((operator_64_false_acc_cse_7_sva(3)) AND COMP_LOOP_nor_257_itm
      AND and_dcpl_265) OR ((operator_64_false_acc_cse_8_sva(3)) AND COMP_LOOP_nor_297_itm
      AND and_dcpl_269) OR ((operator_64_false_acc_cse_9_sva(3)) AND COMP_LOOP_nor_337_itm
      AND and_dcpl_271) OR ((operator_64_false_acc_cse_10_sva(3)) AND COMP_LOOP_nor_377_itm
      AND and_dcpl_273) OR ((operator_64_false_acc_cse_11_sva(3)) AND COMP_LOOP_nor_417_itm
      AND and_dcpl_276) OR ((operator_64_false_acc_cse_12_sva(3)) AND COMP_LOOP_nor_457_itm
      AND and_dcpl_278) OR ((operator_64_false_acc_cse_13_sva(3)) AND COMP_LOOP_nor_497_itm
      AND and_dcpl_283) OR ((operator_64_false_acc_cse_14_sva(3)) AND COMP_LOOP_nor_537_itm
      AND and_dcpl_285) OR ((operator_64_false_acc_cse_15_sva(3)) AND COMP_LOOP_nor_577_itm
      AND and_dcpl_287) OR ((operator_64_false_acc_cse_sva(3)) AND COMP_LOOP_nor_617_itm
      AND and_dcpl_289);
  COMP_LOOP_or_27_nl <= (COMP_LOOP_COMP_LOOP_and_23_itm AND tmp_1_lpi_4_dfm_mx0c0)
      OR (COMP_LOOP_COMP_LOOP_and_83_itm AND and_dcpl_245) OR (COMP_LOOP_COMP_LOOP_and_143_itm
      AND and_dcpl_249) OR (COMP_LOOP_COMP_LOOP_and_203_itm AND and_dcpl_254) OR
      (COMP_LOOP_COMP_LOOP_and_263_itm AND and_dcpl_258) OR (COMP_LOOP_COMP_LOOP_and_323_itm
      AND and_dcpl_262) OR (COMP_LOOP_COMP_LOOP_and_383_itm AND and_dcpl_265) OR
      (COMP_LOOP_COMP_LOOP_and_443_itm AND and_dcpl_269) OR (COMP_LOOP_COMP_LOOP_and_503_itm
      AND and_dcpl_271) OR (COMP_LOOP_COMP_LOOP_and_563_itm AND and_dcpl_273) OR
      (COMP_LOOP_COMP_LOOP_and_623_itm AND and_dcpl_276) OR (COMP_LOOP_COMP_LOOP_and_683_itm
      AND and_dcpl_278) OR (COMP_LOOP_COMP_LOOP_and_743_itm AND and_dcpl_283) OR
      (COMP_LOOP_COMP_LOOP_and_803_itm AND and_dcpl_285) OR (COMP_LOOP_COMP_LOOP_and_863_itm
      AND and_dcpl_287) OR (COMP_LOOP_COMP_LOOP_and_923_itm AND and_dcpl_289);
  COMP_LOOP_or_28_nl <= (COMP_LOOP_COMP_LOOP_and_24_itm AND tmp_1_lpi_4_dfm_mx0c0)
      OR (COMP_LOOP_COMP_LOOP_and_84_itm AND and_dcpl_245) OR (COMP_LOOP_COMP_LOOP_and_144_itm
      AND and_dcpl_249) OR (COMP_LOOP_COMP_LOOP_and_204_itm AND and_dcpl_254) OR
      (COMP_LOOP_COMP_LOOP_and_264_itm AND and_dcpl_258) OR (COMP_LOOP_COMP_LOOP_and_324_itm
      AND and_dcpl_262) OR (COMP_LOOP_COMP_LOOP_and_384_itm AND and_dcpl_265) OR
      (COMP_LOOP_COMP_LOOP_and_444_itm AND and_dcpl_269) OR (COMP_LOOP_COMP_LOOP_and_504_itm
      AND and_dcpl_271) OR (COMP_LOOP_COMP_LOOP_and_564_itm AND and_dcpl_273) OR
      (COMP_LOOP_COMP_LOOP_and_624_itm AND and_dcpl_276) OR (COMP_LOOP_COMP_LOOP_and_684_itm
      AND and_dcpl_278) OR (COMP_LOOP_COMP_LOOP_and_744_itm AND and_dcpl_283) OR
      (COMP_LOOP_COMP_LOOP_and_804_itm AND and_dcpl_285) OR (COMP_LOOP_COMP_LOOP_and_864_itm
      AND and_dcpl_287) OR (COMP_LOOP_COMP_LOOP_and_924_itm AND and_dcpl_289);
  COMP_LOOP_or_29_nl <= (COMP_LOOP_COMP_LOOP_and_25_itm AND tmp_1_lpi_4_dfm_mx0c0)
      OR (COMP_LOOP_COMP_LOOP_and_85_itm AND and_dcpl_245) OR (COMP_LOOP_COMP_LOOP_and_145_itm
      AND and_dcpl_249) OR (COMP_LOOP_COMP_LOOP_and_205_itm AND and_dcpl_254) OR
      (COMP_LOOP_COMP_LOOP_and_265_itm AND and_dcpl_258) OR (COMP_LOOP_COMP_LOOP_and_325_itm
      AND and_dcpl_262) OR (COMP_LOOP_COMP_LOOP_and_385_itm AND and_dcpl_265) OR
      (COMP_LOOP_COMP_LOOP_and_445_itm AND and_dcpl_269) OR (COMP_LOOP_COMP_LOOP_and_505_itm
      AND and_dcpl_271) OR (COMP_LOOP_COMP_LOOP_and_565_itm AND and_dcpl_273) OR
      (COMP_LOOP_COMP_LOOP_and_625_itm AND and_dcpl_276) OR (COMP_LOOP_COMP_LOOP_and_685_itm
      AND and_dcpl_278) OR (COMP_LOOP_COMP_LOOP_and_745_itm AND and_dcpl_283) OR
      (COMP_LOOP_COMP_LOOP_and_805_itm AND and_dcpl_285) OR (COMP_LOOP_COMP_LOOP_and_865_itm
      AND and_dcpl_287) OR (COMP_LOOP_COMP_LOOP_and_925_itm AND and_dcpl_289);
  COMP_LOOP_or_30_nl <= (COMP_LOOP_COMP_LOOP_and_26_itm AND tmp_1_lpi_4_dfm_mx0c0)
      OR (COMP_LOOP_COMP_LOOP_and_86_itm AND and_dcpl_245) OR (COMP_LOOP_COMP_LOOP_and_146_itm
      AND and_dcpl_249) OR (COMP_LOOP_COMP_LOOP_and_206_itm AND and_dcpl_254) OR
      (COMP_LOOP_COMP_LOOP_and_266_itm AND and_dcpl_258) OR (COMP_LOOP_COMP_LOOP_and_326_itm
      AND and_dcpl_262) OR (COMP_LOOP_COMP_LOOP_and_386_itm AND and_dcpl_265) OR
      (COMP_LOOP_COMP_LOOP_and_446_itm AND and_dcpl_269) OR (COMP_LOOP_COMP_LOOP_and_506_itm
      AND and_dcpl_271) OR (COMP_LOOP_COMP_LOOP_and_566_itm AND and_dcpl_273) OR
      (COMP_LOOP_COMP_LOOP_and_626_itm AND and_dcpl_276) OR (COMP_LOOP_COMP_LOOP_and_686_itm
      AND and_dcpl_278) OR (COMP_LOOP_COMP_LOOP_and_746_itm AND and_dcpl_283) OR
      (COMP_LOOP_COMP_LOOP_and_806_itm AND and_dcpl_285) OR (COMP_LOOP_COMP_LOOP_and_866_itm
      AND and_dcpl_287) OR (COMP_LOOP_COMP_LOOP_and_926_itm AND and_dcpl_289);
  COMP_LOOP_or_31_nl <= (COMP_LOOP_COMP_LOOP_and_27_itm AND tmp_1_lpi_4_dfm_mx0c0)
      OR (COMP_LOOP_COMP_LOOP_and_87_itm AND and_dcpl_245) OR (COMP_LOOP_COMP_LOOP_and_147_itm
      AND and_dcpl_249) OR (COMP_LOOP_COMP_LOOP_and_207_itm AND and_dcpl_254) OR
      (COMP_LOOP_COMP_LOOP_and_267_itm AND and_dcpl_258) OR (COMP_LOOP_COMP_LOOP_and_327_itm
      AND and_dcpl_262) OR (COMP_LOOP_COMP_LOOP_and_387_itm AND and_dcpl_265) OR
      (COMP_LOOP_COMP_LOOP_and_447_itm AND and_dcpl_269) OR (COMP_LOOP_COMP_LOOP_and_507_itm
      AND and_dcpl_271) OR (COMP_LOOP_COMP_LOOP_and_567_itm AND and_dcpl_273) OR
      (COMP_LOOP_COMP_LOOP_and_627_itm AND and_dcpl_276) OR (COMP_LOOP_COMP_LOOP_and_687_itm
      AND and_dcpl_278) OR (COMP_LOOP_COMP_LOOP_and_747_itm AND and_dcpl_283) OR
      (COMP_LOOP_COMP_LOOP_and_807_itm AND and_dcpl_285) OR (COMP_LOOP_COMP_LOOP_and_867_itm
      AND and_dcpl_287) OR (COMP_LOOP_COMP_LOOP_and_927_itm AND and_dcpl_289);
  COMP_LOOP_or_32_nl <= (COMP_LOOP_COMP_LOOP_and_28_itm AND tmp_1_lpi_4_dfm_mx0c0)
      OR (COMP_LOOP_COMP_LOOP_and_88_itm AND and_dcpl_245) OR (COMP_LOOP_COMP_LOOP_and_148_itm
      AND and_dcpl_249) OR (COMP_LOOP_COMP_LOOP_and_208_itm AND and_dcpl_254) OR
      (COMP_LOOP_COMP_LOOP_and_268_itm AND and_dcpl_258) OR (COMP_LOOP_COMP_LOOP_and_328_itm
      AND and_dcpl_262) OR (COMP_LOOP_COMP_LOOP_and_388_itm AND and_dcpl_265) OR
      (COMP_LOOP_COMP_LOOP_and_448_itm AND and_dcpl_269) OR (COMP_LOOP_COMP_LOOP_and_508_itm
      AND and_dcpl_271) OR (COMP_LOOP_COMP_LOOP_and_568_itm AND and_dcpl_273) OR
      (COMP_LOOP_COMP_LOOP_and_628_itm AND and_dcpl_276) OR (COMP_LOOP_COMP_LOOP_and_688_itm
      AND and_dcpl_278) OR (COMP_LOOP_COMP_LOOP_and_748_itm AND and_dcpl_283) OR
      (COMP_LOOP_COMP_LOOP_and_808_itm AND and_dcpl_285) OR (COMP_LOOP_COMP_LOOP_and_868_itm
      AND and_dcpl_287) OR (COMP_LOOP_COMP_LOOP_and_928_itm AND and_dcpl_289);
  COMP_LOOP_or_33_nl <= (COMP_LOOP_COMP_LOOP_and_29_itm AND tmp_1_lpi_4_dfm_mx0c0)
      OR (COMP_LOOP_COMP_LOOP_and_89_itm AND and_dcpl_245) OR (COMP_LOOP_COMP_LOOP_and_149_itm
      AND and_dcpl_249) OR (COMP_LOOP_COMP_LOOP_and_209_itm AND and_dcpl_254) OR
      (COMP_LOOP_COMP_LOOP_and_269_itm AND and_dcpl_258) OR (COMP_LOOP_COMP_LOOP_and_329_itm
      AND and_dcpl_262) OR (COMP_LOOP_COMP_LOOP_and_389_itm AND and_dcpl_265) OR
      (COMP_LOOP_COMP_LOOP_and_449_itm AND and_dcpl_269) OR (COMP_LOOP_COMP_LOOP_and_509_itm
      AND and_dcpl_271) OR (COMP_LOOP_COMP_LOOP_and_569_itm AND and_dcpl_273) OR
      (COMP_LOOP_COMP_LOOP_and_629_itm AND and_dcpl_276) OR (COMP_LOOP_COMP_LOOP_and_689_itm
      AND and_dcpl_278) OR (COMP_LOOP_COMP_LOOP_and_749_itm AND and_dcpl_283) OR
      (COMP_LOOP_COMP_LOOP_and_809_itm AND and_dcpl_285) OR (COMP_LOOP_COMP_LOOP_and_869_itm
      AND and_dcpl_287) OR (COMP_LOOP_COMP_LOOP_and_929_itm AND and_dcpl_289);
  not_7089_nl <= NOT not_tmp_597;
  nand_nl <= NOT((fsm_output(7)) AND (fsm_output(1)) AND (fsm_output(0)) AND (NOT
      (fsm_output(9))) AND nor_tmp_1);
  nor_1035_nl <= NOT((NOT (fsm_output(0))) OR (fsm_output(9)) OR (NOT nor_tmp_1));
  mux_2890_nl <= MUX_s_1_2_2(nor_1035_nl, nor_tmp_1, fsm_output(1));
  mux_2896_nl <= MUX_s_1_2_2(mux_tmp_2815, mux_tmp_2823, nor_1040_cse);
  mux_2889_nl <= MUX_s_1_2_2(mux_tmp_2823, mux_2896_nl, fsm_output(1));
  mux_2891_nl <= MUX_s_1_2_2((NOT mux_2890_nl), mux_2889_nl, fsm_output(7));
  mux_2892_nl <= MUX_s_1_2_2(nand_nl, mux_2891_nl, fsm_output(4));
  mux_2895_nl <= MUX_s_1_2_2(mux_tmp_2815, mux_tmp_2823, nor_1040_cse);
  mux_2885_nl <= MUX_s_1_2_2(mux_tmp_2813, mux_tmp_2815, or_3018_cse);
  mux_2887_nl <= MUX_s_1_2_2(mux_2895_nl, mux_2885_nl, fsm_output(1));
  or_3017_nl <= (fsm_output(1)) OR (NOT((NOT (fsm_output(0))) OR (fsm_output(9))))
      OR (fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(6));
  mux_2888_nl <= MUX_s_1_2_2(mux_2887_nl, or_3017_nl, fsm_output(7));
  or_3019_nl <= (fsm_output(4)) OR mux_2888_nl;
  mux_2893_nl <= MUX_s_1_2_2(mux_2892_nl, or_3019_nl, fsm_output(5));
  mux_2879_nl <= MUX_s_1_2_2(mux_tmp_2824, (NOT mux_tmp_2812), fsm_output(9));
  mux_2878_nl <= MUX_s_1_2_2(mux_tmp_2823, mux_tmp_2824, fsm_output(9));
  mux_2880_nl <= MUX_s_1_2_2(mux_2879_nl, mux_2878_nl, fsm_output(0));
  mux_2881_nl <= MUX_s_1_2_2(mux_2880_nl, mux_tmp_2823, fsm_output(1));
  mux_2874_nl <= MUX_s_1_2_2(or_307_cse, or_165_cse, or_3018_cse);
  mux_2875_nl <= MUX_s_1_2_2(mux_2874_nl, or_307_cse, fsm_output(1));
  mux_2882_nl <= MUX_s_1_2_2(mux_2881_nl, mux_2875_nl, fsm_output(7));
  or_3011_nl <= (fsm_output(7)) OR (NOT((NOT (fsm_output(1))) OR (NOT (fsm_output(0)))
      OR (fsm_output(9)))) OR (fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(6));
  mux_2883_nl <= MUX_s_1_2_2(mux_2882_nl, or_3011_nl, fsm_output(4));
  or_3008_nl <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (NOT nor_tmp_1);
  mux_2870_nl <= MUX_s_1_2_2(and_711_cse, nor_tmp_1, nor_1040_cse);
  mux_2871_nl <= MUX_s_1_2_2(nor_tmp_1, mux_2870_nl, fsm_output(1));
  or_3006_nl <= (fsm_output(9)) OR mux_tmp_2815;
  or_3005_nl <= (fsm_output(9)) OR mux_tmp_2813;
  or_3004_nl <= (fsm_output(9)) OR mux_tmp_2812;
  mux_2867_nl <= MUX_s_1_2_2(or_3005_nl, or_3004_nl, fsm_output(0));
  mux_2869_nl <= MUX_s_1_2_2(or_3006_nl, mux_2867_nl, fsm_output(1));
  mux_2872_nl <= MUX_s_1_2_2((NOT mux_2871_nl), mux_2869_nl, fsm_output(7));
  mux_2873_nl <= MUX_s_1_2_2(or_3008_nl, mux_2872_nl, fsm_output(4));
  mux_2884_nl <= MUX_s_1_2_2(mux_2883_nl, mux_2873_nl, fsm_output(5));
  COMP_LOOP_mux_291_nl <= MUX_v_64_2_2(COMP_LOOP_10_modExp_dev_1_while_mul_mut, modExp_dev_result_sva,
      and_dcpl_402);
  or_3024_nl <= (fsm_output(1)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(5))
      OR (fsm_output(3)) OR (fsm_output(8)) OR (NOT (fsm_output(2)));
  or_3025_nl <= (NOT (fsm_output(7))) OR (fsm_output(4)) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(3))) OR (fsm_output(8)) OR (fsm_output(2));
  mux_2900_nl <= MUX_s_1_2_2(or_3025_nl, nand_tmp_150, fsm_output(1));
  mux_2899_nl <= MUX_s_1_2_2(or_3024_nl, mux_2900_nl, fsm_output(6));
  mux_2898_nl <= MUX_s_1_2_2(or_tmp_2743, mux_2899_nl, fsm_output(9));
  or_3026_nl <= (NOT (fsm_output(7))) OR (fsm_output(4)) OR mux_tmp_2749;
  mux_2902_nl <= MUX_s_1_2_2(nand_tmp_150, or_3026_nl, fsm_output(1));
  nand_491_nl <= NOT((fsm_output(6)) AND (NOT mux_2902_nl));
  mux_2901_nl <= MUX_s_1_2_2(nand_491_nl, or_tmp_2743, fsm_output(9));
  mux_2897_nl <= MUX_s_1_2_2(mux_2898_nl, mux_2901_nl, fsm_output(0));
  COMP_LOOP_mux1h_842_nl <= MUX1HOT_v_64_3_2(COMP_LOOP_1_modulo_dev_cmp_return_rsc_z,
      r_sva, modExp_dev_result_sva, STD_LOGIC_VECTOR'( (NOT mux_2897_nl) & and_dcpl_402
      & (NOT mux_2835_cse)));
  z_out <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( UNSIGNED(COMP_LOOP_mux_291_nl)
      * UNSIGNED(COMP_LOOP_mux1h_842_nl)), 64));
  COMP_LOOP_mux_292_nl <= MUX_v_10_2_2((STD_LOGIC_VECTOR'( "0000") & (STAGE_VEC_LOOP_j_sva_9_0(9
      DOWNTO 4))), STAGE_VEC_LOOP_j_sva_9_0, and_dcpl_418);
  COMP_LOOP_mux_293_nl <= MUX_v_10_2_2((STD_LOGIC_VECTOR'( "00000") & COMP_LOOP_k_9_4_sva_4_0),
      STAGE_MAIN_LOOP_lshift_psp_1_sva, and_dcpl_418);
  z_out_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_292_nl),
      11) + CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_293_nl), 11), 11));
  operator_64_false_operator_64_false_or_58_nl <= (NOT(and_dcpl_427 OR and_dcpl_435
      OR and_dcpl_442 OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464
      OR and_dcpl_468 OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_478
      OR and_dcpl_481 OR and_dcpl_484 OR and_dcpl_487 OR and_dcpl_489 OR and_dcpl_496
      OR and_dcpl_498)) OR (NOT mux_2835_cse) OR and_dcpl_493 OR and_dcpl_495;
  operator_64_false_operator_64_false_mux_58_nl <= MUX_s_1_2_2((z_out_3(63)), (STAGE_MAIN_LOOP_div_cmp_z(63)),
      and_dcpl_493);
  operator_64_false_or_130_nl <= (NOT(operator_64_false_operator_64_false_mux_58_nl
      OR and_dcpl_478 OR and_dcpl_481 OR and_dcpl_484 OR and_dcpl_487 OR and_dcpl_489))
      OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442 OR and_dcpl_449 OR and_dcpl_454
      OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468 OR and_dcpl_471 OR and_dcpl_474
      OR and_dcpl_476 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_59_nl <= MUX_s_1_2_2((z_out_3(62)), (STAGE_MAIN_LOOP_div_cmp_z(62)),
      and_dcpl_493);
  operator_64_false_or_131_nl <= (NOT(operator_64_false_operator_64_false_mux_59_nl
      OR and_dcpl_478 OR and_dcpl_481 OR and_dcpl_484 OR and_dcpl_487 OR and_dcpl_489))
      OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442 OR and_dcpl_449 OR and_dcpl_454
      OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468 OR and_dcpl_471 OR and_dcpl_474
      OR and_dcpl_476 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_60_nl <= MUX_s_1_2_2((z_out_3(61)), (STAGE_MAIN_LOOP_div_cmp_z(61)),
      and_dcpl_493);
  operator_64_false_or_132_nl <= (NOT(operator_64_false_operator_64_false_mux_60_nl
      OR and_dcpl_478 OR and_dcpl_487 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435
      OR and_dcpl_442 OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464
      OR and_dcpl_468 OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481
      OR and_dcpl_484 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_61_nl <= MUX_s_1_2_2((z_out_3(60)), (STAGE_MAIN_LOOP_div_cmp_z(60)),
      and_dcpl_493);
  operator_64_false_or_133_nl <= (NOT(operator_64_false_operator_64_false_mux_61_nl
      OR and_dcpl_478 OR and_dcpl_487 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435
      OR and_dcpl_442 OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464
      OR and_dcpl_468 OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481
      OR and_dcpl_484 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_62_nl <= MUX_s_1_2_2((z_out_3(59)), (STAGE_MAIN_LOOP_div_cmp_z(59)),
      and_dcpl_493);
  operator_64_false_or_134_nl <= (NOT(operator_64_false_operator_64_false_mux_62_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_63_nl <= MUX_s_1_2_2((z_out_3(58)), (STAGE_MAIN_LOOP_div_cmp_z(58)),
      and_dcpl_493);
  operator_64_false_or_135_nl <= (NOT(operator_64_false_operator_64_false_mux_63_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_64_nl <= MUX_s_1_2_2((z_out_3(57)), (STAGE_MAIN_LOOP_div_cmp_z(57)),
      and_dcpl_493);
  operator_64_false_or_136_nl <= (NOT(operator_64_false_operator_64_false_mux_64_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_65_nl <= MUX_s_1_2_2((z_out_3(56)), (STAGE_MAIN_LOOP_div_cmp_z(56)),
      and_dcpl_493);
  operator_64_false_or_137_nl <= (NOT(operator_64_false_operator_64_false_mux_65_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_66_nl <= MUX_s_1_2_2((z_out_3(55)), (STAGE_MAIN_LOOP_div_cmp_z(55)),
      and_dcpl_493);
  operator_64_false_or_138_nl <= (NOT(operator_64_false_operator_64_false_mux_66_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_67_nl <= MUX_s_1_2_2((z_out_3(54)), (STAGE_MAIN_LOOP_div_cmp_z(54)),
      and_dcpl_493);
  operator_64_false_or_139_nl <= (NOT(operator_64_false_operator_64_false_mux_67_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_68_nl <= MUX_s_1_2_2((z_out_3(53)), (STAGE_MAIN_LOOP_div_cmp_z(53)),
      and_dcpl_493);
  operator_64_false_or_140_nl <= (NOT(operator_64_false_operator_64_false_mux_68_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_69_nl <= MUX_s_1_2_2((z_out_3(52)), (STAGE_MAIN_LOOP_div_cmp_z(52)),
      and_dcpl_493);
  operator_64_false_or_141_nl <= (NOT(operator_64_false_operator_64_false_mux_69_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_70_nl <= MUX_s_1_2_2((z_out_3(51)), (STAGE_MAIN_LOOP_div_cmp_z(51)),
      and_dcpl_493);
  operator_64_false_or_142_nl <= (NOT(operator_64_false_operator_64_false_mux_70_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_71_nl <= MUX_s_1_2_2((z_out_3(50)), (STAGE_MAIN_LOOP_div_cmp_z(50)),
      and_dcpl_493);
  operator_64_false_or_143_nl <= (NOT(operator_64_false_operator_64_false_mux_71_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_72_nl <= MUX_s_1_2_2((z_out_3(49)), (STAGE_MAIN_LOOP_div_cmp_z(49)),
      and_dcpl_493);
  operator_64_false_or_144_nl <= (NOT(operator_64_false_operator_64_false_mux_72_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_73_nl <= MUX_s_1_2_2((z_out_3(48)), (STAGE_MAIN_LOOP_div_cmp_z(48)),
      and_dcpl_493);
  operator_64_false_or_145_nl <= (NOT(operator_64_false_operator_64_false_mux_73_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_74_nl <= MUX_s_1_2_2((z_out_3(47)), (STAGE_MAIN_LOOP_div_cmp_z(47)),
      and_dcpl_493);
  operator_64_false_or_146_nl <= (NOT(operator_64_false_operator_64_false_mux_74_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_75_nl <= MUX_s_1_2_2((z_out_3(46)), (STAGE_MAIN_LOOP_div_cmp_z(46)),
      and_dcpl_493);
  operator_64_false_or_147_nl <= (NOT(operator_64_false_operator_64_false_mux_75_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_76_nl <= MUX_s_1_2_2((z_out_3(45)), (STAGE_MAIN_LOOP_div_cmp_z(45)),
      and_dcpl_493);
  operator_64_false_or_148_nl <= (NOT(operator_64_false_operator_64_false_mux_76_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_77_nl <= MUX_s_1_2_2((z_out_3(44)), (STAGE_MAIN_LOOP_div_cmp_z(44)),
      and_dcpl_493);
  operator_64_false_or_149_nl <= (NOT(operator_64_false_operator_64_false_mux_77_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_78_nl <= MUX_s_1_2_2((z_out_3(43)), (STAGE_MAIN_LOOP_div_cmp_z(43)),
      and_dcpl_493);
  operator_64_false_or_150_nl <= (NOT(operator_64_false_operator_64_false_mux_78_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_79_nl <= MUX_s_1_2_2((z_out_3(42)), (STAGE_MAIN_LOOP_div_cmp_z(42)),
      and_dcpl_493);
  operator_64_false_or_151_nl <= (NOT(operator_64_false_operator_64_false_mux_79_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_80_nl <= MUX_s_1_2_2((z_out_3(41)), (STAGE_MAIN_LOOP_div_cmp_z(41)),
      and_dcpl_493);
  operator_64_false_or_152_nl <= (NOT(operator_64_false_operator_64_false_mux_80_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_81_nl <= MUX_s_1_2_2((z_out_3(40)), (STAGE_MAIN_LOOP_div_cmp_z(40)),
      and_dcpl_493);
  operator_64_false_or_153_nl <= (NOT(operator_64_false_operator_64_false_mux_81_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_82_nl <= MUX_s_1_2_2((z_out_3(39)), (STAGE_MAIN_LOOP_div_cmp_z(39)),
      and_dcpl_493);
  operator_64_false_or_154_nl <= (NOT(operator_64_false_operator_64_false_mux_82_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_83_nl <= MUX_s_1_2_2((z_out_3(38)), (STAGE_MAIN_LOOP_div_cmp_z(38)),
      and_dcpl_493);
  operator_64_false_or_155_nl <= (NOT(operator_64_false_operator_64_false_mux_83_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_84_nl <= MUX_s_1_2_2((z_out_3(37)), (STAGE_MAIN_LOOP_div_cmp_z(37)),
      and_dcpl_493);
  operator_64_false_or_156_nl <= (NOT(operator_64_false_operator_64_false_mux_84_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_85_nl <= MUX_s_1_2_2((z_out_3(36)), (STAGE_MAIN_LOOP_div_cmp_z(36)),
      and_dcpl_493);
  operator_64_false_or_157_nl <= (NOT(operator_64_false_operator_64_false_mux_85_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_86_nl <= MUX_s_1_2_2((z_out_3(35)), (STAGE_MAIN_LOOP_div_cmp_z(35)),
      and_dcpl_493);
  operator_64_false_or_158_nl <= (NOT(operator_64_false_operator_64_false_mux_86_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_87_nl <= MUX_s_1_2_2((z_out_3(34)), (STAGE_MAIN_LOOP_div_cmp_z(34)),
      and_dcpl_493);
  operator_64_false_or_159_nl <= (NOT(operator_64_false_operator_64_false_mux_87_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_88_nl <= MUX_s_1_2_2((z_out_3(33)), (STAGE_MAIN_LOOP_div_cmp_z(33)),
      and_dcpl_493);
  operator_64_false_or_160_nl <= (NOT(operator_64_false_operator_64_false_mux_88_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_89_nl <= MUX_s_1_2_2((z_out_3(32)), (STAGE_MAIN_LOOP_div_cmp_z(32)),
      and_dcpl_493);
  operator_64_false_or_161_nl <= (NOT(operator_64_false_operator_64_false_mux_89_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_90_nl <= MUX_s_1_2_2((z_out_3(31)), (STAGE_MAIN_LOOP_div_cmp_z(31)),
      and_dcpl_493);
  operator_64_false_or_162_nl <= (NOT(operator_64_false_operator_64_false_mux_90_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_91_nl <= MUX_s_1_2_2((z_out_3(30)), (STAGE_MAIN_LOOP_div_cmp_z(30)),
      and_dcpl_493);
  operator_64_false_or_163_nl <= (NOT(operator_64_false_operator_64_false_mux_91_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_92_nl <= MUX_s_1_2_2((z_out_3(29)), (STAGE_MAIN_LOOP_div_cmp_z(29)),
      and_dcpl_493);
  operator_64_false_or_164_nl <= (NOT(operator_64_false_operator_64_false_mux_92_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_93_nl <= MUX_s_1_2_2((z_out_3(28)), (STAGE_MAIN_LOOP_div_cmp_z(28)),
      and_dcpl_493);
  operator_64_false_or_165_nl <= (NOT(operator_64_false_operator_64_false_mux_93_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_94_nl <= MUX_s_1_2_2((z_out_3(27)), (STAGE_MAIN_LOOP_div_cmp_z(27)),
      and_dcpl_493);
  operator_64_false_or_166_nl <= (NOT(operator_64_false_operator_64_false_mux_94_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_95_nl <= MUX_s_1_2_2((z_out_3(26)), (STAGE_MAIN_LOOP_div_cmp_z(26)),
      and_dcpl_493);
  operator_64_false_or_167_nl <= (NOT(operator_64_false_operator_64_false_mux_95_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_96_nl <= MUX_s_1_2_2((z_out_3(25)), (STAGE_MAIN_LOOP_div_cmp_z(25)),
      and_dcpl_493);
  operator_64_false_or_168_nl <= (NOT(operator_64_false_operator_64_false_mux_96_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_97_nl <= MUX_s_1_2_2((z_out_3(24)), (STAGE_MAIN_LOOP_div_cmp_z(24)),
      and_dcpl_493);
  operator_64_false_or_169_nl <= (NOT(operator_64_false_operator_64_false_mux_97_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_98_nl <= MUX_s_1_2_2((z_out_3(23)), (STAGE_MAIN_LOOP_div_cmp_z(23)),
      and_dcpl_493);
  operator_64_false_or_170_nl <= (NOT(operator_64_false_operator_64_false_mux_98_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_99_nl <= MUX_s_1_2_2((z_out_3(22)), (STAGE_MAIN_LOOP_div_cmp_z(22)),
      and_dcpl_493);
  operator_64_false_or_171_nl <= (NOT(operator_64_false_operator_64_false_mux_99_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_100_nl <= MUX_s_1_2_2((z_out_3(21)), (STAGE_MAIN_LOOP_div_cmp_z(21)),
      and_dcpl_493);
  operator_64_false_or_172_nl <= (NOT(operator_64_false_operator_64_false_mux_100_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_101_nl <= MUX_s_1_2_2((z_out_3(20)), (STAGE_MAIN_LOOP_div_cmp_z(20)),
      and_dcpl_493);
  operator_64_false_or_173_nl <= (NOT(operator_64_false_operator_64_false_mux_101_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_102_nl <= MUX_s_1_2_2((z_out_3(19)), (STAGE_MAIN_LOOP_div_cmp_z(19)),
      and_dcpl_493);
  operator_64_false_or_174_nl <= (NOT(operator_64_false_operator_64_false_mux_102_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_103_nl <= MUX_s_1_2_2((z_out_3(18)), (STAGE_MAIN_LOOP_div_cmp_z(18)),
      and_dcpl_493);
  operator_64_false_or_175_nl <= (NOT(operator_64_false_operator_64_false_mux_103_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_104_nl <= MUX_s_1_2_2((z_out_3(17)), (STAGE_MAIN_LOOP_div_cmp_z(17)),
      and_dcpl_493);
  operator_64_false_or_176_nl <= (NOT(operator_64_false_operator_64_false_mux_104_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_105_nl <= MUX_s_1_2_2((z_out_3(16)), (STAGE_MAIN_LOOP_div_cmp_z(16)),
      and_dcpl_493);
  operator_64_false_or_177_nl <= (NOT(operator_64_false_operator_64_false_mux_105_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_106_nl <= MUX_s_1_2_2((z_out_3(15)), (STAGE_MAIN_LOOP_div_cmp_z(15)),
      and_dcpl_493);
  operator_64_false_or_178_nl <= (NOT(operator_64_false_operator_64_false_mux_106_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_107_nl <= MUX_s_1_2_2((z_out_3(14)), (STAGE_MAIN_LOOP_div_cmp_z(14)),
      and_dcpl_493);
  operator_64_false_or_179_nl <= (NOT(operator_64_false_operator_64_false_mux_107_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_108_nl <= MUX_s_1_2_2((z_out_3(13)), (STAGE_MAIN_LOOP_div_cmp_z(13)),
      and_dcpl_493);
  operator_64_false_or_180_nl <= (NOT(operator_64_false_operator_64_false_mux_108_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_109_nl <= MUX_s_1_2_2((z_out_3(12)), (STAGE_MAIN_LOOP_div_cmp_z(12)),
      and_dcpl_493);
  operator_64_false_or_181_nl <= (NOT(operator_64_false_operator_64_false_mux_109_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_110_nl <= MUX_s_1_2_2((z_out_3(11)), (STAGE_MAIN_LOOP_div_cmp_z(11)),
      and_dcpl_493);
  operator_64_false_or_182_nl <= (NOT(operator_64_false_operator_64_false_mux_110_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_111_nl <= MUX_s_1_2_2((z_out_3(10)), (STAGE_MAIN_LOOP_div_cmp_z(10)),
      and_dcpl_493);
  operator_64_false_or_183_nl <= (NOT(operator_64_false_operator_64_false_mux_111_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_operator_64_false_mux_112_nl <= MUX_s_1_2_2((z_out_3(9)), (STAGE_MAIN_LOOP_div_cmp_z(9)),
      and_dcpl_493);
  operator_64_false_or_184_nl <= (NOT(operator_64_false_operator_64_false_mux_112_nl
      OR and_dcpl_478 OR and_dcpl_489)) OR and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442
      OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR and_dcpl_496 OR and_dcpl_498;
  operator_64_false_mux1h_62_nl <= MUX1HOT_v_2_4_2((STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 8)), STD_LOGIC_VECTOR'( '1' & (NOT (STAGE_VEC_LOOP_j_sva_9_0(9)))),
      (z_out_3(8 DOWNTO 7)), (STAGE_MAIN_LOOP_div_cmp_z(8 DOWNTO 7)), STD_LOGIC_VECTOR'(
      operator_64_false_or_120_itm & and_dcpl_478 & operator_64_false_or_121_cse
      & and_dcpl_493));
  operator_64_false_operator_64_false_nor_111_nl <= NOT(MUX_v_2_2_2(operator_64_false_mux1h_62_nl,
      STD_LOGIC_VECTOR'("11"), and_dcpl_489));
  operator_64_false_or_186_nl <= and_dcpl_481 OR and_dcpl_484 OR and_dcpl_487;
  operator_64_false_or_185_nl <= MUX_v_2_2_2(operator_64_false_operator_64_false_nor_111_nl,
      STD_LOGIC_VECTOR'("11"), operator_64_false_or_186_nl);
  operator_64_false_or_187_nl <= and_dcpl_481 OR and_dcpl_484;
  operator_64_false_mux1h_63_nl <= MUX1HOT_v_7_7_2((NOT (STAGE_MAIN_LOOP_lshift_psp_1_sva(7
      DOWNTO 1))), (STAGE_VEC_LOOP_j_sva_9_0(8 DOWNTO 2)), (NOT (STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 3))), (STD_LOGIC_VECTOR'( "11") & (NOT (STAGE_MAIN_LOOP_lshift_psp_1_sva(9
      DOWNTO 5)))), (NOT (z_out_3(6 DOWNTO 0))), (STD_LOGIC_VECTOR'( "000") & STAGE_MAIN_LOOP_acc_1_psp_sva),
      (NOT (STAGE_MAIN_LOOP_div_cmp_z(6 DOWNTO 0))), STD_LOGIC_VECTOR'( operator_64_false_or_120_itm
      & and_dcpl_478 & operator_64_false_or_187_nl & and_dcpl_487 & operator_64_false_or_121_cse
      & and_dcpl_489 & and_dcpl_493));
  operator_64_false_or_188_nl <= (NOT(and_dcpl_478 OR (NOT mux_2835_cse) OR and_dcpl_489
      OR and_dcpl_493 OR and_dcpl_495 OR and_dcpl_496)) OR and_dcpl_427 OR and_dcpl_435
      OR and_dcpl_442 OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464
      OR and_dcpl_468 OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476 OR and_dcpl_481
      OR and_dcpl_484 OR and_dcpl_487 OR and_dcpl_498;
  operator_64_false_operator_64_false_or_59_nl <= ((COMP_LOOP_slc_acc_3_12_1_slc(5))
      AND (NOT(and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442 OR and_dcpl_449 OR and_dcpl_454
      OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468 OR and_dcpl_471 OR and_dcpl_474
      OR and_dcpl_476 OR and_dcpl_478 OR and_dcpl_481 OR and_dcpl_484 OR and_dcpl_487
      OR (NOT mux_2835_cse) OR and_dcpl_493 OR and_dcpl_495 OR and_dcpl_496))) OR
      and_dcpl_489;
  operator_64_false_operator_64_false_mux_113_nl <= MUX_v_2_2_2((COMP_LOOP_k_9_4_sva_4_0(4
      DOWNTO 3)), (COMP_LOOP_slc_acc_3_12_1_slc(4 DOWNTO 3)), and_dcpl_498);
  operator_64_false_nor_121_nl <= NOT(and_dcpl_478 OR and_dcpl_481 OR and_dcpl_484
      OR and_dcpl_487 OR (NOT mux_2835_cse) OR and_dcpl_493 OR and_dcpl_495 OR and_dcpl_496);
  operator_64_false_and_65_nl <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), operator_64_false_operator_64_false_mux_113_nl,
      operator_64_false_nor_121_nl);
  operator_64_false_or_189_nl <= MUX_v_2_2_2(operator_64_false_and_65_nl, STD_LOGIC_VECTOR'("11"),
      and_dcpl_489);
  operator_64_false_or_191_nl <= and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442 OR
      and_dcpl_449 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_476;
  operator_64_false_or_192_nl <= and_dcpl_478 OR and_dcpl_481 OR and_dcpl_484;
  operator_64_false_mux1h_64_nl <= MUX1HOT_v_3_4_2((COMP_LOOP_k_9_4_sva_4_0(2 DOWNTO
      0)), (COMP_LOOP_k_9_4_sva_4_0(4 DOWNTO 2)), (STD_LOGIC_VECTOR'( "00") & (COMP_LOOP_k_9_4_sva_4_0(4))),
      (COMP_LOOP_slc_acc_3_12_1_slc(2 DOWNTO 0)), STD_LOGIC_VECTOR'( operator_64_false_or_191_nl
      & operator_64_false_or_192_nl & and_dcpl_487 & and_dcpl_498));
  operator_64_false_nor_122_nl <= NOT((NOT mux_2835_cse) OR and_dcpl_493 OR and_dcpl_495
      OR and_dcpl_496);
  operator_64_false_and_66_nl <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), operator_64_false_mux1h_64_nl,
      operator_64_false_nor_122_nl);
  operator_64_false_or_190_nl <= MUX_v_3_2_2(operator_64_false_and_66_nl, STD_LOGIC_VECTOR'("111"),
      and_dcpl_489);
  operator_64_false_operator_64_false_mux_114_nl <= MUX_s_1_2_2((COMP_LOOP_k_9_4_sva_4_0(1)),
      (COMP_LOOP_k_9_4_sva_4_0(3)), and_dcpl_487);
  operator_64_false_or_193_nl <= (operator_64_false_operator_64_false_mux_114_nl
      AND (NOT(and_dcpl_427 OR and_dcpl_435 OR and_dcpl_442 OR and_dcpl_449 OR and_dcpl_454
      OR (NOT mux_2835_cse) OR and_dcpl_493 OR and_dcpl_495 OR and_dcpl_496 OR and_dcpl_498)))
      OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468 OR and_dcpl_471 OR and_dcpl_474
      OR and_dcpl_476 OR and_dcpl_489;
  operator_64_false_operator_64_false_mux_115_nl <= MUX_s_1_2_2((COMP_LOOP_k_9_4_sva_4_0(0)),
      (COMP_LOOP_k_9_4_sva_4_0(2)), and_dcpl_487);
  operator_64_false_or_194_nl <= (operator_64_false_operator_64_false_mux_115_nl
      AND (NOT(and_dcpl_427 OR and_dcpl_435 OR and_dcpl_458 OR and_dcpl_464 OR and_dcpl_468
      OR (NOT mux_2835_cse) OR and_dcpl_493 OR and_dcpl_495 OR and_dcpl_496 OR and_dcpl_498)))
      OR and_dcpl_442 OR and_dcpl_449 OR and_dcpl_454 OR and_dcpl_471 OR and_dcpl_474
      OR and_dcpl_476 OR and_dcpl_489;
  operator_64_false_operator_64_false_or_60_nl <= ((COMP_LOOP_k_9_4_sva_4_0(1)) AND
      (NOT(and_dcpl_427 OR and_dcpl_442 OR and_dcpl_449 OR and_dcpl_458 OR and_dcpl_464
      OR and_dcpl_471 OR and_dcpl_474 OR and_dcpl_481 OR (NOT mux_2835_cse) OR and_dcpl_493
      OR and_dcpl_495 OR and_dcpl_496 OR and_dcpl_498))) OR and_dcpl_435 OR and_dcpl_454
      OR and_dcpl_468 OR and_dcpl_476 OR and_dcpl_478 OR and_dcpl_484 OR and_dcpl_489;
  operator_64_false_operator_64_false_or_61_nl <= ((COMP_LOOP_k_9_4_sva_4_0(0)) AND
      (NOT(and_dcpl_435 OR and_dcpl_442 OR and_dcpl_454 OR and_dcpl_458 OR and_dcpl_468
      OR and_dcpl_471 OR and_dcpl_476 OR and_dcpl_481 OR and_dcpl_484 OR and_dcpl_498)))
      OR and_dcpl_427 OR and_dcpl_449 OR and_dcpl_464 OR and_dcpl_474 OR and_dcpl_478
      OR (NOT mux_2835_cse) OR and_dcpl_489 OR and_dcpl_493 OR and_dcpl_495 OR and_dcpl_496;
  acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(operator_64_false_operator_64_false_or_58_nl
      & operator_64_false_or_130_nl & operator_64_false_or_131_nl & operator_64_false_or_132_nl
      & operator_64_false_or_133_nl & operator_64_false_or_134_nl & operator_64_false_or_135_nl
      & operator_64_false_or_136_nl & operator_64_false_or_137_nl & operator_64_false_or_138_nl
      & operator_64_false_or_139_nl & operator_64_false_or_140_nl & operator_64_false_or_141_nl
      & operator_64_false_or_142_nl & operator_64_false_or_143_nl & operator_64_false_or_144_nl
      & operator_64_false_or_145_nl & operator_64_false_or_146_nl & operator_64_false_or_147_nl
      & operator_64_false_or_148_nl & operator_64_false_or_149_nl & operator_64_false_or_150_nl
      & operator_64_false_or_151_nl & operator_64_false_or_152_nl & operator_64_false_or_153_nl
      & operator_64_false_or_154_nl & operator_64_false_or_155_nl & operator_64_false_or_156_nl
      & operator_64_false_or_157_nl & operator_64_false_or_158_nl & operator_64_false_or_159_nl
      & operator_64_false_or_160_nl & operator_64_false_or_161_nl & operator_64_false_or_162_nl
      & operator_64_false_or_163_nl & operator_64_false_or_164_nl & operator_64_false_or_165_nl
      & operator_64_false_or_166_nl & operator_64_false_or_167_nl & operator_64_false_or_168_nl
      & operator_64_false_or_169_nl & operator_64_false_or_170_nl & operator_64_false_or_171_nl
      & operator_64_false_or_172_nl & operator_64_false_or_173_nl & operator_64_false_or_174_nl
      & operator_64_false_or_175_nl & operator_64_false_or_176_nl & operator_64_false_or_177_nl
      & operator_64_false_or_178_nl & operator_64_false_or_179_nl & operator_64_false_or_180_nl
      & operator_64_false_or_181_nl & operator_64_false_or_182_nl & operator_64_false_or_183_nl
      & operator_64_false_or_184_nl & operator_64_false_or_185_nl & operator_64_false_mux1h_63_nl
      & operator_64_false_or_188_nl) + CONV_UNSIGNED(CONV_SIGNED(SIGNED(operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_1_cse
      & operator_64_false_operator_64_false_or_1_cse & operator_64_false_operator_64_false_or_59_nl
      & operator_64_false_or_189_nl & operator_64_false_or_190_nl & operator_64_false_or_193_nl
      & operator_64_false_or_194_nl & operator_64_false_operator_64_false_or_60_nl
      & operator_64_false_operator_64_false_or_61_nl & '1'), 65), 66), 66));
  z_out_2 <= acc_1_nl(65 DOWNTO 1);
  operator_64_false_or_7_nl <= and_dcpl_511 OR (NOT mux_2863_itm) OR and_925_cse
      OR and_dcpl_525 OR and_936_cse OR and_940_cse OR and_945_cse OR and_950_cse
      OR and_953_cse OR and_957_cse OR and_960_cse OR and_964_cse OR and_966_cse
      OR and_970_cse OR and_973_cse OR and_975_cse OR and_978_cse;
  operator_64_false_mux1h_3_nl <= MUX1HOT_v_64_4_2(p_sva, tmp_10_lpi_4_dfm, (modExp_dev_exp_1_sva_63_9
      & modExp_dev_exp_1_sva_8_4 & (COMP_LOOP_acc_psp_sva(3 DOWNTO 0))), z_out_5,
      STD_LOGIC_VECTOR'( and_dcpl_507 & operator_64_false_or_7_nl & (NOT mux_2835_cse)
      & and_920_cse));
  operator_64_false_operator_64_false_nand_1_nl <= NOT((and_dcpl_507 OR and_dcpl_511
      OR (NOT mux_2835_cse) OR and_920_cse OR and_925_cse OR and_dcpl_525 OR and_936_cse
      OR and_940_cse OR and_945_cse OR and_950_cse OR and_953_cse OR and_957_cse
      OR and_960_cse OR and_964_cse OR and_966_cse OR and_970_cse OR and_973_cse
      OR and_975_cse OR and_978_cse) AND mux_2863_itm);
  operator_64_false_or_10_nl <= and_925_cse OR and_dcpl_525 OR and_936_cse OR and_940_cse
      OR and_945_cse OR and_950_cse OR and_953_cse OR and_957_cse OR and_960_cse
      OR and_964_cse OR and_966_cse OR and_970_cse OR and_973_cse OR and_975_cse
      OR and_978_cse;
  operator_64_false_mux1h_4_nl <= MUX1HOT_v_64_3_2(tmp_1_lpi_4_dfm, (NOT tmp_1_lpi_4_dfm),
      z_out_5, STD_LOGIC_VECTOR'( and_920_cse & (NOT mux_2863_itm) & operator_64_false_or_10_nl));
  operator_64_false_or_11_nl <= and_dcpl_507 OR and_dcpl_511 OR (NOT mux_2835_cse);
  operator_64_false_or_9_nl <= MUX_v_64_2_2(operator_64_false_mux1h_4_nl, STD_LOGIC_VECTOR'("1111111111111111111111111111111111111111111111111111111111111111"),
      operator_64_false_or_11_nl);
  acc_2_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(operator_64_false_mux1h_3_nl
      & operator_64_false_operator_64_false_nand_1_nl) + UNSIGNED(operator_64_false_or_9_nl
      & '1'), 65));
  z_out_3 <= acc_2_nl(64 DOWNTO 1);
  COMP_LOOP_COMP_LOOP_or_3_nl <= (NOT(and_dcpl_582 OR and_dcpl_599)) OR and_dcpl_589
      OR and_dcpl_593;
  not_7303_nl <= NOT and_dcpl_599;
  COMP_LOOP_and_451_nl <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), (STAGE_VEC_LOOP_j_sva_9_0(9
      DOWNTO 6)), not_7303_nl);
  COMP_LOOP_or_41_nl <= and_dcpl_589 OR and_dcpl_593;
  COMP_LOOP_COMP_LOOP_or_4_nl <= MUX_v_4_2_2(COMP_LOOP_and_451_nl, STD_LOGIC_VECTOR'("1111"),
      COMP_LOOP_or_41_nl);
  COMP_LOOP_mux1h_843_nl <= MUX1HOT_v_6_3_2((STAGE_VEC_LOOP_j_sva_9_0(5 DOWNTO 0)),
      (NOT (STAGE_MAIN_LOOP_lshift_psp_1_sva(9 DOWNTO 4))), ('0' & COMP_LOOP_k_9_4_sva_4_0),
      STD_LOGIC_VECTOR'( and_dcpl_582 & and_dcpl_589 & and_dcpl_599));
  COMP_LOOP_or_42_nl <= MUX_v_6_2_2(COMP_LOOP_mux1h_843_nl, STD_LOGIC_VECTOR'("111111"),
      and_dcpl_593);
  COMP_LOOP_or_43_nl <= (NOT(and_dcpl_582 OR and_dcpl_593 OR and_dcpl_599)) OR and_dcpl_589;
  COMP_LOOP_nor_626_nl <= NOT(and_dcpl_589 OR and_dcpl_593 OR and_dcpl_599);
  COMP_LOOP_COMP_LOOP_and_992_nl <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), (COMP_LOOP_k_9_4_sva_4_0(4
      DOWNTO 2)), COMP_LOOP_nor_626_nl);
  COMP_LOOP_mux_294_nl <= MUX_v_2_2_2((COMP_LOOP_k_9_4_sva_4_0(1 DOWNTO 0)), (COMP_LOOP_k_9_4_sva_4_0(4
      DOWNTO 3)), and_dcpl_589);
  COMP_LOOP_nor_627_nl <= NOT(and_dcpl_593 OR and_dcpl_599);
  COMP_LOOP_COMP_LOOP_and_993_nl <= MUX_v_2_2_2(STD_LOGIC_VECTOR'("00"), COMP_LOOP_mux_294_nl,
      COMP_LOOP_nor_627_nl);
  COMP_LOOP_mux1h_844_nl <= MUX1HOT_v_3_3_2(STD_LOGIC_VECTOR'( "010"), (COMP_LOOP_k_9_4_sva_4_0(2
      DOWNTO 0)), (STAGE_MAIN_LOOP_acc_1_psp_sva(3 DOWNTO 1)), STD_LOGIC_VECTOR'(
      and_dcpl_582 & and_dcpl_589 & and_dcpl_593));
  not_7304_nl <= NOT and_dcpl_599;
  COMP_LOOP_and_452_nl <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), COMP_LOOP_mux1h_844_nl,
      not_7304_nl);
  COMP_LOOP_COMP_LOOP_or_5_nl <= ((STAGE_MAIN_LOOP_acc_1_psp_sva(0)) AND (NOT and_dcpl_589))
      OR and_dcpl_582 OR and_dcpl_599;
  acc_3_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_SIGNED(SIGNED(COMP_LOOP_COMP_LOOP_or_3_nl
      & COMP_LOOP_COMP_LOOP_or_4_nl & COMP_LOOP_or_42_nl & COMP_LOOP_or_43_nl), 12),
      13) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_and_992_nl & COMP_LOOP_COMP_LOOP_and_993_nl
      & COMP_LOOP_and_452_nl & COMP_LOOP_COMP_LOOP_or_5_nl & '1'), 10), 13), 13));
  COMP_LOOP_slc_acc_3_12_1_slc <= acc_3_nl(12 DOWNTO 1);
  COMP_LOOP_mux1h_845_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_nor_itm, COMP_LOOP_COMP_LOOP_nor_5_itm,
      COMP_LOOP_COMP_LOOP_nor_9_itm, COMP_LOOP_COMP_LOOP_nor_13_itm, COMP_LOOP_COMP_LOOP_nor_17_itm,
      COMP_LOOP_COMP_LOOP_nor_21_itm, COMP_LOOP_COMP_LOOP_nor_25_itm, COMP_LOOP_COMP_LOOP_nor_29_itm,
      COMP_LOOP_COMP_LOOP_nor_33_itm, COMP_LOOP_COMP_LOOP_nor_37_itm, COMP_LOOP_COMP_LOOP_nor_41_itm,
      COMP_LOOP_COMP_LOOP_nor_45_itm, COMP_LOOP_COMP_LOOP_nor_49_itm, COMP_LOOP_COMP_LOOP_nor_53_itm,
      COMP_LOOP_COMP_LOOP_nor_57_itm, COMP_LOOP_COMP_LOOP_nor_61_itm, STD_LOGIC_VECTOR'(
      and_920_cse & and_925_cse & and_dcpl_621 & and_936_cse & and_940_cse & and_945_cse
      & and_950_cse & and_953_cse & and_957_cse & and_960_cse & and_964_cse & and_966_cse
      & and_970_cse & and_973_cse & and_975_cse & and_978_cse));
  COMP_LOOP_COMP_LOOP_and_994_nl <= (operator_64_false_acc_cse_2_sva(0)) AND COMP_LOOP_nor_51_itm;
  COMP_LOOP_COMP_LOOP_and_995_nl <= (operator_64_false_acc_cse_3_sva(0)) AND COMP_LOOP_nor_91_itm;
  COMP_LOOP_COMP_LOOP_and_996_nl <= (operator_64_false_acc_cse_4_sva(0)) AND COMP_LOOP_nor_131_itm;
  COMP_LOOP_COMP_LOOP_and_997_nl <= (operator_64_false_acc_cse_5_sva(0)) AND COMP_LOOP_nor_171_itm;
  COMP_LOOP_COMP_LOOP_and_998_nl <= (operator_64_false_acc_cse_6_sva(0)) AND COMP_LOOP_nor_211_itm;
  COMP_LOOP_COMP_LOOP_and_999_nl <= (operator_64_false_acc_cse_7_sva(0)) AND COMP_LOOP_nor_251_itm;
  COMP_LOOP_COMP_LOOP_and_1000_nl <= (operator_64_false_acc_cse_8_sva(0)) AND COMP_LOOP_nor_291_itm;
  COMP_LOOP_COMP_LOOP_and_1001_nl <= (operator_64_false_acc_cse_9_sva(0)) AND COMP_LOOP_nor_331_itm;
  COMP_LOOP_COMP_LOOP_and_1002_nl <= (operator_64_false_acc_cse_10_sva(0)) AND COMP_LOOP_nor_371_itm;
  COMP_LOOP_COMP_LOOP_and_1003_nl <= (operator_64_false_acc_cse_11_sva(0)) AND COMP_LOOP_nor_411_itm;
  COMP_LOOP_COMP_LOOP_and_1004_nl <= (operator_64_false_acc_cse_12_sva(0)) AND COMP_LOOP_nor_451_itm;
  COMP_LOOP_COMP_LOOP_and_1005_nl <= (operator_64_false_acc_cse_13_sva(0)) AND COMP_LOOP_nor_491_itm;
  COMP_LOOP_COMP_LOOP_and_1006_nl <= (operator_64_false_acc_cse_14_sva(0)) AND COMP_LOOP_nor_531_itm;
  COMP_LOOP_COMP_LOOP_and_1007_nl <= (operator_64_false_acc_cse_15_sva(0)) AND COMP_LOOP_nor_571_itm;
  COMP_LOOP_COMP_LOOP_and_1008_nl <= (operator_64_false_acc_cse_sva(0)) AND COMP_LOOP_nor_611_itm;
  COMP_LOOP_mux1h_846_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_244_itm, COMP_LOOP_COMP_LOOP_and_994_nl,
      COMP_LOOP_COMP_LOOP_and_995_nl, COMP_LOOP_COMP_LOOP_and_996_nl, COMP_LOOP_COMP_LOOP_and_997_nl,
      COMP_LOOP_COMP_LOOP_and_998_nl, COMP_LOOP_COMP_LOOP_and_999_nl, COMP_LOOP_COMP_LOOP_and_1000_nl,
      COMP_LOOP_COMP_LOOP_and_1001_nl, COMP_LOOP_COMP_LOOP_and_1002_nl, COMP_LOOP_COMP_LOOP_and_1003_nl,
      COMP_LOOP_COMP_LOOP_and_1004_nl, COMP_LOOP_COMP_LOOP_and_1005_nl, COMP_LOOP_COMP_LOOP_and_1006_nl,
      COMP_LOOP_COMP_LOOP_and_1007_nl, COMP_LOOP_COMP_LOOP_and_1008_nl, STD_LOGIC_VECTOR'(
      and_920_cse & and_925_cse & and_dcpl_621 & and_936_cse & and_940_cse & and_945_cse
      & and_950_cse & and_953_cse & and_957_cse & and_960_cse & and_964_cse & and_966_cse
      & and_970_cse & and_973_cse & and_975_cse & and_978_cse));
  COMP_LOOP_COMP_LOOP_and_1009_nl <= (operator_64_false_acc_cse_2_sva(1)) AND COMP_LOOP_nor_52_itm;
  COMP_LOOP_COMP_LOOP_and_1010_nl <= (operator_64_false_acc_cse_3_sva(1)) AND COMP_LOOP_nor_92_itm;
  COMP_LOOP_COMP_LOOP_and_1011_nl <= (operator_64_false_acc_cse_4_sva(1)) AND COMP_LOOP_nor_132_itm;
  COMP_LOOP_COMP_LOOP_and_1012_nl <= (operator_64_false_acc_cse_5_sva(1)) AND COMP_LOOP_nor_172_itm;
  COMP_LOOP_COMP_LOOP_and_1013_nl <= (operator_64_false_acc_cse_6_sva(1)) AND COMP_LOOP_nor_212_itm;
  COMP_LOOP_COMP_LOOP_and_1014_nl <= (operator_64_false_acc_cse_7_sva(1)) AND COMP_LOOP_nor_252_itm;
  COMP_LOOP_COMP_LOOP_and_1015_nl <= (operator_64_false_acc_cse_8_sva(1)) AND COMP_LOOP_nor_292_itm;
  COMP_LOOP_COMP_LOOP_and_1016_nl <= (operator_64_false_acc_cse_9_sva(1)) AND COMP_LOOP_nor_332_itm;
  COMP_LOOP_COMP_LOOP_and_1017_nl <= (operator_64_false_acc_cse_10_sva(1)) AND COMP_LOOP_nor_372_itm;
  COMP_LOOP_COMP_LOOP_and_1018_nl <= (operator_64_false_acc_cse_11_sva(1)) AND COMP_LOOP_nor_412_itm;
  COMP_LOOP_COMP_LOOP_and_1019_nl <= (operator_64_false_acc_cse_12_sva(1)) AND COMP_LOOP_nor_452_itm;
  COMP_LOOP_COMP_LOOP_and_1020_nl <= (operator_64_false_acc_cse_13_sva(1)) AND COMP_LOOP_nor_492_itm;
  COMP_LOOP_COMP_LOOP_and_1021_nl <= (operator_64_false_acc_cse_14_sva(1)) AND COMP_LOOP_nor_532_itm;
  COMP_LOOP_COMP_LOOP_and_1022_nl <= (operator_64_false_acc_cse_15_sva(1)) AND COMP_LOOP_nor_572_itm;
  COMP_LOOP_COMP_LOOP_and_1023_nl <= (operator_64_false_acc_cse_sva(1)) AND COMP_LOOP_nor_612_itm;
  COMP_LOOP_mux1h_847_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_62_itm, COMP_LOOP_COMP_LOOP_and_1009_nl,
      COMP_LOOP_COMP_LOOP_and_1010_nl, COMP_LOOP_COMP_LOOP_and_1011_nl, COMP_LOOP_COMP_LOOP_and_1012_nl,
      COMP_LOOP_COMP_LOOP_and_1013_nl, COMP_LOOP_COMP_LOOP_and_1014_nl, COMP_LOOP_COMP_LOOP_and_1015_nl,
      COMP_LOOP_COMP_LOOP_and_1016_nl, COMP_LOOP_COMP_LOOP_and_1017_nl, COMP_LOOP_COMP_LOOP_and_1018_nl,
      COMP_LOOP_COMP_LOOP_and_1019_nl, COMP_LOOP_COMP_LOOP_and_1020_nl, COMP_LOOP_COMP_LOOP_and_1021_nl,
      COMP_LOOP_COMP_LOOP_and_1022_nl, COMP_LOOP_COMP_LOOP_and_1023_nl, STD_LOGIC_VECTOR'(
      and_920_cse & and_925_cse & and_dcpl_621 & and_936_cse & and_940_cse & and_945_cse
      & and_950_cse & and_953_cse & and_957_cse & and_960_cse & and_964_cse & and_966_cse
      & and_970_cse & and_973_cse & and_975_cse & and_978_cse));
  COMP_LOOP_mux1h_848_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_185_itm, COMP_LOOP_COMP_LOOP_and_77_itm,
      COMP_LOOP_COMP_LOOP_and_137_itm, COMP_LOOP_COMP_LOOP_and_197_itm, COMP_LOOP_COMP_LOOP_and_257_itm,
      COMP_LOOP_COMP_LOOP_and_317_itm, COMP_LOOP_COMP_LOOP_and_377_itm, COMP_LOOP_COMP_LOOP_and_437_itm,
      COMP_LOOP_COMP_LOOP_and_497_itm, COMP_LOOP_COMP_LOOP_and_557_itm, COMP_LOOP_COMP_LOOP_and_617_itm,
      COMP_LOOP_COMP_LOOP_and_677_itm, COMP_LOOP_COMP_LOOP_and_737_itm, COMP_LOOP_COMP_LOOP_and_797_itm,
      COMP_LOOP_COMP_LOOP_and_857_itm, COMP_LOOP_COMP_LOOP_and_917_itm, STD_LOGIC_VECTOR'(
      and_920_cse & and_925_cse & and_dcpl_621 & and_936_cse & and_940_cse & and_945_cse
      & and_950_cse & and_953_cse & and_957_cse & and_960_cse & and_964_cse & and_966_cse
      & and_970_cse & and_973_cse & and_975_cse & and_978_cse));
  COMP_LOOP_COMP_LOOP_and_1024_nl <= (operator_64_false_acc_cse_2_sva(2)) AND COMP_LOOP_nor_54_itm;
  COMP_LOOP_COMP_LOOP_and_1025_nl <= (operator_64_false_acc_cse_3_sva(2)) AND COMP_LOOP_nor_94_itm;
  COMP_LOOP_COMP_LOOP_and_1026_nl <= (operator_64_false_acc_cse_4_sva(2)) AND COMP_LOOP_nor_134_itm;
  COMP_LOOP_COMP_LOOP_and_1027_nl <= (operator_64_false_acc_cse_5_sva(2)) AND COMP_LOOP_nor_174_itm;
  COMP_LOOP_COMP_LOOP_and_1028_nl <= (operator_64_false_acc_cse_6_sva(2)) AND COMP_LOOP_nor_214_itm;
  COMP_LOOP_COMP_LOOP_and_1029_nl <= (operator_64_false_acc_cse_7_sva(2)) AND COMP_LOOP_nor_254_itm;
  COMP_LOOP_COMP_LOOP_and_1030_nl <= (operator_64_false_acc_cse_8_sva(2)) AND COMP_LOOP_nor_294_itm;
  COMP_LOOP_COMP_LOOP_and_1031_nl <= (operator_64_false_acc_cse_9_sva(2)) AND COMP_LOOP_nor_334_itm;
  COMP_LOOP_COMP_LOOP_and_1032_nl <= (operator_64_false_acc_cse_10_sva(2)) AND COMP_LOOP_nor_374_itm;
  COMP_LOOP_COMP_LOOP_and_1033_nl <= (operator_64_false_acc_cse_11_sva(2)) AND COMP_LOOP_nor_414_itm;
  COMP_LOOP_COMP_LOOP_and_1034_nl <= (operator_64_false_acc_cse_12_sva(2)) AND COMP_LOOP_nor_454_itm;
  COMP_LOOP_COMP_LOOP_and_1035_nl <= (operator_64_false_acc_cse_13_sva(2)) AND COMP_LOOP_nor_494_itm;
  COMP_LOOP_COMP_LOOP_and_1036_nl <= (operator_64_false_acc_cse_14_sva(2)) AND COMP_LOOP_nor_534_itm;
  COMP_LOOP_COMP_LOOP_and_1037_nl <= (operator_64_false_acc_cse_15_sva(2)) AND COMP_LOOP_nor_574_itm;
  COMP_LOOP_COMP_LOOP_and_1038_nl <= (operator_64_false_acc_cse_sva(2)) AND COMP_LOOP_nor_614_itm;
  COMP_LOOP_mux1h_849_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_64_itm, COMP_LOOP_COMP_LOOP_and_1024_nl,
      COMP_LOOP_COMP_LOOP_and_1025_nl, COMP_LOOP_COMP_LOOP_and_1026_nl, COMP_LOOP_COMP_LOOP_and_1027_nl,
      COMP_LOOP_COMP_LOOP_and_1028_nl, COMP_LOOP_COMP_LOOP_and_1029_nl, COMP_LOOP_COMP_LOOP_and_1030_nl,
      COMP_LOOP_COMP_LOOP_and_1031_nl, COMP_LOOP_COMP_LOOP_and_1032_nl, COMP_LOOP_COMP_LOOP_and_1033_nl,
      COMP_LOOP_COMP_LOOP_and_1034_nl, COMP_LOOP_COMP_LOOP_and_1035_nl, COMP_LOOP_COMP_LOOP_and_1036_nl,
      COMP_LOOP_COMP_LOOP_and_1037_nl, COMP_LOOP_COMP_LOOP_and_1038_nl, STD_LOGIC_VECTOR'(
      and_920_cse & and_925_cse & and_dcpl_621 & and_936_cse & and_940_cse & and_945_cse
      & and_950_cse & and_953_cse & and_957_cse & and_960_cse & and_964_cse & and_966_cse
      & and_970_cse & and_973_cse & and_975_cse & and_978_cse));
  COMP_LOOP_mux1h_850_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_65_itm, COMP_LOOP_COMP_LOOP_and_79_itm,
      COMP_LOOP_COMP_LOOP_and_139_itm, COMP_LOOP_COMP_LOOP_and_199_itm, COMP_LOOP_COMP_LOOP_and_259_itm,
      COMP_LOOP_COMP_LOOP_and_319_itm, COMP_LOOP_COMP_LOOP_and_379_itm, COMP_LOOP_COMP_LOOP_and_439_itm,
      COMP_LOOP_COMP_LOOP_and_499_itm, COMP_LOOP_COMP_LOOP_and_559_itm, COMP_LOOP_COMP_LOOP_and_619_itm,
      COMP_LOOP_COMP_LOOP_and_679_itm, COMP_LOOP_COMP_LOOP_and_739_itm, COMP_LOOP_COMP_LOOP_and_799_itm,
      COMP_LOOP_COMP_LOOP_and_859_itm, COMP_LOOP_COMP_LOOP_and_919_itm, STD_LOGIC_VECTOR'(
      and_920_cse & and_925_cse & and_dcpl_621 & and_936_cse & and_940_cse & and_945_cse
      & and_950_cse & and_953_cse & and_957_cse & and_960_cse & and_964_cse & and_966_cse
      & and_970_cse & and_973_cse & and_975_cse & and_978_cse));
  COMP_LOOP_mux1h_851_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_66_itm, COMP_LOOP_COMP_LOOP_and_80_itm,
      COMP_LOOP_COMP_LOOP_and_140_itm, COMP_LOOP_COMP_LOOP_and_200_itm, COMP_LOOP_COMP_LOOP_and_260_itm,
      COMP_LOOP_COMP_LOOP_and_320_itm, COMP_LOOP_COMP_LOOP_and_380_itm, COMP_LOOP_COMP_LOOP_and_440_itm,
      COMP_LOOP_COMP_LOOP_and_500_itm, COMP_LOOP_COMP_LOOP_and_560_itm, COMP_LOOP_COMP_LOOP_and_620_itm,
      COMP_LOOP_COMP_LOOP_and_680_itm, COMP_LOOP_COMP_LOOP_and_740_itm, COMP_LOOP_COMP_LOOP_and_800_itm,
      COMP_LOOP_COMP_LOOP_and_860_itm, COMP_LOOP_COMP_LOOP_and_920_itm, STD_LOGIC_VECTOR'(
      and_920_cse & and_925_cse & and_dcpl_621 & and_936_cse & and_940_cse & and_945_cse
      & and_950_cse & and_953_cse & and_957_cse & and_960_cse & and_964_cse & and_966_cse
      & and_970_cse & and_973_cse & and_975_cse & and_978_cse));
  COMP_LOOP_mux1h_852_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_6_itm, COMP_LOOP_COMP_LOOP_and_81_itm,
      COMP_LOOP_COMP_LOOP_and_141_itm, COMP_LOOP_COMP_LOOP_and_201_itm, COMP_LOOP_COMP_LOOP_and_261_itm,
      COMP_LOOP_COMP_LOOP_and_321_itm, COMP_LOOP_COMP_LOOP_and_381_itm, COMP_LOOP_COMP_LOOP_and_441_itm,
      COMP_LOOP_COMP_LOOP_and_501_itm, COMP_LOOP_COMP_LOOP_and_561_itm, COMP_LOOP_COMP_LOOP_and_621_itm,
      COMP_LOOP_COMP_LOOP_and_681_itm, COMP_LOOP_COMP_LOOP_and_741_itm, COMP_LOOP_COMP_LOOP_and_801_itm,
      COMP_LOOP_COMP_LOOP_and_861_itm, COMP_LOOP_COMP_LOOP_and_921_itm, STD_LOGIC_VECTOR'(
      and_920_cse & and_925_cse & and_dcpl_621 & and_936_cse & and_940_cse & and_945_cse
      & and_950_cse & and_953_cse & and_957_cse & and_960_cse & and_964_cse & and_966_cse
      & and_970_cse & and_973_cse & and_975_cse & and_978_cse));
  COMP_LOOP_COMP_LOOP_and_1039_nl <= (operator_64_false_acc_cse_2_sva(3)) AND COMP_LOOP_nor_57_itm;
  COMP_LOOP_COMP_LOOP_and_1040_nl <= (operator_64_false_acc_cse_3_sva(3)) AND COMP_LOOP_nor_97_itm;
  COMP_LOOP_COMP_LOOP_and_1041_nl <= (operator_64_false_acc_cse_4_sva(3)) AND COMP_LOOP_nor_137_itm;
  COMP_LOOP_COMP_LOOP_and_1042_nl <= (operator_64_false_acc_cse_5_sva(3)) AND COMP_LOOP_nor_177_itm;
  COMP_LOOP_COMP_LOOP_and_1043_nl <= (operator_64_false_acc_cse_6_sva(3)) AND COMP_LOOP_nor_217_itm;
  COMP_LOOP_COMP_LOOP_and_1044_nl <= (operator_64_false_acc_cse_7_sva(3)) AND COMP_LOOP_nor_257_itm;
  COMP_LOOP_COMP_LOOP_and_1045_nl <= (operator_64_false_acc_cse_8_sva(3)) AND COMP_LOOP_nor_297_itm;
  COMP_LOOP_COMP_LOOP_and_1046_nl <= (operator_64_false_acc_cse_9_sva(3)) AND COMP_LOOP_nor_337_itm;
  COMP_LOOP_COMP_LOOP_and_1047_nl <= (operator_64_false_acc_cse_10_sva(3)) AND COMP_LOOP_nor_377_itm;
  COMP_LOOP_COMP_LOOP_and_1048_nl <= (operator_64_false_acc_cse_11_sva(3)) AND COMP_LOOP_nor_417_itm;
  COMP_LOOP_COMP_LOOP_and_1049_nl <= (operator_64_false_acc_cse_12_sva(3)) AND COMP_LOOP_nor_457_itm;
  COMP_LOOP_COMP_LOOP_and_1050_nl <= (operator_64_false_acc_cse_13_sva(3)) AND COMP_LOOP_nor_497_itm;
  COMP_LOOP_COMP_LOOP_and_1051_nl <= (operator_64_false_acc_cse_14_sva(3)) AND COMP_LOOP_nor_537_itm;
  COMP_LOOP_COMP_LOOP_and_1052_nl <= (operator_64_false_acc_cse_15_sva(3)) AND COMP_LOOP_nor_577_itm;
  COMP_LOOP_COMP_LOOP_and_1053_nl <= (operator_64_false_acc_cse_sva(3)) AND COMP_LOOP_nor_617_itm;
  COMP_LOOP_mux1h_853_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_68_itm, COMP_LOOP_COMP_LOOP_and_1039_nl,
      COMP_LOOP_COMP_LOOP_and_1040_nl, COMP_LOOP_COMP_LOOP_and_1041_nl, COMP_LOOP_COMP_LOOP_and_1042_nl,
      COMP_LOOP_COMP_LOOP_and_1043_nl, COMP_LOOP_COMP_LOOP_and_1044_nl, COMP_LOOP_COMP_LOOP_and_1045_nl,
      COMP_LOOP_COMP_LOOP_and_1046_nl, COMP_LOOP_COMP_LOOP_and_1047_nl, COMP_LOOP_COMP_LOOP_and_1048_nl,
      COMP_LOOP_COMP_LOOP_and_1049_nl, COMP_LOOP_COMP_LOOP_and_1050_nl, COMP_LOOP_COMP_LOOP_and_1051_nl,
      COMP_LOOP_COMP_LOOP_and_1052_nl, COMP_LOOP_COMP_LOOP_and_1053_nl, STD_LOGIC_VECTOR'(
      and_920_cse & and_925_cse & and_dcpl_621 & and_936_cse & and_940_cse & and_945_cse
      & and_950_cse & and_953_cse & and_957_cse & and_960_cse & and_964_cse & and_966_cse
      & and_970_cse & and_973_cse & and_975_cse & and_978_cse));
  COMP_LOOP_mux1h_854_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_69_itm, COMP_LOOP_COMP_LOOP_and_83_itm,
      COMP_LOOP_COMP_LOOP_and_143_itm, COMP_LOOP_COMP_LOOP_and_203_itm, COMP_LOOP_COMP_LOOP_and_263_itm,
      COMP_LOOP_COMP_LOOP_and_323_itm, COMP_LOOP_COMP_LOOP_and_383_itm, COMP_LOOP_COMP_LOOP_and_443_itm,
      COMP_LOOP_COMP_LOOP_and_503_itm, COMP_LOOP_COMP_LOOP_and_563_itm, COMP_LOOP_COMP_LOOP_and_623_itm,
      COMP_LOOP_COMP_LOOP_and_683_itm, COMP_LOOP_COMP_LOOP_and_743_itm, COMP_LOOP_COMP_LOOP_and_803_itm,
      COMP_LOOP_COMP_LOOP_and_863_itm, COMP_LOOP_COMP_LOOP_and_923_itm, STD_LOGIC_VECTOR'(
      and_920_cse & and_925_cse & and_dcpl_621 & and_936_cse & and_940_cse & and_945_cse
      & and_950_cse & and_953_cse & and_957_cse & and_960_cse & and_964_cse & and_966_cse
      & and_970_cse & and_973_cse & and_975_cse & and_978_cse));
  COMP_LOOP_mux1h_855_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_70_itm, COMP_LOOP_COMP_LOOP_and_84_itm,
      COMP_LOOP_COMP_LOOP_and_144_itm, COMP_LOOP_COMP_LOOP_and_204_itm, COMP_LOOP_COMP_LOOP_and_264_itm,
      COMP_LOOP_COMP_LOOP_and_324_itm, COMP_LOOP_COMP_LOOP_and_384_itm, COMP_LOOP_COMP_LOOP_and_444_itm,
      COMP_LOOP_COMP_LOOP_and_504_itm, COMP_LOOP_COMP_LOOP_and_564_itm, COMP_LOOP_COMP_LOOP_and_624_itm,
      COMP_LOOP_COMP_LOOP_and_684_itm, COMP_LOOP_COMP_LOOP_and_744_itm, COMP_LOOP_COMP_LOOP_and_804_itm,
      COMP_LOOP_COMP_LOOP_and_864_itm, COMP_LOOP_COMP_LOOP_and_924_itm, STD_LOGIC_VECTOR'(
      and_920_cse & and_925_cse & and_dcpl_621 & and_936_cse & and_940_cse & and_945_cse
      & and_950_cse & and_953_cse & and_957_cse & and_960_cse & and_964_cse & and_966_cse
      & and_970_cse & and_973_cse & and_975_cse & and_978_cse));
  COMP_LOOP_mux1h_856_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_10_itm, COMP_LOOP_COMP_LOOP_and_85_itm,
      COMP_LOOP_COMP_LOOP_and_145_itm, COMP_LOOP_COMP_LOOP_and_205_itm, COMP_LOOP_COMP_LOOP_and_265_itm,
      COMP_LOOP_COMP_LOOP_and_325_itm, COMP_LOOP_COMP_LOOP_and_385_itm, COMP_LOOP_COMP_LOOP_and_445_itm,
      COMP_LOOP_COMP_LOOP_and_505_itm, COMP_LOOP_COMP_LOOP_and_565_itm, COMP_LOOP_COMP_LOOP_and_625_itm,
      COMP_LOOP_COMP_LOOP_and_685_itm, COMP_LOOP_COMP_LOOP_and_745_itm, COMP_LOOP_COMP_LOOP_and_805_itm,
      COMP_LOOP_COMP_LOOP_and_865_itm, COMP_LOOP_COMP_LOOP_and_925_itm, STD_LOGIC_VECTOR'(
      and_920_cse & and_925_cse & and_dcpl_621 & and_936_cse & and_940_cse & and_945_cse
      & and_950_cse & and_953_cse & and_957_cse & and_960_cse & and_964_cse & and_966_cse
      & and_970_cse & and_973_cse & and_975_cse & and_978_cse));
  COMP_LOOP_mux1h_857_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_72_itm, COMP_LOOP_COMP_LOOP_and_86_itm,
      COMP_LOOP_COMP_LOOP_and_146_itm, COMP_LOOP_COMP_LOOP_and_206_itm, COMP_LOOP_COMP_LOOP_and_266_itm,
      COMP_LOOP_COMP_LOOP_and_326_itm, COMP_LOOP_COMP_LOOP_and_386_itm, COMP_LOOP_COMP_LOOP_and_446_itm,
      COMP_LOOP_COMP_LOOP_and_506_itm, COMP_LOOP_COMP_LOOP_and_566_itm, COMP_LOOP_COMP_LOOP_and_626_itm,
      COMP_LOOP_COMP_LOOP_and_686_itm, COMP_LOOP_COMP_LOOP_and_746_itm, COMP_LOOP_COMP_LOOP_and_806_itm,
      COMP_LOOP_COMP_LOOP_and_866_itm, COMP_LOOP_COMP_LOOP_and_926_itm, STD_LOGIC_VECTOR'(
      and_920_cse & and_925_cse & and_dcpl_621 & and_936_cse & and_940_cse & and_945_cse
      & and_950_cse & and_953_cse & and_957_cse & and_960_cse & and_964_cse & and_966_cse
      & and_970_cse & and_973_cse & and_975_cse & and_978_cse));
  COMP_LOOP_mux1h_858_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_12_itm, COMP_LOOP_COMP_LOOP_and_87_itm,
      COMP_LOOP_COMP_LOOP_and_147_itm, COMP_LOOP_COMP_LOOP_and_207_itm, COMP_LOOP_COMP_LOOP_and_267_itm,
      COMP_LOOP_COMP_LOOP_and_327_itm, COMP_LOOP_COMP_LOOP_and_387_itm, COMP_LOOP_COMP_LOOP_and_447_itm,
      COMP_LOOP_COMP_LOOP_and_507_itm, COMP_LOOP_COMP_LOOP_and_567_itm, COMP_LOOP_COMP_LOOP_and_627_itm,
      COMP_LOOP_COMP_LOOP_and_687_itm, COMP_LOOP_COMP_LOOP_and_747_itm, COMP_LOOP_COMP_LOOP_and_807_itm,
      COMP_LOOP_COMP_LOOP_and_867_itm, COMP_LOOP_COMP_LOOP_and_927_itm, STD_LOGIC_VECTOR'(
      and_920_cse & and_925_cse & and_dcpl_621 & and_936_cse & and_940_cse & and_945_cse
      & and_950_cse & and_953_cse & and_957_cse & and_960_cse & and_964_cse & and_966_cse
      & and_970_cse & and_973_cse & and_975_cse & and_978_cse));
  COMP_LOOP_mux1h_859_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_13_itm, COMP_LOOP_COMP_LOOP_and_88_itm,
      COMP_LOOP_COMP_LOOP_and_148_itm, COMP_LOOP_COMP_LOOP_and_208_itm, COMP_LOOP_COMP_LOOP_and_268_itm,
      COMP_LOOP_COMP_LOOP_and_328_itm, COMP_LOOP_COMP_LOOP_and_388_itm, COMP_LOOP_COMP_LOOP_and_448_itm,
      COMP_LOOP_COMP_LOOP_and_508_itm, COMP_LOOP_COMP_LOOP_and_568_itm, COMP_LOOP_COMP_LOOP_and_628_itm,
      COMP_LOOP_COMP_LOOP_and_688_itm, COMP_LOOP_COMP_LOOP_and_748_itm, COMP_LOOP_COMP_LOOP_and_808_itm,
      COMP_LOOP_COMP_LOOP_and_868_itm, COMP_LOOP_COMP_LOOP_and_928_itm, STD_LOGIC_VECTOR'(
      and_920_cse & and_925_cse & and_dcpl_621 & and_936_cse & and_940_cse & and_945_cse
      & and_950_cse & and_953_cse & and_957_cse & and_960_cse & and_964_cse & and_966_cse
      & and_970_cse & and_973_cse & and_975_cse & and_978_cse));
  COMP_LOOP_mux1h_860_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_14_itm, COMP_LOOP_COMP_LOOP_and_89_itm,
      COMP_LOOP_COMP_LOOP_and_149_itm, COMP_LOOP_COMP_LOOP_and_209_itm, COMP_LOOP_COMP_LOOP_and_269_itm,
      COMP_LOOP_COMP_LOOP_and_329_itm, COMP_LOOP_COMP_LOOP_and_389_itm, COMP_LOOP_COMP_LOOP_and_449_itm,
      COMP_LOOP_COMP_LOOP_and_509_itm, COMP_LOOP_COMP_LOOP_and_569_itm, COMP_LOOP_COMP_LOOP_and_629_itm,
      COMP_LOOP_COMP_LOOP_and_689_itm, COMP_LOOP_COMP_LOOP_and_749_itm, COMP_LOOP_COMP_LOOP_and_809_itm,
      COMP_LOOP_COMP_LOOP_and_869_itm, COMP_LOOP_COMP_LOOP_and_929_itm, STD_LOGIC_VECTOR'(
      and_920_cse & and_925_cse & and_dcpl_621 & and_936_cse & and_940_cse & and_945_cse
      & and_950_cse & and_953_cse & and_957_cse & and_960_cse & and_964_cse & and_966_cse
      & and_970_cse & and_973_cse & and_975_cse & and_978_cse));
  z_out_5 <= MUX1HOT_v_64_16_2(vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d,
      vec_rsc_0_3_i_qa_d, vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_6_i_qa_d,
      vec_rsc_0_7_i_qa_d, vec_rsc_0_8_i_qa_d, vec_rsc_0_9_i_qa_d, vec_rsc_0_10_i_qa_d,
      vec_rsc_0_11_i_qa_d, vec_rsc_0_12_i_qa_d, vec_rsc_0_13_i_qa_d, vec_rsc_0_14_i_qa_d,
      vec_rsc_0_15_i_qa_d, STD_LOGIC_VECTOR'( COMP_LOOP_mux1h_845_nl & COMP_LOOP_mux1h_846_nl
      & COMP_LOOP_mux1h_847_nl & COMP_LOOP_mux1h_848_nl & COMP_LOOP_mux1h_849_nl
      & COMP_LOOP_mux1h_850_nl & COMP_LOOP_mux1h_851_nl & COMP_LOOP_mux1h_852_nl
      & COMP_LOOP_mux1h_853_nl & COMP_LOOP_mux1h_854_nl & COMP_LOOP_mux1h_855_nl
      & COMP_LOOP_mux1h_856_nl & COMP_LOOP_mux1h_857_nl & COMP_LOOP_mux1h_858_nl
      & COMP_LOOP_mux1h_859_nl & COMP_LOOP_mux1h_860_nl));
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_0_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_0_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_wea : OUT STD_LOGIC;
    vec_rsc_0_0_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_0_1_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_1_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_wea : OUT STD_LOGIC;
    vec_rsc_0_1_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_0_2_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_2_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_wea : OUT STD_LOGIC;
    vec_rsc_0_2_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_0_3_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_3_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_wea : OUT STD_LOGIC;
    vec_rsc_0_3_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_0_4_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_4_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_wea : OUT STD_LOGIC;
    vec_rsc_0_4_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_0_5_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_5_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_wea : OUT STD_LOGIC;
    vec_rsc_0_5_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_0_6_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_6_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_wea : OUT STD_LOGIC;
    vec_rsc_0_6_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_0_7_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_7_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_wea : OUT STD_LOGIC;
    vec_rsc_0_7_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    vec_rsc_0_8_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_8_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_8_wea : OUT STD_LOGIC;
    vec_rsc_0_8_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    vec_rsc_0_9_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_9_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_9_wea : OUT STD_LOGIC;
    vec_rsc_0_9_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    vec_rsc_0_10_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_10_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_10_wea : OUT STD_LOGIC;
    vec_rsc_0_10_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    vec_rsc_0_11_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_11_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_11_wea : OUT STD_LOGIC;
    vec_rsc_0_11_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    vec_rsc_0_12_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_12_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_12_wea : OUT STD_LOGIC;
    vec_rsc_0_12_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    vec_rsc_0_13_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_13_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_13_wea : OUT STD_LOGIC;
    vec_rsc_0_13_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    vec_rsc_0_14_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_14_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_14_wea : OUT STD_LOGIC;
    vec_rsc_0_14_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    vec_rsc_0_15_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_15_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_15_wea : OUT STD_LOGIC;
    vec_rsc_0_15_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC
  );
END inPlaceNTT_DIF;

ARCHITECTURE v7 OF inPlaceNTT_DIF IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_adra_d_iff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da_d_iff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_8_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_9_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_10_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_11_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_12_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_13_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_14_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_15_i_wea_d_iff : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_6_64_64_64_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_0_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_6_64_64_64_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_1_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_6_64_64_64_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_2_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_6_64_64_64_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_3_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_6_64_64_64_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_4_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_6_64_64_64_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_5_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_6_64_64_64_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_6_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_6_64_64_64_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_7_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_6_64_64_64_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_8_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_6_64_64_64_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_9_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_6_64_64_64_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_10_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_6_64_64_64_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_11_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_20_6_64_64_64_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_12_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_21_6_64_64_64_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_13_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_22_6_64_64_64_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_14_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_23_6_64_64_64_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_15_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      p_rsc_triosy_lz : OUT STD_LOGIC;
      r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      r_rsc_triosy_lz : OUT STD_LOGIC;
      vec_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_0_i_adra_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      vec_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_1_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_2_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_3_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_4_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_5_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_6_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_7_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_8_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_9_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_10_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_11_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_12_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_13_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_14_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_15_i_wea_d_pff : OUT STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_core_inst_p_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_r_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_adra_d_pff : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_da_d_pff : STD_LOGIC_VECTOR (63 DOWNTO
      0);

BEGIN
  vec_rsc_0_0_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_6_64_64_64_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_0_i_qa,
      wea => vec_rsc_0_0_wea,
      da => vec_rsc_0_0_i_da,
      adra => vec_rsc_0_0_i_adra,
      adra_d => vec_rsc_0_0_i_adra_d,
      da_d => vec_rsc_0_0_i_da_d,
      qa_d => vec_rsc_0_0_i_qa_d_1,
      wea_d => vec_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_0_i_wea_d_iff
    );
  vec_rsc_0_0_i_qa <= vec_rsc_0_0_qa;
  vec_rsc_0_0_da <= vec_rsc_0_0_i_da;
  vec_rsc_0_0_adra <= vec_rsc_0_0_i_adra;
  vec_rsc_0_0_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_0_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_0_i_qa_d <= vec_rsc_0_0_i_qa_d_1;

  vec_rsc_0_1_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_6_64_64_64_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_1_i_qa,
      wea => vec_rsc_0_1_wea,
      da => vec_rsc_0_1_i_da,
      adra => vec_rsc_0_1_i_adra,
      adra_d => vec_rsc_0_1_i_adra_d,
      da_d => vec_rsc_0_1_i_da_d,
      qa_d => vec_rsc_0_1_i_qa_d_1,
      wea_d => vec_rsc_0_1_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_1_i_wea_d_iff
    );
  vec_rsc_0_1_i_qa <= vec_rsc_0_1_qa;
  vec_rsc_0_1_da <= vec_rsc_0_1_i_da;
  vec_rsc_0_1_adra <= vec_rsc_0_1_i_adra;
  vec_rsc_0_1_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_1_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_1_i_qa_d <= vec_rsc_0_1_i_qa_d_1;

  vec_rsc_0_2_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_6_64_64_64_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_2_i_qa,
      wea => vec_rsc_0_2_wea,
      da => vec_rsc_0_2_i_da,
      adra => vec_rsc_0_2_i_adra,
      adra_d => vec_rsc_0_2_i_adra_d,
      da_d => vec_rsc_0_2_i_da_d,
      qa_d => vec_rsc_0_2_i_qa_d_1,
      wea_d => vec_rsc_0_2_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_2_i_wea_d_iff
    );
  vec_rsc_0_2_i_qa <= vec_rsc_0_2_qa;
  vec_rsc_0_2_da <= vec_rsc_0_2_i_da;
  vec_rsc_0_2_adra <= vec_rsc_0_2_i_adra;
  vec_rsc_0_2_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_2_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_2_i_qa_d <= vec_rsc_0_2_i_qa_d_1;

  vec_rsc_0_3_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_6_64_64_64_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_3_i_qa,
      wea => vec_rsc_0_3_wea,
      da => vec_rsc_0_3_i_da,
      adra => vec_rsc_0_3_i_adra,
      adra_d => vec_rsc_0_3_i_adra_d,
      da_d => vec_rsc_0_3_i_da_d,
      qa_d => vec_rsc_0_3_i_qa_d_1,
      wea_d => vec_rsc_0_3_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_3_i_wea_d_iff
    );
  vec_rsc_0_3_i_qa <= vec_rsc_0_3_qa;
  vec_rsc_0_3_da <= vec_rsc_0_3_i_da;
  vec_rsc_0_3_adra <= vec_rsc_0_3_i_adra;
  vec_rsc_0_3_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_3_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_3_i_qa_d <= vec_rsc_0_3_i_qa_d_1;

  vec_rsc_0_4_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_6_64_64_64_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_4_i_qa,
      wea => vec_rsc_0_4_wea,
      da => vec_rsc_0_4_i_da,
      adra => vec_rsc_0_4_i_adra,
      adra_d => vec_rsc_0_4_i_adra_d,
      da_d => vec_rsc_0_4_i_da_d,
      qa_d => vec_rsc_0_4_i_qa_d_1,
      wea_d => vec_rsc_0_4_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_4_i_wea_d_iff
    );
  vec_rsc_0_4_i_qa <= vec_rsc_0_4_qa;
  vec_rsc_0_4_da <= vec_rsc_0_4_i_da;
  vec_rsc_0_4_adra <= vec_rsc_0_4_i_adra;
  vec_rsc_0_4_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_4_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_4_i_qa_d <= vec_rsc_0_4_i_qa_d_1;

  vec_rsc_0_5_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_6_64_64_64_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_5_i_qa,
      wea => vec_rsc_0_5_wea,
      da => vec_rsc_0_5_i_da,
      adra => vec_rsc_0_5_i_adra,
      adra_d => vec_rsc_0_5_i_adra_d,
      da_d => vec_rsc_0_5_i_da_d,
      qa_d => vec_rsc_0_5_i_qa_d_1,
      wea_d => vec_rsc_0_5_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_5_i_wea_d_iff
    );
  vec_rsc_0_5_i_qa <= vec_rsc_0_5_qa;
  vec_rsc_0_5_da <= vec_rsc_0_5_i_da;
  vec_rsc_0_5_adra <= vec_rsc_0_5_i_adra;
  vec_rsc_0_5_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_5_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_5_i_qa_d <= vec_rsc_0_5_i_qa_d_1;

  vec_rsc_0_6_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_6_64_64_64_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_6_i_qa,
      wea => vec_rsc_0_6_wea,
      da => vec_rsc_0_6_i_da,
      adra => vec_rsc_0_6_i_adra,
      adra_d => vec_rsc_0_6_i_adra_d,
      da_d => vec_rsc_0_6_i_da_d,
      qa_d => vec_rsc_0_6_i_qa_d_1,
      wea_d => vec_rsc_0_6_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_6_i_wea_d_iff
    );
  vec_rsc_0_6_i_qa <= vec_rsc_0_6_qa;
  vec_rsc_0_6_da <= vec_rsc_0_6_i_da;
  vec_rsc_0_6_adra <= vec_rsc_0_6_i_adra;
  vec_rsc_0_6_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_6_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_6_i_qa_d <= vec_rsc_0_6_i_qa_d_1;

  vec_rsc_0_7_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_6_64_64_64_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_7_i_qa,
      wea => vec_rsc_0_7_wea,
      da => vec_rsc_0_7_i_da,
      adra => vec_rsc_0_7_i_adra,
      adra_d => vec_rsc_0_7_i_adra_d,
      da_d => vec_rsc_0_7_i_da_d,
      qa_d => vec_rsc_0_7_i_qa_d_1,
      wea_d => vec_rsc_0_7_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_7_i_wea_d_iff
    );
  vec_rsc_0_7_i_qa <= vec_rsc_0_7_qa;
  vec_rsc_0_7_da <= vec_rsc_0_7_i_da;
  vec_rsc_0_7_adra <= vec_rsc_0_7_i_adra;
  vec_rsc_0_7_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_7_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_7_i_qa_d <= vec_rsc_0_7_i_qa_d_1;

  vec_rsc_0_8_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_6_64_64_64_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_8_i_qa,
      wea => vec_rsc_0_8_wea,
      da => vec_rsc_0_8_i_da,
      adra => vec_rsc_0_8_i_adra,
      adra_d => vec_rsc_0_8_i_adra_d,
      da_d => vec_rsc_0_8_i_da_d,
      qa_d => vec_rsc_0_8_i_qa_d_1,
      wea_d => vec_rsc_0_8_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_8_i_wea_d_iff
    );
  vec_rsc_0_8_i_qa <= vec_rsc_0_8_qa;
  vec_rsc_0_8_da <= vec_rsc_0_8_i_da;
  vec_rsc_0_8_adra <= vec_rsc_0_8_i_adra;
  vec_rsc_0_8_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_8_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_8_i_qa_d <= vec_rsc_0_8_i_qa_d_1;

  vec_rsc_0_9_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_6_64_64_64_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_9_i_qa,
      wea => vec_rsc_0_9_wea,
      da => vec_rsc_0_9_i_da,
      adra => vec_rsc_0_9_i_adra,
      adra_d => vec_rsc_0_9_i_adra_d,
      da_d => vec_rsc_0_9_i_da_d,
      qa_d => vec_rsc_0_9_i_qa_d_1,
      wea_d => vec_rsc_0_9_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_9_i_wea_d_iff
    );
  vec_rsc_0_9_i_qa <= vec_rsc_0_9_qa;
  vec_rsc_0_9_da <= vec_rsc_0_9_i_da;
  vec_rsc_0_9_adra <= vec_rsc_0_9_i_adra;
  vec_rsc_0_9_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_9_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_9_i_qa_d <= vec_rsc_0_9_i_qa_d_1;

  vec_rsc_0_10_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_6_64_64_64_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_10_i_qa,
      wea => vec_rsc_0_10_wea,
      da => vec_rsc_0_10_i_da,
      adra => vec_rsc_0_10_i_adra,
      adra_d => vec_rsc_0_10_i_adra_d,
      da_d => vec_rsc_0_10_i_da_d,
      qa_d => vec_rsc_0_10_i_qa_d_1,
      wea_d => vec_rsc_0_10_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_10_i_wea_d_iff
    );
  vec_rsc_0_10_i_qa <= vec_rsc_0_10_qa;
  vec_rsc_0_10_da <= vec_rsc_0_10_i_da;
  vec_rsc_0_10_adra <= vec_rsc_0_10_i_adra;
  vec_rsc_0_10_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_10_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_10_i_qa_d <= vec_rsc_0_10_i_qa_d_1;

  vec_rsc_0_11_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_6_64_64_64_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_11_i_qa,
      wea => vec_rsc_0_11_wea,
      da => vec_rsc_0_11_i_da,
      adra => vec_rsc_0_11_i_adra,
      adra_d => vec_rsc_0_11_i_adra_d,
      da_d => vec_rsc_0_11_i_da_d,
      qa_d => vec_rsc_0_11_i_qa_d_1,
      wea_d => vec_rsc_0_11_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_11_i_wea_d_iff
    );
  vec_rsc_0_11_i_qa <= vec_rsc_0_11_qa;
  vec_rsc_0_11_da <= vec_rsc_0_11_i_da;
  vec_rsc_0_11_adra <= vec_rsc_0_11_i_adra;
  vec_rsc_0_11_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_11_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_11_i_qa_d <= vec_rsc_0_11_i_qa_d_1;

  vec_rsc_0_12_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_20_6_64_64_64_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_12_i_qa,
      wea => vec_rsc_0_12_wea,
      da => vec_rsc_0_12_i_da,
      adra => vec_rsc_0_12_i_adra,
      adra_d => vec_rsc_0_12_i_adra_d,
      da_d => vec_rsc_0_12_i_da_d,
      qa_d => vec_rsc_0_12_i_qa_d_1,
      wea_d => vec_rsc_0_12_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_12_i_wea_d_iff
    );
  vec_rsc_0_12_i_qa <= vec_rsc_0_12_qa;
  vec_rsc_0_12_da <= vec_rsc_0_12_i_da;
  vec_rsc_0_12_adra <= vec_rsc_0_12_i_adra;
  vec_rsc_0_12_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_12_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_12_i_qa_d <= vec_rsc_0_12_i_qa_d_1;

  vec_rsc_0_13_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_21_6_64_64_64_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_13_i_qa,
      wea => vec_rsc_0_13_wea,
      da => vec_rsc_0_13_i_da,
      adra => vec_rsc_0_13_i_adra,
      adra_d => vec_rsc_0_13_i_adra_d,
      da_d => vec_rsc_0_13_i_da_d,
      qa_d => vec_rsc_0_13_i_qa_d_1,
      wea_d => vec_rsc_0_13_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_13_i_wea_d_iff
    );
  vec_rsc_0_13_i_qa <= vec_rsc_0_13_qa;
  vec_rsc_0_13_da <= vec_rsc_0_13_i_da;
  vec_rsc_0_13_adra <= vec_rsc_0_13_i_adra;
  vec_rsc_0_13_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_13_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_13_i_qa_d <= vec_rsc_0_13_i_qa_d_1;

  vec_rsc_0_14_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_22_6_64_64_64_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_14_i_qa,
      wea => vec_rsc_0_14_wea,
      da => vec_rsc_0_14_i_da,
      adra => vec_rsc_0_14_i_adra,
      adra_d => vec_rsc_0_14_i_adra_d,
      da_d => vec_rsc_0_14_i_da_d,
      qa_d => vec_rsc_0_14_i_qa_d_1,
      wea_d => vec_rsc_0_14_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_14_i_wea_d_iff
    );
  vec_rsc_0_14_i_qa <= vec_rsc_0_14_qa;
  vec_rsc_0_14_da <= vec_rsc_0_14_i_da;
  vec_rsc_0_14_adra <= vec_rsc_0_14_i_adra;
  vec_rsc_0_14_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_14_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_14_i_qa_d <= vec_rsc_0_14_i_qa_d_1;

  vec_rsc_0_15_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_23_6_64_64_64_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_15_i_qa,
      wea => vec_rsc_0_15_wea,
      da => vec_rsc_0_15_i_da,
      adra => vec_rsc_0_15_i_adra,
      adra_d => vec_rsc_0_15_i_adra_d,
      da_d => vec_rsc_0_15_i_da_d,
      qa_d => vec_rsc_0_15_i_qa_d_1,
      wea_d => vec_rsc_0_15_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_15_i_wea_d_iff
    );
  vec_rsc_0_15_i_qa <= vec_rsc_0_15_qa;
  vec_rsc_0_15_da <= vec_rsc_0_15_i_da;
  vec_rsc_0_15_adra <= vec_rsc_0_15_i_adra;
  vec_rsc_0_15_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_15_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_15_i_qa_d <= vec_rsc_0_15_i_qa_d_1;

  inPlaceNTT_DIF_core_inst : inPlaceNTT_DIF_core
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_triosy_0_0_lz => vec_rsc_triosy_0_0_lz,
      vec_rsc_triosy_0_1_lz => vec_rsc_triosy_0_1_lz,
      vec_rsc_triosy_0_2_lz => vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz => vec_rsc_triosy_0_3_lz,
      vec_rsc_triosy_0_4_lz => vec_rsc_triosy_0_4_lz,
      vec_rsc_triosy_0_5_lz => vec_rsc_triosy_0_5_lz,
      vec_rsc_triosy_0_6_lz => vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz => vec_rsc_triosy_0_7_lz,
      vec_rsc_triosy_0_8_lz => vec_rsc_triosy_0_8_lz,
      vec_rsc_triosy_0_9_lz => vec_rsc_triosy_0_9_lz,
      vec_rsc_triosy_0_10_lz => vec_rsc_triosy_0_10_lz,
      vec_rsc_triosy_0_11_lz => vec_rsc_triosy_0_11_lz,
      vec_rsc_triosy_0_12_lz => vec_rsc_triosy_0_12_lz,
      vec_rsc_triosy_0_13_lz => vec_rsc_triosy_0_13_lz,
      vec_rsc_triosy_0_14_lz => vec_rsc_triosy_0_14_lz,
      vec_rsc_triosy_0_15_lz => vec_rsc_triosy_0_15_lz,
      p_rsc_dat => inPlaceNTT_DIF_core_inst_p_rsc_dat,
      p_rsc_triosy_lz => p_rsc_triosy_lz,
      r_rsc_dat => inPlaceNTT_DIF_core_inst_r_rsc_dat,
      r_rsc_triosy_lz => r_rsc_triosy_lz,
      vec_rsc_0_0_i_qa_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_qa_d,
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_1_i_qa_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_1_i_qa_d,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_2_i_qa_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_2_i_qa_d,
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_qa_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_3_i_qa_d,
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_4_i_qa_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_4_i_qa_d,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_5_i_qa_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_5_i_qa_d,
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_qa_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_6_i_qa_d,
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_7_i_qa_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_7_i_qa_d,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_8_i_qa_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_8_i_qa_d,
      vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_9_i_qa_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_9_i_qa_d,
      vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_10_i_qa_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_10_i_qa_d,
      vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_11_i_qa_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_11_i_qa_d,
      vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_12_i_qa_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_12_i_qa_d,
      vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_13_i_qa_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_13_i_qa_d,
      vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_14_i_qa_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_14_i_qa_d,
      vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_15_i_qa_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_15_i_qa_d,
      vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_0_i_adra_d_pff => inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_adra_d_pff,
      vec_rsc_0_0_i_da_d_pff => inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_da_d_pff,
      vec_rsc_0_0_i_wea_d_pff => vec_rsc_0_0_i_wea_d_iff,
      vec_rsc_0_1_i_wea_d_pff => vec_rsc_0_1_i_wea_d_iff,
      vec_rsc_0_2_i_wea_d_pff => vec_rsc_0_2_i_wea_d_iff,
      vec_rsc_0_3_i_wea_d_pff => vec_rsc_0_3_i_wea_d_iff,
      vec_rsc_0_4_i_wea_d_pff => vec_rsc_0_4_i_wea_d_iff,
      vec_rsc_0_5_i_wea_d_pff => vec_rsc_0_5_i_wea_d_iff,
      vec_rsc_0_6_i_wea_d_pff => vec_rsc_0_6_i_wea_d_iff,
      vec_rsc_0_7_i_wea_d_pff => vec_rsc_0_7_i_wea_d_iff,
      vec_rsc_0_8_i_wea_d_pff => vec_rsc_0_8_i_wea_d_iff,
      vec_rsc_0_9_i_wea_d_pff => vec_rsc_0_9_i_wea_d_iff,
      vec_rsc_0_10_i_wea_d_pff => vec_rsc_0_10_i_wea_d_iff,
      vec_rsc_0_11_i_wea_d_pff => vec_rsc_0_11_i_wea_d_iff,
      vec_rsc_0_12_i_wea_d_pff => vec_rsc_0_12_i_wea_d_iff,
      vec_rsc_0_13_i_wea_d_pff => vec_rsc_0_13_i_wea_d_iff,
      vec_rsc_0_14_i_wea_d_pff => vec_rsc_0_14_i_wea_d_iff,
      vec_rsc_0_15_i_wea_d_pff => vec_rsc_0_15_i_wea_d_iff
    );
  inPlaceNTT_DIF_core_inst_p_rsc_dat <= p_rsc_dat;
  inPlaceNTT_DIF_core_inst_r_rsc_dat <= r_rsc_dat;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_qa_d <= vec_rsc_0_0_i_qa_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_1_i_qa_d <= vec_rsc_0_1_i_qa_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_2_i_qa_d <= vec_rsc_0_2_i_qa_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_3_i_qa_d <= vec_rsc_0_3_i_qa_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_4_i_qa_d <= vec_rsc_0_4_i_qa_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_5_i_qa_d <= vec_rsc_0_5_i_qa_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_6_i_qa_d <= vec_rsc_0_6_i_qa_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_7_i_qa_d <= vec_rsc_0_7_i_qa_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_8_i_qa_d <= vec_rsc_0_8_i_qa_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_9_i_qa_d <= vec_rsc_0_9_i_qa_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_10_i_qa_d <= vec_rsc_0_10_i_qa_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_11_i_qa_d <= vec_rsc_0_11_i_qa_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_12_i_qa_d <= vec_rsc_0_12_i_qa_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_13_i_qa_d <= vec_rsc_0_13_i_qa_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_14_i_qa_d <= vec_rsc_0_14_i_qa_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_15_i_qa_d <= vec_rsc_0_15_i_qa_d;
  vec_rsc_0_0_i_adra_d_iff <= inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_adra_d_pff;
  vec_rsc_0_0_i_da_d_iff <= inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_da_d_pff;

END v7;



