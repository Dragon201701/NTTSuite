
--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_pkg_v1 IS

COMPONENT ccs_in_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    dat    : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_in_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    dat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_in_v1;

ARCHITECTURE beh OF ccs_in_v1 IS
BEGIN

  idat <= dat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_out_dreg_pkg_v2 IS

COMPONENT mgc_out_dreg_v2
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    d        : IN  std_logic_vector(width-1 DOWNTO 0);
    z        : OUT std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_out_dreg_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_out_dreg_v2 IS
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    d        : IN  std_logic_vector(width-1 DOWNTO 0);
    z        : OUT std_logic_vector(width-1 DOWNTO 0)
  );
END mgc_out_dreg_v2;

ARCHITECTURE beh OF mgc_out_dreg_v2 IS
BEGIN

  z <= d;

END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/src/funcs.vhd 

-- a package of attributes that give verification tools a hint about
-- the function being implemented
PACKAGE attributes IS
  ATTRIBUTE CALYPTO_FUNC : string;
  ATTRIBUTE CALYPTO_DATA_ORDER : string;
end attributes;

-----------------------------------------------------------------------
-- Package that declares synthesizable functions needed for RTL output
-----------------------------------------------------------------------

LIBRARY ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

PACKAGE funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

   FUNCTION maximum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION minimum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2 : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;
   
-----------------------------------------------------------------
-- logic functions
-----------------------------------------------------------------

   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION or_v (inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- mux functions
-----------------------------------------------------------------

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC_VECTOR;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- latch functions
-----------------------------------------------------------------
   FUNCTION lat_s(dinput: STD_LOGIC       ; clk: STD_LOGIC; doutput: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- tristate functions
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC       ; control: STD_LOGIC) RETURN STD_LOGIC;
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: SIGNED  ) RETURN STD_LOGIC;

   -- RETURN 2 bits (left => lt, right => eq)
   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED;
 
   FUNCTION fabs(arg1: SIGNED  ) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "**" (l, r: UNSIGNED) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "**" (l, r: SIGNED  ) RETURN SIGNED  ;

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-- *_stdar functions use shift functions from std_logic_arith
-----------------------------------------------------------------

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;

   -----------------------------------------------------------------
   -- *_stdar functions use shift functions from std_logic_arith
   -----------------------------------------------------------------
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC;
   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE;
   --FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR ;

   FUNCTION ceil_log2(size : NATURAL) return NATURAL;
   FUNCTION bits(size : NATURAL) return NATURAL;    

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   
END funcs;


--------------------------- B O D Y ----------------------------


PACKAGE BODY funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC IS
     BEGIN IF arg1 THEN RETURN '1'; ELSE RETURN '0'; END IF; END;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
--     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;

   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
     VARIABLE result: STD_LOGIC_VECTOR(0 DOWNTO 0);
   BEGIN
     result := (0 => arg1);
     RETURN result;
   END;

   FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 > arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION minimum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 < arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;

   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := input1'LENGTH;
     ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
     ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     --synopsys translate_off
     FOR i IN len-1 DOWNTO 0 LOOP
       result(i) := resolved(input1a(i) & input2a(i));
     END LOOP;
     --synopsys translate_on
     RETURN result;
   END;

   FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED) RETURN UNSIGNED IS
   BEGIN RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

   FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED) RETURN SIGNED IS
   BEGIN RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

-----------------------------------------------------------------
-- Logic Functions
-----------------------------------------------------------------

   FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;
   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(and_v(inputs, 1)); END;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(or_v(inputs, 1)); END;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(xor_v(inputs, 1)); END;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result AND inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

   FUNCTION or_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     -- this if is added as a quick fix for a bug in catapult evaluating the loop even if inputs'LENGTH==1
     -- see dts0100971279
     IF icnt2 > 1 THEN
       FOR i IN icnt2-1 DOWNTO 1 LOOP
         inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
         result := result OR inputsx(olenM1 DOWNTO 0);
       END LOOP;
     END IF;
     RETURN result;
   END;

   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result XOR inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

-----------------------------------------------------------------
-- Muxes
-----------------------------------------------------------------
   
   FUNCTION mux_sel2_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(1 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 4;
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector( size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "01" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "10" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "11" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel3_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(2 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 8;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "001" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "010" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "011" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN "100" =>
       result := inputs0(5*size-1 DOWNTO 4*size);
     WHEN "101" =>
       result := inputs0(6*size-1 DOWNTO 5*size);
     WHEN "110" =>
       result := inputs0(7*size-1 DOWNTO 6*size);
     WHEN "111" =>
       result := inputs0(8*size-1 DOWNTO 7*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel4_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(3 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 16;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "0000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "0001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "0010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "0011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "0100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "0101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "0110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "0111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "1000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "1001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "1010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "1011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "1100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "1101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "1110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "1111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel5_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(4 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 32;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0 );
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "00001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "00010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "00011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "00100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "00101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "00110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "00111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "01000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "01001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "01010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "01011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "01100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "01101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "01110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "01111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "10000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "10001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "10010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "10011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "10100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "10101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "10110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "10111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "11000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "11001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "11010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "11011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "11100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "11101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "11110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "11111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel6_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(5 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 64;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "000001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "000010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "000011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "000100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "000101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "000110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "000111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "001000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "001001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "001010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "001011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "001100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "001101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "001110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "001111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "010000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "010001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "010010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "010011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "010100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "010101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "010110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "010111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "011000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "011001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "011010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "011011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "011100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "011101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "011110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "011111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN "100000" =>
       result := inputs0( 33*size-1 DOWNTO 32*size);
     WHEN "100001" =>
       result := inputs0( 34*size-1 DOWNTO 33*size);
     WHEN "100010" =>
       result := inputs0( 35*size-1 DOWNTO 34*size);
     WHEN "100011" =>
       result := inputs0( 36*size-1 DOWNTO 35*size);
     WHEN "100100" =>
       result := inputs0( 37*size-1 DOWNTO 36*size);
     WHEN "100101" =>
       result := inputs0( 38*size-1 DOWNTO 37*size);
     WHEN "100110" =>
       result := inputs0( 39*size-1 DOWNTO 38*size);
     WHEN "100111" =>
       result := inputs0( 40*size-1 DOWNTO 39*size);
     WHEN "101000" =>
       result := inputs0( 41*size-1 DOWNTO 40*size);
     WHEN "101001" =>
       result := inputs0( 42*size-1 DOWNTO 41*size);
     WHEN "101010" =>
       result := inputs0( 43*size-1 DOWNTO 42*size);
     WHEN "101011" =>
       result := inputs0( 44*size-1 DOWNTO 43*size);
     WHEN "101100" =>
       result := inputs0( 45*size-1 DOWNTO 44*size);
     WHEN "101101" =>
       result := inputs0( 46*size-1 DOWNTO 45*size);
     WHEN "101110" =>
       result := inputs0( 47*size-1 DOWNTO 46*size);
     WHEN "101111" =>
       result := inputs0( 48*size-1 DOWNTO 47*size);
     WHEN "110000" =>
       result := inputs0( 49*size-1 DOWNTO 48*size);
     WHEN "110001" =>
       result := inputs0( 50*size-1 DOWNTO 49*size);
     WHEN "110010" =>
       result := inputs0( 51*size-1 DOWNTO 50*size);
     WHEN "110011" =>
       result := inputs0( 52*size-1 DOWNTO 51*size);
     WHEN "110100" =>
       result := inputs0( 53*size-1 DOWNTO 52*size);
     WHEN "110101" =>
       result := inputs0( 54*size-1 DOWNTO 53*size);
     WHEN "110110" =>
       result := inputs0( 55*size-1 DOWNTO 54*size);
     WHEN "110111" =>
       result := inputs0( 56*size-1 DOWNTO 55*size);
     WHEN "111000" =>
       result := inputs0( 57*size-1 DOWNTO 56*size);
     WHEN "111001" =>
       result := inputs0( 58*size-1 DOWNTO 57*size);
     WHEN "111010" =>
       result := inputs0( 59*size-1 DOWNTO 58*size);
     WHEN "111011" =>
       result := inputs0( 60*size-1 DOWNTO 59*size);
     WHEN "111100" =>
       result := inputs0( 61*size-1 DOWNTO 60*size);
     WHEN "111101" =>
       result := inputs0( 62*size-1 DOWNTO 61*size);
     WHEN "111110" =>
       result := inputs0( 63*size-1 DOWNTO 62*size);
     WHEN "111111" =>
       result := inputs0( 64*size-1 DOWNTO 63*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS  --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2 SEVERITY FAILURE;
     --synopsys translate_on
       CASE sel IS
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0( size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1  DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0(size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
       RETURN result;
   END;
--   BEGIN RETURN mux_v(inputs, TO_STDLOGICVECTOR(sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     ALIAS    sel0   : STD_LOGIC_VECTOR( sel'LENGTH-1 DOWNTO 0 ) IS sel;

     VARIABLE sellen : INTEGER RANGE 2-sel'LENGTH TO sel'LENGTH;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2**sel'LENGTH;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
     TYPE inputs_array_type is array(natural range <>) of std_logic_vector( olen - 1 DOWNTO 0);
     VARIABLE inputs_array : inputs_array_type( 2**sel'LENGTH - 1 DOWNTO 0);
   BEGIN
     sellen := sel'LENGTH;
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2**sellen SEVERITY FAILURE;
     sellen := 2-sellen;
     --synopsys translate_on
     CASE sellen IS
     WHEN 1 =>
       CASE sel0(0) IS

       WHEN '1' 
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0(  size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1 DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0( size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
     WHEN 2 =>
       result := mux_sel2_v(inputs, not sel);
     WHEN 3 =>
       result := mux_sel3_v(inputs, not sel);
     WHEN 4 =>
       result := mux_sel4_v(inputs, not sel);
     WHEN 5 =>
       result := mux_sel5_v(inputs, not sel);
     WHEN 6 =>
       result := mux_sel6_v(inputs, not sel);
     WHEN others =>
       -- synopsys translate_off
       IF(Is_X(sel0)) THEN
         result := (others => 'X');
       ELSE
       -- synopsys translate_on
         FOR i in 0 to 2**sel'LENGTH - 1 LOOP
           inputs_array(i) := inputs0( ((i + 1) * olen) - 1  DOWNTO i*olen);
         END LOOP;
         result := inputs_array(CONV_INTEGER( (UNSIGNED(NOT sel0)) ));
       -- synopsys translate_off
       END IF;
       -- synopsys translate_on
     END CASE;
     RETURN result;
   END;

 
-----------------------------------------------------------------
-- Latches
-----------------------------------------------------------------

   FUNCTION lat_s(dinput: STD_LOGIC; clk: STD_LOGIC; doutput: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN mux_s(STD_LOGIC_VECTOR'(doutput & dinput), clk); END;

   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR ; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR ) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     --synopsys translate_off
     ASSERT dinput'LENGTH = doutput'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN mux_v(doutput & dinput, clk);
   END;

-----------------------------------------------------------------
-- Tri-States
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC; control: STD_LOGIC) RETURN STD_LOGIC IS
--   BEGIN RETURN TO_STDLOGIC(tri_v(TO_STDLOGICVECTOR(dinput), control)); END;
--
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR ; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
--     VARIABLE result: STD_LOGIC_VECTOR(dinput'range);
--   BEGIN
--     CASE control IS
--     WHEN '0' | 'L' =>
--       result := (others => 'Z');
--     WHEN '1' | 'H' =>
--       FOR i IN dinput'range LOOP
--         result(i) := to_UX01(dinput(i));
--       END LOOP;
--     WHEN others =>
--       -- synopsys translate_off
--       result := (others => 'X');
--       -- synopsys translate_on
--     END CASE;
--     RETURN result;
--   END;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;

   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     VARIABLE diff: UNSIGNED(l'LENGTH DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     diff := ('0'&l) - ('0'&r);
     RETURN diff(l'LENGTH);
   END;
   FUNCTION "<"(l, r: SIGNED  ) RETURN STD_LOGIC IS
   BEGIN
     RETURN (UNSIGNED(l) < UNSIGNED(r)) xor (l(l'LEFT) xor r(r'LEFT));
   END;

   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION "<=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">"(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;
   FUNCTION ">=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;

   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN not or_s(l xor r);
   END;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   --some functions to placate spyglass
   FUNCTION mult_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a*b;
   END mult_natural;

   FUNCTION div_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a/b;
   END div_natural;

   FUNCTION mod_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a mod b;
   END mod_natural;

   FUNCTION add_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a+b;
   END add_unsigned;

   FUNCTION sub_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a-b;
   END sub_unsigned;

   FUNCTION sub_int(a,b : INTEGER) RETURN INTEGER IS
   BEGIN
     return a-b;
   END sub_int;

   FUNCTION concat_0(b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return '0' & b;
   END concat_0;

   FUNCTION concat_uns(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a&b;
   END concat_uns;

   FUNCTION concat_vect(a,b : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     return a&b;
   END concat_vect;





   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED IS
     CONSTANT ninps : NATURAL := arg'LENGTH / width;
     ALIAS    arg0  : UNSIGNED(arg'LENGTH-1 DOWNTO 0) IS arg;
     VARIABLE result: UNSIGNED(width-1 DOWNTO 0);
     VARIABLE from  : INTEGER;
     VARIABLE dto   : INTEGER;
   BEGIN
     --synopsys translate_off
     ASSERT arg'LENGTH = width * ninps SEVERITY FAILURE;
     --synopsys translate_on
     result := (OTHERS => '0');
     FOR i IN ninps-1 DOWNTO 0 LOOP
       --result := result + arg0((i+1)*width-1 DOWNTO i*width);
       from := mult_natural((i+1), width)-1; --2.1.6.3
       dto  := mult_natural(i,width); --2.1.6.3
       result := add_unsigned(result , arg0(from DOWNTO dto) );
     END LOOP;
     RETURN result;
   END faccu;

   FUNCTION  fabs (arg1: SIGNED) RETURN UNSIGNED IS
   BEGIN
     CASE arg1(arg1'LEFT) IS
     WHEN '1'
     --synopsys translate_off
          | 'H'
     --synopsys translate_on
       =>
       RETURN UNSIGNED'("0") - UNSIGNED(arg1);
     WHEN '0'
     --synopsys translate_off
          | 'L'
     --synopsys translate_on
       =>
       RETURN UNSIGNED(arg1);
     WHEN others =>
       RETURN resolve_unsigned(UNSIGNED(arg1), UNSIGNED'("0") - UNSIGNED(arg1));
     END CASE;
   END;

   PROCEDURE divmod(l, r: UNSIGNED; rdiv, rmod: OUT UNSIGNED) IS
     CONSTANT llen: INTEGER := l'LENGTH;
     CONSTANT rlen: INTEGER := r'LENGTH;
     CONSTANT llen_plus_rlen: INTEGER := llen + rlen;
     VARIABLE lbuf: UNSIGNED(llen+rlen-1 DOWNTO 0);
     VARIABLE diff: UNSIGNED(rlen DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT rdiv'LENGTH = llen AND rmod'LENGTH = rlen SEVERITY FAILURE;
     --synopsys translate_on
     lbuf := (others => '0');
     lbuf(llen-1 DOWNTO 0) := l;
     FOR i IN rdiv'range LOOP
       diff := sub_unsigned(lbuf(llen_plus_rlen-1 DOWNTO llen-1) ,(concat_0(r)));
       rdiv(i) := not diff(rlen);
       IF diff(rlen) = '0' THEN
         lbuf(llen_plus_rlen-1 DOWNTO llen-1) := diff;
       END IF;
       lbuf(llen_plus_rlen-1 DOWNTO 1) := lbuf(llen_plus_rlen-2 DOWNTO 0);
     END LOOP;
     rmod := lbuf(llen_plus_rlen-1 DOWNTO llen);
   END divmod;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rdiv;
   END "/";

   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rmod;
   END;

   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN l MOD r; END;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rdiv := UNSIGNED'("0") - rdiv;
     END IF;
     RETURN SIGNED(rdiv); -- overflow problem "1000" / "11"
   END "/";

   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
     CONSTANT rnul: UNSIGNED(r'LENGTH-1 DOWNTO 0) := (others => '0');
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     IF rmod /= rnul AND to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rmod := UNSIGNED(r) + rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "MOD";

   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "REM";

   FUNCTION mult_unsigned(l,r : UNSIGNED) return UNSIGNED is
   BEGIN
     return l*r; 
   END mult_unsigned;

   FUNCTION "**" (l, r : UNSIGNED) RETURN UNSIGNED IS
     CONSTANT llen  : NATURAL := l'LENGTH;
     VARIABLE result: UNSIGNED(llen-1 DOWNTO 0);
     VARIABLE fak   : UNSIGNED(llen-1 DOWNTO 0);
   BEGIN
     fak := l;
     result := (others => '0'); result(0) := '1';
     FOR i IN r'reverse_range LOOP
       --was:result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(result & (result*fak)), r(i)));
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR( concat_uns(result , mult_unsigned(result,fak) )), r(i)));

       fak := mult_unsigned(fak , fak);
     END LOOP;
     RETURN result;
   END "**";

   FUNCTION "**" (l, r : SIGNED) RETURN SIGNED IS
     CONSTANT rlen  : NATURAL := r'LENGTH;
     ALIAS    r0    : SIGNED(0 TO r'LENGTH-1) IS r;
     VARIABLE result: SIGNED(l'range);
   BEGIN
     CASE r(r'LEFT) IS
     WHEN '0'
   --synopsys translate_off
          | 'L'
   --synopsys translate_on
     =>
       result := SIGNED(UNSIGNED(l) ** UNSIGNED(r0(1 TO r'LENGTH-1)));
     WHEN '1'
   --synopsys translate_off
          | 'H'
   --synopsys translate_on
     =>
       result := (others => '0');
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END "**";

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-----------------------------------------------------------------

   FUNCTION add_nat(arg1 : NATURAL; arg2 : NATURAL ) RETURN NATURAL IS
   BEGIN
     return (arg1 + arg2);
   END;
   
--   FUNCTION UNSIGNED_2_BIT_VECTOR(arg1 : NATURAL; arg2 : NATURAL ) RETURN BIT_VECTOR IS
--   BEGIN
--     return (arg1 + arg2);
--   END;
   
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(SIGNED(result), arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
        =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
        =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;


   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     --SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: NATURAL range 1 TO len;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => '0');
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         --was:temp(i2+sw) := result(i2);
         temp_idx := add_nat(i2,sw);
         temp(temp_idx) := result(i2);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: sw_range;
     VARIABLE result_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => sbit);
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         -- was: temp(i2) := result(i2+sw);
         result_idx := add_nat(i2,sw);
         temp(i2) := result(result_idx);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;


   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := arg1'LENGTH;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     VARIABLE temp: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     SUBTYPE sw_range IS NATURAL range 0 TO len-1;
     VARIABLE sw: sw_range;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     result := (others=>'0');
     result := arg1;
     sw := sdir MOD len;
     FOR i IN arg2'reverse_range LOOP
       EXIT WHEN sw = 0;
       IF signd2 AND i = arg2'LEFT THEN 
         sw := sub_int(len,sw); 
       END IF;
       -- temp := result(len-sw-1 DOWNTO 0) & result(len-1 DOWNTO len-sw)
       FOR i2 IN len-1 DOWNTO 0 LOOP
         --was: temp((i2+sw) MOD len) := result(i2);
         temp_idx := add_nat(i2,sw) MOD len;
         temp(temp_idx) := result(i2);
       END LOOP;
       result := mux_v(STD_LOGIC_VECTOR(concat_vect(result,temp)), arg2(i));
       sw := mod_natural(mult_natural(sw,2), len);
     END LOOP;
     RETURN result;
   END frot;

   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, -1); END;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, -1); END;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC IS
     CONSTANT len : INTEGER := vec'LENGTH;
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
   BEGIN
     IF index >= len OR index < 0 THEN
       RETURN 'X';
     END IF;
     RETURN vec0(index);
   END;

   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     CONSTANT indexPwidthM1 : INTEGER := index+width-1; --2.1.6.3
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
     CONSTANT xxx : STD_LOGIC_VECTOR(width-1 DOWNTO 0) := (others => 'X');
   BEGIN
     IF index+width > len OR index < 0 THEN
       RETURN xxx;
     END IF;
     RETURN vec0(indexPwidthM1 DOWNTO index);
   END;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     VARIABLE vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     CONSTANT xxx : STD_LOGIC_VECTOR(len-1 DOWNTO 0) := (others => 'X');
   BEGIN
     vec0 := vec;
     IF index >= len OR index < 0 THEN
       RETURN xxx;
     END IF;
     vec0(index) := dinput;
     RETURN vec0;
   END;

   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE IS
     VARIABLE n_b : POSITIVE;
     VARIABLE p_v : NATURAL;
   BEGIN
     p_v := p;
     FOR i IN 1 TO 32 LOOP
       p_v := div_natural(p_v,2);
       n_b := i;
       EXIT WHEN (p_v = 0);
     END LOOP;
     RETURN n_b;
   END;


--   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
--
--     CONSTANT vlen: INTEGER := vec'LENGTH;
--     CONSTANT ilen: INTEGER := dinput'LENGTH;
--     CONSTANT max_shift: INTEGER := vlen-ilen;
--     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
--     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
--     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
--     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
--     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
--     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
--   BEGIN
--     inp := (others => '0');
--     mask := (others => '0');
--
--     IF index > max_shift OR index < 0 THEN
--       RETURN xxx;
--     END IF;
--
--     shift := CONV_UNSIGNED(index, shift'LENGTH);
--     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
--     mask(ilen-1 DOWNTO 0) := ones;
--     inp := fshl(inp, shift, vlen);
--     mask := fshl(mask, shift, vlen);
--     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
--     RETURN vec0;
--   END;

   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR IS

     type enable_matrix is array (0 to enable'LENGTH-1 ) of std_logic_vector(byte_width-1 downto 0);
     CONSTANT vlen: INTEGER := vec'LENGTH;
     CONSTANT ilen: INTEGER := dinput'LENGTH;
     CONSTANT max_shift: INTEGER := vlen-ilen;
     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask2: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE enables: enable_matrix;
     VARIABLE cat_enables: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0 );
     VARIABLE lsbi : INTEGER;
     VARIABLE msbi : INTEGER;

   BEGIN
     cat_enables := (others => '0');
     lsbi := 0;
     msbi := byte_width-1;
     inp := (others => '0');
     mask := (others => '0');

     IF index > max_shift OR index < 0 THEN
       RETURN xxx;
     END IF;

     --initialize enables
     for i in 0 TO (enable'LENGTH-1) loop
       enables(i)  := (others => enable(i));
       cat_enables(msbi downto lsbi) := enables(i) ;
       lsbi := msbi+1;
       msbi := msbi+byte_width;
     end loop;


     shift := CONV_UNSIGNED(index, shift'LENGTH);
     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
     mask(ilen-1 DOWNTO 0) := UNSIGNED((STD_LOGIC_VECTOR(ones) AND cat_enables));
     inp := fshl(inp, shift, vlen);
     mask := fshl(mask, shift, vlen);
     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
     RETURN vec0;
   END;


   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;
   
   FUNCTION bits(size : NATURAL) return NATURAL is
   begin
     return ceil_log2(size);
   END;

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH) xor conv_std_logic_vector(c, s'LENGTH);
     cout := ( (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH)) or (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) or (conv_std_logic_vector(b, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) );
   END PROCEDURE csa;

   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH);
     cout := (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH));
   END PROCEDURE csha;

END funcs;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_comps.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_comps IS
 
FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
FUNCTION ceil_log2(size : NATURAL) return NATURAL;
 

COMPONENT mgc_not
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_and
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nand
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_or
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xnor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux
  GENERIC (
    width  :  NATURAL;
    ctrlw  :  NATURAL;
    p2ctrlw : NATURAL := 0
  );
  PORT (
    a: in  std_logic_vector(width*(2**ctrlw) - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw            - 1 DOWNTO 0);
    z: out std_logic_vector(width            - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux1hot
  GENERIC (
    width  : NATURAL;
    ctrlw  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ctrlw - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw       - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_reg_pos
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;  -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL  -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_reg_neg
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;   -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_generic_reg
  GENERIC(
   width: natural := 8;
   ph_clk: integer range 0 to 1 := 1; -- clock polarity, 1=rising_edge
   ph_en: integer range 0 to 1 := 1;
   ph_a_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   ph_s_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   a_rst_used: integer range 0 to 1 := 1;
   s_rst_used: integer range 0 to 1 := 0;
   en_used: integer range 0 to 1 := 1
  );
  PORT(
   d: std_logic_vector(width-1 downto 0);
   clk: in std_logic;
   en: in std_logic;
   a_rst: in std_logic;
   s_rst: in std_logic;
   q: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_equal
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a : in  std_logic_vector(width-1 DOWNTO 0);
    b : in  std_logic_vector(width-1 DOWNTO 0);
    eq: out std_logic;
    ne: out std_logic
  );
END COMPONENT;

COMPONENT mgc_shift_l
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rot
  GENERIC (
    width  : NATURAL;
    width_s: NATURAL;
    signd_s: NATURAL;      -- 0:unsigned 1:signed
    sleft  : NATURAL;      -- 0:right 1:left;
    log2w  : NATURAL := 0; -- LOG2(width)
    l2wp2  : NATURAL := 0  --2**LOG2(width)
  );
  PORT (
    a : in  std_logic_vector(width  -1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width  -1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_sub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_ci
  GENERIC (
    width_a : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width_a, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width_a, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width_a,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width_a,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_addc
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add3
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_c : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_c : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(ifeqsel(width_c,0,width,width_c)-1 DOWNTO 0);
    d: in  std_logic_vector(0 DOWNTO 0);
    e: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_sub_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addc_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     c: in std_logic_vector(0 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addsub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    add: in  std_logic;
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_accu
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_abs
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_fast
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_pipe
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2  : NATURAL;
    add_d2  : NATURAL
  );
  PORT (
    a   : in  std_logic_vector(width_a-1 DOWNTO 0);
    b   : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2  : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c   : in  std_logic_vector(width_c-1 DOWNTO 0);
    d   : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2  : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst : in  std_logic_vector(width_e-1 DOWNTO 0);
    z   : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1_pipe
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2   : NATURAL;
    add_d2   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2     : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2     : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_e-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL
  );
  PORT (
    a:   in  std_logic_vector(width_a-1 DOWNTO 0);
    b:   in  std_logic_vector(width_b-1 DOWNTO 0);
    c:   in  std_logic_vector(width_c-1 DOWNTO 0);
    cst: in  std_logic_vector(width_cst-1 DOWNTO 0);
    d:   in  std_logic_vector(width_d-1 DOWNTO 0);
    z:   out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1_pipe
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_cst-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mulacc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2acc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    add_cxd : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    d         : in  std_logic_vector(width_d-1 DOWNTO 0);
    e         : in  std_logic_vector(width_e-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_div
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mod
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rem
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_csa
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     c: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_csha
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_rom
    GENERIC (
      rom_id : natural := 1;
      size : natural := 33;
      width : natural := 32
      );
    PORT (
      data_in : std_logic_vector((size*width)-1 downto 0);
      addr : std_logic_vector(ceil_log2(size)-1 downto 0);
      data_out : out std_logic_vector(width-1 downto 0)
    );
END COMPONENT;

END mgc_comps;

PACKAGE BODY mgc_comps IS
 
   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;
 
END mgc_comps;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_rem IS
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END mgc_rem;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

USE work.funcs.all;

ARCHITECTURE beh OF mgc_rem IS
BEGIN
  z <= std_logic_vector(unsigned(a) rem unsigned(b)) WHEN signd = 0 ELSE
       std_logic_vector(  signed(a) rem   signed(b));
END beh;

--------> ../td_ccore_solutions/modulo_7c916ad59326b02df02b1a80099f3e2761bb_0/rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Mon Aug  2 16:56:58 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    modulo_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;
USE work.mgc_comps.ALL;


ENTITY modulo_core IS
  PORT(
    base_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    m_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    return_rsc_z : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    ccs_ccore_start_rsc_dat : IN STD_LOGIC;
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_srst : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC
  );
END modulo_core;

ARCHITECTURE v1 OF modulo_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL base_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL return_rsci_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL ccs_ccore_start_rsci_idat : STD_LOGIC;
  SIGNAL rem_12_cmp_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_1_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_2_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_3_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_4_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_5_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_6_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_7_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_8_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_9_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_10_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_11_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_1_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_2_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_3_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_4_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_5_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_6_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_7_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_8_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_9_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_10_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_11_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_1_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_2_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_3_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_4_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_5_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_6_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_7_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_8_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_9_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_10_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12_cmp_11_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_tmp : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_tmp : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL and_dcpl_1 : STD_LOGIC;
  SIGNAL and_dcpl_2 : STD_LOGIC;
  SIGNAL and_dcpl_3 : STD_LOGIC;
  SIGNAL and_dcpl_4 : STD_LOGIC;
  SIGNAL and_dcpl_6 : STD_LOGIC;
  SIGNAL and_dcpl_8 : STD_LOGIC;
  SIGNAL and_dcpl_9 : STD_LOGIC;
  SIGNAL and_dcpl_11 : STD_LOGIC;
  SIGNAL and_dcpl_13 : STD_LOGIC;
  SIGNAL and_dcpl_18 : STD_LOGIC;
  SIGNAL and_dcpl_23 : STD_LOGIC;
  SIGNAL and_dcpl_28 : STD_LOGIC;
  SIGNAL and_dcpl_29 : STD_LOGIC;
  SIGNAL and_dcpl_30 : STD_LOGIC;
  SIGNAL and_dcpl_31 : STD_LOGIC;
  SIGNAL and_dcpl_33 : STD_LOGIC;
  SIGNAL and_dcpl_35 : STD_LOGIC;
  SIGNAL and_dcpl_36 : STD_LOGIC;
  SIGNAL and_dcpl_38 : STD_LOGIC;
  SIGNAL and_dcpl_40 : STD_LOGIC;
  SIGNAL and_dcpl_45 : STD_LOGIC;
  SIGNAL and_dcpl_50 : STD_LOGIC;
  SIGNAL and_dcpl_55 : STD_LOGIC;
  SIGNAL and_dcpl_56 : STD_LOGIC;
  SIGNAL and_dcpl_57 : STD_LOGIC;
  SIGNAL and_dcpl_58 : STD_LOGIC;
  SIGNAL and_dcpl_60 : STD_LOGIC;
  SIGNAL and_dcpl_62 : STD_LOGIC;
  SIGNAL and_dcpl_63 : STD_LOGIC;
  SIGNAL and_dcpl_65 : STD_LOGIC;
  SIGNAL and_dcpl_67 : STD_LOGIC;
  SIGNAL and_dcpl_72 : STD_LOGIC;
  SIGNAL and_dcpl_77 : STD_LOGIC;
  SIGNAL and_dcpl_82 : STD_LOGIC;
  SIGNAL and_dcpl_83 : STD_LOGIC;
  SIGNAL and_dcpl_84 : STD_LOGIC;
  SIGNAL and_dcpl_85 : STD_LOGIC;
  SIGNAL and_dcpl_87 : STD_LOGIC;
  SIGNAL and_dcpl_89 : STD_LOGIC;
  SIGNAL and_dcpl_90 : STD_LOGIC;
  SIGNAL and_dcpl_92 : STD_LOGIC;
  SIGNAL and_dcpl_94 : STD_LOGIC;
  SIGNAL and_dcpl_99 : STD_LOGIC;
  SIGNAL and_dcpl_104 : STD_LOGIC;
  SIGNAL and_dcpl_109 : STD_LOGIC;
  SIGNAL and_dcpl_110 : STD_LOGIC;
  SIGNAL and_dcpl_111 : STD_LOGIC;
  SIGNAL and_dcpl_112 : STD_LOGIC;
  SIGNAL and_dcpl_114 : STD_LOGIC;
  SIGNAL and_dcpl_115 : STD_LOGIC;
  SIGNAL and_dcpl_117 : STD_LOGIC;
  SIGNAL and_dcpl_119 : STD_LOGIC;
  SIGNAL and_dcpl_121 : STD_LOGIC;
  SIGNAL and_dcpl_126 : STD_LOGIC;
  SIGNAL and_dcpl_129 : STD_LOGIC;
  SIGNAL and_dcpl_136 : STD_LOGIC;
  SIGNAL and_dcpl_137 : STD_LOGIC;
  SIGNAL and_dcpl_138 : STD_LOGIC;
  SIGNAL and_dcpl_139 : STD_LOGIC;
  SIGNAL and_dcpl_141 : STD_LOGIC;
  SIGNAL and_dcpl_143 : STD_LOGIC;
  SIGNAL and_dcpl_144 : STD_LOGIC;
  SIGNAL and_dcpl_146 : STD_LOGIC;
  SIGNAL and_dcpl_148 : STD_LOGIC;
  SIGNAL and_dcpl_153 : STD_LOGIC;
  SIGNAL and_dcpl_158 : STD_LOGIC;
  SIGNAL and_dcpl_163 : STD_LOGIC;
  SIGNAL and_dcpl_164 : STD_LOGIC;
  SIGNAL and_dcpl_165 : STD_LOGIC;
  SIGNAL and_dcpl_166 : STD_LOGIC;
  SIGNAL and_dcpl_168 : STD_LOGIC;
  SIGNAL and_dcpl_170 : STD_LOGIC;
  SIGNAL and_dcpl_171 : STD_LOGIC;
  SIGNAL and_dcpl_173 : STD_LOGIC;
  SIGNAL and_dcpl_175 : STD_LOGIC;
  SIGNAL and_dcpl_180 : STD_LOGIC;
  SIGNAL and_dcpl_185 : STD_LOGIC;
  SIGNAL and_dcpl_190 : STD_LOGIC;
  SIGNAL and_dcpl_191 : STD_LOGIC;
  SIGNAL and_dcpl_192 : STD_LOGIC;
  SIGNAL and_dcpl_193 : STD_LOGIC;
  SIGNAL and_dcpl_195 : STD_LOGIC;
  SIGNAL and_dcpl_197 : STD_LOGIC;
  SIGNAL and_dcpl_198 : STD_LOGIC;
  SIGNAL and_dcpl_200 : STD_LOGIC;
  SIGNAL and_dcpl_202 : STD_LOGIC;
  SIGNAL and_dcpl_207 : STD_LOGIC;
  SIGNAL and_dcpl_212 : STD_LOGIC;
  SIGNAL and_dcpl_217 : STD_LOGIC;
  SIGNAL and_dcpl_218 : STD_LOGIC;
  SIGNAL and_dcpl_219 : STD_LOGIC;
  SIGNAL and_dcpl_220 : STD_LOGIC;
  SIGNAL and_dcpl_222 : STD_LOGIC;
  SIGNAL and_dcpl_224 : STD_LOGIC;
  SIGNAL and_dcpl_225 : STD_LOGIC;
  SIGNAL and_dcpl_227 : STD_LOGIC;
  SIGNAL and_dcpl_229 : STD_LOGIC;
  SIGNAL and_dcpl_234 : STD_LOGIC;
  SIGNAL and_dcpl_239 : STD_LOGIC;
  SIGNAL and_dcpl_244 : STD_LOGIC;
  SIGNAL and_dcpl_245 : STD_LOGIC;
  SIGNAL and_dcpl_246 : STD_LOGIC;
  SIGNAL and_dcpl_247 : STD_LOGIC;
  SIGNAL and_dcpl_249 : STD_LOGIC;
  SIGNAL and_dcpl_251 : STD_LOGIC;
  SIGNAL and_dcpl_252 : STD_LOGIC;
  SIGNAL and_dcpl_254 : STD_LOGIC;
  SIGNAL and_dcpl_256 : STD_LOGIC;
  SIGNAL and_dcpl_261 : STD_LOGIC;
  SIGNAL and_dcpl_266 : STD_LOGIC;
  SIGNAL and_dcpl_271 : STD_LOGIC;
  SIGNAL and_dcpl_272 : STD_LOGIC;
  SIGNAL and_dcpl_274 : STD_LOGIC;
  SIGNAL and_dcpl_276 : STD_LOGIC;
  SIGNAL and_dcpl_278 : STD_LOGIC;
  SIGNAL and_dcpl_280 : STD_LOGIC;
  SIGNAL and_dcpl_285 : STD_LOGIC;
  SIGNAL and_dcpl_291 : STD_LOGIC;
  SIGNAL and_dcpl_292 : STD_LOGIC;
  SIGNAL and_dcpl_293 : STD_LOGIC;
  SIGNAL and_dcpl_294 : STD_LOGIC;
  SIGNAL and_dcpl_295 : STD_LOGIC;
  SIGNAL and_dcpl_296 : STD_LOGIC;
  SIGNAL and_dcpl_298 : STD_LOGIC;
  SIGNAL not_tmp_54 : STD_LOGIC;
  SIGNAL or_tmp_2 : STD_LOGIC;
  SIGNAL and_dcpl_300 : STD_LOGIC;
  SIGNAL and_dcpl_301 : STD_LOGIC;
  SIGNAL and_dcpl_302 : STD_LOGIC;
  SIGNAL and_dcpl_304 : STD_LOGIC;
  SIGNAL and_tmp : STD_LOGIC;
  SIGNAL and_dcpl_306 : STD_LOGIC;
  SIGNAL and_dcpl_307 : STD_LOGIC;
  SIGNAL and_dcpl_308 : STD_LOGIC;
  SIGNAL and_dcpl_310 : STD_LOGIC;
  SIGNAL and_tmp_2 : STD_LOGIC;
  SIGNAL and_dcpl_312 : STD_LOGIC;
  SIGNAL and_dcpl_313 : STD_LOGIC;
  SIGNAL and_dcpl_314 : STD_LOGIC;
  SIGNAL and_dcpl_316 : STD_LOGIC;
  SIGNAL and_tmp_5 : STD_LOGIC;
  SIGNAL and_dcpl_318 : STD_LOGIC;
  SIGNAL and_tmp_9 : STD_LOGIC;
  SIGNAL and_dcpl_324 : STD_LOGIC;
  SIGNAL and_tmp_13 : STD_LOGIC;
  SIGNAL and_dcpl_330 : STD_LOGIC;
  SIGNAL mux_tmp_19 : STD_LOGIC;
  SIGNAL and_tmp_17 : STD_LOGIC;
  SIGNAL and_dcpl_336 : STD_LOGIC;
  SIGNAL mux_tmp_22 : STD_LOGIC;
  SIGNAL mux_tmp_23 : STD_LOGIC;
  SIGNAL and_tmp_21 : STD_LOGIC;
  SIGNAL and_dcpl_342 : STD_LOGIC;
  SIGNAL mux_tmp_26 : STD_LOGIC;
  SIGNAL mux_tmp_27 : STD_LOGIC;
  SIGNAL mux_tmp_28 : STD_LOGIC;
  SIGNAL and_tmp_25 : STD_LOGIC;
  SIGNAL and_dcpl_348 : STD_LOGIC;
  SIGNAL and_tmp_35 : STD_LOGIC;
  SIGNAL and_dcpl_355 : STD_LOGIC;
  SIGNAL and_dcpl_356 : STD_LOGIC;
  SIGNAL and_dcpl_358 : STD_LOGIC;
  SIGNAL or_tmp_80 : STD_LOGIC;
  SIGNAL and_dcpl_360 : STD_LOGIC;
  SIGNAL and_dcpl_362 : STD_LOGIC;
  SIGNAL mux_tmp_32 : STD_LOGIC;
  SIGNAL and_dcpl_364 : STD_LOGIC;
  SIGNAL and_dcpl_366 : STD_LOGIC;
  SIGNAL mux_tmp_34 : STD_LOGIC;
  SIGNAL mux_tmp_35 : STD_LOGIC;
  SIGNAL and_dcpl_368 : STD_LOGIC;
  SIGNAL and_dcpl_370 : STD_LOGIC;
  SIGNAL mux_tmp_37 : STD_LOGIC;
  SIGNAL mux_tmp_38 : STD_LOGIC;
  SIGNAL mux_tmp_39 : STD_LOGIC;
  SIGNAL and_dcpl_372 : STD_LOGIC;
  SIGNAL mux_tmp_41 : STD_LOGIC;
  SIGNAL mux_tmp_42 : STD_LOGIC;
  SIGNAL mux_tmp_43 : STD_LOGIC;
  SIGNAL mux_tmp_44 : STD_LOGIC;
  SIGNAL and_dcpl_376 : STD_LOGIC;
  SIGNAL mux_tmp_46 : STD_LOGIC;
  SIGNAL mux_tmp_47 : STD_LOGIC;
  SIGNAL mux_tmp_48 : STD_LOGIC;
  SIGNAL mux_tmp_49 : STD_LOGIC;
  SIGNAL mux_tmp_50 : STD_LOGIC;
  SIGNAL and_dcpl_379 : STD_LOGIC;
  SIGNAL mux_tmp_52 : STD_LOGIC;
  SIGNAL mux_tmp_53 : STD_LOGIC;
  SIGNAL mux_tmp_54 : STD_LOGIC;
  SIGNAL mux_tmp_55 : STD_LOGIC;
  SIGNAL mux_tmp_56 : STD_LOGIC;
  SIGNAL mux_tmp_57 : STD_LOGIC;
  SIGNAL and_dcpl_382 : STD_LOGIC;
  SIGNAL mux_tmp_59 : STD_LOGIC;
  SIGNAL mux_tmp_60 : STD_LOGIC;
  SIGNAL mux_tmp_61 : STD_LOGIC;
  SIGNAL mux_tmp_62 : STD_LOGIC;
  SIGNAL mux_tmp_63 : STD_LOGIC;
  SIGNAL mux_tmp_64 : STD_LOGIC;
  SIGNAL mux_tmp_65 : STD_LOGIC;
  SIGNAL and_dcpl_385 : STD_LOGIC;
  SIGNAL mux_tmp_67 : STD_LOGIC;
  SIGNAL mux_tmp_68 : STD_LOGIC;
  SIGNAL mux_tmp_69 : STD_LOGIC;
  SIGNAL mux_tmp_70 : STD_LOGIC;
  SIGNAL mux_tmp_71 : STD_LOGIC;
  SIGNAL mux_tmp_72 : STD_LOGIC;
  SIGNAL mux_tmp_73 : STD_LOGIC;
  SIGNAL mux_tmp_74 : STD_LOGIC;
  SIGNAL and_dcpl_388 : STD_LOGIC;
  SIGNAL and_tmp_44 : STD_LOGIC;
  SIGNAL mux_tmp_76 : STD_LOGIC;
  SIGNAL and_dcpl_393 : STD_LOGIC;
  SIGNAL and_dcpl_394 : STD_LOGIC;
  SIGNAL and_dcpl_395 : STD_LOGIC;
  SIGNAL or_tmp_185 : STD_LOGIC;
  SIGNAL and_dcpl_397 : STD_LOGIC;
  SIGNAL and_dcpl_398 : STD_LOGIC;
  SIGNAL and_tmp_45 : STD_LOGIC;
  SIGNAL and_dcpl_400 : STD_LOGIC;
  SIGNAL and_dcpl_401 : STD_LOGIC;
  SIGNAL and_tmp_47 : STD_LOGIC;
  SIGNAL and_dcpl_403 : STD_LOGIC;
  SIGNAL and_dcpl_404 : STD_LOGIC;
  SIGNAL and_tmp_50 : STD_LOGIC;
  SIGNAL and_dcpl_406 : STD_LOGIC;
  SIGNAL and_tmp_54 : STD_LOGIC;
  SIGNAL and_dcpl_409 : STD_LOGIC;
  SIGNAL and_tmp_58 : STD_LOGIC;
  SIGNAL and_dcpl_413 : STD_LOGIC;
  SIGNAL mux_tmp_84 : STD_LOGIC;
  SIGNAL and_tmp_62 : STD_LOGIC;
  SIGNAL and_dcpl_417 : STD_LOGIC;
  SIGNAL mux_tmp_87 : STD_LOGIC;
  SIGNAL mux_tmp_88 : STD_LOGIC;
  SIGNAL and_tmp_66 : STD_LOGIC;
  SIGNAL and_dcpl_421 : STD_LOGIC;
  SIGNAL mux_tmp_91 : STD_LOGIC;
  SIGNAL mux_tmp_92 : STD_LOGIC;
  SIGNAL mux_tmp_93 : STD_LOGIC;
  SIGNAL and_tmp_70 : STD_LOGIC;
  SIGNAL and_dcpl_425 : STD_LOGIC;
  SIGNAL and_tmp_80 : STD_LOGIC;
  SIGNAL and_dcpl_430 : STD_LOGIC;
  SIGNAL and_dcpl_431 : STD_LOGIC;
  SIGNAL or_tmp_263 : STD_LOGIC;
  SIGNAL and_dcpl_433 : STD_LOGIC;
  SIGNAL mux_tmp_97 : STD_LOGIC;
  SIGNAL and_dcpl_435 : STD_LOGIC;
  SIGNAL mux_tmp_99 : STD_LOGIC;
  SIGNAL mux_tmp_100 : STD_LOGIC;
  SIGNAL and_dcpl_437 : STD_LOGIC;
  SIGNAL mux_tmp_102 : STD_LOGIC;
  SIGNAL mux_tmp_103 : STD_LOGIC;
  SIGNAL mux_tmp_104 : STD_LOGIC;
  SIGNAL and_dcpl_439 : STD_LOGIC;
  SIGNAL mux_tmp_106 : STD_LOGIC;
  SIGNAL mux_tmp_107 : STD_LOGIC;
  SIGNAL mux_tmp_108 : STD_LOGIC;
  SIGNAL mux_tmp_109 : STD_LOGIC;
  SIGNAL and_dcpl_442 : STD_LOGIC;
  SIGNAL mux_tmp_111 : STD_LOGIC;
  SIGNAL mux_tmp_112 : STD_LOGIC;
  SIGNAL mux_tmp_113 : STD_LOGIC;
  SIGNAL mux_tmp_114 : STD_LOGIC;
  SIGNAL mux_tmp_115 : STD_LOGIC;
  SIGNAL and_dcpl_445 : STD_LOGIC;
  SIGNAL mux_tmp_117 : STD_LOGIC;
  SIGNAL mux_tmp_118 : STD_LOGIC;
  SIGNAL mux_tmp_119 : STD_LOGIC;
  SIGNAL mux_tmp_120 : STD_LOGIC;
  SIGNAL mux_tmp_121 : STD_LOGIC;
  SIGNAL mux_tmp_122 : STD_LOGIC;
  SIGNAL and_dcpl_448 : STD_LOGIC;
  SIGNAL mux_tmp_124 : STD_LOGIC;
  SIGNAL mux_tmp_125 : STD_LOGIC;
  SIGNAL mux_tmp_126 : STD_LOGIC;
  SIGNAL mux_tmp_127 : STD_LOGIC;
  SIGNAL mux_tmp_128 : STD_LOGIC;
  SIGNAL mux_tmp_129 : STD_LOGIC;
  SIGNAL mux_tmp_130 : STD_LOGIC;
  SIGNAL and_dcpl_451 : STD_LOGIC;
  SIGNAL mux_tmp_132 : STD_LOGIC;
  SIGNAL mux_tmp_133 : STD_LOGIC;
  SIGNAL mux_tmp_134 : STD_LOGIC;
  SIGNAL mux_tmp_135 : STD_LOGIC;
  SIGNAL mux_tmp_136 : STD_LOGIC;
  SIGNAL mux_tmp_137 : STD_LOGIC;
  SIGNAL mux_tmp_138 : STD_LOGIC;
  SIGNAL mux_tmp_139 : STD_LOGIC;
  SIGNAL and_dcpl_454 : STD_LOGIC;
  SIGNAL and_tmp_89 : STD_LOGIC;
  SIGNAL mux_tmp_141 : STD_LOGIC;
  SIGNAL and_dcpl_460 : STD_LOGIC;
  SIGNAL and_dcpl_461 : STD_LOGIC;
  SIGNAL and_dcpl_462 : STD_LOGIC;
  SIGNAL and_dcpl_463 : STD_LOGIC;
  SIGNAL not_tmp_332 : STD_LOGIC;
  SIGNAL or_tmp_368 : STD_LOGIC;
  SIGNAL and_dcpl_465 : STD_LOGIC;
  SIGNAL and_dcpl_466 : STD_LOGIC;
  SIGNAL and_dcpl_467 : STD_LOGIC;
  SIGNAL and_tmp_90 : STD_LOGIC;
  SIGNAL and_dcpl_469 : STD_LOGIC;
  SIGNAL and_dcpl_470 : STD_LOGIC;
  SIGNAL and_dcpl_471 : STD_LOGIC;
  SIGNAL and_tmp_92 : STD_LOGIC;
  SIGNAL and_dcpl_473 : STD_LOGIC;
  SIGNAL and_dcpl_474 : STD_LOGIC;
  SIGNAL and_dcpl_475 : STD_LOGIC;
  SIGNAL and_tmp_95 : STD_LOGIC;
  SIGNAL and_dcpl_477 : STD_LOGIC;
  SIGNAL and_tmp_99 : STD_LOGIC;
  SIGNAL and_dcpl_480 : STD_LOGIC;
  SIGNAL and_tmp_103 : STD_LOGIC;
  SIGNAL and_dcpl_483 : STD_LOGIC;
  SIGNAL mux_tmp_149 : STD_LOGIC;
  SIGNAL and_tmp_107 : STD_LOGIC;
  SIGNAL and_dcpl_486 : STD_LOGIC;
  SIGNAL mux_tmp_152 : STD_LOGIC;
  SIGNAL mux_tmp_153 : STD_LOGIC;
  SIGNAL and_tmp_111 : STD_LOGIC;
  SIGNAL and_dcpl_489 : STD_LOGIC;
  SIGNAL mux_tmp_156 : STD_LOGIC;
  SIGNAL mux_tmp_157 : STD_LOGIC;
  SIGNAL mux_tmp_158 : STD_LOGIC;
  SIGNAL and_tmp_115 : STD_LOGIC;
  SIGNAL and_dcpl_492 : STD_LOGIC;
  SIGNAL and_tmp_125 : STD_LOGIC;
  SIGNAL and_dcpl_498 : STD_LOGIC;
  SIGNAL or_tmp_446 : STD_LOGIC;
  SIGNAL and_dcpl_500 : STD_LOGIC;
  SIGNAL mux_tmp_162 : STD_LOGIC;
  SIGNAL and_dcpl_502 : STD_LOGIC;
  SIGNAL mux_tmp_164 : STD_LOGIC;
  SIGNAL mux_tmp_165 : STD_LOGIC;
  SIGNAL and_dcpl_504 : STD_LOGIC;
  SIGNAL mux_tmp_167 : STD_LOGIC;
  SIGNAL mux_tmp_168 : STD_LOGIC;
  SIGNAL mux_tmp_169 : STD_LOGIC;
  SIGNAL and_dcpl_506 : STD_LOGIC;
  SIGNAL mux_tmp_171 : STD_LOGIC;
  SIGNAL mux_tmp_172 : STD_LOGIC;
  SIGNAL mux_tmp_173 : STD_LOGIC;
  SIGNAL mux_tmp_174 : STD_LOGIC;
  SIGNAL and_dcpl_508 : STD_LOGIC;
  SIGNAL mux_tmp_176 : STD_LOGIC;
  SIGNAL mux_tmp_177 : STD_LOGIC;
  SIGNAL mux_tmp_178 : STD_LOGIC;
  SIGNAL mux_tmp_179 : STD_LOGIC;
  SIGNAL mux_tmp_180 : STD_LOGIC;
  SIGNAL and_dcpl_510 : STD_LOGIC;
  SIGNAL mux_tmp_182 : STD_LOGIC;
  SIGNAL mux_tmp_183 : STD_LOGIC;
  SIGNAL mux_tmp_184 : STD_LOGIC;
  SIGNAL mux_tmp_185 : STD_LOGIC;
  SIGNAL mux_tmp_186 : STD_LOGIC;
  SIGNAL mux_tmp_187 : STD_LOGIC;
  SIGNAL and_dcpl_512 : STD_LOGIC;
  SIGNAL mux_tmp_189 : STD_LOGIC;
  SIGNAL mux_tmp_190 : STD_LOGIC;
  SIGNAL mux_tmp_191 : STD_LOGIC;
  SIGNAL mux_tmp_192 : STD_LOGIC;
  SIGNAL mux_tmp_193 : STD_LOGIC;
  SIGNAL mux_tmp_194 : STD_LOGIC;
  SIGNAL mux_tmp_195 : STD_LOGIC;
  SIGNAL and_dcpl_514 : STD_LOGIC;
  SIGNAL mux_tmp_197 : STD_LOGIC;
  SIGNAL mux_tmp_198 : STD_LOGIC;
  SIGNAL mux_tmp_199 : STD_LOGIC;
  SIGNAL mux_tmp_200 : STD_LOGIC;
  SIGNAL mux_tmp_201 : STD_LOGIC;
  SIGNAL mux_tmp_202 : STD_LOGIC;
  SIGNAL mux_tmp_203 : STD_LOGIC;
  SIGNAL mux_tmp_204 : STD_LOGIC;
  SIGNAL and_dcpl_516 : STD_LOGIC;
  SIGNAL and_tmp_134 : STD_LOGIC;
  SIGNAL mux_tmp_206 : STD_LOGIC;
  SIGNAL and_dcpl_520 : STD_LOGIC;
  SIGNAL and_dcpl_521 : STD_LOGIC;
  SIGNAL or_tmp_551 : STD_LOGIC;
  SIGNAL and_dcpl_523 : STD_LOGIC;
  SIGNAL and_dcpl_524 : STD_LOGIC;
  SIGNAL and_tmp_135 : STD_LOGIC;
  SIGNAL and_dcpl_526 : STD_LOGIC;
  SIGNAL and_dcpl_527 : STD_LOGIC;
  SIGNAL and_tmp_137 : STD_LOGIC;
  SIGNAL and_dcpl_529 : STD_LOGIC;
  SIGNAL and_dcpl_530 : STD_LOGIC;
  SIGNAL and_tmp_140 : STD_LOGIC;
  SIGNAL and_dcpl_532 : STD_LOGIC;
  SIGNAL and_tmp_144 : STD_LOGIC;
  SIGNAL and_dcpl_534 : STD_LOGIC;
  SIGNAL and_tmp_148 : STD_LOGIC;
  SIGNAL and_dcpl_536 : STD_LOGIC;
  SIGNAL mux_tmp_214 : STD_LOGIC;
  SIGNAL and_tmp_152 : STD_LOGIC;
  SIGNAL and_dcpl_538 : STD_LOGIC;
  SIGNAL mux_tmp_217 : STD_LOGIC;
  SIGNAL mux_tmp_218 : STD_LOGIC;
  SIGNAL and_tmp_156 : STD_LOGIC;
  SIGNAL and_dcpl_540 : STD_LOGIC;
  SIGNAL mux_tmp_221 : STD_LOGIC;
  SIGNAL mux_tmp_222 : STD_LOGIC;
  SIGNAL mux_tmp_223 : STD_LOGIC;
  SIGNAL and_tmp_160 : STD_LOGIC;
  SIGNAL and_dcpl_542 : STD_LOGIC;
  SIGNAL and_tmp_170 : STD_LOGIC;
  SIGNAL and_dcpl_546 : STD_LOGIC;
  SIGNAL or_tmp_629 : STD_LOGIC;
  SIGNAL and_dcpl_548 : STD_LOGIC;
  SIGNAL mux_tmp_227 : STD_LOGIC;
  SIGNAL and_dcpl_550 : STD_LOGIC;
  SIGNAL mux_tmp_229 : STD_LOGIC;
  SIGNAL mux_tmp_230 : STD_LOGIC;
  SIGNAL and_dcpl_552 : STD_LOGIC;
  SIGNAL mux_tmp_232 : STD_LOGIC;
  SIGNAL mux_tmp_233 : STD_LOGIC;
  SIGNAL mux_tmp_234 : STD_LOGIC;
  SIGNAL and_dcpl_554 : STD_LOGIC;
  SIGNAL mux_tmp_236 : STD_LOGIC;
  SIGNAL mux_tmp_237 : STD_LOGIC;
  SIGNAL mux_tmp_238 : STD_LOGIC;
  SIGNAL mux_tmp_239 : STD_LOGIC;
  SIGNAL and_dcpl_556 : STD_LOGIC;
  SIGNAL mux_tmp_241 : STD_LOGIC;
  SIGNAL mux_tmp_242 : STD_LOGIC;
  SIGNAL mux_tmp_243 : STD_LOGIC;
  SIGNAL mux_tmp_244 : STD_LOGIC;
  SIGNAL mux_tmp_245 : STD_LOGIC;
  SIGNAL and_dcpl_558 : STD_LOGIC;
  SIGNAL mux_tmp_247 : STD_LOGIC;
  SIGNAL mux_tmp_248 : STD_LOGIC;
  SIGNAL mux_tmp_249 : STD_LOGIC;
  SIGNAL mux_tmp_250 : STD_LOGIC;
  SIGNAL mux_tmp_251 : STD_LOGIC;
  SIGNAL mux_tmp_252 : STD_LOGIC;
  SIGNAL and_dcpl_560 : STD_LOGIC;
  SIGNAL mux_tmp_254 : STD_LOGIC;
  SIGNAL mux_tmp_255 : STD_LOGIC;
  SIGNAL mux_tmp_256 : STD_LOGIC;
  SIGNAL mux_tmp_257 : STD_LOGIC;
  SIGNAL mux_tmp_258 : STD_LOGIC;
  SIGNAL mux_tmp_259 : STD_LOGIC;
  SIGNAL mux_tmp_260 : STD_LOGIC;
  SIGNAL and_dcpl_562 : STD_LOGIC;
  SIGNAL mux_tmp_262 : STD_LOGIC;
  SIGNAL mux_tmp_263 : STD_LOGIC;
  SIGNAL mux_tmp_264 : STD_LOGIC;
  SIGNAL mux_tmp_265 : STD_LOGIC;
  SIGNAL mux_tmp_266 : STD_LOGIC;
  SIGNAL mux_tmp_267 : STD_LOGIC;
  SIGNAL mux_tmp_268 : STD_LOGIC;
  SIGNAL mux_tmp_269 : STD_LOGIC;
  SIGNAL and_dcpl_564 : STD_LOGIC;
  SIGNAL and_tmp_179 : STD_LOGIC;
  SIGNAL mux_tmp_271 : STD_LOGIC;
  SIGNAL and_dcpl_568 : STD_LOGIC;
  SIGNAL and_dcpl_569 : STD_LOGIC;
  SIGNAL and_dcpl_570 : STD_LOGIC;
  SIGNAL and_dcpl_571 : STD_LOGIC;
  SIGNAL or_tmp_733 : STD_LOGIC;
  SIGNAL and_dcpl_573 : STD_LOGIC;
  SIGNAL and_dcpl_574 : STD_LOGIC;
  SIGNAL and_dcpl_575 : STD_LOGIC;
  SIGNAL and_tmp_180 : STD_LOGIC;
  SIGNAL and_dcpl_577 : STD_LOGIC;
  SIGNAL and_dcpl_578 : STD_LOGIC;
  SIGNAL and_dcpl_579 : STD_LOGIC;
  SIGNAL and_tmp_182 : STD_LOGIC;
  SIGNAL and_dcpl_581 : STD_LOGIC;
  SIGNAL and_dcpl_582 : STD_LOGIC;
  SIGNAL and_dcpl_583 : STD_LOGIC;
  SIGNAL and_tmp_185 : STD_LOGIC;
  SIGNAL and_dcpl_585 : STD_LOGIC;
  SIGNAL and_tmp_189 : STD_LOGIC;
  SIGNAL and_dcpl_589 : STD_LOGIC;
  SIGNAL and_tmp_193 : STD_LOGIC;
  SIGNAL and_dcpl_593 : STD_LOGIC;
  SIGNAL mux_tmp_279 : STD_LOGIC;
  SIGNAL and_tmp_197 : STD_LOGIC;
  SIGNAL and_dcpl_597 : STD_LOGIC;
  SIGNAL mux_tmp_282 : STD_LOGIC;
  SIGNAL mux_tmp_283 : STD_LOGIC;
  SIGNAL and_tmp_201 : STD_LOGIC;
  SIGNAL and_dcpl_601 : STD_LOGIC;
  SIGNAL mux_tmp_286 : STD_LOGIC;
  SIGNAL mux_tmp_287 : STD_LOGIC;
  SIGNAL mux_tmp_288 : STD_LOGIC;
  SIGNAL and_tmp_205 : STD_LOGIC;
  SIGNAL and_dcpl_605 : STD_LOGIC;
  SIGNAL or_tmp_808 : STD_LOGIC;
  SIGNAL mux_tmp_291 : STD_LOGIC;
  SIGNAL mux_tmp_292 : STD_LOGIC;
  SIGNAL mux_tmp_293 : STD_LOGIC;
  SIGNAL mux_tmp_294 : STD_LOGIC;
  SIGNAL mux_tmp_295 : STD_LOGIC;
  SIGNAL mux_tmp_296 : STD_LOGIC;
  SIGNAL mux_tmp_297 : STD_LOGIC;
  SIGNAL mux_tmp_298 : STD_LOGIC;
  SIGNAL and_tmp_206 : STD_LOGIC;
  SIGNAL and_dcpl_610 : STD_LOGIC;
  SIGNAL or_tmp_820 : STD_LOGIC;
  SIGNAL and_dcpl_612 : STD_LOGIC;
  SIGNAL mux_tmp_301 : STD_LOGIC;
  SIGNAL and_dcpl_614 : STD_LOGIC;
  SIGNAL mux_tmp_303 : STD_LOGIC;
  SIGNAL mux_tmp_304 : STD_LOGIC;
  SIGNAL and_dcpl_616 : STD_LOGIC;
  SIGNAL mux_tmp_306 : STD_LOGIC;
  SIGNAL mux_tmp_307 : STD_LOGIC;
  SIGNAL mux_tmp_308 : STD_LOGIC;
  SIGNAL and_dcpl_618 : STD_LOGIC;
  SIGNAL mux_tmp_310 : STD_LOGIC;
  SIGNAL mux_tmp_311 : STD_LOGIC;
  SIGNAL mux_tmp_312 : STD_LOGIC;
  SIGNAL mux_tmp_313 : STD_LOGIC;
  SIGNAL and_dcpl_622 : STD_LOGIC;
  SIGNAL mux_tmp_315 : STD_LOGIC;
  SIGNAL mux_tmp_316 : STD_LOGIC;
  SIGNAL mux_tmp_317 : STD_LOGIC;
  SIGNAL mux_tmp_318 : STD_LOGIC;
  SIGNAL mux_tmp_319 : STD_LOGIC;
  SIGNAL and_dcpl_625 : STD_LOGIC;
  SIGNAL mux_tmp_321 : STD_LOGIC;
  SIGNAL mux_tmp_322 : STD_LOGIC;
  SIGNAL mux_tmp_323 : STD_LOGIC;
  SIGNAL mux_tmp_324 : STD_LOGIC;
  SIGNAL mux_tmp_325 : STD_LOGIC;
  SIGNAL mux_tmp_326 : STD_LOGIC;
  SIGNAL and_dcpl_628 : STD_LOGIC;
  SIGNAL mux_tmp_328 : STD_LOGIC;
  SIGNAL mux_tmp_329 : STD_LOGIC;
  SIGNAL mux_tmp_330 : STD_LOGIC;
  SIGNAL mux_tmp_331 : STD_LOGIC;
  SIGNAL mux_tmp_332 : STD_LOGIC;
  SIGNAL mux_tmp_333 : STD_LOGIC;
  SIGNAL mux_tmp_334 : STD_LOGIC;
  SIGNAL and_dcpl_631 : STD_LOGIC;
  SIGNAL mux_tmp_336 : STD_LOGIC;
  SIGNAL mux_tmp_337 : STD_LOGIC;
  SIGNAL mux_tmp_338 : STD_LOGIC;
  SIGNAL mux_tmp_339 : STD_LOGIC;
  SIGNAL mux_tmp_340 : STD_LOGIC;
  SIGNAL mux_tmp_341 : STD_LOGIC;
  SIGNAL mux_tmp_342 : STD_LOGIC;
  SIGNAL mux_tmp_343 : STD_LOGIC;
  SIGNAL and_dcpl_634 : STD_LOGIC;
  SIGNAL or_tmp_921 : STD_LOGIC;
  SIGNAL mux_tmp_345 : STD_LOGIC;
  SIGNAL mux_tmp_346 : STD_LOGIC;
  SIGNAL mux_tmp_347 : STD_LOGIC;
  SIGNAL mux_tmp_348 : STD_LOGIC;
  SIGNAL mux_tmp_349 : STD_LOGIC;
  SIGNAL mux_tmp_350 : STD_LOGIC;
  SIGNAL mux_tmp_351 : STD_LOGIC;
  SIGNAL mux_tmp_352 : STD_LOGIC;
  SIGNAL mux_tmp_353 : STD_LOGIC;
  SIGNAL mux_tmp_354 : STD_LOGIC;
  SIGNAL and_dcpl_638 : STD_LOGIC;
  SIGNAL and_dcpl_639 : STD_LOGIC;
  SIGNAL or_tmp_934 : STD_LOGIC;
  SIGNAL and_dcpl_641 : STD_LOGIC;
  SIGNAL and_dcpl_642 : STD_LOGIC;
  SIGNAL and_tmp_207 : STD_LOGIC;
  SIGNAL and_dcpl_644 : STD_LOGIC;
  SIGNAL and_dcpl_645 : STD_LOGIC;
  SIGNAL and_tmp_209 : STD_LOGIC;
  SIGNAL and_dcpl_647 : STD_LOGIC;
  SIGNAL and_dcpl_648 : STD_LOGIC;
  SIGNAL and_tmp_212 : STD_LOGIC;
  SIGNAL and_dcpl_650 : STD_LOGIC;
  SIGNAL and_tmp_216 : STD_LOGIC;
  SIGNAL and_dcpl_653 : STD_LOGIC;
  SIGNAL and_tmp_220 : STD_LOGIC;
  SIGNAL and_dcpl_657 : STD_LOGIC;
  SIGNAL mux_tmp_362 : STD_LOGIC;
  SIGNAL and_tmp_224 : STD_LOGIC;
  SIGNAL and_dcpl_661 : STD_LOGIC;
  SIGNAL mux_tmp_365 : STD_LOGIC;
  SIGNAL mux_tmp_366 : STD_LOGIC;
  SIGNAL and_tmp_228 : STD_LOGIC;
  SIGNAL and_dcpl_665 : STD_LOGIC;
  SIGNAL mux_tmp_369 : STD_LOGIC;
  SIGNAL mux_tmp_370 : STD_LOGIC;
  SIGNAL mux_tmp_371 : STD_LOGIC;
  SIGNAL and_tmp_232 : STD_LOGIC;
  SIGNAL and_dcpl_669 : STD_LOGIC;
  SIGNAL or_tmp_1009 : STD_LOGIC;
  SIGNAL mux_tmp_374 : STD_LOGIC;
  SIGNAL mux_tmp_375 : STD_LOGIC;
  SIGNAL mux_tmp_376 : STD_LOGIC;
  SIGNAL mux_tmp_377 : STD_LOGIC;
  SIGNAL mux_tmp_378 : STD_LOGIC;
  SIGNAL mux_tmp_379 : STD_LOGIC;
  SIGNAL mux_tmp_380 : STD_LOGIC;
  SIGNAL mux_tmp_381 : STD_LOGIC;
  SIGNAL and_tmp_233 : STD_LOGIC;
  SIGNAL and_dcpl_673 : STD_LOGIC;
  SIGNAL or_tmp_1021 : STD_LOGIC;
  SIGNAL and_dcpl_675 : STD_LOGIC;
  SIGNAL mux_tmp_384 : STD_LOGIC;
  SIGNAL and_dcpl_677 : STD_LOGIC;
  SIGNAL mux_tmp_386 : STD_LOGIC;
  SIGNAL mux_tmp_387 : STD_LOGIC;
  SIGNAL and_dcpl_679 : STD_LOGIC;
  SIGNAL mux_tmp_389 : STD_LOGIC;
  SIGNAL mux_tmp_390 : STD_LOGIC;
  SIGNAL mux_tmp_391 : STD_LOGIC;
  SIGNAL and_dcpl_681 : STD_LOGIC;
  SIGNAL mux_tmp_393 : STD_LOGIC;
  SIGNAL mux_tmp_394 : STD_LOGIC;
  SIGNAL mux_tmp_395 : STD_LOGIC;
  SIGNAL mux_tmp_396 : STD_LOGIC;
  SIGNAL and_dcpl_684 : STD_LOGIC;
  SIGNAL mux_tmp_398 : STD_LOGIC;
  SIGNAL mux_tmp_399 : STD_LOGIC;
  SIGNAL mux_tmp_400 : STD_LOGIC;
  SIGNAL mux_tmp_401 : STD_LOGIC;
  SIGNAL mux_tmp_402 : STD_LOGIC;
  SIGNAL and_dcpl_687 : STD_LOGIC;
  SIGNAL mux_tmp_404 : STD_LOGIC;
  SIGNAL mux_tmp_405 : STD_LOGIC;
  SIGNAL mux_tmp_406 : STD_LOGIC;
  SIGNAL mux_tmp_407 : STD_LOGIC;
  SIGNAL mux_tmp_408 : STD_LOGIC;
  SIGNAL mux_tmp_409 : STD_LOGIC;
  SIGNAL and_dcpl_690 : STD_LOGIC;
  SIGNAL mux_tmp_411 : STD_LOGIC;
  SIGNAL mux_tmp_412 : STD_LOGIC;
  SIGNAL mux_tmp_413 : STD_LOGIC;
  SIGNAL mux_tmp_414 : STD_LOGIC;
  SIGNAL mux_tmp_415 : STD_LOGIC;
  SIGNAL mux_tmp_416 : STD_LOGIC;
  SIGNAL mux_tmp_417 : STD_LOGIC;
  SIGNAL and_dcpl_693 : STD_LOGIC;
  SIGNAL mux_tmp_419 : STD_LOGIC;
  SIGNAL mux_tmp_420 : STD_LOGIC;
  SIGNAL mux_tmp_421 : STD_LOGIC;
  SIGNAL mux_tmp_422 : STD_LOGIC;
  SIGNAL mux_tmp_423 : STD_LOGIC;
  SIGNAL mux_tmp_424 : STD_LOGIC;
  SIGNAL mux_tmp_425 : STD_LOGIC;
  SIGNAL mux_tmp_426 : STD_LOGIC;
  SIGNAL and_dcpl_696 : STD_LOGIC;
  SIGNAL or_tmp_1122 : STD_LOGIC;
  SIGNAL mux_tmp_428 : STD_LOGIC;
  SIGNAL mux_tmp_429 : STD_LOGIC;
  SIGNAL mux_tmp_430 : STD_LOGIC;
  SIGNAL mux_tmp_431 : STD_LOGIC;
  SIGNAL mux_tmp_432 : STD_LOGIC;
  SIGNAL mux_tmp_433 : STD_LOGIC;
  SIGNAL mux_tmp_434 : STD_LOGIC;
  SIGNAL mux_tmp_435 : STD_LOGIC;
  SIGNAL mux_tmp_436 : STD_LOGIC;
  SIGNAL mux_tmp_437 : STD_LOGIC;
  SIGNAL rem_12cyc_st_10_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_10_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_9_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_9_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_8_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_8_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_7_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_7_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_6_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_6_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_5_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_5_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_4_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_4_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_3_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_3_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_2_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_2_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_12_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL result_sva_duc : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12cyc_st_12_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL COMP_LOOP_asn_itm_12 : STD_LOGIC;
  SIGNAL main_stage_0_13 : STD_LOGIC;
  SIGNAL main_stage_0_3 : STD_LOGIC;
  SIGNAL COMP_LOOP_asn_itm_1 : STD_LOGIC;
  SIGNAL main_stage_0_2 : STD_LOGIC;
  SIGNAL main_stage_0_4 : STD_LOGIC;
  SIGNAL COMP_LOOP_asn_itm_2 : STD_LOGIC;
  SIGNAL main_stage_0_5 : STD_LOGIC;
  SIGNAL COMP_LOOP_asn_itm_3 : STD_LOGIC;
  SIGNAL main_stage_0_6 : STD_LOGIC;
  SIGNAL COMP_LOOP_asn_itm_4 : STD_LOGIC;
  SIGNAL COMP_LOOP_asn_itm_5 : STD_LOGIC;
  SIGNAL main_stage_0_8 : STD_LOGIC;
  SIGNAL COMP_LOOP_asn_itm_7 : STD_LOGIC;
  SIGNAL main_stage_0_9 : STD_LOGIC;
  SIGNAL COMP_LOOP_asn_itm_8 : STD_LOGIC;
  SIGNAL main_stage_0_10 : STD_LOGIC;
  SIGNAL COMP_LOOP_asn_itm_9 : STD_LOGIC;
  SIGNAL main_stage_0_7 : STD_LOGIC;
  SIGNAL COMP_LOOP_asn_itm_6 : STD_LOGIC;
  SIGNAL main_stage_0_11 : STD_LOGIC;
  SIGNAL COMP_LOOP_asn_itm_10 : STD_LOGIC;
  SIGNAL COMP_LOOP_and_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_2_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_4_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_6_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_8_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_10_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_12_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_14_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_16_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_18_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_20_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_22_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_24_cse : STD_LOGIC;
  SIGNAL or_1_cse : STD_LOGIC;
  SIGNAL or_6_cse : STD_LOGIC;
  SIGNAL or_10_cse : STD_LOGIC;
  SIGNAL or_15_cse : STD_LOGIC;
  SIGNAL or_21_cse : STD_LOGIC;
  SIGNAL or_28_cse : STD_LOGIC;
  SIGNAL or_37_cse : STD_LOGIC;
  SIGNAL or_48_cse : STD_LOGIC;
  SIGNAL or_83_cse : STD_LOGIC;
  SIGNAL nand_276_cse : STD_LOGIC;
  SIGNAL or_88_cse : STD_LOGIC;
  SIGNAL nand_274_cse : STD_LOGIC;
  SIGNAL or_93_cse : STD_LOGIC;
  SIGNAL nand_271_cse : STD_LOGIC;
  SIGNAL or_100_cse : STD_LOGIC;
  SIGNAL nand_267_cse : STD_LOGIC;
  SIGNAL or_109_cse : STD_LOGIC;
  SIGNAL or_120_cse : STD_LOGIC;
  SIGNAL or_133_cse : STD_LOGIC;
  SIGNAL or_148_cse : STD_LOGIC;
  SIGNAL or_190_cse : STD_LOGIC;
  SIGNAL or_195_cse : STD_LOGIC;
  SIGNAL or_199_cse : STD_LOGIC;
  SIGNAL or_204_cse : STD_LOGIC;
  SIGNAL or_210_cse : STD_LOGIC;
  SIGNAL or_217_cse : STD_LOGIC;
  SIGNAL or_226_cse : STD_LOGIC;
  SIGNAL or_237_cse : STD_LOGIC;
  SIGNAL or_270_cse : STD_LOGIC;
  SIGNAL or_275_cse : STD_LOGIC;
  SIGNAL or_280_cse : STD_LOGIC;
  SIGNAL or_287_cse : STD_LOGIC;
  SIGNAL or_296_cse : STD_LOGIC;
  SIGNAL or_307_cse : STD_LOGIC;
  SIGNAL or_320_cse : STD_LOGIC;
  SIGNAL or_335_cse : STD_LOGIC;
  SIGNAL nand_281_cse : STD_LOGIC;
  SIGNAL or_377_cse : STD_LOGIC;
  SIGNAL or_382_cse : STD_LOGIC;
  SIGNAL or_386_cse : STD_LOGIC;
  SIGNAL or_391_cse : STD_LOGIC;
  SIGNAL or_397_cse : STD_LOGIC;
  SIGNAL nand_215_cse : STD_LOGIC;
  SIGNAL or_404_cse : STD_LOGIC;
  SIGNAL nand_212_cse : STD_LOGIC;
  SIGNAL or_413_cse : STD_LOGIC;
  SIGNAL nand_208_cse : STD_LOGIC;
  SIGNAL or_424_cse : STD_LOGIC;
  SIGNAL or_458_cse : STD_LOGIC;
  SIGNAL or_463_cse : STD_LOGIC;
  SIGNAL nand_198_cse : STD_LOGIC;
  SIGNAL or_468_cse : STD_LOGIC;
  SIGNAL or_475_cse : STD_LOGIC;
  SIGNAL nand_189_cse : STD_LOGIC;
  SIGNAL or_484_cse : STD_LOGIC;
  SIGNAL or_495_cse : STD_LOGIC;
  SIGNAL or_508_cse : STD_LOGIC;
  SIGNAL nand_203_cse : STD_LOGIC;
  SIGNAL or_523_cse : STD_LOGIC;
  SIGNAL nand_250_cse : STD_LOGIC;
  SIGNAL or_564_cse : STD_LOGIC;
  SIGNAL or_569_cse : STD_LOGIC;
  SIGNAL or_573_cse : STD_LOGIC;
  SIGNAL or_578_cse : STD_LOGIC;
  SIGNAL or_584_cse : STD_LOGIC;
  SIGNAL or_591_cse : STD_LOGIC;
  SIGNAL or_600_cse : STD_LOGIC;
  SIGNAL or_611_cse : STD_LOGIC;
  SIGNAL or_643_cse : STD_LOGIC;
  SIGNAL or_648_cse : STD_LOGIC;
  SIGNAL or_653_cse : STD_LOGIC;
  SIGNAL or_660_cse : STD_LOGIC;
  SIGNAL or_669_cse : STD_LOGIC;
  SIGNAL or_680_cse : STD_LOGIC;
  SIGNAL or_693_cse : STD_LOGIC;
  SIGNAL or_708_cse : STD_LOGIC;
  SIGNAL or_748_cse : STD_LOGIC;
  SIGNAL or_753_cse : STD_LOGIC;
  SIGNAL or_757_cse : STD_LOGIC;
  SIGNAL or_762_cse : STD_LOGIC;
  SIGNAL or_768_cse : STD_LOGIC;
  SIGNAL or_775_cse : STD_LOGIC;
  SIGNAL or_784_cse : STD_LOGIC;
  SIGNAL or_795_cse : STD_LOGIC;
  SIGNAL or_837_cse : STD_LOGIC;
  SIGNAL nand_84_cse : STD_LOGIC;
  SIGNAL or_842_cse : STD_LOGIC;
  SIGNAL or_847_cse : STD_LOGIC;
  SIGNAL nand_79_cse : STD_LOGIC;
  SIGNAL or_854_cse : STD_LOGIC;
  SIGNAL or_863_cse : STD_LOGIC;
  SIGNAL or_874_cse : STD_LOGIC;
  SIGNAL or_887_cse : STD_LOGIC;
  SIGNAL or_902_cse : STD_LOGIC;
  SIGNAL or_952_cse : STD_LOGIC;
  SIGNAL or_957_cse : STD_LOGIC;
  SIGNAL or_961_cse : STD_LOGIC;
  SIGNAL or_966_cse : STD_LOGIC;
  SIGNAL or_972_cse : STD_LOGIC;
  SIGNAL or_979_cse : STD_LOGIC;
  SIGNAL or_988_cse : STD_LOGIC;
  SIGNAL or_999_cse : STD_LOGIC;
  SIGNAL nand_57_cse : STD_LOGIC;
  SIGNAL or_1045_cse : STD_LOGIC;
  SIGNAL or_1050_cse : STD_LOGIC;
  SIGNAL or_1057_cse : STD_LOGIC;
  SIGNAL or_1066_cse : STD_LOGIC;
  SIGNAL nand_36_cse : STD_LOGIC;
  SIGNAL nand_29_cse : STD_LOGIC;
  SIGNAL nand_21_cse : STD_LOGIC;
  SIGNAL nand_222_cse : STD_LOGIC;
  SIGNAL nand_223_cse : STD_LOGIC;
  SIGNAL main_stage_0_12 : STD_LOGIC;
  SIGNAL m_buf_sva_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_11 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_12 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_asn_itm_11 : STD_LOGIC;
  SIGNAL mut_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12cyc_st_11_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_11_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL result_sva_duc_mx0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_and_26_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_28_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_30_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_32_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_34_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_36_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_38_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_40_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_42_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_44_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_46_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_48_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_50_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_52_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_54_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_56_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_58_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_60_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_62_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_64_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_66_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_68_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_70_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_72_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_74_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_76_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_78_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_80_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_82_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_84_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_86_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_88_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_90_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_92_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_94_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_96_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_98_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_100_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_102_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_104_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_106_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_108_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_110_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_112_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_114_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_116_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_118_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_120_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_122_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_124_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_126_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_128_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_130_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_132_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_134_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_136_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_138_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_140_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_142_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_144_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_146_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_148_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_150_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_152_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_154_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_156_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_158_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_160_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_162_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_164_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_166_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_168_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_170_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_172_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_174_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_176_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_178_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_180_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_182_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_184_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_186_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_188_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_190_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_192_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_194_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_196_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_198_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_200_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_202_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_204_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_206_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_208_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_210_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_212_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_214_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_216_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_218_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_220_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_222_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_224_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_226_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_228_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_230_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_232_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_234_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_236_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_238_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_240_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_242_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_244_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_246_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_248_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_250_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_252_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_254_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_256_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_258_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_260_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_262_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_264_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_266_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_268_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_270_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_272_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_274_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_276_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_278_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_280_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_282_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_284_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_and_286_cse : STD_LOGIC;

  SIGNAL qelse_acc_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mux_11_nl : STD_LOGIC;
  SIGNAL mux_10_nl : STD_LOGIC;
  SIGNAL mux_9_nl : STD_LOGIC;
  SIGNAL mux_8_nl : STD_LOGIC;
  SIGNAL mux_7_nl : STD_LOGIC;
  SIGNAL mux_6_nl : STD_LOGIC;
  SIGNAL mux_5_nl : STD_LOGIC;
  SIGNAL mux_4_nl : STD_LOGIC;
  SIGNAL mux_3_nl : STD_LOGIC;
  SIGNAL mux_2_nl : STD_LOGIC;
  SIGNAL mux_1_nl : STD_LOGIC;
  SIGNAL mux_nl : STD_LOGIC;
  SIGNAL and_273_nl : STD_LOGIC;
  SIGNAL and_275_nl : STD_LOGIC;
  SIGNAL and_277_nl : STD_LOGIC;
  SIGNAL and_279_nl : STD_LOGIC;
  SIGNAL and_281_nl : STD_LOGIC;
  SIGNAL and_282_nl : STD_LOGIC;
  SIGNAL and_283_nl : STD_LOGIC;
  SIGNAL and_284_nl : STD_LOGIC;
  SIGNAL and_286_nl : STD_LOGIC;
  SIGNAL and_287_nl : STD_LOGIC;
  SIGNAL and_288_nl : STD_LOGIC;
  SIGNAL and_289_nl : STD_LOGIC;
  SIGNAL and_290_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_xor_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_nl : STD_LOGIC;
  SIGNAL mux_12_nl : STD_LOGIC;
  SIGNAL nor_nl : STD_LOGIC;
  SIGNAL mux_13_nl : STD_LOGIC;
  SIGNAL nor_516_nl : STD_LOGIC;
  SIGNAL mux_14_nl : STD_LOGIC;
  SIGNAL nor_515_nl : STD_LOGIC;
  SIGNAL mux_15_nl : STD_LOGIC;
  SIGNAL nor_514_nl : STD_LOGIC;
  SIGNAL mux_16_nl : STD_LOGIC;
  SIGNAL nor_513_nl : STD_LOGIC;
  SIGNAL mux_17_nl : STD_LOGIC;
  SIGNAL nor_511_nl : STD_LOGIC;
  SIGNAL mux_18_nl : STD_LOGIC;
  SIGNAL nor_512_nl : STD_LOGIC;
  SIGNAL nor_508_nl : STD_LOGIC;
  SIGNAL mux_20_nl : STD_LOGIC;
  SIGNAL nor_509_nl : STD_LOGIC;
  SIGNAL mux_21_nl : STD_LOGIC;
  SIGNAL nor_510_nl : STD_LOGIC;
  SIGNAL nor_504_nl : STD_LOGIC;
  SIGNAL nor_505_nl : STD_LOGIC;
  SIGNAL mux_24_nl : STD_LOGIC;
  SIGNAL nor_506_nl : STD_LOGIC;
  SIGNAL mux_25_nl : STD_LOGIC;
  SIGNAL nor_507_nl : STD_LOGIC;
  SIGNAL nor_499_nl : STD_LOGIC;
  SIGNAL or_61_nl : STD_LOGIC;
  SIGNAL nor_500_nl : STD_LOGIC;
  SIGNAL nor_501_nl : STD_LOGIC;
  SIGNAL mux_29_nl : STD_LOGIC;
  SIGNAL nor_502_nl : STD_LOGIC;
  SIGNAL mux_30_nl : STD_LOGIC;
  SIGNAL nor_503_nl : STD_LOGIC;
  SIGNAL mux_31_nl : STD_LOGIC;
  SIGNAL nor_498_nl : STD_LOGIC;
  SIGNAL and_1168_nl : STD_LOGIC;
  SIGNAL mux_33_nl : STD_LOGIC;
  SIGNAL nor_497_nl : STD_LOGIC;
  SIGNAL and_1166_nl : STD_LOGIC;
  SIGNAL and_1167_nl : STD_LOGIC;
  SIGNAL mux_36_nl : STD_LOGIC;
  SIGNAL nor_496_nl : STD_LOGIC;
  SIGNAL and_1163_nl : STD_LOGIC;
  SIGNAL and_1164_nl : STD_LOGIC;
  SIGNAL and_1165_nl : STD_LOGIC;
  SIGNAL mux_40_nl : STD_LOGIC;
  SIGNAL nor_495_nl : STD_LOGIC;
  SIGNAL and_1159_nl : STD_LOGIC;
  SIGNAL and_1160_nl : STD_LOGIC;
  SIGNAL and_1161_nl : STD_LOGIC;
  SIGNAL and_1162_nl : STD_LOGIC;
  SIGNAL mux_45_nl : STD_LOGIC;
  SIGNAL nor_494_nl : STD_LOGIC;
  SIGNAL nor_492_nl : STD_LOGIC;
  SIGNAL and_1155_nl : STD_LOGIC;
  SIGNAL and_1156_nl : STD_LOGIC;
  SIGNAL and_1157_nl : STD_LOGIC;
  SIGNAL and_1158_nl : STD_LOGIC;
  SIGNAL mux_51_nl : STD_LOGIC;
  SIGNAL nor_493_nl : STD_LOGIC;
  SIGNAL nor_489_nl : STD_LOGIC;
  SIGNAL nor_490_nl : STD_LOGIC;
  SIGNAL and_1151_nl : STD_LOGIC;
  SIGNAL and_1152_nl : STD_LOGIC;
  SIGNAL and_1153_nl : STD_LOGIC;
  SIGNAL and_1154_nl : STD_LOGIC;
  SIGNAL mux_58_nl : STD_LOGIC;
  SIGNAL nor_491_nl : STD_LOGIC;
  SIGNAL nor_485_nl : STD_LOGIC;
  SIGNAL nor_486_nl : STD_LOGIC;
  SIGNAL nor_487_nl : STD_LOGIC;
  SIGNAL and_1147_nl : STD_LOGIC;
  SIGNAL and_1148_nl : STD_LOGIC;
  SIGNAL and_1149_nl : STD_LOGIC;
  SIGNAL and_1150_nl : STD_LOGIC;
  SIGNAL mux_66_nl : STD_LOGIC;
  SIGNAL nor_488_nl : STD_LOGIC;
  SIGNAL nor_480_nl : STD_LOGIC;
  SIGNAL or_165_nl : STD_LOGIC;
  SIGNAL nor_481_nl : STD_LOGIC;
  SIGNAL nor_482_nl : STD_LOGIC;
  SIGNAL nor_483_nl : STD_LOGIC;
  SIGNAL and_1143_nl : STD_LOGIC;
  SIGNAL and_1144_nl : STD_LOGIC;
  SIGNAL and_1145_nl : STD_LOGIC;
  SIGNAL and_1146_nl : STD_LOGIC;
  SIGNAL mux_75_nl : STD_LOGIC;
  SIGNAL nor_484_nl : STD_LOGIC;
  SIGNAL nor_479_nl : STD_LOGIC;
  SIGNAL or_175_nl : STD_LOGIC;
  SIGNAL mux_77_nl : STD_LOGIC;
  SIGNAL nor_478_nl : STD_LOGIC;
  SIGNAL mux_78_nl : STD_LOGIC;
  SIGNAL nor_477_nl : STD_LOGIC;
  SIGNAL mux_79_nl : STD_LOGIC;
  SIGNAL nor_476_nl : STD_LOGIC;
  SIGNAL mux_80_nl : STD_LOGIC;
  SIGNAL nor_475_nl : STD_LOGIC;
  SIGNAL mux_81_nl : STD_LOGIC;
  SIGNAL nor_474_nl : STD_LOGIC;
  SIGNAL mux_82_nl : STD_LOGIC;
  SIGNAL nor_472_nl : STD_LOGIC;
  SIGNAL mux_83_nl : STD_LOGIC;
  SIGNAL nor_473_nl : STD_LOGIC;
  SIGNAL nor_469_nl : STD_LOGIC;
  SIGNAL mux_85_nl : STD_LOGIC;
  SIGNAL nor_470_nl : STD_LOGIC;
  SIGNAL mux_86_nl : STD_LOGIC;
  SIGNAL nor_471_nl : STD_LOGIC;
  SIGNAL nor_465_nl : STD_LOGIC;
  SIGNAL nor_466_nl : STD_LOGIC;
  SIGNAL mux_89_nl : STD_LOGIC;
  SIGNAL nor_467_nl : STD_LOGIC;
  SIGNAL mux_90_nl : STD_LOGIC;
  SIGNAL nor_468_nl : STD_LOGIC;
  SIGNAL nor_460_nl : STD_LOGIC;
  SIGNAL or_250_nl : STD_LOGIC;
  SIGNAL nor_461_nl : STD_LOGIC;
  SIGNAL nor_462_nl : STD_LOGIC;
  SIGNAL mux_94_nl : STD_LOGIC;
  SIGNAL nor_463_nl : STD_LOGIC;
  SIGNAL mux_95_nl : STD_LOGIC;
  SIGNAL nor_464_nl : STD_LOGIC;
  SIGNAL mux_96_nl : STD_LOGIC;
  SIGNAL nor_459_nl : STD_LOGIC;
  SIGNAL and_1142_nl : STD_LOGIC;
  SIGNAL mux_98_nl : STD_LOGIC;
  SIGNAL nor_458_nl : STD_LOGIC;
  SIGNAL and_1140_nl : STD_LOGIC;
  SIGNAL and_1141_nl : STD_LOGIC;
  SIGNAL mux_101_nl : STD_LOGIC;
  SIGNAL nor_457_nl : STD_LOGIC;
  SIGNAL and_1137_nl : STD_LOGIC;
  SIGNAL and_1138_nl : STD_LOGIC;
  SIGNAL and_1139_nl : STD_LOGIC;
  SIGNAL mux_105_nl : STD_LOGIC;
  SIGNAL nor_456_nl : STD_LOGIC;
  SIGNAL and_1133_nl : STD_LOGIC;
  SIGNAL and_1134_nl : STD_LOGIC;
  SIGNAL and_1135_nl : STD_LOGIC;
  SIGNAL and_1136_nl : STD_LOGIC;
  SIGNAL mux_110_nl : STD_LOGIC;
  SIGNAL nor_455_nl : STD_LOGIC;
  SIGNAL nor_453_nl : STD_LOGIC;
  SIGNAL and_1129_nl : STD_LOGIC;
  SIGNAL and_1130_nl : STD_LOGIC;
  SIGNAL and_1131_nl : STD_LOGIC;
  SIGNAL and_1132_nl : STD_LOGIC;
  SIGNAL mux_116_nl : STD_LOGIC;
  SIGNAL nor_454_nl : STD_LOGIC;
  SIGNAL nor_450_nl : STD_LOGIC;
  SIGNAL nor_451_nl : STD_LOGIC;
  SIGNAL and_1125_nl : STD_LOGIC;
  SIGNAL and_1126_nl : STD_LOGIC;
  SIGNAL and_1127_nl : STD_LOGIC;
  SIGNAL and_1128_nl : STD_LOGIC;
  SIGNAL mux_123_nl : STD_LOGIC;
  SIGNAL nor_452_nl : STD_LOGIC;
  SIGNAL nor_446_nl : STD_LOGIC;
  SIGNAL nor_447_nl : STD_LOGIC;
  SIGNAL nor_448_nl : STD_LOGIC;
  SIGNAL and_1121_nl : STD_LOGIC;
  SIGNAL and_1122_nl : STD_LOGIC;
  SIGNAL and_1123_nl : STD_LOGIC;
  SIGNAL and_1124_nl : STD_LOGIC;
  SIGNAL mux_131_nl : STD_LOGIC;
  SIGNAL nor_449_nl : STD_LOGIC;
  SIGNAL nor_441_nl : STD_LOGIC;
  SIGNAL or_352_nl : STD_LOGIC;
  SIGNAL nor_442_nl : STD_LOGIC;
  SIGNAL nor_443_nl : STD_LOGIC;
  SIGNAL nor_444_nl : STD_LOGIC;
  SIGNAL and_1117_nl : STD_LOGIC;
  SIGNAL and_1118_nl : STD_LOGIC;
  SIGNAL and_1119_nl : STD_LOGIC;
  SIGNAL and_1120_nl : STD_LOGIC;
  SIGNAL mux_140_nl : STD_LOGIC;
  SIGNAL nor_445_nl : STD_LOGIC;
  SIGNAL and_1116_nl : STD_LOGIC;
  SIGNAL or_362_nl : STD_LOGIC;
  SIGNAL mux_142_nl : STD_LOGIC;
  SIGNAL and_1172_nl : STD_LOGIC;
  SIGNAL mux_143_nl : STD_LOGIC;
  SIGNAL and_1114_nl : STD_LOGIC;
  SIGNAL mux_144_nl : STD_LOGIC;
  SIGNAL and_1113_nl : STD_LOGIC;
  SIGNAL mux_145_nl : STD_LOGIC;
  SIGNAL and_1112_nl : STD_LOGIC;
  SIGNAL mux_146_nl : STD_LOGIC;
  SIGNAL and_1111_nl : STD_LOGIC;
  SIGNAL mux_147_nl : STD_LOGIC;
  SIGNAL and_1109_nl : STD_LOGIC;
  SIGNAL mux_148_nl : STD_LOGIC;
  SIGNAL and_1110_nl : STD_LOGIC;
  SIGNAL and_1106_nl : STD_LOGIC;
  SIGNAL mux_150_nl : STD_LOGIC;
  SIGNAL and_1107_nl : STD_LOGIC;
  SIGNAL mux_151_nl : STD_LOGIC;
  SIGNAL and_1108_nl : STD_LOGIC;
  SIGNAL and_1102_nl : STD_LOGIC;
  SIGNAL and_1103_nl : STD_LOGIC;
  SIGNAL mux_154_nl : STD_LOGIC;
  SIGNAL and_1104_nl : STD_LOGIC;
  SIGNAL mux_155_nl : STD_LOGIC;
  SIGNAL and_1105_nl : STD_LOGIC;
  SIGNAL and_1097_nl : STD_LOGIC;
  SIGNAL or_437_nl : STD_LOGIC;
  SIGNAL and_1098_nl : STD_LOGIC;
  SIGNAL and_1099_nl : STD_LOGIC;
  SIGNAL mux_159_nl : STD_LOGIC;
  SIGNAL and_1100_nl : STD_LOGIC;
  SIGNAL mux_160_nl : STD_LOGIC;
  SIGNAL and_1101_nl : STD_LOGIC;
  SIGNAL mux_161_nl : STD_LOGIC;
  SIGNAL and_1171_nl : STD_LOGIC;
  SIGNAL and_1094_nl : STD_LOGIC;
  SIGNAL mux_163_nl : STD_LOGIC;
  SIGNAL and_1095_nl : STD_LOGIC;
  SIGNAL and_1091_nl : STD_LOGIC;
  SIGNAL and_1092_nl : STD_LOGIC;
  SIGNAL mux_166_nl : STD_LOGIC;
  SIGNAL and_1093_nl : STD_LOGIC;
  SIGNAL and_1087_nl : STD_LOGIC;
  SIGNAL and_1088_nl : STD_LOGIC;
  SIGNAL and_1089_nl : STD_LOGIC;
  SIGNAL mux_170_nl : STD_LOGIC;
  SIGNAL and_1090_nl : STD_LOGIC;
  SIGNAL and_1082_nl : STD_LOGIC;
  SIGNAL and_1083_nl : STD_LOGIC;
  SIGNAL and_1084_nl : STD_LOGIC;
  SIGNAL and_1085_nl : STD_LOGIC;
  SIGNAL mux_175_nl : STD_LOGIC;
  SIGNAL and_1086_nl : STD_LOGIC;
  SIGNAL and_1076_nl : STD_LOGIC;
  SIGNAL and_1077_nl : STD_LOGIC;
  SIGNAL and_1078_nl : STD_LOGIC;
  SIGNAL and_1079_nl : STD_LOGIC;
  SIGNAL and_1080_nl : STD_LOGIC;
  SIGNAL mux_181_nl : STD_LOGIC;
  SIGNAL and_1081_nl : STD_LOGIC;
  SIGNAL and_1069_nl : STD_LOGIC;
  SIGNAL and_1070_nl : STD_LOGIC;
  SIGNAL and_1071_nl : STD_LOGIC;
  SIGNAL and_1072_nl : STD_LOGIC;
  SIGNAL and_1073_nl : STD_LOGIC;
  SIGNAL and_1074_nl : STD_LOGIC;
  SIGNAL mux_188_nl : STD_LOGIC;
  SIGNAL and_1075_nl : STD_LOGIC;
  SIGNAL and_1061_nl : STD_LOGIC;
  SIGNAL and_1062_nl : STD_LOGIC;
  SIGNAL and_1063_nl : STD_LOGIC;
  SIGNAL and_1064_nl : STD_LOGIC;
  SIGNAL and_1065_nl : STD_LOGIC;
  SIGNAL and_1066_nl : STD_LOGIC;
  SIGNAL and_1067_nl : STD_LOGIC;
  SIGNAL mux_196_nl : STD_LOGIC;
  SIGNAL and_1068_nl : STD_LOGIC;
  SIGNAL and_1052_nl : STD_LOGIC;
  SIGNAL or_540_nl : STD_LOGIC;
  SIGNAL and_1053_nl : STD_LOGIC;
  SIGNAL and_1054_nl : STD_LOGIC;
  SIGNAL and_1055_nl : STD_LOGIC;
  SIGNAL and_1056_nl : STD_LOGIC;
  SIGNAL and_1057_nl : STD_LOGIC;
  SIGNAL and_1058_nl : STD_LOGIC;
  SIGNAL and_1059_nl : STD_LOGIC;
  SIGNAL mux_205_nl : STD_LOGIC;
  SIGNAL and_1060_nl : STD_LOGIC;
  SIGNAL nor_438_nl : STD_LOGIC;
  SIGNAL or_550_nl : STD_LOGIC;
  SIGNAL mux_207_nl : STD_LOGIC;
  SIGNAL and_1170_nl : STD_LOGIC;
  SIGNAL mux_208_nl : STD_LOGIC;
  SIGNAL and_1050_nl : STD_LOGIC;
  SIGNAL mux_209_nl : STD_LOGIC;
  SIGNAL and_1049_nl : STD_LOGIC;
  SIGNAL mux_210_nl : STD_LOGIC;
  SIGNAL and_1048_nl : STD_LOGIC;
  SIGNAL mux_211_nl : STD_LOGIC;
  SIGNAL and_1047_nl : STD_LOGIC;
  SIGNAL mux_212_nl : STD_LOGIC;
  SIGNAL and_1045_nl : STD_LOGIC;
  SIGNAL mux_213_nl : STD_LOGIC;
  SIGNAL and_1046_nl : STD_LOGIC;
  SIGNAL and_1042_nl : STD_LOGIC;
  SIGNAL mux_215_nl : STD_LOGIC;
  SIGNAL and_1043_nl : STD_LOGIC;
  SIGNAL mux_216_nl : STD_LOGIC;
  SIGNAL and_1044_nl : STD_LOGIC;
  SIGNAL and_1038_nl : STD_LOGIC;
  SIGNAL and_1039_nl : STD_LOGIC;
  SIGNAL mux_219_nl : STD_LOGIC;
  SIGNAL and_1040_nl : STD_LOGIC;
  SIGNAL mux_220_nl : STD_LOGIC;
  SIGNAL and_1041_nl : STD_LOGIC;
  SIGNAL and_1033_nl : STD_LOGIC;
  SIGNAL or_624_nl : STD_LOGIC;
  SIGNAL and_1034_nl : STD_LOGIC;
  SIGNAL and_1035_nl : STD_LOGIC;
  SIGNAL mux_224_nl : STD_LOGIC;
  SIGNAL and_1036_nl : STD_LOGIC;
  SIGNAL mux_225_nl : STD_LOGIC;
  SIGNAL and_1037_nl : STD_LOGIC;
  SIGNAL mux_226_nl : STD_LOGIC;
  SIGNAL and_1169_nl : STD_LOGIC;
  SIGNAL and_1030_nl : STD_LOGIC;
  SIGNAL mux_228_nl : STD_LOGIC;
  SIGNAL and_1031_nl : STD_LOGIC;
  SIGNAL and_1027_nl : STD_LOGIC;
  SIGNAL and_1028_nl : STD_LOGIC;
  SIGNAL mux_231_nl : STD_LOGIC;
  SIGNAL and_1029_nl : STD_LOGIC;
  SIGNAL and_1023_nl : STD_LOGIC;
  SIGNAL and_1024_nl : STD_LOGIC;
  SIGNAL and_1025_nl : STD_LOGIC;
  SIGNAL mux_235_nl : STD_LOGIC;
  SIGNAL and_1026_nl : STD_LOGIC;
  SIGNAL and_1018_nl : STD_LOGIC;
  SIGNAL and_1019_nl : STD_LOGIC;
  SIGNAL and_1020_nl : STD_LOGIC;
  SIGNAL and_1021_nl : STD_LOGIC;
  SIGNAL mux_240_nl : STD_LOGIC;
  SIGNAL and_1022_nl : STD_LOGIC;
  SIGNAL and_1012_nl : STD_LOGIC;
  SIGNAL and_1013_nl : STD_LOGIC;
  SIGNAL and_1014_nl : STD_LOGIC;
  SIGNAL and_1015_nl : STD_LOGIC;
  SIGNAL and_1016_nl : STD_LOGIC;
  SIGNAL mux_246_nl : STD_LOGIC;
  SIGNAL and_1017_nl : STD_LOGIC;
  SIGNAL and_1005_nl : STD_LOGIC;
  SIGNAL and_1006_nl : STD_LOGIC;
  SIGNAL and_1007_nl : STD_LOGIC;
  SIGNAL and_1008_nl : STD_LOGIC;
  SIGNAL and_1009_nl : STD_LOGIC;
  SIGNAL and_1010_nl : STD_LOGIC;
  SIGNAL mux_253_nl : STD_LOGIC;
  SIGNAL and_1011_nl : STD_LOGIC;
  SIGNAL and_997_nl : STD_LOGIC;
  SIGNAL and_998_nl : STD_LOGIC;
  SIGNAL and_999_nl : STD_LOGIC;
  SIGNAL and_1000_nl : STD_LOGIC;
  SIGNAL and_1001_nl : STD_LOGIC;
  SIGNAL and_1002_nl : STD_LOGIC;
  SIGNAL and_1003_nl : STD_LOGIC;
  SIGNAL mux_261_nl : STD_LOGIC;
  SIGNAL and_1004_nl : STD_LOGIC;
  SIGNAL and_988_nl : STD_LOGIC;
  SIGNAL or_725_nl : STD_LOGIC;
  SIGNAL and_989_nl : STD_LOGIC;
  SIGNAL and_990_nl : STD_LOGIC;
  SIGNAL and_991_nl : STD_LOGIC;
  SIGNAL and_992_nl : STD_LOGIC;
  SIGNAL and_993_nl : STD_LOGIC;
  SIGNAL and_994_nl : STD_LOGIC;
  SIGNAL and_995_nl : STD_LOGIC;
  SIGNAL mux_270_nl : STD_LOGIC;
  SIGNAL and_996_nl : STD_LOGIC;
  SIGNAL and_987_nl : STD_LOGIC;
  SIGNAL or_735_nl : STD_LOGIC;
  SIGNAL mux_272_nl : STD_LOGIC;
  SIGNAL nor_435_nl : STD_LOGIC;
  SIGNAL mux_273_nl : STD_LOGIC;
  SIGNAL nor_434_nl : STD_LOGIC;
  SIGNAL mux_274_nl : STD_LOGIC;
  SIGNAL nor_433_nl : STD_LOGIC;
  SIGNAL mux_275_nl : STD_LOGIC;
  SIGNAL nor_432_nl : STD_LOGIC;
  SIGNAL mux_276_nl : STD_LOGIC;
  SIGNAL nor_431_nl : STD_LOGIC;
  SIGNAL mux_277_nl : STD_LOGIC;
  SIGNAL nor_429_nl : STD_LOGIC;
  SIGNAL mux_278_nl : STD_LOGIC;
  SIGNAL nor_430_nl : STD_LOGIC;
  SIGNAL nor_426_nl : STD_LOGIC;
  SIGNAL mux_280_nl : STD_LOGIC;
  SIGNAL nor_427_nl : STD_LOGIC;
  SIGNAL mux_281_nl : STD_LOGIC;
  SIGNAL nor_428_nl : STD_LOGIC;
  SIGNAL nor_422_nl : STD_LOGIC;
  SIGNAL nor_423_nl : STD_LOGIC;
  SIGNAL mux_284_nl : STD_LOGIC;
  SIGNAL nor_424_nl : STD_LOGIC;
  SIGNAL mux_285_nl : STD_LOGIC;
  SIGNAL nor_425_nl : STD_LOGIC;
  SIGNAL nor_417_nl : STD_LOGIC;
  SIGNAL or_808_nl : STD_LOGIC;
  SIGNAL nor_418_nl : STD_LOGIC;
  SIGNAL nor_419_nl : STD_LOGIC;
  SIGNAL mux_289_nl : STD_LOGIC;
  SIGNAL nor_420_nl : STD_LOGIC;
  SIGNAL mux_290_nl : STD_LOGIC;
  SIGNAL nor_421_nl : STD_LOGIC;
  SIGNAL nor_408_nl : STD_LOGIC;
  SIGNAL or_823_nl : STD_LOGIC;
  SIGNAL nor_409_nl : STD_LOGIC;
  SIGNAL or_822_nl : STD_LOGIC;
  SIGNAL nor_410_nl : STD_LOGIC;
  SIGNAL or_821_nl : STD_LOGIC;
  SIGNAL nor_411_nl : STD_LOGIC;
  SIGNAL or_820_nl : STD_LOGIC;
  SIGNAL nor_412_nl : STD_LOGIC;
  SIGNAL or_819_nl : STD_LOGIC;
  SIGNAL nor_413_nl : STD_LOGIC;
  SIGNAL or_818_nl : STD_LOGIC;
  SIGNAL nor_414_nl : STD_LOGIC;
  SIGNAL or_817_nl : STD_LOGIC;
  SIGNAL nor_415_nl : STD_LOGIC;
  SIGNAL or_816_nl : STD_LOGIC;
  SIGNAL mux_299_nl : STD_LOGIC;
  SIGNAL nor_416_nl : STD_LOGIC;
  SIGNAL or_815_nl : STD_LOGIC;
  SIGNAL mux_300_nl : STD_LOGIC;
  SIGNAL nor_407_nl : STD_LOGIC;
  SIGNAL and_986_nl : STD_LOGIC;
  SIGNAL mux_302_nl : STD_LOGIC;
  SIGNAL nor_406_nl : STD_LOGIC;
  SIGNAL and_984_nl : STD_LOGIC;
  SIGNAL and_985_nl : STD_LOGIC;
  SIGNAL mux_305_nl : STD_LOGIC;
  SIGNAL nor_405_nl : STD_LOGIC;
  SIGNAL and_981_nl : STD_LOGIC;
  SIGNAL and_982_nl : STD_LOGIC;
  SIGNAL and_983_nl : STD_LOGIC;
  SIGNAL mux_309_nl : STD_LOGIC;
  SIGNAL nor_404_nl : STD_LOGIC;
  SIGNAL and_977_nl : STD_LOGIC;
  SIGNAL and_978_nl : STD_LOGIC;
  SIGNAL and_979_nl : STD_LOGIC;
  SIGNAL and_980_nl : STD_LOGIC;
  SIGNAL mux_314_nl : STD_LOGIC;
  SIGNAL nor_403_nl : STD_LOGIC;
  SIGNAL nor_401_nl : STD_LOGIC;
  SIGNAL and_973_nl : STD_LOGIC;
  SIGNAL and_974_nl : STD_LOGIC;
  SIGNAL and_975_nl : STD_LOGIC;
  SIGNAL and_976_nl : STD_LOGIC;
  SIGNAL mux_320_nl : STD_LOGIC;
  SIGNAL nor_402_nl : STD_LOGIC;
  SIGNAL nor_398_nl : STD_LOGIC;
  SIGNAL nor_399_nl : STD_LOGIC;
  SIGNAL and_969_nl : STD_LOGIC;
  SIGNAL and_970_nl : STD_LOGIC;
  SIGNAL and_971_nl : STD_LOGIC;
  SIGNAL and_972_nl : STD_LOGIC;
  SIGNAL mux_327_nl : STD_LOGIC;
  SIGNAL nor_400_nl : STD_LOGIC;
  SIGNAL nor_394_nl : STD_LOGIC;
  SIGNAL nor_395_nl : STD_LOGIC;
  SIGNAL nor_396_nl : STD_LOGIC;
  SIGNAL and_965_nl : STD_LOGIC;
  SIGNAL and_966_nl : STD_LOGIC;
  SIGNAL and_967_nl : STD_LOGIC;
  SIGNAL and_968_nl : STD_LOGIC;
  SIGNAL mux_335_nl : STD_LOGIC;
  SIGNAL nor_397_nl : STD_LOGIC;
  SIGNAL nor_389_nl : STD_LOGIC;
  SIGNAL or_919_nl : STD_LOGIC;
  SIGNAL nor_390_nl : STD_LOGIC;
  SIGNAL nor_391_nl : STD_LOGIC;
  SIGNAL nor_392_nl : STD_LOGIC;
  SIGNAL and_961_nl : STD_LOGIC;
  SIGNAL and_962_nl : STD_LOGIC;
  SIGNAL and_963_nl : STD_LOGIC;
  SIGNAL and_964_nl : STD_LOGIC;
  SIGNAL mux_344_nl : STD_LOGIC;
  SIGNAL nor_393_nl : STD_LOGIC;
  SIGNAL nor_379_nl : STD_LOGIC;
  SIGNAL or_938_nl : STD_LOGIC;
  SIGNAL nor_380_nl : STD_LOGIC;
  SIGNAL or_937_nl : STD_LOGIC;
  SIGNAL nor_381_nl : STD_LOGIC;
  SIGNAL or_936_nl : STD_LOGIC;
  SIGNAL nor_382_nl : STD_LOGIC;
  SIGNAL or_935_nl : STD_LOGIC;
  SIGNAL nor_383_nl : STD_LOGIC;
  SIGNAL or_934_nl : STD_LOGIC;
  SIGNAL nor_384_nl : STD_LOGIC;
  SIGNAL or_933_nl : STD_LOGIC;
  SIGNAL nor_385_nl : STD_LOGIC;
  SIGNAL or_932_nl : STD_LOGIC;
  SIGNAL nor_386_nl : STD_LOGIC;
  SIGNAL or_931_nl : STD_LOGIC;
  SIGNAL nor_387_nl : STD_LOGIC;
  SIGNAL or_930_nl : STD_LOGIC;
  SIGNAL nor_388_nl : STD_LOGIC;
  SIGNAL or_929_nl : STD_LOGIC;
  SIGNAL mux_355_nl : STD_LOGIC;
  SIGNAL nor_378_nl : STD_LOGIC;
  SIGNAL mux_356_nl : STD_LOGIC;
  SIGNAL nor_377_nl : STD_LOGIC;
  SIGNAL mux_357_nl : STD_LOGIC;
  SIGNAL nor_376_nl : STD_LOGIC;
  SIGNAL mux_358_nl : STD_LOGIC;
  SIGNAL nor_375_nl : STD_LOGIC;
  SIGNAL mux_359_nl : STD_LOGIC;
  SIGNAL nor_374_nl : STD_LOGIC;
  SIGNAL mux_360_nl : STD_LOGIC;
  SIGNAL nor_372_nl : STD_LOGIC;
  SIGNAL mux_361_nl : STD_LOGIC;
  SIGNAL nor_373_nl : STD_LOGIC;
  SIGNAL nor_369_nl : STD_LOGIC;
  SIGNAL mux_363_nl : STD_LOGIC;
  SIGNAL nor_370_nl : STD_LOGIC;
  SIGNAL mux_364_nl : STD_LOGIC;
  SIGNAL nor_371_nl : STD_LOGIC;
  SIGNAL nor_365_nl : STD_LOGIC;
  SIGNAL nor_366_nl : STD_LOGIC;
  SIGNAL mux_367_nl : STD_LOGIC;
  SIGNAL nor_367_nl : STD_LOGIC;
  SIGNAL mux_368_nl : STD_LOGIC;
  SIGNAL nor_368_nl : STD_LOGIC;
  SIGNAL nor_360_nl : STD_LOGIC;
  SIGNAL or_1012_nl : STD_LOGIC;
  SIGNAL nor_361_nl : STD_LOGIC;
  SIGNAL nor_362_nl : STD_LOGIC;
  SIGNAL mux_372_nl : STD_LOGIC;
  SIGNAL nor_363_nl : STD_LOGIC;
  SIGNAL mux_373_nl : STD_LOGIC;
  SIGNAL nor_364_nl : STD_LOGIC;
  SIGNAL nor_351_nl : STD_LOGIC;
  SIGNAL or_1027_nl : STD_LOGIC;
  SIGNAL nor_352_nl : STD_LOGIC;
  SIGNAL or_1026_nl : STD_LOGIC;
  SIGNAL nor_353_nl : STD_LOGIC;
  SIGNAL or_1025_nl : STD_LOGIC;
  SIGNAL nor_354_nl : STD_LOGIC;
  SIGNAL or_1024_nl : STD_LOGIC;
  SIGNAL nor_355_nl : STD_LOGIC;
  SIGNAL or_1023_nl : STD_LOGIC;
  SIGNAL nor_356_nl : STD_LOGIC;
  SIGNAL or_1022_nl : STD_LOGIC;
  SIGNAL nor_357_nl : STD_LOGIC;
  SIGNAL or_1021_nl : STD_LOGIC;
  SIGNAL nor_358_nl : STD_LOGIC;
  SIGNAL or_1020_nl : STD_LOGIC;
  SIGNAL mux_382_nl : STD_LOGIC;
  SIGNAL nor_359_nl : STD_LOGIC;
  SIGNAL or_1019_nl : STD_LOGIC;
  SIGNAL mux_383_nl : STD_LOGIC;
  SIGNAL nor_350_nl : STD_LOGIC;
  SIGNAL and_960_nl : STD_LOGIC;
  SIGNAL mux_385_nl : STD_LOGIC;
  SIGNAL nor_349_nl : STD_LOGIC;
  SIGNAL and_958_nl : STD_LOGIC;
  SIGNAL and_959_nl : STD_LOGIC;
  SIGNAL mux_388_nl : STD_LOGIC;
  SIGNAL nor_348_nl : STD_LOGIC;
  SIGNAL and_955_nl : STD_LOGIC;
  SIGNAL and_956_nl : STD_LOGIC;
  SIGNAL and_957_nl : STD_LOGIC;
  SIGNAL mux_392_nl : STD_LOGIC;
  SIGNAL nor_347_nl : STD_LOGIC;
  SIGNAL and_951_nl : STD_LOGIC;
  SIGNAL and_952_nl : STD_LOGIC;
  SIGNAL and_953_nl : STD_LOGIC;
  SIGNAL and_954_nl : STD_LOGIC;
  SIGNAL mux_397_nl : STD_LOGIC;
  SIGNAL nor_346_nl : STD_LOGIC;
  SIGNAL nor_344_nl : STD_LOGIC;
  SIGNAL and_947_nl : STD_LOGIC;
  SIGNAL and_948_nl : STD_LOGIC;
  SIGNAL and_949_nl : STD_LOGIC;
  SIGNAL and_950_nl : STD_LOGIC;
  SIGNAL mux_403_nl : STD_LOGIC;
  SIGNAL nor_345_nl : STD_LOGIC;
  SIGNAL nor_341_nl : STD_LOGIC;
  SIGNAL nor_342_nl : STD_LOGIC;
  SIGNAL and_943_nl : STD_LOGIC;
  SIGNAL and_944_nl : STD_LOGIC;
  SIGNAL and_945_nl : STD_LOGIC;
  SIGNAL and_946_nl : STD_LOGIC;
  SIGNAL mux_410_nl : STD_LOGIC;
  SIGNAL nor_343_nl : STD_LOGIC;
  SIGNAL nor_337_nl : STD_LOGIC;
  SIGNAL nor_338_nl : STD_LOGIC;
  SIGNAL nor_339_nl : STD_LOGIC;
  SIGNAL and_939_nl : STD_LOGIC;
  SIGNAL and_940_nl : STD_LOGIC;
  SIGNAL and_941_nl : STD_LOGIC;
  SIGNAL and_942_nl : STD_LOGIC;
  SIGNAL mux_418_nl : STD_LOGIC;
  SIGNAL nor_340_nl : STD_LOGIC;
  SIGNAL nor_332_nl : STD_LOGIC;
  SIGNAL nand_12_nl : STD_LOGIC;
  SIGNAL nor_333_nl : STD_LOGIC;
  SIGNAL nor_334_nl : STD_LOGIC;
  SIGNAL nor_335_nl : STD_LOGIC;
  SIGNAL and_935_nl : STD_LOGIC;
  SIGNAL and_936_nl : STD_LOGIC;
  SIGNAL and_937_nl : STD_LOGIC;
  SIGNAL and_938_nl : STD_LOGIC;
  SIGNAL mux_427_nl : STD_LOGIC;
  SIGNAL nor_336_nl : STD_LOGIC;
  SIGNAL nor_323_nl : STD_LOGIC;
  SIGNAL nand_1_nl : STD_LOGIC;
  SIGNAL nor_324_nl : STD_LOGIC;
  SIGNAL nand_2_nl : STD_LOGIC;
  SIGNAL nor_325_nl : STD_LOGIC;
  SIGNAL nand_3_nl : STD_LOGIC;
  SIGNAL nor_326_nl : STD_LOGIC;
  SIGNAL nand_4_nl : STD_LOGIC;
  SIGNAL nor_327_nl : STD_LOGIC;
  SIGNAL nand_5_nl : STD_LOGIC;
  SIGNAL nor_328_nl : STD_LOGIC;
  SIGNAL nand_6_nl : STD_LOGIC;
  SIGNAL nor_329_nl : STD_LOGIC;
  SIGNAL nand_7_nl : STD_LOGIC;
  SIGNAL nor_330_nl : STD_LOGIC;
  SIGNAL nand_8_nl : STD_LOGIC;
  SIGNAL nor_331_nl : STD_LOGIC;
  SIGNAL nand_9_nl : STD_LOGIC;
  SIGNAL and_934_nl : STD_LOGIC;
  SIGNAL nand_11_nl : STD_LOGIC;
  SIGNAL base_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL m_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL return_rsci_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL return_rsci_z : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL ccs_ccore_start_rsci_dat : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL ccs_ccore_start_rsci_idat_1 : STD_LOGIC_VECTOR (0 DOWNTO 0);

  SIGNAL rem_12_cmp_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_12_cmp_1_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_1_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_1_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_12_cmp_2_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_2_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_2_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_12_cmp_3_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_3_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_3_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_12_cmp_4_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_4_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_4_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_12_cmp_5_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_5_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_5_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_12_cmp_6_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_6_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_6_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_12_cmp_7_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_7_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_7_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_12_cmp_8_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_8_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_8_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_12_cmp_9_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_9_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_9_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_12_cmp_10_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_10_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_10_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_12_cmp_11_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_11_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_12_cmp_11_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_v_64_11_2(input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(10 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_13_2(input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(12 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_64_2_2(input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  base_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 1,
      width => 64
      )
    PORT MAP(
      dat => base_rsci_dat,
      idat => base_rsci_idat_1
    );
  base_rsci_dat <= base_rsc_dat;
  base_rsci_idat <= base_rsci_idat_1;

  m_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 2,
      width => 64
      )
    PORT MAP(
      dat => m_rsci_dat,
      idat => m_rsci_idat_1
    );
  m_rsci_dat <= m_rsc_dat;
  m_rsci_idat <= m_rsci_idat_1;

  return_rsci : work.mgc_out_dreg_pkg_v2.mgc_out_dreg_v2
    GENERIC MAP(
      rscid => 3,
      width => 64
      )
    PORT MAP(
      d => return_rsci_d_1,
      z => return_rsci_z
    );
  return_rsci_d_1 <= return_rsci_d;
  return_rsc_z <= return_rsci_z;

  ccs_ccore_start_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 8,
      width => 1
      )
    PORT MAP(
      dat => ccs_ccore_start_rsci_dat,
      idat => ccs_ccore_start_rsci_idat_1
    );
  ccs_ccore_start_rsci_dat(0) <= ccs_ccore_start_rsc_dat;
  ccs_ccore_start_rsci_idat <= ccs_ccore_start_rsci_idat_1(0);

  rem_12_cmp : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_12_cmp_a,
      b => rem_12_cmp_b,
      z => rem_12_cmp_z_1
    );
  rem_12_cmp_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_12_cmp_a_63_0),65));
  rem_12_cmp_b <= '0' & rem_12_cmp_b_63_0;
  rem_12_cmp_z <= rem_12_cmp_z_1;

  rem_12_cmp_1 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_12_cmp_1_a,
      b => rem_12_cmp_1_b,
      z => rem_12_cmp_1_z_1
    );
  rem_12_cmp_1_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_12_cmp_1_a_63_0),65));
  rem_12_cmp_1_b <= '0' & rem_12_cmp_1_b_63_0;
  rem_12_cmp_1_z <= rem_12_cmp_1_z_1;

  rem_12_cmp_2 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_12_cmp_2_a,
      b => rem_12_cmp_2_b,
      z => rem_12_cmp_2_z_1
    );
  rem_12_cmp_2_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_12_cmp_2_a_63_0),65));
  rem_12_cmp_2_b <= '0' & rem_12_cmp_2_b_63_0;
  rem_12_cmp_2_z <= rem_12_cmp_2_z_1;

  rem_12_cmp_3 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_12_cmp_3_a,
      b => rem_12_cmp_3_b,
      z => rem_12_cmp_3_z_1
    );
  rem_12_cmp_3_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_12_cmp_3_a_63_0),65));
  rem_12_cmp_3_b <= '0' & rem_12_cmp_3_b_63_0;
  rem_12_cmp_3_z <= rem_12_cmp_3_z_1;

  rem_12_cmp_4 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_12_cmp_4_a,
      b => rem_12_cmp_4_b,
      z => rem_12_cmp_4_z_1
    );
  rem_12_cmp_4_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_12_cmp_4_a_63_0),65));
  rem_12_cmp_4_b <= '0' & rem_12_cmp_4_b_63_0;
  rem_12_cmp_4_z <= rem_12_cmp_4_z_1;

  rem_12_cmp_5 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_12_cmp_5_a,
      b => rem_12_cmp_5_b,
      z => rem_12_cmp_5_z_1
    );
  rem_12_cmp_5_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_12_cmp_5_a_63_0),65));
  rem_12_cmp_5_b <= '0' & rem_12_cmp_5_b_63_0;
  rem_12_cmp_5_z <= rem_12_cmp_5_z_1;

  rem_12_cmp_6 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_12_cmp_6_a,
      b => rem_12_cmp_6_b,
      z => rem_12_cmp_6_z_1
    );
  rem_12_cmp_6_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_12_cmp_6_a_63_0),65));
  rem_12_cmp_6_b <= '0' & rem_12_cmp_6_b_63_0;
  rem_12_cmp_6_z <= rem_12_cmp_6_z_1;

  rem_12_cmp_7 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_12_cmp_7_a,
      b => rem_12_cmp_7_b,
      z => rem_12_cmp_7_z_1
    );
  rem_12_cmp_7_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_12_cmp_7_a_63_0),65));
  rem_12_cmp_7_b <= '0' & rem_12_cmp_7_b_63_0;
  rem_12_cmp_7_z <= rem_12_cmp_7_z_1;

  rem_12_cmp_8 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_12_cmp_8_a,
      b => rem_12_cmp_8_b,
      z => rem_12_cmp_8_z_1
    );
  rem_12_cmp_8_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_12_cmp_8_a_63_0),65));
  rem_12_cmp_8_b <= '0' & rem_12_cmp_8_b_63_0;
  rem_12_cmp_8_z <= rem_12_cmp_8_z_1;

  rem_12_cmp_9 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_12_cmp_9_a,
      b => rem_12_cmp_9_b,
      z => rem_12_cmp_9_z_1
    );
  rem_12_cmp_9_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_12_cmp_9_a_63_0),65));
  rem_12_cmp_9_b <= '0' & rem_12_cmp_9_b_63_0;
  rem_12_cmp_9_z <= rem_12_cmp_9_z_1;

  rem_12_cmp_10 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_12_cmp_10_a,
      b => rem_12_cmp_10_b,
      z => rem_12_cmp_10_z_1
    );
  rem_12_cmp_10_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_12_cmp_10_a_63_0),65));
  rem_12_cmp_10_b <= '0' & rem_12_cmp_10_b_63_0;
  rem_12_cmp_10_z <= rem_12_cmp_10_z_1;

  rem_12_cmp_11 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_12_cmp_11_a,
      b => rem_12_cmp_11_b,
      z => rem_12_cmp_11_z_1
    );
  rem_12_cmp_11_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_12_cmp_11_a_63_0),65));
  rem_12_cmp_11_b <= '0' & rem_12_cmp_11_b_63_0;
  rem_12_cmp_11_z <= rem_12_cmp_11_z_1;

  COMP_LOOP_and_26_cse <= ccs_ccore_en AND main_stage_0_12 AND COMP_LOOP_asn_itm_11;
  COMP_LOOP_and_cse <= ccs_ccore_en AND (and_dcpl_294 OR and_dcpl_300 OR and_dcpl_306
      OR and_dcpl_312 OR and_dcpl_318 OR and_dcpl_324 OR and_dcpl_330 OR and_dcpl_336
      OR and_dcpl_342 OR and_dcpl_348 OR and_tmp_35);
  COMP_LOOP_and_2_cse <= ccs_ccore_en AND (and_dcpl_356 OR and_dcpl_360 OR and_dcpl_364
      OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_376 OR and_dcpl_379 OR and_dcpl_382
      OR and_dcpl_385 OR and_dcpl_388 OR mux_tmp_76);
  COMP_LOOP_and_4_cse <= ccs_ccore_en AND (and_dcpl_394 OR and_dcpl_397 OR and_dcpl_400
      OR and_dcpl_403 OR and_dcpl_406 OR and_dcpl_409 OR and_dcpl_413 OR and_dcpl_417
      OR and_dcpl_421 OR and_dcpl_425 OR and_tmp_80);
  COMP_LOOP_and_6_cse <= ccs_ccore_en AND (and_dcpl_431 OR and_dcpl_433 OR and_dcpl_435
      OR and_dcpl_437 OR and_dcpl_439 OR and_dcpl_442 OR and_dcpl_445 OR and_dcpl_448
      OR and_dcpl_451 OR and_dcpl_454 OR mux_tmp_141);
  COMP_LOOP_and_8_cse <= ccs_ccore_en AND (and_dcpl_461 OR and_dcpl_465 OR and_dcpl_469
      OR and_dcpl_473 OR and_dcpl_477 OR and_dcpl_480 OR and_dcpl_483 OR and_dcpl_486
      OR and_dcpl_489 OR and_dcpl_492 OR and_tmp_125);
  COMP_LOOP_and_10_cse <= ccs_ccore_en AND (and_dcpl_498 OR and_dcpl_500 OR and_dcpl_502
      OR and_dcpl_504 OR and_dcpl_506 OR and_dcpl_508 OR and_dcpl_510 OR and_dcpl_512
      OR and_dcpl_514 OR and_dcpl_516 OR mux_tmp_206);
  COMP_LOOP_and_12_cse <= ccs_ccore_en AND (and_dcpl_520 OR and_dcpl_523 OR and_dcpl_526
      OR and_dcpl_529 OR and_dcpl_532 OR and_dcpl_534 OR and_dcpl_536 OR and_dcpl_538
      OR and_dcpl_540 OR and_dcpl_542 OR and_tmp_170);
  COMP_LOOP_and_14_cse <= ccs_ccore_en AND (and_dcpl_546 OR and_dcpl_548 OR and_dcpl_550
      OR and_dcpl_552 OR and_dcpl_554 OR and_dcpl_556 OR and_dcpl_558 OR and_dcpl_560
      OR and_dcpl_562 OR and_dcpl_564 OR mux_tmp_271);
  COMP_LOOP_and_16_cse <= ccs_ccore_en AND (and_dcpl_569 OR and_dcpl_573 OR and_dcpl_577
      OR and_dcpl_581 OR and_dcpl_585 OR and_dcpl_589 OR and_dcpl_593 OR and_dcpl_597
      OR and_dcpl_601 OR and_dcpl_605 OR and_tmp_206);
  COMP_LOOP_and_18_cse <= ccs_ccore_en AND (and_dcpl_610 OR and_dcpl_612 OR and_dcpl_614
      OR and_dcpl_616 OR and_dcpl_618 OR and_dcpl_622 OR and_dcpl_625 OR and_dcpl_628
      OR and_dcpl_631 OR and_dcpl_634 OR mux_tmp_354);
  COMP_LOOP_and_20_cse <= ccs_ccore_en AND (and_dcpl_638 OR and_dcpl_641 OR and_dcpl_644
      OR and_dcpl_647 OR and_dcpl_650 OR and_dcpl_653 OR and_dcpl_657 OR and_dcpl_661
      OR and_dcpl_665 OR and_dcpl_669 OR and_tmp_233);
  COMP_LOOP_and_22_cse <= ccs_ccore_en AND (and_dcpl_673 OR and_dcpl_675 OR and_dcpl_677
      OR and_dcpl_679 OR and_dcpl_681 OR and_dcpl_684 OR and_dcpl_687 OR and_dcpl_690
      OR and_dcpl_693 OR and_dcpl_696 OR mux_tmp_437);
  COMP_LOOP_and_28_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_2;
  COMP_LOOP_and_30_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_6;
  COMP_LOOP_and_32_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_9;
  COMP_LOOP_and_34_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_11;
  COMP_LOOP_and_36_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_2;
  COMP_LOOP_and_38_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_6;
  COMP_LOOP_and_40_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_9;
  COMP_LOOP_and_42_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_11;
  COMP_LOOP_and_44_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_18 AND (NOT (rem_12cyc_st_10_1_0(0)));
  COMP_LOOP_and_46_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_18 AND (rem_12cyc_st_10_1_0(0));
  COMP_LOOP_and_48_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_23 AND (NOT (rem_12cyc_st_10_1_0(0)));
  COMP_LOOP_and_50_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_23 AND (rem_12cyc_st_10_1_0(0));
  COMP_LOOP_and_52_cse <= ccs_ccore_en AND and_dcpl_3;
  COMP_LOOP_and_54_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_29;
  COMP_LOOP_and_56_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_33;
  COMP_LOOP_and_58_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_36;
  COMP_LOOP_and_60_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_38;
  COMP_LOOP_and_62_cse <= ccs_ccore_en AND and_dcpl_40 AND and_dcpl_29;
  COMP_LOOP_and_64_cse <= ccs_ccore_en AND and_dcpl_40 AND and_dcpl_33;
  COMP_LOOP_and_66_cse <= ccs_ccore_en AND and_dcpl_40 AND and_dcpl_36;
  COMP_LOOP_and_68_cse <= ccs_ccore_en AND and_dcpl_40 AND and_dcpl_38;
  COMP_LOOP_and_70_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_45 AND (NOT (rem_12cyc_st_9_1_0(0)));
  COMP_LOOP_and_72_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_45 AND (rem_12cyc_st_9_1_0(0));
  COMP_LOOP_and_74_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_50 AND (NOT (rem_12cyc_st_9_1_0(0)));
  COMP_LOOP_and_76_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_50 AND (rem_12cyc_st_9_1_0(0));
  COMP_LOOP_and_78_cse <= ccs_ccore_en AND and_dcpl_30;
  COMP_LOOP_and_80_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_56;
  COMP_LOOP_and_82_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_60;
  COMP_LOOP_and_84_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_63;
  COMP_LOOP_and_86_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_65;
  COMP_LOOP_and_88_cse <= ccs_ccore_en AND and_dcpl_67 AND and_dcpl_56;
  COMP_LOOP_and_90_cse <= ccs_ccore_en AND and_dcpl_67 AND and_dcpl_60;
  COMP_LOOP_and_92_cse <= ccs_ccore_en AND and_dcpl_67 AND and_dcpl_63;
  COMP_LOOP_and_94_cse <= ccs_ccore_en AND and_dcpl_67 AND and_dcpl_65;
  COMP_LOOP_and_96_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_72 AND (NOT (rem_12cyc_st_8_1_0(0)));
  COMP_LOOP_and_98_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_72 AND (rem_12cyc_st_8_1_0(0));
  COMP_LOOP_and_100_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_77 AND (NOT
      (rem_12cyc_st_8_1_0(0)));
  COMP_LOOP_and_102_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_77 AND (rem_12cyc_st_8_1_0(0));
  COMP_LOOP_and_104_cse <= ccs_ccore_en AND and_dcpl_57;
  COMP_LOOP_and_106_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_83;
  COMP_LOOP_and_108_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_87;
  COMP_LOOP_and_110_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_90;
  COMP_LOOP_and_112_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_92;
  COMP_LOOP_and_114_cse <= ccs_ccore_en AND and_dcpl_94 AND and_dcpl_83;
  COMP_LOOP_and_116_cse <= ccs_ccore_en AND and_dcpl_94 AND and_dcpl_87;
  COMP_LOOP_and_118_cse <= ccs_ccore_en AND and_dcpl_94 AND and_dcpl_90;
  COMP_LOOP_and_120_cse <= ccs_ccore_en AND and_dcpl_94 AND and_dcpl_92;
  COMP_LOOP_and_122_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_99 AND (NOT
      (rem_12cyc_st_7_1_0(0)));
  COMP_LOOP_and_124_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_99 AND (rem_12cyc_st_7_1_0(0));
  COMP_LOOP_and_126_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_104 AND (NOT
      (rem_12cyc_st_7_1_0(0)));
  COMP_LOOP_and_128_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_104 AND (rem_12cyc_st_7_1_0(0));
  COMP_LOOP_and_130_cse <= ccs_ccore_en AND and_dcpl_84;
  COMP_LOOP_and_132_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_110;
  COMP_LOOP_and_134_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_115;
  COMP_LOOP_and_136_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_117;
  COMP_LOOP_and_138_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_119;
  COMP_LOOP_and_140_cse <= ccs_ccore_en AND and_dcpl_121 AND and_dcpl_110;
  COMP_LOOP_and_142_cse <= ccs_ccore_en AND and_dcpl_121 AND and_dcpl_115;
  COMP_LOOP_and_144_cse <= ccs_ccore_en AND and_dcpl_121 AND and_dcpl_117;
  COMP_LOOP_and_146_cse <= ccs_ccore_en AND and_dcpl_121 AND and_dcpl_119;
  COMP_LOOP_and_148_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_126 AND (NOT
      (rem_12cyc_st_6_1_0(1)));
  COMP_LOOP_and_150_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_129 AND (NOT
      (rem_12cyc_st_6_1_0(1)));
  COMP_LOOP_and_152_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_126 AND (rem_12cyc_st_6_1_0(1));
  COMP_LOOP_and_154_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_129 AND (rem_12cyc_st_6_1_0(1));
  COMP_LOOP_and_156_cse <= ccs_ccore_en AND and_dcpl_111;
  COMP_LOOP_and_158_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_137;
  COMP_LOOP_and_160_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_141;
  COMP_LOOP_and_162_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_144;
  COMP_LOOP_and_164_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_146;
  COMP_LOOP_and_166_cse <= ccs_ccore_en AND and_dcpl_148 AND and_dcpl_137;
  COMP_LOOP_and_168_cse <= ccs_ccore_en AND and_dcpl_148 AND and_dcpl_141;
  COMP_LOOP_and_170_cse <= ccs_ccore_en AND and_dcpl_148 AND and_dcpl_144;
  COMP_LOOP_and_172_cse <= ccs_ccore_en AND and_dcpl_148 AND and_dcpl_146;
  COMP_LOOP_and_174_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_153 AND (NOT
      (rem_12cyc_st_5_1_0(0)));
  COMP_LOOP_and_176_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_153 AND (rem_12cyc_st_5_1_0(0));
  COMP_LOOP_and_178_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_158 AND (NOT
      (rem_12cyc_st_5_1_0(0)));
  COMP_LOOP_and_180_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_158 AND (rem_12cyc_st_5_1_0(0));
  COMP_LOOP_and_182_cse <= ccs_ccore_en AND and_dcpl_138;
  COMP_LOOP_and_184_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_164;
  COMP_LOOP_and_186_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_168;
  COMP_LOOP_and_188_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_171;
  COMP_LOOP_and_190_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_173;
  COMP_LOOP_and_192_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_175 AND (NOT
      (rem_12cyc_st_4_1_0(0)));
  COMP_LOOP_and_194_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_175 AND (rem_12cyc_st_4_1_0(0));
  COMP_LOOP_and_196_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_180 AND (NOT
      (rem_12cyc_st_4_1_0(0)));
  COMP_LOOP_and_198_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_180 AND (rem_12cyc_st_4_1_0(0));
  COMP_LOOP_and_200_cse <= ccs_ccore_en AND and_dcpl_185 AND and_dcpl_164;
  COMP_LOOP_and_202_cse <= ccs_ccore_en AND and_dcpl_185 AND and_dcpl_168;
  COMP_LOOP_and_204_cse <= ccs_ccore_en AND and_dcpl_185 AND and_dcpl_171;
  COMP_LOOP_and_206_cse <= ccs_ccore_en AND and_dcpl_185 AND and_dcpl_173;
  COMP_LOOP_and_208_cse <= ccs_ccore_en AND and_dcpl_165;
  COMP_LOOP_and_210_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_191;
  COMP_LOOP_and_212_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_195;
  COMP_LOOP_and_214_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_198;
  COMP_LOOP_and_216_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_200;
  COMP_LOOP_and_218_cse <= ccs_ccore_en AND and_dcpl_202 AND and_dcpl_191;
  COMP_LOOP_and_220_cse <= ccs_ccore_en AND and_dcpl_202 AND and_dcpl_195;
  COMP_LOOP_and_222_cse <= ccs_ccore_en AND and_dcpl_202 AND and_dcpl_198;
  COMP_LOOP_and_224_cse <= ccs_ccore_en AND and_dcpl_202 AND and_dcpl_200;
  COMP_LOOP_and_226_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_207 AND (NOT
      (rem_12cyc_st_3_1_0(0)));
  COMP_LOOP_and_228_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_207 AND (rem_12cyc_st_3_1_0(0));
  COMP_LOOP_and_230_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_212 AND (NOT
      (rem_12cyc_st_3_1_0(0)));
  COMP_LOOP_and_232_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_212 AND (rem_12cyc_st_3_1_0(0));
  COMP_LOOP_and_234_cse <= ccs_ccore_en AND and_dcpl_192;
  COMP_LOOP_and_236_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_218;
  COMP_LOOP_and_238_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_222;
  COMP_LOOP_and_240_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_225;
  COMP_LOOP_and_242_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_227;
  COMP_LOOP_and_244_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_229 AND (NOT
      (rem_12cyc_st_2_1_0(0)));
  COMP_LOOP_and_246_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_229 AND (rem_12cyc_st_2_1_0(0));
  COMP_LOOP_and_248_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_234 AND (NOT
      (rem_12cyc_st_2_1_0(0)));
  COMP_LOOP_and_250_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_234 AND (rem_12cyc_st_2_1_0(0));
  COMP_LOOP_and_252_cse <= ccs_ccore_en AND and_dcpl_239 AND and_dcpl_218;
  COMP_LOOP_and_254_cse <= ccs_ccore_en AND and_dcpl_239 AND and_dcpl_222;
  COMP_LOOP_and_256_cse <= ccs_ccore_en AND and_dcpl_239 AND and_dcpl_225;
  COMP_LOOP_and_258_cse <= ccs_ccore_en AND and_dcpl_239 AND and_dcpl_227;
  COMP_LOOP_and_260_cse <= ccs_ccore_en AND and_dcpl_219;
  COMP_LOOP_and_262_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_245;
  COMP_LOOP_and_264_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_249;
  COMP_LOOP_and_266_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_252;
  COMP_LOOP_and_268_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_254;
  COMP_LOOP_and_270_cse <= ccs_ccore_en AND and_dcpl_256 AND and_dcpl_245;
  COMP_LOOP_and_272_cse <= ccs_ccore_en AND and_dcpl_256 AND and_dcpl_249;
  COMP_LOOP_and_274_cse <= ccs_ccore_en AND and_dcpl_256 AND and_dcpl_252;
  COMP_LOOP_and_276_cse <= ccs_ccore_en AND and_dcpl_256 AND and_dcpl_254;
  COMP_LOOP_and_278_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_261 AND (NOT
      (rem_12cyc_1_0(0)));
  COMP_LOOP_and_280_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_261 AND (rem_12cyc_1_0(0));
  COMP_LOOP_and_282_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_266 AND (NOT
      (rem_12cyc_1_0(0)));
  COMP_LOOP_and_284_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_266 AND (rem_12cyc_1_0(0));
  COMP_LOOP_and_286_cse <= ccs_ccore_en AND and_dcpl_246;
  COMP_LOOP_and_24_cse <= ccs_ccore_en AND ccs_ccore_start_rsci_idat;
  and_273_nl <= and_dcpl_272 AND and_dcpl_271;
  and_275_nl <= and_dcpl_272 AND and_dcpl_274;
  and_277_nl <= and_dcpl_272 AND and_dcpl_276;
  and_279_nl <= and_dcpl_272 AND and_dcpl_278;
  and_281_nl <= and_dcpl_280 AND and_dcpl_271;
  and_282_nl <= and_dcpl_280 AND and_dcpl_274;
  and_283_nl <= and_dcpl_280 AND and_dcpl_276;
  and_284_nl <= and_dcpl_280 AND and_dcpl_278;
  and_286_nl <= and_dcpl_285 AND and_dcpl_271;
  and_287_nl <= and_dcpl_285 AND and_dcpl_274;
  and_288_nl <= and_dcpl_285 AND and_dcpl_276;
  and_289_nl <= and_dcpl_285 AND and_dcpl_278;
  and_290_nl <= CONV_SL_1_1(rem_12cyc_st_12_3_2=STD_LOGIC_VECTOR'("11"));
  result_sva_duc_mx0 <= MUX1HOT_v_64_13_2((rem_12_cmp_1_z(63 DOWNTO 0)), (rem_12_cmp_2_z(63
      DOWNTO 0)), (rem_12_cmp_3_z(63 DOWNTO 0)), (rem_12_cmp_4_z(63 DOWNTO 0)), (rem_12_cmp_5_z(63
      DOWNTO 0)), (rem_12_cmp_6_z(63 DOWNTO 0)), (rem_12_cmp_7_z(63 DOWNTO 0)), (rem_12_cmp_8_z(63
      DOWNTO 0)), (rem_12_cmp_9_z(63 DOWNTO 0)), (rem_12_cmp_10_z(63 DOWNTO 0)),
      (rem_12_cmp_11_z(63 DOWNTO 0)), (rem_12_cmp_z(63 DOWNTO 0)), result_sva_duc,
      STD_LOGIC_VECTOR'( and_273_nl & and_275_nl & and_277_nl & and_279_nl & and_281_nl
      & and_282_nl & and_283_nl & and_284_nl & and_286_nl & and_287_nl & and_288_nl
      & and_289_nl & and_290_nl));
  COMP_LOOP_acc_1_tmp <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(rem_12cyc_3_2 &
      rem_12cyc_1_0) + UNSIGNED'( "0001"), 4));
  COMP_LOOP_COMP_LOOP_xor_nl <= (COMP_LOOP_acc_1_tmp(2)) XOR (COMP_LOOP_acc_1_tmp(3));
  COMP_LOOP_nor_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_tmp(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10")));
  COMP_LOOP_acc_tmp <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(COMP_LOOP_COMP_LOOP_xor_nl,
      1), 2) + CONV_UNSIGNED(CONV_UNSIGNED(COMP_LOOP_nor_nl, 1), 2), 2));
  and_dcpl_1 <= NOT((rem_12cyc_st_10_3_2(1)) OR (rem_12cyc_st_10_1_0(1)));
  and_dcpl_2 <= and_dcpl_1 AND (NOT (rem_12cyc_st_10_1_0(0)));
  and_dcpl_3 <= main_stage_0_11 AND COMP_LOOP_asn_itm_10;
  and_dcpl_4 <= and_dcpl_3 AND (NOT (rem_12cyc_st_10_3_2(0)));
  and_dcpl_6 <= and_dcpl_1 AND (rem_12cyc_st_10_1_0(0));
  and_dcpl_8 <= (NOT (rem_12cyc_st_10_3_2(1))) AND (rem_12cyc_st_10_1_0(1));
  and_dcpl_9 <= and_dcpl_8 AND (NOT (rem_12cyc_st_10_1_0(0)));
  and_dcpl_11 <= and_dcpl_8 AND (rem_12cyc_st_10_1_0(0));
  and_dcpl_13 <= and_dcpl_3 AND (rem_12cyc_st_10_3_2(0));
  and_dcpl_18 <= (rem_12cyc_st_10_3_2(1)) AND (NOT (rem_12cyc_st_10_1_0(1)));
  and_dcpl_23 <= (rem_12cyc_st_10_3_2(1)) AND (rem_12cyc_st_10_1_0(1));
  and_dcpl_28 <= NOT((rem_12cyc_st_9_3_2(1)) OR (rem_12cyc_st_9_1_0(1)));
  and_dcpl_29 <= and_dcpl_28 AND (NOT (rem_12cyc_st_9_1_0(0)));
  and_dcpl_30 <= main_stage_0_10 AND COMP_LOOP_asn_itm_9;
  and_dcpl_31 <= and_dcpl_30 AND (NOT (rem_12cyc_st_9_3_2(0)));
  and_dcpl_33 <= and_dcpl_28 AND (rem_12cyc_st_9_1_0(0));
  and_dcpl_35 <= (NOT (rem_12cyc_st_9_3_2(1))) AND (rem_12cyc_st_9_1_0(1));
  and_dcpl_36 <= and_dcpl_35 AND (NOT (rem_12cyc_st_9_1_0(0)));
  and_dcpl_38 <= and_dcpl_35 AND (rem_12cyc_st_9_1_0(0));
  and_dcpl_40 <= and_dcpl_30 AND (rem_12cyc_st_9_3_2(0));
  and_dcpl_45 <= (rem_12cyc_st_9_3_2(1)) AND (NOT (rem_12cyc_st_9_1_0(1)));
  and_dcpl_50 <= (rem_12cyc_st_9_3_2(1)) AND (rem_12cyc_st_9_1_0(1));
  and_dcpl_55 <= NOT((rem_12cyc_st_8_3_2(1)) OR (rem_12cyc_st_8_1_0(1)));
  and_dcpl_56 <= and_dcpl_55 AND (NOT (rem_12cyc_st_8_1_0(0)));
  and_dcpl_57 <= main_stage_0_9 AND COMP_LOOP_asn_itm_8;
  and_dcpl_58 <= and_dcpl_57 AND (NOT (rem_12cyc_st_8_3_2(0)));
  and_dcpl_60 <= and_dcpl_55 AND (rem_12cyc_st_8_1_0(0));
  and_dcpl_62 <= (NOT (rem_12cyc_st_8_3_2(1))) AND (rem_12cyc_st_8_1_0(1));
  and_dcpl_63 <= and_dcpl_62 AND (NOT (rem_12cyc_st_8_1_0(0)));
  and_dcpl_65 <= and_dcpl_62 AND (rem_12cyc_st_8_1_0(0));
  and_dcpl_67 <= and_dcpl_57 AND (rem_12cyc_st_8_3_2(0));
  and_dcpl_72 <= (rem_12cyc_st_8_3_2(1)) AND (NOT (rem_12cyc_st_8_1_0(1)));
  and_dcpl_77 <= (rem_12cyc_st_8_3_2(1)) AND (rem_12cyc_st_8_1_0(1));
  and_dcpl_82 <= NOT((rem_12cyc_st_7_3_2(1)) OR (rem_12cyc_st_7_1_0(1)));
  and_dcpl_83 <= and_dcpl_82 AND (NOT (rem_12cyc_st_7_1_0(0)));
  and_dcpl_84 <= main_stage_0_8 AND COMP_LOOP_asn_itm_7;
  and_dcpl_85 <= and_dcpl_84 AND (NOT (rem_12cyc_st_7_3_2(0)));
  and_dcpl_87 <= and_dcpl_82 AND (rem_12cyc_st_7_1_0(0));
  and_dcpl_89 <= (NOT (rem_12cyc_st_7_3_2(1))) AND (rem_12cyc_st_7_1_0(1));
  and_dcpl_90 <= and_dcpl_89 AND (NOT (rem_12cyc_st_7_1_0(0)));
  and_dcpl_92 <= and_dcpl_89 AND (rem_12cyc_st_7_1_0(0));
  and_dcpl_94 <= and_dcpl_84 AND (rem_12cyc_st_7_3_2(0));
  and_dcpl_99 <= (rem_12cyc_st_7_3_2(1)) AND (NOT (rem_12cyc_st_7_1_0(1)));
  and_dcpl_104 <= (rem_12cyc_st_7_3_2(1)) AND (rem_12cyc_st_7_1_0(1));
  and_dcpl_109 <= NOT((rem_12cyc_st_6_3_2(1)) OR (rem_12cyc_st_6_1_0(0)));
  and_dcpl_110 <= and_dcpl_109 AND (NOT (rem_12cyc_st_6_1_0(1)));
  and_dcpl_111 <= main_stage_0_7 AND COMP_LOOP_asn_itm_6;
  and_dcpl_112 <= and_dcpl_111 AND (NOT (rem_12cyc_st_6_3_2(0)));
  and_dcpl_114 <= (NOT (rem_12cyc_st_6_3_2(1))) AND (rem_12cyc_st_6_1_0(0));
  and_dcpl_115 <= and_dcpl_114 AND (NOT (rem_12cyc_st_6_1_0(1)));
  and_dcpl_117 <= and_dcpl_109 AND (rem_12cyc_st_6_1_0(1));
  and_dcpl_119 <= and_dcpl_114 AND (rem_12cyc_st_6_1_0(1));
  and_dcpl_121 <= and_dcpl_111 AND (rem_12cyc_st_6_3_2(0));
  and_dcpl_126 <= (rem_12cyc_st_6_3_2(1)) AND (NOT (rem_12cyc_st_6_1_0(0)));
  and_dcpl_129 <= (rem_12cyc_st_6_3_2(1)) AND (rem_12cyc_st_6_1_0(0));
  and_dcpl_136 <= NOT((rem_12cyc_st_5_3_2(1)) OR (rem_12cyc_st_5_1_0(1)));
  and_dcpl_137 <= and_dcpl_136 AND (NOT (rem_12cyc_st_5_1_0(0)));
  and_dcpl_138 <= main_stage_0_6 AND COMP_LOOP_asn_itm_5;
  and_dcpl_139 <= and_dcpl_138 AND (NOT (rem_12cyc_st_5_3_2(0)));
  and_dcpl_141 <= and_dcpl_136 AND (rem_12cyc_st_5_1_0(0));
  and_dcpl_143 <= (NOT (rem_12cyc_st_5_3_2(1))) AND (rem_12cyc_st_5_1_0(1));
  and_dcpl_144 <= and_dcpl_143 AND (NOT (rem_12cyc_st_5_1_0(0)));
  and_dcpl_146 <= and_dcpl_143 AND (rem_12cyc_st_5_1_0(0));
  and_dcpl_148 <= and_dcpl_138 AND (rem_12cyc_st_5_3_2(0));
  and_dcpl_153 <= (rem_12cyc_st_5_3_2(1)) AND (NOT (rem_12cyc_st_5_1_0(1)));
  and_dcpl_158 <= (rem_12cyc_st_5_3_2(1)) AND (rem_12cyc_st_5_1_0(1));
  and_dcpl_163 <= NOT((rem_12cyc_st_4_3_2(0)) OR (rem_12cyc_st_4_1_0(1)));
  and_dcpl_164 <= and_dcpl_163 AND (NOT (rem_12cyc_st_4_1_0(0)));
  and_dcpl_165 <= main_stage_0_5 AND COMP_LOOP_asn_itm_4;
  and_dcpl_166 <= and_dcpl_165 AND (NOT (rem_12cyc_st_4_3_2(1)));
  and_dcpl_168 <= and_dcpl_163 AND (rem_12cyc_st_4_1_0(0));
  and_dcpl_170 <= (NOT (rem_12cyc_st_4_3_2(0))) AND (rem_12cyc_st_4_1_0(1));
  and_dcpl_171 <= and_dcpl_170 AND (NOT (rem_12cyc_st_4_1_0(0)));
  and_dcpl_173 <= and_dcpl_170 AND (rem_12cyc_st_4_1_0(0));
  and_dcpl_175 <= (rem_12cyc_st_4_3_2(0)) AND (NOT (rem_12cyc_st_4_1_0(1)));
  and_dcpl_180 <= (rem_12cyc_st_4_3_2(0)) AND (rem_12cyc_st_4_1_0(1));
  and_dcpl_185 <= and_dcpl_165 AND (rem_12cyc_st_4_3_2(1));
  and_dcpl_190 <= NOT((rem_12cyc_st_3_3_2(1)) OR (rem_12cyc_st_3_1_0(1)));
  and_dcpl_191 <= and_dcpl_190 AND (NOT (rem_12cyc_st_3_1_0(0)));
  and_dcpl_192 <= main_stage_0_4 AND COMP_LOOP_asn_itm_3;
  and_dcpl_193 <= and_dcpl_192 AND (NOT (rem_12cyc_st_3_3_2(0)));
  and_dcpl_195 <= and_dcpl_190 AND (rem_12cyc_st_3_1_0(0));
  and_dcpl_197 <= (NOT (rem_12cyc_st_3_3_2(1))) AND (rem_12cyc_st_3_1_0(1));
  and_dcpl_198 <= and_dcpl_197 AND (NOT (rem_12cyc_st_3_1_0(0)));
  and_dcpl_200 <= and_dcpl_197 AND (rem_12cyc_st_3_1_0(0));
  and_dcpl_202 <= and_dcpl_192 AND (rem_12cyc_st_3_3_2(0));
  and_dcpl_207 <= (rem_12cyc_st_3_3_2(1)) AND (NOT (rem_12cyc_st_3_1_0(1)));
  and_dcpl_212 <= (rem_12cyc_st_3_3_2(1)) AND (rem_12cyc_st_3_1_0(1));
  and_dcpl_217 <= NOT((rem_12cyc_st_2_3_2(0)) OR (rem_12cyc_st_2_1_0(1)));
  and_dcpl_218 <= and_dcpl_217 AND (NOT (rem_12cyc_st_2_1_0(0)));
  and_dcpl_219 <= main_stage_0_3 AND COMP_LOOP_asn_itm_2;
  and_dcpl_220 <= and_dcpl_219 AND (NOT (rem_12cyc_st_2_3_2(1)));
  and_dcpl_222 <= and_dcpl_217 AND (rem_12cyc_st_2_1_0(0));
  and_dcpl_224 <= (NOT (rem_12cyc_st_2_3_2(0))) AND (rem_12cyc_st_2_1_0(1));
  and_dcpl_225 <= and_dcpl_224 AND (NOT (rem_12cyc_st_2_1_0(0)));
  and_dcpl_227 <= and_dcpl_224 AND (rem_12cyc_st_2_1_0(0));
  and_dcpl_229 <= (rem_12cyc_st_2_3_2(0)) AND (NOT (rem_12cyc_st_2_1_0(1)));
  and_dcpl_234 <= (rem_12cyc_st_2_3_2(0)) AND (rem_12cyc_st_2_1_0(1));
  and_dcpl_239 <= and_dcpl_219 AND (rem_12cyc_st_2_3_2(1));
  and_dcpl_244 <= NOT((rem_12cyc_3_2(1)) OR (rem_12cyc_1_0(1)));
  and_dcpl_245 <= and_dcpl_244 AND (NOT (rem_12cyc_1_0(0)));
  and_dcpl_246 <= main_stage_0_2 AND COMP_LOOP_asn_itm_1;
  and_dcpl_247 <= and_dcpl_246 AND (NOT (rem_12cyc_3_2(0)));
  and_dcpl_249 <= and_dcpl_244 AND (rem_12cyc_1_0(0));
  and_dcpl_251 <= (NOT (rem_12cyc_3_2(1))) AND (rem_12cyc_1_0(1));
  and_dcpl_252 <= and_dcpl_251 AND (NOT (rem_12cyc_1_0(0)));
  and_dcpl_254 <= and_dcpl_251 AND (rem_12cyc_1_0(0));
  and_dcpl_256 <= and_dcpl_246 AND (rem_12cyc_3_2(0));
  and_dcpl_261 <= (rem_12cyc_3_2(1)) AND (NOT (rem_12cyc_1_0(1)));
  and_dcpl_266 <= (rem_12cyc_3_2(1)) AND (rem_12cyc_1_0(1));
  and_dcpl_271 <= NOT(CONV_SL_1_1(rem_12cyc_st_12_1_0/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_272 <= NOT(CONV_SL_1_1(rem_12cyc_st_12_3_2/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_274 <= CONV_SL_1_1(rem_12cyc_st_12_1_0=STD_LOGIC_VECTOR'("01"));
  and_dcpl_276 <= CONV_SL_1_1(rem_12cyc_st_12_1_0=STD_LOGIC_VECTOR'("10"));
  and_dcpl_278 <= CONV_SL_1_1(rem_12cyc_st_12_1_0=STD_LOGIC_VECTOR'("11"));
  and_dcpl_280 <= CONV_SL_1_1(rem_12cyc_st_12_3_2=STD_LOGIC_VECTOR'("01"));
  and_dcpl_285 <= CONV_SL_1_1(rem_12cyc_st_12_3_2=STD_LOGIC_VECTOR'("10"));
  and_dcpl_291 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_292 <= ccs_ccore_start_rsci_idat AND (NOT (COMP_LOOP_acc_tmp(0)));
  and_dcpl_293 <= and_dcpl_292 AND (NOT (COMP_LOOP_acc_tmp(1)));
  and_dcpl_294 <= and_dcpl_293 AND and_dcpl_291;
  and_dcpl_295 <= NOT(CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_296 <= and_dcpl_295 AND (NOT (rem_12cyc_st_2_1_0(1)));
  and_dcpl_298 <= (NOT (rem_12cyc_st_2_1_0(0))) AND main_stage_0_3 AND COMP_LOOP_asn_itm_2;
  not_tmp_54 <= NOT(COMP_LOOP_asn_itm_1 AND main_stage_0_2);
  or_tmp_2 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_54;
  or_1_cse <= CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("00"));
  nor_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_2));
  mux_12_nl <= MUX_s_1_2_2(nor_nl, or_tmp_2, or_1_cse);
  and_dcpl_300 <= mux_12_nl AND and_dcpl_298 AND and_dcpl_296;
  and_dcpl_301 <= NOT(CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_302 <= and_dcpl_301 AND (NOT (rem_12cyc_st_3_1_0(1)));
  and_dcpl_304 <= (NOT (rem_12cyc_st_3_1_0(0))) AND main_stage_0_4 AND COMP_LOOP_asn_itm_3;
  or_6_cse <= (rem_12cyc_st_2_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp <= or_6_cse AND or_tmp_2;
  nor_516_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp));
  mux_13_nl <= MUX_s_1_2_2(nor_516_nl, and_tmp, or_1_cse);
  and_dcpl_306 <= mux_13_nl AND and_dcpl_304 AND and_dcpl_302;
  and_dcpl_307 <= NOT(CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_308 <= and_dcpl_307 AND (NOT (rem_12cyc_st_4_1_0(1)));
  and_dcpl_310 <= (NOT (rem_12cyc_st_4_1_0(0))) AND main_stage_0_5 AND COMP_LOOP_asn_itm_4;
  or_10_cse <= (rem_12cyc_st_3_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_2 <= or_6_cse AND or_10_cse AND or_tmp_2;
  nor_515_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_2));
  mux_14_nl <= MUX_s_1_2_2(nor_515_nl, and_tmp_2, or_1_cse);
  and_dcpl_312 <= mux_14_nl AND and_dcpl_310 AND and_dcpl_308;
  and_dcpl_313 <= NOT(CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_314 <= and_dcpl_313 AND (NOT (rem_12cyc_st_5_1_0(1)));
  and_dcpl_316 <= (NOT (rem_12cyc_st_5_1_0(0))) AND main_stage_0_6 AND COMP_LOOP_asn_itm_5;
  or_15_cse <= (rem_12cyc_st_4_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_5 <= or_6_cse AND or_10_cse AND or_15_cse AND or_tmp_2;
  nor_514_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_5));
  mux_15_nl <= MUX_s_1_2_2(nor_514_nl, and_tmp_5, or_1_cse);
  and_dcpl_318 <= mux_15_nl AND and_dcpl_316 AND and_dcpl_314;
  or_21_cse <= (rem_12cyc_st_5_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_9 <= or_6_cse AND or_10_cse AND or_15_cse AND or_21_cse AND or_tmp_2;
  nor_513_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_9));
  mux_16_nl <= MUX_s_1_2_2(nor_513_nl, and_tmp_9, or_1_cse);
  and_dcpl_324 <= mux_16_nl AND and_dcpl_112 AND and_dcpl_110;
  or_28_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_511_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_2));
  mux_17_nl <= MUX_s_1_2_2(nor_511_nl, or_tmp_2, or_28_cse);
  and_tmp_13 <= or_6_cse AND or_10_cse AND or_15_cse AND or_21_cse AND mux_17_nl;
  nor_512_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_13));
  mux_18_nl <= MUX_s_1_2_2(nor_512_nl, and_tmp_13, or_1_cse);
  and_dcpl_330 <= mux_18_nl AND and_dcpl_85 AND and_dcpl_83;
  or_37_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_508_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_2));
  mux_tmp_19 <= MUX_s_1_2_2(nor_508_nl, or_tmp_2, or_37_cse);
  nor_509_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_19));
  mux_20_nl <= MUX_s_1_2_2(nor_509_nl, mux_tmp_19, or_28_cse);
  and_tmp_17 <= or_6_cse AND or_10_cse AND or_15_cse AND or_21_cse AND mux_20_nl;
  nor_510_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_17));
  mux_21_nl <= MUX_s_1_2_2(nor_510_nl, and_tmp_17, or_1_cse);
  and_dcpl_336 <= mux_21_nl AND and_dcpl_58 AND and_dcpl_56;
  or_48_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_504_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_2));
  mux_tmp_22 <= MUX_s_1_2_2(nor_504_nl, or_tmp_2, or_48_cse);
  nor_505_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_22));
  mux_tmp_23 <= MUX_s_1_2_2(nor_505_nl, mux_tmp_22, or_37_cse);
  nor_506_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_23));
  mux_24_nl <= MUX_s_1_2_2(nor_506_nl, mux_tmp_23, or_28_cse);
  and_tmp_21 <= or_6_cse AND or_10_cse AND or_15_cse AND or_21_cse AND mux_24_nl;
  nor_507_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_21));
  mux_25_nl <= MUX_s_1_2_2(nor_507_nl, and_tmp_21, or_1_cse);
  and_dcpl_342 <= mux_25_nl AND and_dcpl_31 AND and_dcpl_29;
  nor_499_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_2));
  or_61_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_26 <= MUX_s_1_2_2(nor_499_nl, or_tmp_2, or_61_nl);
  nor_500_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_26));
  mux_tmp_27 <= MUX_s_1_2_2(nor_500_nl, mux_tmp_26, or_48_cse);
  nor_501_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_27));
  mux_tmp_28 <= MUX_s_1_2_2(nor_501_nl, mux_tmp_27, or_37_cse);
  nor_502_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_28));
  mux_29_nl <= MUX_s_1_2_2(nor_502_nl, mux_tmp_28, or_28_cse);
  and_tmp_25 <= or_6_cse AND or_10_cse AND or_15_cse AND or_21_cse AND mux_29_nl;
  nor_503_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_25));
  mux_30_nl <= MUX_s_1_2_2(nor_503_nl, and_tmp_25, or_1_cse);
  and_dcpl_348 <= mux_30_nl AND and_dcpl_4 AND and_dcpl_2;
  and_tmp_35 <= ((NOT main_stage_0_2) OR (NOT COMP_LOOP_asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_8)
      OR (NOT COMP_LOOP_asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_9)
      OR (NOT COMP_LOOP_asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_10)
      OR (NOT COMP_LOOP_asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"))) AND or_6_cse AND
      or_10_cse AND or_15_cse AND or_21_cse AND ((NOT main_stage_0_7) OR (NOT COMP_LOOP_asn_itm_6)
      OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00")))
      AND ((NOT main_stage_0_11) OR (NOT COMP_LOOP_asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("00"))) AND (CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT ccs_ccore_start_rsci_idat));
  and_dcpl_355 <= CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_356 <= and_dcpl_293 AND and_dcpl_355;
  and_dcpl_358 <= (rem_12cyc_st_2_1_0(0)) AND main_stage_0_3 AND COMP_LOOP_asn_itm_2;
  or_tmp_80 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_54;
  or_83_cse <= CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("00"));
  nor_498_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_80));
  mux_31_nl <= MUX_s_1_2_2(nor_498_nl, or_tmp_80, or_83_cse);
  and_dcpl_360 <= mux_31_nl AND and_dcpl_358 AND and_dcpl_296;
  and_dcpl_362 <= (rem_12cyc_st_3_1_0(0)) AND main_stage_0_4 AND COMP_LOOP_asn_itm_3;
  nand_276_cse <= NOT(COMP_LOOP_asn_itm_2 AND main_stage_0_3 AND (rem_12cyc_st_2_1_0(0)));
  or_88_cse <= (rem_12cyc_st_2_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1168_nl <= nand_276_cse AND or_tmp_80;
  mux_tmp_32 <= MUX_s_1_2_2(and_1168_nl, or_tmp_80, or_88_cse);
  nor_497_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_32));
  mux_33_nl <= MUX_s_1_2_2(nor_497_nl, mux_tmp_32, or_83_cse);
  and_dcpl_364 <= mux_33_nl AND and_dcpl_362 AND and_dcpl_302;
  and_dcpl_366 <= (rem_12cyc_st_4_1_0(0)) AND main_stage_0_5 AND COMP_LOOP_asn_itm_4;
  nand_274_cse <= NOT(COMP_LOOP_asn_itm_3 AND main_stage_0_4 AND (rem_12cyc_st_3_1_0(0)));
  or_93_cse <= (rem_12cyc_st_3_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1166_nl <= nand_274_cse AND or_tmp_80;
  mux_tmp_34 <= MUX_s_1_2_2(and_1166_nl, or_tmp_80, or_93_cse);
  and_1167_nl <= nand_276_cse AND mux_tmp_34;
  mux_tmp_35 <= MUX_s_1_2_2(and_1167_nl, mux_tmp_34, or_88_cse);
  nor_496_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_35));
  mux_36_nl <= MUX_s_1_2_2(nor_496_nl, mux_tmp_35, or_83_cse);
  and_dcpl_368 <= mux_36_nl AND and_dcpl_366 AND and_dcpl_308;
  and_dcpl_370 <= (rem_12cyc_st_5_1_0(0)) AND main_stage_0_6 AND COMP_LOOP_asn_itm_5;
  nand_271_cse <= NOT(COMP_LOOP_asn_itm_4 AND main_stage_0_5 AND (rem_12cyc_st_4_1_0(0)));
  or_100_cse <= (rem_12cyc_st_4_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1163_nl <= nand_271_cse AND or_tmp_80;
  mux_tmp_37 <= MUX_s_1_2_2(and_1163_nl, or_tmp_80, or_100_cse);
  and_1164_nl <= nand_274_cse AND mux_tmp_37;
  mux_tmp_38 <= MUX_s_1_2_2(and_1164_nl, mux_tmp_37, or_93_cse);
  and_1165_nl <= nand_276_cse AND mux_tmp_38;
  mux_tmp_39 <= MUX_s_1_2_2(and_1165_nl, mux_tmp_38, or_88_cse);
  nor_495_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_39));
  mux_40_nl <= MUX_s_1_2_2(nor_495_nl, mux_tmp_39, or_83_cse);
  and_dcpl_372 <= mux_40_nl AND and_dcpl_370 AND and_dcpl_314;
  nand_267_cse <= NOT(COMP_LOOP_asn_itm_5 AND main_stage_0_6 AND (rem_12cyc_st_5_1_0(0)));
  or_109_cse <= (rem_12cyc_st_5_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1159_nl <= nand_267_cse AND or_tmp_80;
  mux_tmp_41 <= MUX_s_1_2_2(and_1159_nl, or_tmp_80, or_109_cse);
  and_1160_nl <= nand_271_cse AND mux_tmp_41;
  mux_tmp_42 <= MUX_s_1_2_2(and_1160_nl, mux_tmp_41, or_100_cse);
  and_1161_nl <= nand_274_cse AND mux_tmp_42;
  mux_tmp_43 <= MUX_s_1_2_2(and_1161_nl, mux_tmp_42, or_93_cse);
  and_1162_nl <= nand_276_cse AND mux_tmp_43;
  mux_tmp_44 <= MUX_s_1_2_2(and_1162_nl, mux_tmp_43, or_88_cse);
  nor_494_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_44));
  mux_45_nl <= MUX_s_1_2_2(nor_494_nl, mux_tmp_44, or_83_cse);
  and_dcpl_376 <= mux_45_nl AND and_dcpl_112 AND and_dcpl_115;
  or_120_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_492_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_80));
  mux_tmp_46 <= MUX_s_1_2_2(nor_492_nl, or_tmp_80, or_120_cse);
  and_1155_nl <= nand_267_cse AND mux_tmp_46;
  mux_tmp_47 <= MUX_s_1_2_2(and_1155_nl, mux_tmp_46, or_109_cse);
  and_1156_nl <= nand_271_cse AND mux_tmp_47;
  mux_tmp_48 <= MUX_s_1_2_2(and_1156_nl, mux_tmp_47, or_100_cse);
  and_1157_nl <= nand_274_cse AND mux_tmp_48;
  mux_tmp_49 <= MUX_s_1_2_2(and_1157_nl, mux_tmp_48, or_93_cse);
  and_1158_nl <= nand_276_cse AND mux_tmp_49;
  mux_tmp_50 <= MUX_s_1_2_2(and_1158_nl, mux_tmp_49, or_88_cse);
  nor_493_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_50));
  mux_51_nl <= MUX_s_1_2_2(nor_493_nl, mux_tmp_50, or_83_cse);
  and_dcpl_379 <= mux_51_nl AND and_dcpl_85 AND and_dcpl_87;
  or_133_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_489_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_80));
  mux_tmp_52 <= MUX_s_1_2_2(nor_489_nl, or_tmp_80, or_133_cse);
  nor_490_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_52));
  mux_tmp_53 <= MUX_s_1_2_2(nor_490_nl, mux_tmp_52, or_120_cse);
  and_1151_nl <= nand_267_cse AND mux_tmp_53;
  mux_tmp_54 <= MUX_s_1_2_2(and_1151_nl, mux_tmp_53, or_109_cse);
  and_1152_nl <= nand_271_cse AND mux_tmp_54;
  mux_tmp_55 <= MUX_s_1_2_2(and_1152_nl, mux_tmp_54, or_100_cse);
  and_1153_nl <= nand_274_cse AND mux_tmp_55;
  mux_tmp_56 <= MUX_s_1_2_2(and_1153_nl, mux_tmp_55, or_93_cse);
  and_1154_nl <= nand_276_cse AND mux_tmp_56;
  mux_tmp_57 <= MUX_s_1_2_2(and_1154_nl, mux_tmp_56, or_88_cse);
  nor_491_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_57));
  mux_58_nl <= MUX_s_1_2_2(nor_491_nl, mux_tmp_57, or_83_cse);
  and_dcpl_382 <= mux_58_nl AND and_dcpl_58 AND and_dcpl_60;
  or_148_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_485_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_80));
  mux_tmp_59 <= MUX_s_1_2_2(nor_485_nl, or_tmp_80, or_148_cse);
  nor_486_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_59));
  mux_tmp_60 <= MUX_s_1_2_2(nor_486_nl, mux_tmp_59, or_133_cse);
  nor_487_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_60));
  mux_tmp_61 <= MUX_s_1_2_2(nor_487_nl, mux_tmp_60, or_120_cse);
  and_1147_nl <= nand_267_cse AND mux_tmp_61;
  mux_tmp_62 <= MUX_s_1_2_2(and_1147_nl, mux_tmp_61, or_109_cse);
  and_1148_nl <= nand_271_cse AND mux_tmp_62;
  mux_tmp_63 <= MUX_s_1_2_2(and_1148_nl, mux_tmp_62, or_100_cse);
  and_1149_nl <= nand_274_cse AND mux_tmp_63;
  mux_tmp_64 <= MUX_s_1_2_2(and_1149_nl, mux_tmp_63, or_93_cse);
  and_1150_nl <= nand_276_cse AND mux_tmp_64;
  mux_tmp_65 <= MUX_s_1_2_2(and_1150_nl, mux_tmp_64, or_88_cse);
  nor_488_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_65));
  mux_66_nl <= MUX_s_1_2_2(nor_488_nl, mux_tmp_65, or_83_cse);
  and_dcpl_385 <= mux_66_nl AND and_dcpl_31 AND and_dcpl_33;
  nor_480_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_80));
  or_165_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_67 <= MUX_s_1_2_2(nor_480_nl, or_tmp_80, or_165_nl);
  nor_481_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_67));
  mux_tmp_68 <= MUX_s_1_2_2(nor_481_nl, mux_tmp_67, or_148_cse);
  nor_482_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_68));
  mux_tmp_69 <= MUX_s_1_2_2(nor_482_nl, mux_tmp_68, or_133_cse);
  nor_483_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_69));
  mux_tmp_70 <= MUX_s_1_2_2(nor_483_nl, mux_tmp_69, or_120_cse);
  and_1143_nl <= nand_267_cse AND mux_tmp_70;
  mux_tmp_71 <= MUX_s_1_2_2(and_1143_nl, mux_tmp_70, or_109_cse);
  and_1144_nl <= nand_271_cse AND mux_tmp_71;
  mux_tmp_72 <= MUX_s_1_2_2(and_1144_nl, mux_tmp_71, or_100_cse);
  and_1145_nl <= nand_274_cse AND mux_tmp_72;
  mux_tmp_73 <= MUX_s_1_2_2(and_1145_nl, mux_tmp_72, or_93_cse);
  and_1146_nl <= nand_276_cse AND mux_tmp_73;
  mux_tmp_74 <= MUX_s_1_2_2(and_1146_nl, mux_tmp_73, or_88_cse);
  nor_484_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_74));
  mux_75_nl <= MUX_s_1_2_2(nor_484_nl, mux_tmp_74, or_83_cse);
  and_dcpl_388 <= mux_75_nl AND and_dcpl_4 AND and_dcpl_6;
  nand_250_cse <= NOT((COMP_LOOP_acc_1_tmp(0)) AND ccs_ccore_start_rsci_idat);
  and_tmp_44 <= ((NOT main_stage_0_8) OR (NOT COMP_LOOP_asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_9)
      OR (NOT COMP_LOOP_asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_10)
      OR (NOT COMP_LOOP_asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_3)
      OR (NOT COMP_LOOP_asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_4)
      OR (NOT COMP_LOOP_asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_5)
      OR (NOT COMP_LOOP_asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_6)
      OR (NOT COMP_LOOP_asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_7)
      OR (NOT COMP_LOOP_asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_11)
      OR (NOT COMP_LOOP_asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("00"))) AND (CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("00"))
      OR (COMP_LOOP_acc_1_tmp(1)) OR nand_250_cse);
  nor_479_nl <= NOT((rem_12cyc_1_0(0)) OR (NOT and_tmp_44));
  or_175_nl <= (NOT main_stage_0_2) OR (NOT COMP_LOOP_asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_1_0(1));
  mux_tmp_76 <= MUX_s_1_2_2(nor_479_nl, and_tmp_44, or_175_nl);
  and_dcpl_393 <= CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_394 <= and_dcpl_293 AND and_dcpl_393;
  and_dcpl_395 <= and_dcpl_295 AND (rem_12cyc_st_2_1_0(1));
  or_tmp_185 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_54;
  or_190_cse <= CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("00"));
  nor_478_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_185));
  mux_77_nl <= MUX_s_1_2_2(nor_478_nl, or_tmp_185, or_190_cse);
  and_dcpl_397 <= mux_77_nl AND and_dcpl_298 AND and_dcpl_395;
  and_dcpl_398 <= and_dcpl_301 AND (rem_12cyc_st_3_1_0(1));
  or_195_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp_45 <= or_195_cse AND or_tmp_185;
  nor_477_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_45));
  mux_78_nl <= MUX_s_1_2_2(nor_477_nl, and_tmp_45, or_190_cse);
  and_dcpl_400 <= mux_78_nl AND and_dcpl_304 AND and_dcpl_398;
  and_dcpl_401 <= and_dcpl_307 AND (rem_12cyc_st_4_1_0(1));
  or_199_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_47 <= or_195_cse AND or_199_cse AND or_tmp_185;
  nor_476_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_47));
  mux_79_nl <= MUX_s_1_2_2(nor_476_nl, and_tmp_47, or_190_cse);
  and_dcpl_403 <= mux_79_nl AND and_dcpl_310 AND and_dcpl_401;
  and_dcpl_404 <= and_dcpl_313 AND (rem_12cyc_st_5_1_0(1));
  or_204_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_50 <= or_195_cse AND or_199_cse AND or_204_cse AND or_tmp_185;
  nor_475_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_50));
  mux_80_nl <= MUX_s_1_2_2(nor_475_nl, and_tmp_50, or_190_cse);
  and_dcpl_406 <= mux_80_nl AND and_dcpl_316 AND and_dcpl_404;
  or_210_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_54 <= or_195_cse AND or_199_cse AND or_204_cse AND or_210_cse AND or_tmp_185;
  nor_474_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_54));
  mux_81_nl <= MUX_s_1_2_2(nor_474_nl, and_tmp_54, or_190_cse);
  and_dcpl_409 <= mux_81_nl AND and_dcpl_112 AND and_dcpl_117;
  or_217_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_472_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_185));
  mux_82_nl <= MUX_s_1_2_2(nor_472_nl, or_tmp_185, or_217_cse);
  and_tmp_58 <= or_195_cse AND or_199_cse AND or_204_cse AND or_210_cse AND mux_82_nl;
  nor_473_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_58));
  mux_83_nl <= MUX_s_1_2_2(nor_473_nl, and_tmp_58, or_190_cse);
  and_dcpl_413 <= mux_83_nl AND and_dcpl_85 AND and_dcpl_90;
  or_226_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_469_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_185));
  mux_tmp_84 <= MUX_s_1_2_2(nor_469_nl, or_tmp_185, or_226_cse);
  nor_470_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_84));
  mux_85_nl <= MUX_s_1_2_2(nor_470_nl, mux_tmp_84, or_217_cse);
  and_tmp_62 <= or_195_cse AND or_199_cse AND or_204_cse AND or_210_cse AND mux_85_nl;
  nor_471_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_62));
  mux_86_nl <= MUX_s_1_2_2(nor_471_nl, and_tmp_62, or_190_cse);
  and_dcpl_417 <= mux_86_nl AND and_dcpl_58 AND and_dcpl_63;
  or_237_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_465_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_185));
  mux_tmp_87 <= MUX_s_1_2_2(nor_465_nl, or_tmp_185, or_237_cse);
  nor_466_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_87));
  mux_tmp_88 <= MUX_s_1_2_2(nor_466_nl, mux_tmp_87, or_226_cse);
  nor_467_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_88));
  mux_89_nl <= MUX_s_1_2_2(nor_467_nl, mux_tmp_88, or_217_cse);
  and_tmp_66 <= or_195_cse AND or_199_cse AND or_204_cse AND or_210_cse AND mux_89_nl;
  nor_468_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_66));
  mux_90_nl <= MUX_s_1_2_2(nor_468_nl, and_tmp_66, or_190_cse);
  and_dcpl_421 <= mux_90_nl AND and_dcpl_31 AND and_dcpl_36;
  nor_460_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_185));
  or_250_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_91 <= MUX_s_1_2_2(nor_460_nl, or_tmp_185, or_250_nl);
  nor_461_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_91));
  mux_tmp_92 <= MUX_s_1_2_2(nor_461_nl, mux_tmp_91, or_237_cse);
  nor_462_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_92));
  mux_tmp_93 <= MUX_s_1_2_2(nor_462_nl, mux_tmp_92, or_226_cse);
  nor_463_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_93));
  mux_94_nl <= MUX_s_1_2_2(nor_463_nl, mux_tmp_93, or_217_cse);
  and_tmp_70 <= or_195_cse AND or_199_cse AND or_204_cse AND or_210_cse AND mux_94_nl;
  nor_464_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_70));
  mux_95_nl <= MUX_s_1_2_2(nor_464_nl, and_tmp_70, or_190_cse);
  and_dcpl_425 <= mux_95_nl AND and_dcpl_4 AND and_dcpl_9;
  and_tmp_80 <= ((NOT main_stage_0_2) OR (NOT COMP_LOOP_asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10"))) AND ((NOT main_stage_0_8)
      OR (NOT COMP_LOOP_asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_9)
      OR (NOT COMP_LOOP_asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_10)
      OR (NOT COMP_LOOP_asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"))) AND or_195_cse
      AND or_199_cse AND or_204_cse AND or_210_cse AND ((NOT main_stage_0_7) OR (NOT
      COMP_LOOP_asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_11)
      OR (NOT COMP_LOOP_asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("00"))) AND (CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT ccs_ccore_start_rsci_idat));
  and_dcpl_430 <= CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_431 <= and_dcpl_293 AND and_dcpl_430;
  or_tmp_263 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_54;
  or_270_cse <= CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("00"));
  nor_459_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_263));
  mux_96_nl <= MUX_s_1_2_2(nor_459_nl, or_tmp_263, or_270_cse);
  and_dcpl_433 <= mux_96_nl AND and_dcpl_358 AND and_dcpl_395;
  or_275_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1142_nl <= nand_276_cse AND or_tmp_263;
  mux_tmp_97 <= MUX_s_1_2_2(and_1142_nl, or_tmp_263, or_275_cse);
  nor_458_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_97));
  mux_98_nl <= MUX_s_1_2_2(nor_458_nl, mux_tmp_97, or_270_cse);
  and_dcpl_435 <= mux_98_nl AND and_dcpl_362 AND and_dcpl_398;
  or_280_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1140_nl <= nand_274_cse AND or_tmp_263;
  mux_tmp_99 <= MUX_s_1_2_2(and_1140_nl, or_tmp_263, or_280_cse);
  and_1141_nl <= nand_276_cse AND mux_tmp_99;
  mux_tmp_100 <= MUX_s_1_2_2(and_1141_nl, mux_tmp_99, or_275_cse);
  nor_457_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_100));
  mux_101_nl <= MUX_s_1_2_2(nor_457_nl, mux_tmp_100, or_270_cse);
  and_dcpl_437 <= mux_101_nl AND and_dcpl_366 AND and_dcpl_401;
  or_287_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1137_nl <= nand_271_cse AND or_tmp_263;
  mux_tmp_102 <= MUX_s_1_2_2(and_1137_nl, or_tmp_263, or_287_cse);
  and_1138_nl <= nand_274_cse AND mux_tmp_102;
  mux_tmp_103 <= MUX_s_1_2_2(and_1138_nl, mux_tmp_102, or_280_cse);
  and_1139_nl <= nand_276_cse AND mux_tmp_103;
  mux_tmp_104 <= MUX_s_1_2_2(and_1139_nl, mux_tmp_103, or_275_cse);
  nor_456_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_104));
  mux_105_nl <= MUX_s_1_2_2(nor_456_nl, mux_tmp_104, or_270_cse);
  and_dcpl_439 <= mux_105_nl AND and_dcpl_370 AND and_dcpl_404;
  or_296_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1133_nl <= nand_267_cse AND or_tmp_263;
  mux_tmp_106 <= MUX_s_1_2_2(and_1133_nl, or_tmp_263, or_296_cse);
  and_1134_nl <= nand_271_cse AND mux_tmp_106;
  mux_tmp_107 <= MUX_s_1_2_2(and_1134_nl, mux_tmp_106, or_287_cse);
  and_1135_nl <= nand_274_cse AND mux_tmp_107;
  mux_tmp_108 <= MUX_s_1_2_2(and_1135_nl, mux_tmp_107, or_280_cse);
  and_1136_nl <= nand_276_cse AND mux_tmp_108;
  mux_tmp_109 <= MUX_s_1_2_2(and_1136_nl, mux_tmp_108, or_275_cse);
  nor_455_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_109));
  mux_110_nl <= MUX_s_1_2_2(nor_455_nl, mux_tmp_109, or_270_cse);
  and_dcpl_442 <= mux_110_nl AND and_dcpl_112 AND and_dcpl_119;
  or_307_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_453_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_263));
  mux_tmp_111 <= MUX_s_1_2_2(nor_453_nl, or_tmp_263, or_307_cse);
  and_1129_nl <= nand_267_cse AND mux_tmp_111;
  mux_tmp_112 <= MUX_s_1_2_2(and_1129_nl, mux_tmp_111, or_296_cse);
  and_1130_nl <= nand_271_cse AND mux_tmp_112;
  mux_tmp_113 <= MUX_s_1_2_2(and_1130_nl, mux_tmp_112, or_287_cse);
  and_1131_nl <= nand_274_cse AND mux_tmp_113;
  mux_tmp_114 <= MUX_s_1_2_2(and_1131_nl, mux_tmp_113, or_280_cse);
  and_1132_nl <= nand_276_cse AND mux_tmp_114;
  mux_tmp_115 <= MUX_s_1_2_2(and_1132_nl, mux_tmp_114, or_275_cse);
  nor_454_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_115));
  mux_116_nl <= MUX_s_1_2_2(nor_454_nl, mux_tmp_115, or_270_cse);
  and_dcpl_445 <= mux_116_nl AND and_dcpl_85 AND and_dcpl_92;
  or_320_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_450_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_263));
  mux_tmp_117 <= MUX_s_1_2_2(nor_450_nl, or_tmp_263, or_320_cse);
  nor_451_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_117));
  mux_tmp_118 <= MUX_s_1_2_2(nor_451_nl, mux_tmp_117, or_307_cse);
  and_1125_nl <= nand_267_cse AND mux_tmp_118;
  mux_tmp_119 <= MUX_s_1_2_2(and_1125_nl, mux_tmp_118, or_296_cse);
  and_1126_nl <= nand_271_cse AND mux_tmp_119;
  mux_tmp_120 <= MUX_s_1_2_2(and_1126_nl, mux_tmp_119, or_287_cse);
  and_1127_nl <= nand_274_cse AND mux_tmp_120;
  mux_tmp_121 <= MUX_s_1_2_2(and_1127_nl, mux_tmp_120, or_280_cse);
  and_1128_nl <= nand_276_cse AND mux_tmp_121;
  mux_tmp_122 <= MUX_s_1_2_2(and_1128_nl, mux_tmp_121, or_275_cse);
  nor_452_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_122));
  mux_123_nl <= MUX_s_1_2_2(nor_452_nl, mux_tmp_122, or_270_cse);
  and_dcpl_448 <= mux_123_nl AND and_dcpl_58 AND and_dcpl_65;
  or_335_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_446_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_263));
  mux_tmp_124 <= MUX_s_1_2_2(nor_446_nl, or_tmp_263, or_335_cse);
  nor_447_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_124));
  mux_tmp_125 <= MUX_s_1_2_2(nor_447_nl, mux_tmp_124, or_320_cse);
  nor_448_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_125));
  mux_tmp_126 <= MUX_s_1_2_2(nor_448_nl, mux_tmp_125, or_307_cse);
  and_1121_nl <= nand_267_cse AND mux_tmp_126;
  mux_tmp_127 <= MUX_s_1_2_2(and_1121_nl, mux_tmp_126, or_296_cse);
  and_1122_nl <= nand_271_cse AND mux_tmp_127;
  mux_tmp_128 <= MUX_s_1_2_2(and_1122_nl, mux_tmp_127, or_287_cse);
  and_1123_nl <= nand_274_cse AND mux_tmp_128;
  mux_tmp_129 <= MUX_s_1_2_2(and_1123_nl, mux_tmp_128, or_280_cse);
  and_1124_nl <= nand_276_cse AND mux_tmp_129;
  mux_tmp_130 <= MUX_s_1_2_2(and_1124_nl, mux_tmp_129, or_275_cse);
  nor_449_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_130));
  mux_131_nl <= MUX_s_1_2_2(nor_449_nl, mux_tmp_130, or_270_cse);
  and_dcpl_451 <= mux_131_nl AND and_dcpl_31 AND and_dcpl_38;
  nor_441_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_263));
  or_352_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_132 <= MUX_s_1_2_2(nor_441_nl, or_tmp_263, or_352_nl);
  nor_442_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_132));
  mux_tmp_133 <= MUX_s_1_2_2(nor_442_nl, mux_tmp_132, or_335_cse);
  nor_443_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_133));
  mux_tmp_134 <= MUX_s_1_2_2(nor_443_nl, mux_tmp_133, or_320_cse);
  nor_444_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_134));
  mux_tmp_135 <= MUX_s_1_2_2(nor_444_nl, mux_tmp_134, or_307_cse);
  and_1117_nl <= nand_267_cse AND mux_tmp_135;
  mux_tmp_136 <= MUX_s_1_2_2(and_1117_nl, mux_tmp_135, or_296_cse);
  and_1118_nl <= nand_271_cse AND mux_tmp_136;
  mux_tmp_137 <= MUX_s_1_2_2(and_1118_nl, mux_tmp_136, or_287_cse);
  and_1119_nl <= nand_274_cse AND mux_tmp_137;
  mux_tmp_138 <= MUX_s_1_2_2(and_1119_nl, mux_tmp_137, or_280_cse);
  and_1120_nl <= nand_276_cse AND mux_tmp_138;
  mux_tmp_139 <= MUX_s_1_2_2(and_1120_nl, mux_tmp_138, or_275_cse);
  nor_445_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_139));
  mux_140_nl <= MUX_s_1_2_2(nor_445_nl, mux_tmp_139, or_270_cse);
  and_dcpl_454 <= mux_140_nl AND and_dcpl_4 AND and_dcpl_11;
  nand_222_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND ccs_ccore_start_rsci_idat);
  and_tmp_89 <= ((NOT main_stage_0_8) OR (NOT COMP_LOOP_asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_9)
      OR (NOT COMP_LOOP_asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_10)
      OR (NOT COMP_LOOP_asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_3)
      OR (NOT COMP_LOOP_asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_4)
      OR (NOT COMP_LOOP_asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_5)
      OR (NOT COMP_LOOP_asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_6)
      OR (NOT COMP_LOOP_asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_7)
      OR (NOT COMP_LOOP_asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_11)
      OR (NOT COMP_LOOP_asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("00"))) AND (CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("00"))
      OR nand_222_cse);
  nand_223_cse <= NOT(CONV_SL_1_1(rem_12cyc_1_0=STD_LOGIC_VECTOR'("11")));
  and_1116_nl <= nand_223_cse AND and_tmp_89;
  or_362_nl <= (NOT main_stage_0_2) OR (NOT COMP_LOOP_asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_141 <= MUX_s_1_2_2(and_1116_nl, and_tmp_89, or_362_nl);
  and_dcpl_460 <= ccs_ccore_start_rsci_idat AND CONV_SL_1_1(COMP_LOOP_acc_tmp=STD_LOGIC_VECTOR'("01"));
  and_dcpl_461 <= and_dcpl_460 AND and_dcpl_291;
  and_dcpl_462 <= CONV_SL_1_1(rem_12cyc_st_2_3_2=STD_LOGIC_VECTOR'("01"));
  and_dcpl_463 <= and_dcpl_462 AND (NOT (rem_12cyc_st_2_1_0(1)));
  not_tmp_332 <= NOT((rem_12cyc_3_2(0)) AND COMP_LOOP_asn_itm_1 AND main_stage_0_2);
  or_tmp_368 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00")) OR (rem_12cyc_3_2(1))
      OR not_tmp_332;
  nand_281_cse <= NOT((COMP_LOOP_acc_tmp(0)) AND ccs_ccore_start_rsci_idat);
  or_377_cse <= CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (COMP_LOOP_acc_tmp(1));
  and_1172_nl <= nand_281_cse AND or_tmp_368;
  mux_142_nl <= MUX_s_1_2_2(and_1172_nl, or_tmp_368, or_377_cse);
  and_dcpl_465 <= mux_142_nl AND and_dcpl_298 AND and_dcpl_463;
  and_dcpl_466 <= CONV_SL_1_1(rem_12cyc_st_3_3_2=STD_LOGIC_VECTOR'("01"));
  and_dcpl_467 <= and_dcpl_466 AND (NOT (rem_12cyc_st_3_1_0(1)));
  or_382_cse <= (rem_12cyc_st_2_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp_90 <= or_382_cse AND or_tmp_368;
  and_1114_nl <= nand_281_cse AND and_tmp_90;
  mux_143_nl <= MUX_s_1_2_2(and_1114_nl, and_tmp_90, or_377_cse);
  and_dcpl_469 <= mux_143_nl AND and_dcpl_304 AND and_dcpl_467;
  and_dcpl_470 <= CONV_SL_1_1(rem_12cyc_st_4_3_2=STD_LOGIC_VECTOR'("01"));
  and_dcpl_471 <= and_dcpl_470 AND (NOT (rem_12cyc_st_4_1_0(1)));
  or_386_cse <= (rem_12cyc_st_3_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_92 <= or_382_cse AND or_386_cse AND or_tmp_368;
  and_1113_nl <= nand_281_cse AND and_tmp_92;
  mux_144_nl <= MUX_s_1_2_2(and_1113_nl, and_tmp_92, or_377_cse);
  and_dcpl_473 <= mux_144_nl AND and_dcpl_310 AND and_dcpl_471;
  and_dcpl_474 <= CONV_SL_1_1(rem_12cyc_st_5_3_2=STD_LOGIC_VECTOR'("01"));
  and_dcpl_475 <= and_dcpl_474 AND (NOT (rem_12cyc_st_5_1_0(1)));
  or_391_cse <= (rem_12cyc_st_4_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_95 <= or_382_cse AND or_386_cse AND or_391_cse AND or_tmp_368;
  and_1112_nl <= nand_281_cse AND and_tmp_95;
  mux_145_nl <= MUX_s_1_2_2(and_1112_nl, and_tmp_95, or_377_cse);
  and_dcpl_477 <= mux_145_nl AND and_dcpl_316 AND and_dcpl_475;
  or_397_cse <= (rem_12cyc_st_5_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_99 <= or_382_cse AND or_386_cse AND or_391_cse AND or_397_cse AND or_tmp_368;
  and_1111_nl <= nand_281_cse AND and_tmp_99;
  mux_146_nl <= MUX_s_1_2_2(and_1111_nl, and_tmp_99, or_377_cse);
  and_dcpl_480 <= mux_146_nl AND and_dcpl_121 AND and_dcpl_110;
  nand_215_cse <= NOT((rem_12cyc_st_6_3_2(0)) AND COMP_LOOP_asn_itm_6 AND main_stage_0_7);
  or_404_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00")) OR (rem_12cyc_st_6_3_2(1));
  and_1109_nl <= nand_215_cse AND or_tmp_368;
  mux_147_nl <= MUX_s_1_2_2(and_1109_nl, or_tmp_368, or_404_cse);
  and_tmp_103 <= or_382_cse AND or_386_cse AND or_391_cse AND or_397_cse AND mux_147_nl;
  and_1110_nl <= nand_281_cse AND and_tmp_103;
  mux_148_nl <= MUX_s_1_2_2(and_1110_nl, and_tmp_103, or_377_cse);
  and_dcpl_483 <= mux_148_nl AND and_dcpl_94 AND and_dcpl_83;
  nand_212_cse <= NOT((rem_12cyc_st_7_3_2(0)) AND COMP_LOOP_asn_itm_7 AND main_stage_0_8);
  or_413_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00")) OR (rem_12cyc_st_7_3_2(1));
  and_1106_nl <= nand_212_cse AND or_tmp_368;
  mux_tmp_149 <= MUX_s_1_2_2(and_1106_nl, or_tmp_368, or_413_cse);
  and_1107_nl <= nand_215_cse AND mux_tmp_149;
  mux_150_nl <= MUX_s_1_2_2(and_1107_nl, mux_tmp_149, or_404_cse);
  and_tmp_107 <= or_382_cse AND or_386_cse AND or_391_cse AND or_397_cse AND mux_150_nl;
  and_1108_nl <= nand_281_cse AND and_tmp_107;
  mux_151_nl <= MUX_s_1_2_2(and_1108_nl, and_tmp_107, or_377_cse);
  and_dcpl_486 <= mux_151_nl AND and_dcpl_67 AND and_dcpl_56;
  nand_208_cse <= NOT((rem_12cyc_st_8_3_2(0)) AND COMP_LOOP_asn_itm_8 AND main_stage_0_9);
  or_424_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00")) OR (rem_12cyc_st_8_3_2(1));
  and_1102_nl <= nand_208_cse AND or_tmp_368;
  mux_tmp_152 <= MUX_s_1_2_2(and_1102_nl, or_tmp_368, or_424_cse);
  and_1103_nl <= nand_212_cse AND mux_tmp_152;
  mux_tmp_153 <= MUX_s_1_2_2(and_1103_nl, mux_tmp_152, or_413_cse);
  and_1104_nl <= nand_215_cse AND mux_tmp_153;
  mux_154_nl <= MUX_s_1_2_2(and_1104_nl, mux_tmp_153, or_404_cse);
  and_tmp_111 <= or_382_cse AND or_386_cse AND or_391_cse AND or_397_cse AND mux_154_nl;
  and_1105_nl <= nand_281_cse AND and_tmp_111;
  mux_155_nl <= MUX_s_1_2_2(and_1105_nl, and_tmp_111, or_377_cse);
  and_dcpl_489 <= mux_155_nl AND and_dcpl_40 AND and_dcpl_29;
  nand_203_cse <= NOT((rem_12cyc_st_9_3_2(0)) AND COMP_LOOP_asn_itm_9 AND main_stage_0_10);
  and_1097_nl <= nand_203_cse AND or_tmp_368;
  or_437_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00")) OR (rem_12cyc_st_9_3_2(1));
  mux_tmp_156 <= MUX_s_1_2_2(and_1097_nl, or_tmp_368, or_437_nl);
  and_1098_nl <= nand_208_cse AND mux_tmp_156;
  mux_tmp_157 <= MUX_s_1_2_2(and_1098_nl, mux_tmp_156, or_424_cse);
  and_1099_nl <= nand_212_cse AND mux_tmp_157;
  mux_tmp_158 <= MUX_s_1_2_2(and_1099_nl, mux_tmp_157, or_413_cse);
  and_1100_nl <= nand_215_cse AND mux_tmp_158;
  mux_159_nl <= MUX_s_1_2_2(and_1100_nl, mux_tmp_158, or_404_cse);
  and_tmp_115 <= or_382_cse AND or_386_cse AND or_391_cse AND or_397_cse AND mux_159_nl;
  and_1101_nl <= nand_281_cse AND and_tmp_115;
  mux_160_nl <= MUX_s_1_2_2(and_1101_nl, and_tmp_115, or_377_cse);
  and_dcpl_492 <= mux_160_nl AND and_dcpl_13 AND and_dcpl_2;
  and_tmp_125 <= ((NOT main_stage_0_2) OR (NOT COMP_LOOP_asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_8)
      OR (NOT COMP_LOOP_asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_9)
      OR (NOT COMP_LOOP_asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_10)
      OR (NOT COMP_LOOP_asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("01"))) AND or_382_cse
      AND or_386_cse AND or_391_cse AND or_397_cse AND ((NOT main_stage_0_7) OR (NOT
      COMP_LOOP_asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_11)
      OR (NOT COMP_LOOP_asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("01"))) AND (CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT ccs_ccore_start_rsci_idat));
  and_dcpl_498 <= and_dcpl_460 AND and_dcpl_355;
  or_tmp_446 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("01")) OR (rem_12cyc_3_2(1))
      OR not_tmp_332;
  or_458_cse <= CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (COMP_LOOP_acc_tmp(1));
  and_1171_nl <= nand_281_cse AND or_tmp_446;
  mux_161_nl <= MUX_s_1_2_2(and_1171_nl, or_tmp_446, or_458_cse);
  and_dcpl_500 <= mux_161_nl AND and_dcpl_358 AND and_dcpl_463;
  or_463_cse <= (rem_12cyc_st_2_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("01"));
  and_1094_nl <= nand_276_cse AND or_tmp_446;
  mux_tmp_162 <= MUX_s_1_2_2(and_1094_nl, or_tmp_446, or_463_cse);
  and_1095_nl <= nand_281_cse AND mux_tmp_162;
  mux_163_nl <= MUX_s_1_2_2(and_1095_nl, mux_tmp_162, or_458_cse);
  and_dcpl_502 <= mux_163_nl AND and_dcpl_362 AND and_dcpl_467;
  nand_198_cse <= NOT((rem_12cyc_st_3_3_2(0)) AND COMP_LOOP_asn_itm_3 AND main_stage_0_4
      AND (rem_12cyc_st_3_1_0(0)));
  or_468_cse <= (rem_12cyc_st_3_1_0(1)) OR (rem_12cyc_st_3_3_2(1));
  and_1091_nl <= nand_198_cse AND or_tmp_446;
  mux_tmp_164 <= MUX_s_1_2_2(and_1091_nl, or_tmp_446, or_468_cse);
  and_1092_nl <= nand_276_cse AND mux_tmp_164;
  mux_tmp_165 <= MUX_s_1_2_2(and_1092_nl, mux_tmp_164, or_463_cse);
  and_1093_nl <= nand_281_cse AND mux_tmp_165;
  mux_166_nl <= MUX_s_1_2_2(and_1093_nl, mux_tmp_165, or_458_cse);
  and_dcpl_504 <= mux_166_nl AND and_dcpl_366 AND and_dcpl_471;
  or_475_cse <= (rem_12cyc_st_4_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("01"));
  and_1087_nl <= nand_271_cse AND or_tmp_446;
  mux_tmp_167 <= MUX_s_1_2_2(and_1087_nl, or_tmp_446, or_475_cse);
  and_1088_nl <= nand_198_cse AND mux_tmp_167;
  mux_tmp_168 <= MUX_s_1_2_2(and_1088_nl, mux_tmp_167, or_468_cse);
  and_1089_nl <= nand_276_cse AND mux_tmp_168;
  mux_tmp_169 <= MUX_s_1_2_2(and_1089_nl, mux_tmp_168, or_463_cse);
  and_1090_nl <= nand_281_cse AND mux_tmp_169;
  mux_170_nl <= MUX_s_1_2_2(and_1090_nl, mux_tmp_169, or_458_cse);
  and_dcpl_506 <= mux_170_nl AND and_dcpl_370 AND and_dcpl_475;
  nand_189_cse <= NOT((rem_12cyc_st_5_3_2(0)) AND COMP_LOOP_asn_itm_5 AND main_stage_0_6
      AND (rem_12cyc_st_5_1_0(0)));
  or_484_cse <= (rem_12cyc_st_5_1_0(1)) OR (rem_12cyc_st_5_3_2(1));
  and_1082_nl <= nand_189_cse AND or_tmp_446;
  mux_tmp_171 <= MUX_s_1_2_2(and_1082_nl, or_tmp_446, or_484_cse);
  and_1083_nl <= nand_271_cse AND mux_tmp_171;
  mux_tmp_172 <= MUX_s_1_2_2(and_1083_nl, mux_tmp_171, or_475_cse);
  and_1084_nl <= nand_198_cse AND mux_tmp_172;
  mux_tmp_173 <= MUX_s_1_2_2(and_1084_nl, mux_tmp_172, or_468_cse);
  and_1085_nl <= nand_276_cse AND mux_tmp_173;
  mux_tmp_174 <= MUX_s_1_2_2(and_1085_nl, mux_tmp_173, or_463_cse);
  and_1086_nl <= nand_281_cse AND mux_tmp_174;
  mux_175_nl <= MUX_s_1_2_2(and_1086_nl, mux_tmp_174, or_458_cse);
  and_dcpl_508 <= mux_175_nl AND and_dcpl_121 AND and_dcpl_115;
  or_495_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01")) OR (rem_12cyc_st_6_3_2(1));
  and_1076_nl <= nand_215_cse AND or_tmp_446;
  mux_tmp_176 <= MUX_s_1_2_2(and_1076_nl, or_tmp_446, or_495_cse);
  and_1077_nl <= nand_189_cse AND mux_tmp_176;
  mux_tmp_177 <= MUX_s_1_2_2(and_1077_nl, mux_tmp_176, or_484_cse);
  and_1078_nl <= nand_271_cse AND mux_tmp_177;
  mux_tmp_178 <= MUX_s_1_2_2(and_1078_nl, mux_tmp_177, or_475_cse);
  and_1079_nl <= nand_198_cse AND mux_tmp_178;
  mux_tmp_179 <= MUX_s_1_2_2(and_1079_nl, mux_tmp_178, or_468_cse);
  and_1080_nl <= nand_276_cse AND mux_tmp_179;
  mux_tmp_180 <= MUX_s_1_2_2(and_1080_nl, mux_tmp_179, or_463_cse);
  and_1081_nl <= nand_281_cse AND mux_tmp_180;
  mux_181_nl <= MUX_s_1_2_2(and_1081_nl, mux_tmp_180, or_458_cse);
  and_dcpl_510 <= mux_181_nl AND and_dcpl_94 AND and_dcpl_87;
  or_508_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01")) OR (rem_12cyc_st_7_3_2(1));
  and_1069_nl <= nand_212_cse AND or_tmp_446;
  mux_tmp_182 <= MUX_s_1_2_2(and_1069_nl, or_tmp_446, or_508_cse);
  and_1070_nl <= nand_215_cse AND mux_tmp_182;
  mux_tmp_183 <= MUX_s_1_2_2(and_1070_nl, mux_tmp_182, or_495_cse);
  and_1071_nl <= nand_189_cse AND mux_tmp_183;
  mux_tmp_184 <= MUX_s_1_2_2(and_1071_nl, mux_tmp_183, or_484_cse);
  and_1072_nl <= nand_271_cse AND mux_tmp_184;
  mux_tmp_185 <= MUX_s_1_2_2(and_1072_nl, mux_tmp_184, or_475_cse);
  and_1073_nl <= nand_198_cse AND mux_tmp_185;
  mux_tmp_186 <= MUX_s_1_2_2(and_1073_nl, mux_tmp_185, or_468_cse);
  and_1074_nl <= nand_276_cse AND mux_tmp_186;
  mux_tmp_187 <= MUX_s_1_2_2(and_1074_nl, mux_tmp_186, or_463_cse);
  and_1075_nl <= nand_281_cse AND mux_tmp_187;
  mux_188_nl <= MUX_s_1_2_2(and_1075_nl, mux_tmp_187, or_458_cse);
  and_dcpl_512 <= mux_188_nl AND and_dcpl_67 AND and_dcpl_60;
  or_523_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01")) OR (rem_12cyc_st_8_3_2(1));
  and_1061_nl <= nand_208_cse AND or_tmp_446;
  mux_tmp_189 <= MUX_s_1_2_2(and_1061_nl, or_tmp_446, or_523_cse);
  and_1062_nl <= nand_212_cse AND mux_tmp_189;
  mux_tmp_190 <= MUX_s_1_2_2(and_1062_nl, mux_tmp_189, or_508_cse);
  and_1063_nl <= nand_215_cse AND mux_tmp_190;
  mux_tmp_191 <= MUX_s_1_2_2(and_1063_nl, mux_tmp_190, or_495_cse);
  and_1064_nl <= nand_189_cse AND mux_tmp_191;
  mux_tmp_192 <= MUX_s_1_2_2(and_1064_nl, mux_tmp_191, or_484_cse);
  and_1065_nl <= nand_271_cse AND mux_tmp_192;
  mux_tmp_193 <= MUX_s_1_2_2(and_1065_nl, mux_tmp_192, or_475_cse);
  and_1066_nl <= nand_198_cse AND mux_tmp_193;
  mux_tmp_194 <= MUX_s_1_2_2(and_1066_nl, mux_tmp_193, or_468_cse);
  and_1067_nl <= nand_276_cse AND mux_tmp_194;
  mux_tmp_195 <= MUX_s_1_2_2(and_1067_nl, mux_tmp_194, or_463_cse);
  and_1068_nl <= nand_281_cse AND mux_tmp_195;
  mux_196_nl <= MUX_s_1_2_2(and_1068_nl, mux_tmp_195, or_458_cse);
  and_dcpl_514 <= mux_196_nl AND and_dcpl_40 AND and_dcpl_33;
  and_1052_nl <= nand_203_cse AND or_tmp_446;
  or_540_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01")) OR (rem_12cyc_st_9_3_2(1));
  mux_tmp_197 <= MUX_s_1_2_2(and_1052_nl, or_tmp_446, or_540_nl);
  and_1053_nl <= nand_208_cse AND mux_tmp_197;
  mux_tmp_198 <= MUX_s_1_2_2(and_1053_nl, mux_tmp_197, or_523_cse);
  and_1054_nl <= nand_212_cse AND mux_tmp_198;
  mux_tmp_199 <= MUX_s_1_2_2(and_1054_nl, mux_tmp_198, or_508_cse);
  and_1055_nl <= nand_215_cse AND mux_tmp_199;
  mux_tmp_200 <= MUX_s_1_2_2(and_1055_nl, mux_tmp_199, or_495_cse);
  and_1056_nl <= nand_189_cse AND mux_tmp_200;
  mux_tmp_201 <= MUX_s_1_2_2(and_1056_nl, mux_tmp_200, or_484_cse);
  and_1057_nl <= nand_271_cse AND mux_tmp_201;
  mux_tmp_202 <= MUX_s_1_2_2(and_1057_nl, mux_tmp_201, or_475_cse);
  and_1058_nl <= nand_198_cse AND mux_tmp_202;
  mux_tmp_203 <= MUX_s_1_2_2(and_1058_nl, mux_tmp_202, or_468_cse);
  and_1059_nl <= nand_276_cse AND mux_tmp_203;
  mux_tmp_204 <= MUX_s_1_2_2(and_1059_nl, mux_tmp_203, or_463_cse);
  and_1060_nl <= nand_281_cse AND mux_tmp_204;
  mux_205_nl <= MUX_s_1_2_2(and_1060_nl, mux_tmp_204, or_458_cse);
  and_dcpl_516 <= mux_205_nl AND and_dcpl_13 AND and_dcpl_6;
  and_tmp_134 <= ((NOT main_stage_0_8) OR (NOT COMP_LOOP_asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_9)
      OR (NOT COMP_LOOP_asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_10)
      OR (NOT COMP_LOOP_asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_3)
      OR (NOT COMP_LOOP_asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_4)
      OR (NOT COMP_LOOP_asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_5)
      OR (NOT COMP_LOOP_asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_6)
      OR (NOT COMP_LOOP_asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_7)
      OR (NOT COMP_LOOP_asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_11)
      OR (NOT COMP_LOOP_asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("01"))) AND (CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("01"))
      OR (COMP_LOOP_acc_1_tmp(1)) OR nand_250_cse);
  nor_438_nl <= NOT((rem_12cyc_1_0(0)) OR (NOT and_tmp_134));
  or_550_nl <= (NOT main_stage_0_2) OR (NOT COMP_LOOP_asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_1_0(1));
  mux_tmp_206 <= MUX_s_1_2_2(nor_438_nl, and_tmp_134, or_550_nl);
  and_dcpl_520 <= and_dcpl_460 AND and_dcpl_393;
  and_dcpl_521 <= and_dcpl_462 AND (rem_12cyc_st_2_1_0(1));
  or_tmp_551 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10")) OR (rem_12cyc_3_2(1))
      OR not_tmp_332;
  or_564_cse <= CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (COMP_LOOP_acc_tmp(1));
  and_1170_nl <= nand_281_cse AND or_tmp_551;
  mux_207_nl <= MUX_s_1_2_2(and_1170_nl, or_tmp_551, or_564_cse);
  and_dcpl_523 <= mux_207_nl AND and_dcpl_298 AND and_dcpl_521;
  and_dcpl_524 <= and_dcpl_466 AND (rem_12cyc_st_3_1_0(1));
  or_569_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp_135 <= or_569_cse AND or_tmp_551;
  and_1050_nl <= nand_281_cse AND and_tmp_135;
  mux_208_nl <= MUX_s_1_2_2(and_1050_nl, and_tmp_135, or_564_cse);
  and_dcpl_526 <= mux_208_nl AND and_dcpl_304 AND and_dcpl_524;
  and_dcpl_527 <= and_dcpl_470 AND (rem_12cyc_st_4_1_0(1));
  or_573_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_137 <= or_569_cse AND or_573_cse AND or_tmp_551;
  and_1049_nl <= nand_281_cse AND and_tmp_137;
  mux_209_nl <= MUX_s_1_2_2(and_1049_nl, and_tmp_137, or_564_cse);
  and_dcpl_529 <= mux_209_nl AND and_dcpl_310 AND and_dcpl_527;
  and_dcpl_530 <= and_dcpl_474 AND (rem_12cyc_st_5_1_0(1));
  or_578_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_140 <= or_569_cse AND or_573_cse AND or_578_cse AND or_tmp_551;
  and_1048_nl <= nand_281_cse AND and_tmp_140;
  mux_210_nl <= MUX_s_1_2_2(and_1048_nl, and_tmp_140, or_564_cse);
  and_dcpl_532 <= mux_210_nl AND and_dcpl_316 AND and_dcpl_530;
  or_584_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_144 <= or_569_cse AND or_573_cse AND or_578_cse AND or_584_cse AND or_tmp_551;
  and_1047_nl <= nand_281_cse AND and_tmp_144;
  mux_211_nl <= MUX_s_1_2_2(and_1047_nl, and_tmp_144, or_564_cse);
  and_dcpl_534 <= mux_211_nl AND and_dcpl_121 AND and_dcpl_117;
  or_591_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10")) OR (rem_12cyc_st_6_3_2(1));
  and_1045_nl <= nand_215_cse AND or_tmp_551;
  mux_212_nl <= MUX_s_1_2_2(and_1045_nl, or_tmp_551, or_591_cse);
  and_tmp_148 <= or_569_cse AND or_573_cse AND or_578_cse AND or_584_cse AND mux_212_nl;
  and_1046_nl <= nand_281_cse AND and_tmp_148;
  mux_213_nl <= MUX_s_1_2_2(and_1046_nl, and_tmp_148, or_564_cse);
  and_dcpl_536 <= mux_213_nl AND and_dcpl_94 AND and_dcpl_90;
  or_600_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10")) OR (rem_12cyc_st_7_3_2(1));
  and_1042_nl <= nand_212_cse AND or_tmp_551;
  mux_tmp_214 <= MUX_s_1_2_2(and_1042_nl, or_tmp_551, or_600_cse);
  and_1043_nl <= nand_215_cse AND mux_tmp_214;
  mux_215_nl <= MUX_s_1_2_2(and_1043_nl, mux_tmp_214, or_591_cse);
  and_tmp_152 <= or_569_cse AND or_573_cse AND or_578_cse AND or_584_cse AND mux_215_nl;
  and_1044_nl <= nand_281_cse AND and_tmp_152;
  mux_216_nl <= MUX_s_1_2_2(and_1044_nl, and_tmp_152, or_564_cse);
  and_dcpl_538 <= mux_216_nl AND and_dcpl_67 AND and_dcpl_63;
  or_611_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10")) OR (rem_12cyc_st_8_3_2(1));
  and_1038_nl <= nand_208_cse AND or_tmp_551;
  mux_tmp_217 <= MUX_s_1_2_2(and_1038_nl, or_tmp_551, or_611_cse);
  and_1039_nl <= nand_212_cse AND mux_tmp_217;
  mux_tmp_218 <= MUX_s_1_2_2(and_1039_nl, mux_tmp_217, or_600_cse);
  and_1040_nl <= nand_215_cse AND mux_tmp_218;
  mux_219_nl <= MUX_s_1_2_2(and_1040_nl, mux_tmp_218, or_591_cse);
  and_tmp_156 <= or_569_cse AND or_573_cse AND or_578_cse AND or_584_cse AND mux_219_nl;
  and_1041_nl <= nand_281_cse AND and_tmp_156;
  mux_220_nl <= MUX_s_1_2_2(and_1041_nl, and_tmp_156, or_564_cse);
  and_dcpl_540 <= mux_220_nl AND and_dcpl_40 AND and_dcpl_36;
  and_1033_nl <= nand_203_cse AND or_tmp_551;
  or_624_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10")) OR (rem_12cyc_st_9_3_2(1));
  mux_tmp_221 <= MUX_s_1_2_2(and_1033_nl, or_tmp_551, or_624_nl);
  and_1034_nl <= nand_208_cse AND mux_tmp_221;
  mux_tmp_222 <= MUX_s_1_2_2(and_1034_nl, mux_tmp_221, or_611_cse);
  and_1035_nl <= nand_212_cse AND mux_tmp_222;
  mux_tmp_223 <= MUX_s_1_2_2(and_1035_nl, mux_tmp_222, or_600_cse);
  and_1036_nl <= nand_215_cse AND mux_tmp_223;
  mux_224_nl <= MUX_s_1_2_2(and_1036_nl, mux_tmp_223, or_591_cse);
  and_tmp_160 <= or_569_cse AND or_573_cse AND or_578_cse AND or_584_cse AND mux_224_nl;
  and_1037_nl <= nand_281_cse AND and_tmp_160;
  mux_225_nl <= MUX_s_1_2_2(and_1037_nl, and_tmp_160, or_564_cse);
  and_dcpl_542 <= mux_225_nl AND and_dcpl_13 AND and_dcpl_9;
  and_tmp_170 <= ((NOT main_stage_0_2) OR (NOT COMP_LOOP_asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10"))) AND ((NOT main_stage_0_8)
      OR (NOT COMP_LOOP_asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_9)
      OR (NOT COMP_LOOP_asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_10)
      OR (NOT COMP_LOOP_asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("01"))) AND or_569_cse
      AND or_573_cse AND or_578_cse AND or_584_cse AND ((NOT main_stage_0_7) OR (NOT
      COMP_LOOP_asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_11)
      OR (NOT COMP_LOOP_asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("01"))) AND (CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT ccs_ccore_start_rsci_idat));
  and_dcpl_546 <= and_dcpl_460 AND and_dcpl_430;
  or_tmp_629 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("11")) OR (rem_12cyc_3_2(1))
      OR not_tmp_332;
  or_643_cse <= CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (COMP_LOOP_acc_tmp(1));
  and_1169_nl <= nand_281_cse AND or_tmp_629;
  mux_226_nl <= MUX_s_1_2_2(and_1169_nl, or_tmp_629, or_643_cse);
  and_dcpl_548 <= mux_226_nl AND and_dcpl_358 AND and_dcpl_521;
  or_648_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("01"));
  and_1030_nl <= nand_276_cse AND or_tmp_629;
  mux_tmp_227 <= MUX_s_1_2_2(and_1030_nl, or_tmp_629, or_648_cse);
  and_1031_nl <= nand_281_cse AND mux_tmp_227;
  mux_228_nl <= MUX_s_1_2_2(and_1031_nl, mux_tmp_227, or_643_cse);
  and_dcpl_550 <= mux_228_nl AND and_dcpl_362 AND and_dcpl_524;
  or_653_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR (rem_12cyc_st_3_3_2(1));
  and_1027_nl <= nand_198_cse AND or_tmp_629;
  mux_tmp_229 <= MUX_s_1_2_2(and_1027_nl, or_tmp_629, or_653_cse);
  and_1028_nl <= nand_276_cse AND mux_tmp_229;
  mux_tmp_230 <= MUX_s_1_2_2(and_1028_nl, mux_tmp_229, or_648_cse);
  and_1029_nl <= nand_281_cse AND mux_tmp_230;
  mux_231_nl <= MUX_s_1_2_2(and_1029_nl, mux_tmp_230, or_643_cse);
  and_dcpl_552 <= mux_231_nl AND and_dcpl_366 AND and_dcpl_527;
  or_660_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("01"));
  and_1023_nl <= nand_271_cse AND or_tmp_629;
  mux_tmp_232 <= MUX_s_1_2_2(and_1023_nl, or_tmp_629, or_660_cse);
  and_1024_nl <= nand_198_cse AND mux_tmp_232;
  mux_tmp_233 <= MUX_s_1_2_2(and_1024_nl, mux_tmp_232, or_653_cse);
  and_1025_nl <= nand_276_cse AND mux_tmp_233;
  mux_tmp_234 <= MUX_s_1_2_2(and_1025_nl, mux_tmp_233, or_648_cse);
  and_1026_nl <= nand_281_cse AND mux_tmp_234;
  mux_235_nl <= MUX_s_1_2_2(and_1026_nl, mux_tmp_234, or_643_cse);
  and_dcpl_554 <= mux_235_nl AND and_dcpl_370 AND and_dcpl_530;
  or_669_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR (rem_12cyc_st_5_3_2(1));
  and_1018_nl <= nand_189_cse AND or_tmp_629;
  mux_tmp_236 <= MUX_s_1_2_2(and_1018_nl, or_tmp_629, or_669_cse);
  and_1019_nl <= nand_271_cse AND mux_tmp_236;
  mux_tmp_237 <= MUX_s_1_2_2(and_1019_nl, mux_tmp_236, or_660_cse);
  and_1020_nl <= nand_198_cse AND mux_tmp_237;
  mux_tmp_238 <= MUX_s_1_2_2(and_1020_nl, mux_tmp_237, or_653_cse);
  and_1021_nl <= nand_276_cse AND mux_tmp_238;
  mux_tmp_239 <= MUX_s_1_2_2(and_1021_nl, mux_tmp_238, or_648_cse);
  and_1022_nl <= nand_281_cse AND mux_tmp_239;
  mux_240_nl <= MUX_s_1_2_2(and_1022_nl, mux_tmp_239, or_643_cse);
  and_dcpl_556 <= mux_240_nl AND and_dcpl_121 AND and_dcpl_119;
  or_680_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("11")) OR (rem_12cyc_st_6_3_2(1));
  and_1012_nl <= nand_215_cse AND or_tmp_629;
  mux_tmp_241 <= MUX_s_1_2_2(and_1012_nl, or_tmp_629, or_680_cse);
  and_1013_nl <= nand_189_cse AND mux_tmp_241;
  mux_tmp_242 <= MUX_s_1_2_2(and_1013_nl, mux_tmp_241, or_669_cse);
  and_1014_nl <= nand_271_cse AND mux_tmp_242;
  mux_tmp_243 <= MUX_s_1_2_2(and_1014_nl, mux_tmp_242, or_660_cse);
  and_1015_nl <= nand_198_cse AND mux_tmp_243;
  mux_tmp_244 <= MUX_s_1_2_2(and_1015_nl, mux_tmp_243, or_653_cse);
  and_1016_nl <= nand_276_cse AND mux_tmp_244;
  mux_tmp_245 <= MUX_s_1_2_2(and_1016_nl, mux_tmp_244, or_648_cse);
  and_1017_nl <= nand_281_cse AND mux_tmp_245;
  mux_246_nl <= MUX_s_1_2_2(and_1017_nl, mux_tmp_245, or_643_cse);
  and_dcpl_558 <= mux_246_nl AND and_dcpl_94 AND and_dcpl_92;
  or_693_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("11")) OR (rem_12cyc_st_7_3_2(1));
  and_1005_nl <= nand_212_cse AND or_tmp_629;
  mux_tmp_247 <= MUX_s_1_2_2(and_1005_nl, or_tmp_629, or_693_cse);
  and_1006_nl <= nand_215_cse AND mux_tmp_247;
  mux_tmp_248 <= MUX_s_1_2_2(and_1006_nl, mux_tmp_247, or_680_cse);
  and_1007_nl <= nand_189_cse AND mux_tmp_248;
  mux_tmp_249 <= MUX_s_1_2_2(and_1007_nl, mux_tmp_248, or_669_cse);
  and_1008_nl <= nand_271_cse AND mux_tmp_249;
  mux_tmp_250 <= MUX_s_1_2_2(and_1008_nl, mux_tmp_249, or_660_cse);
  and_1009_nl <= nand_198_cse AND mux_tmp_250;
  mux_tmp_251 <= MUX_s_1_2_2(and_1009_nl, mux_tmp_250, or_653_cse);
  and_1010_nl <= nand_276_cse AND mux_tmp_251;
  mux_tmp_252 <= MUX_s_1_2_2(and_1010_nl, mux_tmp_251, or_648_cse);
  and_1011_nl <= nand_281_cse AND mux_tmp_252;
  mux_253_nl <= MUX_s_1_2_2(and_1011_nl, mux_tmp_252, or_643_cse);
  and_dcpl_560 <= mux_253_nl AND and_dcpl_67 AND and_dcpl_65;
  or_708_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("11")) OR (rem_12cyc_st_8_3_2(1));
  and_997_nl <= nand_208_cse AND or_tmp_629;
  mux_tmp_254 <= MUX_s_1_2_2(and_997_nl, or_tmp_629, or_708_cse);
  and_998_nl <= nand_212_cse AND mux_tmp_254;
  mux_tmp_255 <= MUX_s_1_2_2(and_998_nl, mux_tmp_254, or_693_cse);
  and_999_nl <= nand_215_cse AND mux_tmp_255;
  mux_tmp_256 <= MUX_s_1_2_2(and_999_nl, mux_tmp_255, or_680_cse);
  and_1000_nl <= nand_189_cse AND mux_tmp_256;
  mux_tmp_257 <= MUX_s_1_2_2(and_1000_nl, mux_tmp_256, or_669_cse);
  and_1001_nl <= nand_271_cse AND mux_tmp_257;
  mux_tmp_258 <= MUX_s_1_2_2(and_1001_nl, mux_tmp_257, or_660_cse);
  and_1002_nl <= nand_198_cse AND mux_tmp_258;
  mux_tmp_259 <= MUX_s_1_2_2(and_1002_nl, mux_tmp_258, or_653_cse);
  and_1003_nl <= nand_276_cse AND mux_tmp_259;
  mux_tmp_260 <= MUX_s_1_2_2(and_1003_nl, mux_tmp_259, or_648_cse);
  and_1004_nl <= nand_281_cse AND mux_tmp_260;
  mux_261_nl <= MUX_s_1_2_2(and_1004_nl, mux_tmp_260, or_643_cse);
  and_dcpl_562 <= mux_261_nl AND and_dcpl_40 AND and_dcpl_38;
  and_988_nl <= nand_203_cse AND or_tmp_629;
  or_725_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("11")) OR (rem_12cyc_st_9_3_2(1));
  mux_tmp_262 <= MUX_s_1_2_2(and_988_nl, or_tmp_629, or_725_nl);
  and_989_nl <= nand_208_cse AND mux_tmp_262;
  mux_tmp_263 <= MUX_s_1_2_2(and_989_nl, mux_tmp_262, or_708_cse);
  and_990_nl <= nand_212_cse AND mux_tmp_263;
  mux_tmp_264 <= MUX_s_1_2_2(and_990_nl, mux_tmp_263, or_693_cse);
  and_991_nl <= nand_215_cse AND mux_tmp_264;
  mux_tmp_265 <= MUX_s_1_2_2(and_991_nl, mux_tmp_264, or_680_cse);
  and_992_nl <= nand_189_cse AND mux_tmp_265;
  mux_tmp_266 <= MUX_s_1_2_2(and_992_nl, mux_tmp_265, or_669_cse);
  and_993_nl <= nand_271_cse AND mux_tmp_266;
  mux_tmp_267 <= MUX_s_1_2_2(and_993_nl, mux_tmp_266, or_660_cse);
  and_994_nl <= nand_198_cse AND mux_tmp_267;
  mux_tmp_268 <= MUX_s_1_2_2(and_994_nl, mux_tmp_267, or_653_cse);
  and_995_nl <= nand_276_cse AND mux_tmp_268;
  mux_tmp_269 <= MUX_s_1_2_2(and_995_nl, mux_tmp_268, or_648_cse);
  and_996_nl <= nand_281_cse AND mux_tmp_269;
  mux_270_nl <= MUX_s_1_2_2(and_996_nl, mux_tmp_269, or_643_cse);
  and_dcpl_564 <= mux_270_nl AND and_dcpl_13 AND and_dcpl_11;
  and_tmp_179 <= (NOT(main_stage_0_8 AND COMP_LOOP_asn_itm_7 AND CONV_SL_1_1(rem_12cyc_st_7_1_0=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(rem_12cyc_st_7_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_9
      AND COMP_LOOP_asn_itm_8 AND CONV_SL_1_1(rem_12cyc_st_8_1_0=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(rem_12cyc_st_8_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_10
      AND COMP_LOOP_asn_itm_9 AND CONV_SL_1_1(rem_12cyc_st_9_1_0=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(rem_12cyc_st_9_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_3
      AND COMP_LOOP_asn_itm_2 AND CONV_SL_1_1(rem_12cyc_st_2_1_0=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(rem_12cyc_st_2_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_4
      AND COMP_LOOP_asn_itm_3 AND CONV_SL_1_1(rem_12cyc_st_3_1_0=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(rem_12cyc_st_3_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_5
      AND COMP_LOOP_asn_itm_4 AND CONV_SL_1_1(rem_12cyc_st_4_1_0=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(rem_12cyc_st_4_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_6
      AND COMP_LOOP_asn_itm_5 AND CONV_SL_1_1(rem_12cyc_st_5_1_0=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(rem_12cyc_st_5_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_7
      AND COMP_LOOP_asn_itm_6 AND CONV_SL_1_1(rem_12cyc_st_6_1_0=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(rem_12cyc_st_6_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_11
      AND COMP_LOOP_asn_itm_10 AND CONV_SL_1_1(rem_12cyc_st_10_1_0=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(rem_12cyc_st_10_3_2=STD_LOGIC_VECTOR'("01")))) AND ((COMP_LOOP_acc_tmp(1))
      OR (NOT((COMP_LOOP_acc_tmp(0)) AND CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO
      0)=STD_LOGIC_VECTOR'("11")) AND ccs_ccore_start_rsci_idat)));
  and_987_nl <= (NOT((rem_12cyc_3_2(0)) AND CONV_SL_1_1(rem_12cyc_1_0=STD_LOGIC_VECTOR'("11"))))
      AND and_tmp_179;
  or_735_nl <= (NOT main_stage_0_2) OR (NOT COMP_LOOP_asn_itm_1) OR (rem_12cyc_3_2(1));
  mux_tmp_271 <= MUX_s_1_2_2(and_987_nl, and_tmp_179, or_735_nl);
  and_dcpl_568 <= and_dcpl_292 AND (COMP_LOOP_acc_tmp(1));
  and_dcpl_569 <= and_dcpl_568 AND and_dcpl_291;
  and_dcpl_570 <= CONV_SL_1_1(rem_12cyc_st_2_3_2=STD_LOGIC_VECTOR'("10"));
  and_dcpl_571 <= and_dcpl_570 AND (NOT (rem_12cyc_st_2_1_0(1)));
  or_tmp_733 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR not_tmp_54;
  or_748_cse <= CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("10"));
  nor_435_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_733));
  mux_272_nl <= MUX_s_1_2_2(nor_435_nl, or_tmp_733, or_748_cse);
  and_dcpl_573 <= mux_272_nl AND and_dcpl_298 AND and_dcpl_571;
  and_dcpl_574 <= CONV_SL_1_1(rem_12cyc_st_3_3_2=STD_LOGIC_VECTOR'("10"));
  and_dcpl_575 <= and_dcpl_574 AND (NOT (rem_12cyc_st_3_1_0(1)));
  or_753_cse <= (rem_12cyc_st_2_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp_180 <= or_753_cse AND or_tmp_733;
  nor_434_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_180));
  mux_273_nl <= MUX_s_1_2_2(nor_434_nl, and_tmp_180, or_748_cse);
  and_dcpl_577 <= mux_273_nl AND and_dcpl_304 AND and_dcpl_575;
  and_dcpl_578 <= CONV_SL_1_1(rem_12cyc_st_4_3_2=STD_LOGIC_VECTOR'("10"));
  and_dcpl_579 <= and_dcpl_578 AND (NOT (rem_12cyc_st_4_1_0(1)));
  or_757_cse <= (rem_12cyc_st_3_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_182 <= or_753_cse AND or_757_cse AND or_tmp_733;
  nor_433_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_182));
  mux_274_nl <= MUX_s_1_2_2(nor_433_nl, and_tmp_182, or_748_cse);
  and_dcpl_581 <= mux_274_nl AND and_dcpl_310 AND and_dcpl_579;
  and_dcpl_582 <= CONV_SL_1_1(rem_12cyc_st_5_3_2=STD_LOGIC_VECTOR'("10"));
  and_dcpl_583 <= and_dcpl_582 AND (NOT (rem_12cyc_st_5_1_0(1)));
  or_762_cse <= (rem_12cyc_st_4_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_185 <= or_753_cse AND or_757_cse AND or_762_cse AND or_tmp_733;
  nor_432_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_185));
  mux_275_nl <= MUX_s_1_2_2(nor_432_nl, and_tmp_185, or_748_cse);
  and_dcpl_585 <= mux_275_nl AND and_dcpl_316 AND and_dcpl_583;
  or_768_cse <= (rem_12cyc_st_5_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_189 <= or_753_cse AND or_757_cse AND or_762_cse AND or_768_cse AND or_tmp_733;
  nor_431_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_189));
  mux_276_nl <= MUX_s_1_2_2(nor_431_nl, and_tmp_189, or_748_cse);
  and_dcpl_589 <= mux_276_nl AND and_dcpl_112 AND and_dcpl_126 AND (NOT (rem_12cyc_st_6_1_0(1)));
  or_775_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_429_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_733));
  mux_277_nl <= MUX_s_1_2_2(nor_429_nl, or_tmp_733, or_775_cse);
  and_tmp_193 <= or_753_cse AND or_757_cse AND or_762_cse AND or_768_cse AND mux_277_nl;
  nor_430_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_193));
  mux_278_nl <= MUX_s_1_2_2(nor_430_nl, and_tmp_193, or_748_cse);
  and_dcpl_593 <= mux_278_nl AND and_dcpl_85 AND and_dcpl_99 AND (NOT (rem_12cyc_st_7_1_0(0)));
  or_784_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_426_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_733));
  mux_tmp_279 <= MUX_s_1_2_2(nor_426_nl, or_tmp_733, or_784_cse);
  nor_427_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_279));
  mux_280_nl <= MUX_s_1_2_2(nor_427_nl, mux_tmp_279, or_775_cse);
  and_tmp_197 <= or_753_cse AND or_757_cse AND or_762_cse AND or_768_cse AND mux_280_nl;
  nor_428_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_197));
  mux_281_nl <= MUX_s_1_2_2(nor_428_nl, and_tmp_197, or_748_cse);
  and_dcpl_597 <= mux_281_nl AND and_dcpl_58 AND and_dcpl_72 AND (NOT (rem_12cyc_st_8_1_0(0)));
  or_795_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_422_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_733));
  mux_tmp_282 <= MUX_s_1_2_2(nor_422_nl, or_tmp_733, or_795_cse);
  nor_423_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_282));
  mux_tmp_283 <= MUX_s_1_2_2(nor_423_nl, mux_tmp_282, or_784_cse);
  nor_424_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_283));
  mux_284_nl <= MUX_s_1_2_2(nor_424_nl, mux_tmp_283, or_775_cse);
  and_tmp_201 <= or_753_cse AND or_757_cse AND or_762_cse AND or_768_cse AND mux_284_nl;
  nor_425_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_201));
  mux_285_nl <= MUX_s_1_2_2(nor_425_nl, and_tmp_201, or_748_cse);
  and_dcpl_601 <= mux_285_nl AND and_dcpl_31 AND and_dcpl_45 AND (NOT (rem_12cyc_st_9_1_0(0)));
  nor_417_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_733));
  or_808_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("10"));
  mux_tmp_286 <= MUX_s_1_2_2(nor_417_nl, or_tmp_733, or_808_nl);
  nor_418_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_286));
  mux_tmp_287 <= MUX_s_1_2_2(nor_418_nl, mux_tmp_286, or_795_cse);
  nor_419_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_287));
  mux_tmp_288 <= MUX_s_1_2_2(nor_419_nl, mux_tmp_287, or_784_cse);
  nor_420_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_288));
  mux_289_nl <= MUX_s_1_2_2(nor_420_nl, mux_tmp_288, or_775_cse);
  and_tmp_205 <= or_753_cse AND or_757_cse AND or_762_cse AND or_768_cse AND mux_289_nl;
  nor_421_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_205));
  mux_290_nl <= MUX_s_1_2_2(nor_421_nl, and_tmp_205, or_748_cse);
  and_dcpl_605 <= mux_290_nl AND and_dcpl_4 AND and_dcpl_18 AND (NOT (rem_12cyc_st_10_1_0(0)));
  or_tmp_808 <= CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT ccs_ccore_start_rsci_idat);
  nor_408_nl <= NOT((rem_12cyc_st_10_3_2(1)) OR (NOT or_tmp_808));
  or_823_nl <= (NOT main_stage_0_11) OR (NOT COMP_LOOP_asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_10_3_2(0));
  mux_tmp_291 <= MUX_s_1_2_2(nor_408_nl, or_tmp_808, or_823_nl);
  nor_409_nl <= NOT((rem_12cyc_st_6_3_2(1)) OR (NOT mux_tmp_291));
  or_822_nl <= (NOT main_stage_0_7) OR (NOT COMP_LOOP_asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_6_3_2(0));
  mux_tmp_292 <= MUX_s_1_2_2(nor_409_nl, mux_tmp_291, or_822_nl);
  nor_410_nl <= NOT((rem_12cyc_st_5_3_2(1)) OR (NOT mux_tmp_292));
  or_821_nl <= (NOT main_stage_0_6) OR (NOT COMP_LOOP_asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_5_3_2(0));
  mux_tmp_293 <= MUX_s_1_2_2(nor_410_nl, mux_tmp_292, or_821_nl);
  nor_411_nl <= NOT((rem_12cyc_st_4_3_2(1)) OR (NOT mux_tmp_293));
  or_820_nl <= (NOT main_stage_0_5) OR (NOT COMP_LOOP_asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_4_3_2(0));
  mux_tmp_294 <= MUX_s_1_2_2(nor_411_nl, mux_tmp_293, or_820_nl);
  nor_412_nl <= NOT((rem_12cyc_st_3_3_2(1)) OR (NOT mux_tmp_294));
  or_819_nl <= (NOT main_stage_0_4) OR (NOT COMP_LOOP_asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_3_3_2(0));
  mux_tmp_295 <= MUX_s_1_2_2(nor_412_nl, mux_tmp_294, or_819_nl);
  nor_413_nl <= NOT((rem_12cyc_st_2_3_2(1)) OR (NOT mux_tmp_295));
  or_818_nl <= (NOT main_stage_0_3) OR (NOT COMP_LOOP_asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_2_3_2(0));
  mux_tmp_296 <= MUX_s_1_2_2(nor_413_nl, mux_tmp_295, or_818_nl);
  nor_414_nl <= NOT((rem_12cyc_st_9_3_2(1)) OR (NOT mux_tmp_296));
  or_817_nl <= (NOT main_stage_0_10) OR (NOT COMP_LOOP_asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_9_3_2(0));
  mux_tmp_297 <= MUX_s_1_2_2(nor_414_nl, mux_tmp_296, or_817_nl);
  nor_415_nl <= NOT((rem_12cyc_st_8_3_2(1)) OR (NOT mux_tmp_297));
  or_816_nl <= (NOT main_stage_0_9) OR (NOT COMP_LOOP_asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_8_3_2(0));
  mux_tmp_298 <= MUX_s_1_2_2(nor_415_nl, mux_tmp_297, or_816_nl);
  nor_416_nl <= NOT((rem_12cyc_st_7_3_2(1)) OR (NOT mux_tmp_298));
  or_815_nl <= (NOT main_stage_0_8) OR (NOT COMP_LOOP_asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_7_3_2(0));
  mux_299_nl <= MUX_s_1_2_2(nor_416_nl, mux_tmp_298, or_815_nl);
  and_tmp_206 <= ((NOT main_stage_0_2) OR (NOT COMP_LOOP_asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00"))) AND mux_299_nl;
  and_dcpl_610 <= and_dcpl_568 AND and_dcpl_355;
  or_tmp_820 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR not_tmp_54;
  or_837_cse <= CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("10"));
  nor_407_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_820));
  mux_300_nl <= MUX_s_1_2_2(nor_407_nl, or_tmp_820, or_837_cse);
  and_dcpl_612 <= mux_300_nl AND and_dcpl_358 AND and_dcpl_571;
  nand_84_cse <= NOT((rem_12cyc_st_2_3_2(1)) AND COMP_LOOP_asn_itm_2 AND main_stage_0_3
      AND (rem_12cyc_st_2_1_0(0)));
  or_842_cse <= (rem_12cyc_st_2_1_0(1)) OR (rem_12cyc_st_2_3_2(0));
  and_986_nl <= nand_84_cse AND or_tmp_820;
  mux_tmp_301 <= MUX_s_1_2_2(and_986_nl, or_tmp_820, or_842_cse);
  nor_406_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_301));
  mux_302_nl <= MUX_s_1_2_2(nor_406_nl, mux_tmp_301, or_837_cse);
  and_dcpl_614 <= mux_302_nl AND and_dcpl_362 AND and_dcpl_575;
  or_847_cse <= (rem_12cyc_st_3_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("10"));
  and_984_nl <= nand_274_cse AND or_tmp_820;
  mux_tmp_303 <= MUX_s_1_2_2(and_984_nl, or_tmp_820, or_847_cse);
  and_985_nl <= nand_84_cse AND mux_tmp_303;
  mux_tmp_304 <= MUX_s_1_2_2(and_985_nl, mux_tmp_303, or_842_cse);
  nor_405_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_304));
  mux_305_nl <= MUX_s_1_2_2(nor_405_nl, mux_tmp_304, or_837_cse);
  and_dcpl_616 <= mux_305_nl AND and_dcpl_366 AND and_dcpl_579;
  nand_79_cse <= NOT((rem_12cyc_st_4_3_2(1)) AND COMP_LOOP_asn_itm_4 AND main_stage_0_5
      AND (rem_12cyc_st_4_1_0(0)));
  or_854_cse <= (rem_12cyc_st_4_1_0(1)) OR (rem_12cyc_st_4_3_2(0));
  and_981_nl <= nand_79_cse AND or_tmp_820;
  mux_tmp_306 <= MUX_s_1_2_2(and_981_nl, or_tmp_820, or_854_cse);
  and_982_nl <= nand_274_cse AND mux_tmp_306;
  mux_tmp_307 <= MUX_s_1_2_2(and_982_nl, mux_tmp_306, or_847_cse);
  and_983_nl <= nand_84_cse AND mux_tmp_307;
  mux_tmp_308 <= MUX_s_1_2_2(and_983_nl, mux_tmp_307, or_842_cse);
  nor_404_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_308));
  mux_309_nl <= MUX_s_1_2_2(nor_404_nl, mux_tmp_308, or_837_cse);
  and_dcpl_618 <= mux_309_nl AND and_dcpl_370 AND and_dcpl_583;
  or_863_cse <= (rem_12cyc_st_5_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("10"));
  and_977_nl <= nand_267_cse AND or_tmp_820;
  mux_tmp_310 <= MUX_s_1_2_2(and_977_nl, or_tmp_820, or_863_cse);
  and_978_nl <= nand_79_cse AND mux_tmp_310;
  mux_tmp_311 <= MUX_s_1_2_2(and_978_nl, mux_tmp_310, or_854_cse);
  and_979_nl <= nand_274_cse AND mux_tmp_311;
  mux_tmp_312 <= MUX_s_1_2_2(and_979_nl, mux_tmp_311, or_847_cse);
  and_980_nl <= nand_84_cse AND mux_tmp_312;
  mux_tmp_313 <= MUX_s_1_2_2(and_980_nl, mux_tmp_312, or_842_cse);
  nor_403_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_313));
  mux_314_nl <= MUX_s_1_2_2(nor_403_nl, mux_tmp_313, or_837_cse);
  and_dcpl_622 <= mux_314_nl AND and_dcpl_112 AND and_dcpl_129 AND (NOT (rem_12cyc_st_6_1_0(1)));
  or_874_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_401_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_820));
  mux_tmp_315 <= MUX_s_1_2_2(nor_401_nl, or_tmp_820, or_874_cse);
  and_973_nl <= nand_267_cse AND mux_tmp_315;
  mux_tmp_316 <= MUX_s_1_2_2(and_973_nl, mux_tmp_315, or_863_cse);
  and_974_nl <= nand_79_cse AND mux_tmp_316;
  mux_tmp_317 <= MUX_s_1_2_2(and_974_nl, mux_tmp_316, or_854_cse);
  and_975_nl <= nand_274_cse AND mux_tmp_317;
  mux_tmp_318 <= MUX_s_1_2_2(and_975_nl, mux_tmp_317, or_847_cse);
  and_976_nl <= nand_84_cse AND mux_tmp_318;
  mux_tmp_319 <= MUX_s_1_2_2(and_976_nl, mux_tmp_318, or_842_cse);
  nor_402_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_319));
  mux_320_nl <= MUX_s_1_2_2(nor_402_nl, mux_tmp_319, or_837_cse);
  and_dcpl_625 <= mux_320_nl AND and_dcpl_85 AND and_dcpl_99 AND (rem_12cyc_st_7_1_0(0));
  or_887_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_398_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_820));
  mux_tmp_321 <= MUX_s_1_2_2(nor_398_nl, or_tmp_820, or_887_cse);
  nor_399_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_321));
  mux_tmp_322 <= MUX_s_1_2_2(nor_399_nl, mux_tmp_321, or_874_cse);
  and_969_nl <= nand_267_cse AND mux_tmp_322;
  mux_tmp_323 <= MUX_s_1_2_2(and_969_nl, mux_tmp_322, or_863_cse);
  and_970_nl <= nand_79_cse AND mux_tmp_323;
  mux_tmp_324 <= MUX_s_1_2_2(and_970_nl, mux_tmp_323, or_854_cse);
  and_971_nl <= nand_274_cse AND mux_tmp_324;
  mux_tmp_325 <= MUX_s_1_2_2(and_971_nl, mux_tmp_324, or_847_cse);
  and_972_nl <= nand_84_cse AND mux_tmp_325;
  mux_tmp_326 <= MUX_s_1_2_2(and_972_nl, mux_tmp_325, or_842_cse);
  nor_400_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_326));
  mux_327_nl <= MUX_s_1_2_2(nor_400_nl, mux_tmp_326, or_837_cse);
  and_dcpl_628 <= mux_327_nl AND and_dcpl_58 AND and_dcpl_72 AND (rem_12cyc_st_8_1_0(0));
  or_902_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_394_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_820));
  mux_tmp_328 <= MUX_s_1_2_2(nor_394_nl, or_tmp_820, or_902_cse);
  nor_395_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_328));
  mux_tmp_329 <= MUX_s_1_2_2(nor_395_nl, mux_tmp_328, or_887_cse);
  nor_396_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_329));
  mux_tmp_330 <= MUX_s_1_2_2(nor_396_nl, mux_tmp_329, or_874_cse);
  and_965_nl <= nand_267_cse AND mux_tmp_330;
  mux_tmp_331 <= MUX_s_1_2_2(and_965_nl, mux_tmp_330, or_863_cse);
  and_966_nl <= nand_79_cse AND mux_tmp_331;
  mux_tmp_332 <= MUX_s_1_2_2(and_966_nl, mux_tmp_331, or_854_cse);
  and_967_nl <= nand_274_cse AND mux_tmp_332;
  mux_tmp_333 <= MUX_s_1_2_2(and_967_nl, mux_tmp_332, or_847_cse);
  and_968_nl <= nand_84_cse AND mux_tmp_333;
  mux_tmp_334 <= MUX_s_1_2_2(and_968_nl, mux_tmp_333, or_842_cse);
  nor_397_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_334));
  mux_335_nl <= MUX_s_1_2_2(nor_397_nl, mux_tmp_334, or_837_cse);
  and_dcpl_631 <= mux_335_nl AND and_dcpl_31 AND and_dcpl_45 AND (rem_12cyc_st_9_1_0(0));
  nor_389_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_820));
  or_919_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("10"));
  mux_tmp_336 <= MUX_s_1_2_2(nor_389_nl, or_tmp_820, or_919_nl);
  nor_390_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_336));
  mux_tmp_337 <= MUX_s_1_2_2(nor_390_nl, mux_tmp_336, or_902_cse);
  nor_391_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_337));
  mux_tmp_338 <= MUX_s_1_2_2(nor_391_nl, mux_tmp_337, or_887_cse);
  nor_392_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_338));
  mux_tmp_339 <= MUX_s_1_2_2(nor_392_nl, mux_tmp_338, or_874_cse);
  and_961_nl <= nand_267_cse AND mux_tmp_339;
  mux_tmp_340 <= MUX_s_1_2_2(and_961_nl, mux_tmp_339, or_863_cse);
  and_962_nl <= nand_79_cse AND mux_tmp_340;
  mux_tmp_341 <= MUX_s_1_2_2(and_962_nl, mux_tmp_340, or_854_cse);
  and_963_nl <= nand_274_cse AND mux_tmp_341;
  mux_tmp_342 <= MUX_s_1_2_2(and_963_nl, mux_tmp_341, or_847_cse);
  and_964_nl <= nand_84_cse AND mux_tmp_342;
  mux_tmp_343 <= MUX_s_1_2_2(and_964_nl, mux_tmp_342, or_842_cse);
  nor_393_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_343));
  mux_344_nl <= MUX_s_1_2_2(nor_393_nl, mux_tmp_343, or_837_cse);
  and_dcpl_634 <= mux_344_nl AND and_dcpl_4 AND and_dcpl_18 AND (rem_12cyc_st_10_1_0(0));
  or_tmp_921 <= CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("10")) OR (COMP_LOOP_acc_1_tmp(1))
      OR nand_250_cse;
  nor_379_nl <= NOT((rem_12cyc_st_10_3_2(1)) OR (NOT or_tmp_921));
  or_938_nl <= (NOT main_stage_0_11) OR (NOT COMP_LOOP_asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_10_3_2(0));
  mux_tmp_345 <= MUX_s_1_2_2(nor_379_nl, or_tmp_921, or_938_nl);
  nor_380_nl <= NOT((rem_12cyc_st_6_3_2(1)) OR (NOT mux_tmp_345));
  or_937_nl <= (NOT main_stage_0_7) OR (NOT COMP_LOOP_asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_6_3_2(0));
  mux_tmp_346 <= MUX_s_1_2_2(nor_380_nl, mux_tmp_345, or_937_nl);
  nor_381_nl <= NOT((rem_12cyc_st_5_3_2(1)) OR (NOT mux_tmp_346));
  or_936_nl <= (NOT main_stage_0_6) OR (NOT COMP_LOOP_asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_5_3_2(0));
  mux_tmp_347 <= MUX_s_1_2_2(nor_381_nl, mux_tmp_346, or_936_nl);
  nor_382_nl <= NOT((rem_12cyc_st_4_3_2(1)) OR (NOT mux_tmp_347));
  or_935_nl <= (NOT main_stage_0_5) OR (NOT COMP_LOOP_asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_4_3_2(0));
  mux_tmp_348 <= MUX_s_1_2_2(nor_382_nl, mux_tmp_347, or_935_nl);
  nor_383_nl <= NOT((rem_12cyc_st_3_3_2(1)) OR (NOT mux_tmp_348));
  or_934_nl <= (NOT main_stage_0_4) OR (NOT COMP_LOOP_asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_3_3_2(0));
  mux_tmp_349 <= MUX_s_1_2_2(nor_383_nl, mux_tmp_348, or_934_nl);
  nor_384_nl <= NOT((rem_12cyc_st_2_3_2(1)) OR (NOT mux_tmp_349));
  or_933_nl <= (NOT main_stage_0_3) OR (NOT COMP_LOOP_asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_2_3_2(0));
  mux_tmp_350 <= MUX_s_1_2_2(nor_384_nl, mux_tmp_349, or_933_nl);
  nor_385_nl <= NOT((rem_12cyc_st_9_3_2(1)) OR (NOT mux_tmp_350));
  or_932_nl <= (NOT main_stage_0_10) OR (NOT COMP_LOOP_asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_9_3_2(0));
  mux_tmp_351 <= MUX_s_1_2_2(nor_385_nl, mux_tmp_350, or_932_nl);
  nor_386_nl <= NOT((rem_12cyc_st_8_3_2(1)) OR (NOT mux_tmp_351));
  or_931_nl <= (NOT main_stage_0_9) OR (NOT COMP_LOOP_asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_8_3_2(0));
  mux_tmp_352 <= MUX_s_1_2_2(nor_386_nl, mux_tmp_351, or_931_nl);
  nor_387_nl <= NOT((rem_12cyc_st_7_3_2(1)) OR (NOT mux_tmp_352));
  or_930_nl <= (NOT main_stage_0_8) OR (NOT COMP_LOOP_asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_7_3_2(0));
  mux_tmp_353 <= MUX_s_1_2_2(nor_387_nl, mux_tmp_352, or_930_nl);
  nor_388_nl <= NOT((rem_12cyc_1_0(0)) OR (NOT mux_tmp_353));
  or_929_nl <= (NOT main_stage_0_2) OR (NOT COMP_LOOP_asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_1_0(1));
  mux_tmp_354 <= MUX_s_1_2_2(nor_388_nl, mux_tmp_353, or_929_nl);
  and_dcpl_638 <= and_dcpl_568 AND and_dcpl_393;
  and_dcpl_639 <= and_dcpl_570 AND (rem_12cyc_st_2_1_0(1));
  or_tmp_934 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR not_tmp_54;
  or_952_cse <= CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("10"));
  nor_378_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_934));
  mux_355_nl <= MUX_s_1_2_2(nor_378_nl, or_tmp_934, or_952_cse);
  and_dcpl_641 <= mux_355_nl AND and_dcpl_298 AND and_dcpl_639;
  and_dcpl_642 <= and_dcpl_574 AND (rem_12cyc_st_3_1_0(1));
  or_957_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp_207 <= or_957_cse AND or_tmp_934;
  nor_377_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_207));
  mux_356_nl <= MUX_s_1_2_2(nor_377_nl, and_tmp_207, or_952_cse);
  and_dcpl_644 <= mux_356_nl AND and_dcpl_304 AND and_dcpl_642;
  and_dcpl_645 <= and_dcpl_578 AND (rem_12cyc_st_4_1_0(1));
  or_961_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_209 <= or_957_cse AND or_961_cse AND or_tmp_934;
  nor_376_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_209));
  mux_357_nl <= MUX_s_1_2_2(nor_376_nl, and_tmp_209, or_952_cse);
  and_dcpl_647 <= mux_357_nl AND and_dcpl_310 AND and_dcpl_645;
  and_dcpl_648 <= and_dcpl_582 AND (rem_12cyc_st_5_1_0(1));
  or_966_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_212 <= or_957_cse AND or_961_cse AND or_966_cse AND or_tmp_934;
  nor_375_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_212));
  mux_358_nl <= MUX_s_1_2_2(nor_375_nl, and_tmp_212, or_952_cse);
  and_dcpl_650 <= mux_358_nl AND and_dcpl_316 AND and_dcpl_648;
  or_972_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_216 <= or_957_cse AND or_961_cse AND or_966_cse AND or_972_cse AND or_tmp_934;
  nor_374_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_216));
  mux_359_nl <= MUX_s_1_2_2(nor_374_nl, and_tmp_216, or_952_cse);
  and_dcpl_653 <= mux_359_nl AND and_dcpl_112 AND and_dcpl_126 AND (rem_12cyc_st_6_1_0(1));
  or_979_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_372_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_934));
  mux_360_nl <= MUX_s_1_2_2(nor_372_nl, or_tmp_934, or_979_cse);
  and_tmp_220 <= or_957_cse AND or_961_cse AND or_966_cse AND or_972_cse AND mux_360_nl;
  nor_373_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_220));
  mux_361_nl <= MUX_s_1_2_2(nor_373_nl, and_tmp_220, or_952_cse);
  and_dcpl_657 <= mux_361_nl AND and_dcpl_85 AND and_dcpl_104 AND (NOT (rem_12cyc_st_7_1_0(0)));
  or_988_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_369_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_934));
  mux_tmp_362 <= MUX_s_1_2_2(nor_369_nl, or_tmp_934, or_988_cse);
  nor_370_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_362));
  mux_363_nl <= MUX_s_1_2_2(nor_370_nl, mux_tmp_362, or_979_cse);
  and_tmp_224 <= or_957_cse AND or_961_cse AND or_966_cse AND or_972_cse AND mux_363_nl;
  nor_371_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_224));
  mux_364_nl <= MUX_s_1_2_2(nor_371_nl, and_tmp_224, or_952_cse);
  and_dcpl_661 <= mux_364_nl AND and_dcpl_58 AND and_dcpl_77 AND (NOT (rem_12cyc_st_8_1_0(0)));
  or_999_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_365_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_934));
  mux_tmp_365 <= MUX_s_1_2_2(nor_365_nl, or_tmp_934, or_999_cse);
  nor_366_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_365));
  mux_tmp_366 <= MUX_s_1_2_2(nor_366_nl, mux_tmp_365, or_988_cse);
  nor_367_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_366));
  mux_367_nl <= MUX_s_1_2_2(nor_367_nl, mux_tmp_366, or_979_cse);
  and_tmp_228 <= or_957_cse AND or_961_cse AND or_966_cse AND or_972_cse AND mux_367_nl;
  nor_368_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_228));
  mux_368_nl <= MUX_s_1_2_2(nor_368_nl, and_tmp_228, or_952_cse);
  and_dcpl_665 <= mux_368_nl AND and_dcpl_31 AND and_dcpl_50 AND (NOT (rem_12cyc_st_9_1_0(0)));
  nor_360_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_934));
  or_1012_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("10"));
  mux_tmp_369 <= MUX_s_1_2_2(nor_360_nl, or_tmp_934, or_1012_nl);
  nor_361_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_369));
  mux_tmp_370 <= MUX_s_1_2_2(nor_361_nl, mux_tmp_369, or_999_cse);
  nor_362_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_370));
  mux_tmp_371 <= MUX_s_1_2_2(nor_362_nl, mux_tmp_370, or_988_cse);
  nor_363_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_371));
  mux_372_nl <= MUX_s_1_2_2(nor_363_nl, mux_tmp_371, or_979_cse);
  and_tmp_232 <= or_957_cse AND or_961_cse AND or_966_cse AND or_972_cse AND mux_372_nl;
  nor_364_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_232));
  mux_373_nl <= MUX_s_1_2_2(nor_364_nl, and_tmp_232, or_952_cse);
  and_dcpl_669 <= mux_373_nl AND and_dcpl_4 AND and_dcpl_23 AND (NOT (rem_12cyc_st_10_1_0(0)));
  or_tmp_1009 <= CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT ccs_ccore_start_rsci_idat);
  nor_351_nl <= NOT((rem_12cyc_st_10_3_2(1)) OR (NOT or_tmp_1009));
  or_1027_nl <= (NOT main_stage_0_11) OR (NOT COMP_LOOP_asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_10_3_2(0));
  mux_tmp_374 <= MUX_s_1_2_2(nor_351_nl, or_tmp_1009, or_1027_nl);
  nor_352_nl <= NOT((rem_12cyc_st_6_3_2(1)) OR (NOT mux_tmp_374));
  or_1026_nl <= (NOT main_stage_0_7) OR (NOT COMP_LOOP_asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_6_3_2(0));
  mux_tmp_375 <= MUX_s_1_2_2(nor_352_nl, mux_tmp_374, or_1026_nl);
  nor_353_nl <= NOT((rem_12cyc_st_5_3_2(1)) OR (NOT mux_tmp_375));
  or_1025_nl <= (NOT main_stage_0_6) OR (NOT COMP_LOOP_asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_5_3_2(0));
  mux_tmp_376 <= MUX_s_1_2_2(nor_353_nl, mux_tmp_375, or_1025_nl);
  nor_354_nl <= NOT((rem_12cyc_st_4_3_2(1)) OR (NOT mux_tmp_376));
  or_1024_nl <= (NOT main_stage_0_5) OR (NOT COMP_LOOP_asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_4_3_2(0));
  mux_tmp_377 <= MUX_s_1_2_2(nor_354_nl, mux_tmp_376, or_1024_nl);
  nor_355_nl <= NOT((rem_12cyc_st_3_3_2(1)) OR (NOT mux_tmp_377));
  or_1023_nl <= (NOT main_stage_0_4) OR (NOT COMP_LOOP_asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_3_3_2(0));
  mux_tmp_378 <= MUX_s_1_2_2(nor_355_nl, mux_tmp_377, or_1023_nl);
  nor_356_nl <= NOT((rem_12cyc_st_2_3_2(1)) OR (NOT mux_tmp_378));
  or_1022_nl <= (NOT main_stage_0_3) OR (NOT COMP_LOOP_asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_2_3_2(0));
  mux_tmp_379 <= MUX_s_1_2_2(nor_356_nl, mux_tmp_378, or_1022_nl);
  nor_357_nl <= NOT((rem_12cyc_st_9_3_2(1)) OR (NOT mux_tmp_379));
  or_1021_nl <= (NOT main_stage_0_10) OR (NOT COMP_LOOP_asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_9_3_2(0));
  mux_tmp_380 <= MUX_s_1_2_2(nor_357_nl, mux_tmp_379, or_1021_nl);
  nor_358_nl <= NOT((rem_12cyc_st_8_3_2(1)) OR (NOT mux_tmp_380));
  or_1020_nl <= (NOT main_stage_0_9) OR (NOT COMP_LOOP_asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_8_3_2(0));
  mux_tmp_381 <= MUX_s_1_2_2(nor_358_nl, mux_tmp_380, or_1020_nl);
  nor_359_nl <= NOT((rem_12cyc_st_7_3_2(1)) OR (NOT mux_tmp_381));
  or_1019_nl <= (NOT main_stage_0_8) OR (NOT COMP_LOOP_asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_7_3_2(0));
  mux_382_nl <= MUX_s_1_2_2(nor_359_nl, mux_tmp_381, or_1019_nl);
  and_tmp_233 <= ((NOT main_stage_0_2) OR (NOT COMP_LOOP_asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10"))) AND mux_382_nl;
  and_dcpl_673 <= and_dcpl_568 AND and_dcpl_430;
  or_tmp_1021 <= (NOT(CONV_SL_1_1(rem_12cyc_1_0=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(rem_12cyc_3_2=STD_LOGIC_VECTOR'("10"))))
      OR not_tmp_54;
  nand_57_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(COMP_LOOP_acc_tmp=STD_LOGIC_VECTOR'("10")));
  nor_350_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_1021));
  mux_383_nl <= MUX_s_1_2_2(nor_350_nl, or_tmp_1021, nand_57_cse);
  and_dcpl_675 <= mux_383_nl AND and_dcpl_358 AND and_dcpl_639;
  or_1045_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR (rem_12cyc_st_2_3_2(0));
  and_960_nl <= nand_84_cse AND or_tmp_1021;
  mux_tmp_384 <= MUX_s_1_2_2(and_960_nl, or_tmp_1021, or_1045_cse);
  nor_349_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_384));
  mux_385_nl <= MUX_s_1_2_2(nor_349_nl, mux_tmp_384, nand_57_cse);
  and_dcpl_677 <= mux_385_nl AND and_dcpl_362 AND and_dcpl_642;
  or_1050_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("10"));
  and_958_nl <= nand_274_cse AND or_tmp_1021;
  mux_tmp_386 <= MUX_s_1_2_2(and_958_nl, or_tmp_1021, or_1050_cse);
  and_959_nl <= nand_84_cse AND mux_tmp_386;
  mux_tmp_387 <= MUX_s_1_2_2(and_959_nl, mux_tmp_386, or_1045_cse);
  nor_348_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_387));
  mux_388_nl <= MUX_s_1_2_2(nor_348_nl, mux_tmp_387, nand_57_cse);
  and_dcpl_679 <= mux_388_nl AND and_dcpl_366 AND and_dcpl_645;
  or_1057_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR (rem_12cyc_st_4_3_2(0));
  and_955_nl <= nand_79_cse AND or_tmp_1021;
  mux_tmp_389 <= MUX_s_1_2_2(and_955_nl, or_tmp_1021, or_1057_cse);
  and_956_nl <= nand_274_cse AND mux_tmp_389;
  mux_tmp_390 <= MUX_s_1_2_2(and_956_nl, mux_tmp_389, or_1050_cse);
  and_957_nl <= nand_84_cse AND mux_tmp_390;
  mux_tmp_391 <= MUX_s_1_2_2(and_957_nl, mux_tmp_390, or_1045_cse);
  nor_347_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_391));
  mux_392_nl <= MUX_s_1_2_2(nor_347_nl, mux_tmp_391, nand_57_cse);
  and_dcpl_681 <= mux_392_nl AND and_dcpl_370 AND and_dcpl_648;
  or_1066_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("10"));
  and_951_nl <= nand_267_cse AND or_tmp_1021;
  mux_tmp_393 <= MUX_s_1_2_2(and_951_nl, or_tmp_1021, or_1066_cse);
  and_952_nl <= nand_79_cse AND mux_tmp_393;
  mux_tmp_394 <= MUX_s_1_2_2(and_952_nl, mux_tmp_393, or_1057_cse);
  and_953_nl <= nand_274_cse AND mux_tmp_394;
  mux_tmp_395 <= MUX_s_1_2_2(and_953_nl, mux_tmp_394, or_1050_cse);
  and_954_nl <= nand_84_cse AND mux_tmp_395;
  mux_tmp_396 <= MUX_s_1_2_2(and_954_nl, mux_tmp_395, or_1045_cse);
  nor_346_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_396));
  mux_397_nl <= MUX_s_1_2_2(nor_346_nl, mux_tmp_396, nand_57_cse);
  and_dcpl_684 <= mux_397_nl AND and_dcpl_112 AND and_dcpl_129 AND (rem_12cyc_st_6_1_0(1));
  nand_36_cse <= NOT(CONV_SL_1_1(rem_12cyc_st_6_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_6_3_2=STD_LOGIC_VECTOR'("10")));
  nor_344_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_1021));
  mux_tmp_398 <= MUX_s_1_2_2(nor_344_nl, or_tmp_1021, nand_36_cse);
  and_947_nl <= nand_267_cse AND mux_tmp_398;
  mux_tmp_399 <= MUX_s_1_2_2(and_947_nl, mux_tmp_398, or_1066_cse);
  and_948_nl <= nand_79_cse AND mux_tmp_399;
  mux_tmp_400 <= MUX_s_1_2_2(and_948_nl, mux_tmp_399, or_1057_cse);
  and_949_nl <= nand_274_cse AND mux_tmp_400;
  mux_tmp_401 <= MUX_s_1_2_2(and_949_nl, mux_tmp_400, or_1050_cse);
  and_950_nl <= nand_84_cse AND mux_tmp_401;
  mux_tmp_402 <= MUX_s_1_2_2(and_950_nl, mux_tmp_401, or_1045_cse);
  nor_345_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_402));
  mux_403_nl <= MUX_s_1_2_2(nor_345_nl, mux_tmp_402, nand_57_cse);
  and_dcpl_687 <= mux_403_nl AND and_dcpl_85 AND and_dcpl_104 AND (rem_12cyc_st_7_1_0(0));
  nand_29_cse <= NOT(CONV_SL_1_1(rem_12cyc_st_7_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_7_3_2=STD_LOGIC_VECTOR'("10")));
  nor_341_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_1021));
  mux_tmp_404 <= MUX_s_1_2_2(nor_341_nl, or_tmp_1021, nand_29_cse);
  nor_342_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_404));
  mux_tmp_405 <= MUX_s_1_2_2(nor_342_nl, mux_tmp_404, nand_36_cse);
  and_943_nl <= nand_267_cse AND mux_tmp_405;
  mux_tmp_406 <= MUX_s_1_2_2(and_943_nl, mux_tmp_405, or_1066_cse);
  and_944_nl <= nand_79_cse AND mux_tmp_406;
  mux_tmp_407 <= MUX_s_1_2_2(and_944_nl, mux_tmp_406, or_1057_cse);
  and_945_nl <= nand_274_cse AND mux_tmp_407;
  mux_tmp_408 <= MUX_s_1_2_2(and_945_nl, mux_tmp_407, or_1050_cse);
  and_946_nl <= nand_84_cse AND mux_tmp_408;
  mux_tmp_409 <= MUX_s_1_2_2(and_946_nl, mux_tmp_408, or_1045_cse);
  nor_343_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_409));
  mux_410_nl <= MUX_s_1_2_2(nor_343_nl, mux_tmp_409, nand_57_cse);
  and_dcpl_690 <= mux_410_nl AND and_dcpl_58 AND and_dcpl_77 AND (rem_12cyc_st_8_1_0(0));
  nand_21_cse <= NOT(CONV_SL_1_1(rem_12cyc_st_8_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_8_3_2=STD_LOGIC_VECTOR'("10")));
  nor_337_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_1021));
  mux_tmp_411 <= MUX_s_1_2_2(nor_337_nl, or_tmp_1021, nand_21_cse);
  nor_338_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_411));
  mux_tmp_412 <= MUX_s_1_2_2(nor_338_nl, mux_tmp_411, nand_29_cse);
  nor_339_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_412));
  mux_tmp_413 <= MUX_s_1_2_2(nor_339_nl, mux_tmp_412, nand_36_cse);
  and_939_nl <= nand_267_cse AND mux_tmp_413;
  mux_tmp_414 <= MUX_s_1_2_2(and_939_nl, mux_tmp_413, or_1066_cse);
  and_940_nl <= nand_79_cse AND mux_tmp_414;
  mux_tmp_415 <= MUX_s_1_2_2(and_940_nl, mux_tmp_414, or_1057_cse);
  and_941_nl <= nand_274_cse AND mux_tmp_415;
  mux_tmp_416 <= MUX_s_1_2_2(and_941_nl, mux_tmp_415, or_1050_cse);
  and_942_nl <= nand_84_cse AND mux_tmp_416;
  mux_tmp_417 <= MUX_s_1_2_2(and_942_nl, mux_tmp_416, or_1045_cse);
  nor_340_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_417));
  mux_418_nl <= MUX_s_1_2_2(nor_340_nl, mux_tmp_417, nand_57_cse);
  and_dcpl_693 <= mux_418_nl AND and_dcpl_31 AND and_dcpl_50 AND (rem_12cyc_st_9_1_0(0));
  nor_332_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_1021));
  nand_12_nl <= NOT(CONV_SL_1_1(rem_12cyc_st_9_1_0=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(rem_12cyc_st_9_3_2=STD_LOGIC_VECTOR'("10")));
  mux_tmp_419 <= MUX_s_1_2_2(nor_332_nl, or_tmp_1021, nand_12_nl);
  nor_333_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_419));
  mux_tmp_420 <= MUX_s_1_2_2(nor_333_nl, mux_tmp_419, nand_21_cse);
  nor_334_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_420));
  mux_tmp_421 <= MUX_s_1_2_2(nor_334_nl, mux_tmp_420, nand_29_cse);
  nor_335_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_421));
  mux_tmp_422 <= MUX_s_1_2_2(nor_335_nl, mux_tmp_421, nand_36_cse);
  and_935_nl <= nand_267_cse AND mux_tmp_422;
  mux_tmp_423 <= MUX_s_1_2_2(and_935_nl, mux_tmp_422, or_1066_cse);
  and_936_nl <= nand_79_cse AND mux_tmp_423;
  mux_tmp_424 <= MUX_s_1_2_2(and_936_nl, mux_tmp_423, or_1057_cse);
  and_937_nl <= nand_274_cse AND mux_tmp_424;
  mux_tmp_425 <= MUX_s_1_2_2(and_937_nl, mux_tmp_424, or_1050_cse);
  and_938_nl <= nand_84_cse AND mux_tmp_425;
  mux_tmp_426 <= MUX_s_1_2_2(and_938_nl, mux_tmp_425, or_1045_cse);
  nor_336_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_426));
  mux_427_nl <= MUX_s_1_2_2(nor_336_nl, mux_tmp_426, nand_57_cse);
  and_dcpl_696 <= mux_427_nl AND and_dcpl_4 AND and_dcpl_23 AND (rem_12cyc_st_10_1_0(0));
  or_tmp_1122 <= CONV_SL_1_1(COMP_LOOP_acc_tmp/=STD_LOGIC_VECTOR'("10")) OR nand_222_cse;
  nor_323_nl <= NOT((rem_12cyc_st_10_3_2(1)) OR (NOT or_tmp_1122));
  nand_1_nl <= NOT(main_stage_0_11 AND COMP_LOOP_asn_itm_10 AND CONV_SL_1_1(rem_12cyc_st_10_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_10_3_2(0))));
  mux_tmp_428 <= MUX_s_1_2_2(nor_323_nl, or_tmp_1122, nand_1_nl);
  nor_324_nl <= NOT((rem_12cyc_st_6_3_2(1)) OR (NOT mux_tmp_428));
  nand_2_nl <= NOT(main_stage_0_7 AND COMP_LOOP_asn_itm_6 AND CONV_SL_1_1(rem_12cyc_st_6_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_6_3_2(0))));
  mux_tmp_429 <= MUX_s_1_2_2(nor_324_nl, mux_tmp_428, nand_2_nl);
  nor_325_nl <= NOT((rem_12cyc_st_5_3_2(1)) OR (NOT mux_tmp_429));
  nand_3_nl <= NOT(main_stage_0_6 AND COMP_LOOP_asn_itm_5 AND CONV_SL_1_1(rem_12cyc_st_5_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_5_3_2(0))));
  mux_tmp_430 <= MUX_s_1_2_2(nor_325_nl, mux_tmp_429, nand_3_nl);
  nor_326_nl <= NOT((rem_12cyc_st_4_3_2(1)) OR (NOT mux_tmp_430));
  nand_4_nl <= NOT(main_stage_0_5 AND COMP_LOOP_asn_itm_4 AND CONV_SL_1_1(rem_12cyc_st_4_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_4_3_2(0))));
  mux_tmp_431 <= MUX_s_1_2_2(nor_326_nl, mux_tmp_430, nand_4_nl);
  nor_327_nl <= NOT((rem_12cyc_st_3_3_2(1)) OR (NOT mux_tmp_431));
  nand_5_nl <= NOT(main_stage_0_4 AND COMP_LOOP_asn_itm_3 AND CONV_SL_1_1(rem_12cyc_st_3_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_3_3_2(0))));
  mux_tmp_432 <= MUX_s_1_2_2(nor_327_nl, mux_tmp_431, nand_5_nl);
  nor_328_nl <= NOT((rem_12cyc_st_2_3_2(1)) OR (NOT mux_tmp_432));
  nand_6_nl <= NOT(main_stage_0_3 AND COMP_LOOP_asn_itm_2 AND CONV_SL_1_1(rem_12cyc_st_2_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_2_3_2(0))));
  mux_tmp_433 <= MUX_s_1_2_2(nor_328_nl, mux_tmp_432, nand_6_nl);
  nor_329_nl <= NOT((rem_12cyc_st_9_3_2(1)) OR (NOT mux_tmp_433));
  nand_7_nl <= NOT(main_stage_0_10 AND COMP_LOOP_asn_itm_9 AND CONV_SL_1_1(rem_12cyc_st_9_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_9_3_2(0))));
  mux_tmp_434 <= MUX_s_1_2_2(nor_329_nl, mux_tmp_433, nand_7_nl);
  nor_330_nl <= NOT((rem_12cyc_st_8_3_2(1)) OR (NOT mux_tmp_434));
  nand_8_nl <= NOT(main_stage_0_9 AND COMP_LOOP_asn_itm_8 AND CONV_SL_1_1(rem_12cyc_st_8_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_8_3_2(0))));
  mux_tmp_435 <= MUX_s_1_2_2(nor_330_nl, mux_tmp_434, nand_8_nl);
  nor_331_nl <= NOT((rem_12cyc_st_7_3_2(1)) OR (NOT mux_tmp_435));
  nand_9_nl <= NOT(main_stage_0_8 AND COMP_LOOP_asn_itm_7 AND CONV_SL_1_1(rem_12cyc_st_7_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_7_3_2(0))));
  mux_tmp_436 <= MUX_s_1_2_2(nor_331_nl, mux_tmp_435, nand_9_nl);
  and_934_nl <= nand_223_cse AND mux_tmp_436;
  nand_11_nl <= NOT(main_stage_0_2 AND COMP_LOOP_asn_itm_1 AND CONV_SL_1_1(rem_12cyc_3_2=STD_LOGIC_VECTOR'("10")));
  mux_tmp_437 <= MUX_s_1_2_2(and_934_nl, mux_tmp_436, nand_11_nl);
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( ccs_ccore_en = '1' ) THEN
        return_rsci_d <= MUX_v_64_2_2(result_sva_duc_mx0, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(qelse_acc_nl),
            64)), mux_11_nl);
        m_buf_sva_12 <= m_buf_sva_11;
        m_buf_sva_11 <= m_buf_sva_10;
        m_buf_sva_10 <= m_buf_sva_9;
        m_buf_sva_9 <= m_buf_sva_8;
        m_buf_sva_8 <= m_buf_sva_7;
        m_buf_sva_7 <= m_buf_sva_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        COMP_LOOP_asn_itm_12 <= '0';
        COMP_LOOP_asn_itm_11 <= '0';
        COMP_LOOP_asn_itm_10 <= '0';
        COMP_LOOP_asn_itm_9 <= '0';
        COMP_LOOP_asn_itm_8 <= '0';
        COMP_LOOP_asn_itm_7 <= '0';
        COMP_LOOP_asn_itm_6 <= '0';
        COMP_LOOP_asn_itm_5 <= '0';
        COMP_LOOP_asn_itm_4 <= '0';
        COMP_LOOP_asn_itm_3 <= '0';
        COMP_LOOP_asn_itm_2 <= '0';
        COMP_LOOP_asn_itm_1 <= '0';
        main_stage_0_2 <= '0';
        main_stage_0_3 <= '0';
        main_stage_0_4 <= '0';
        main_stage_0_5 <= '0';
        main_stage_0_6 <= '0';
        main_stage_0_7 <= '0';
        main_stage_0_8 <= '0';
        main_stage_0_9 <= '0';
        main_stage_0_10 <= '0';
        main_stage_0_11 <= '0';
        main_stage_0_12 <= '0';
        main_stage_0_13 <= '0';
      ELSIF ( ccs_ccore_en = '1' ) THEN
        COMP_LOOP_asn_itm_12 <= COMP_LOOP_asn_itm_11;
        COMP_LOOP_asn_itm_11 <= COMP_LOOP_asn_itm_10;
        COMP_LOOP_asn_itm_10 <= COMP_LOOP_asn_itm_9;
        COMP_LOOP_asn_itm_9 <= COMP_LOOP_asn_itm_8;
        COMP_LOOP_asn_itm_8 <= COMP_LOOP_asn_itm_7;
        COMP_LOOP_asn_itm_7 <= COMP_LOOP_asn_itm_6;
        COMP_LOOP_asn_itm_6 <= COMP_LOOP_asn_itm_5;
        COMP_LOOP_asn_itm_5 <= COMP_LOOP_asn_itm_4;
        COMP_LOOP_asn_itm_4 <= COMP_LOOP_asn_itm_3;
        COMP_LOOP_asn_itm_3 <= COMP_LOOP_asn_itm_2;
        COMP_LOOP_asn_itm_2 <= COMP_LOOP_asn_itm_1;
        COMP_LOOP_asn_itm_1 <= ccs_ccore_start_rsci_idat;
        main_stage_0_2 <= '1';
        main_stage_0_3 <= main_stage_0_2;
        main_stage_0_4 <= main_stage_0_3;
        main_stage_0_5 <= main_stage_0_4;
        main_stage_0_6 <= main_stage_0_5;
        main_stage_0_7 <= main_stage_0_6;
        main_stage_0_8 <= main_stage_0_7;
        main_stage_0_9 <= main_stage_0_8;
        main_stage_0_10 <= main_stage_0_9;
        main_stage_0_11 <= main_stage_0_10;
        main_stage_0_12 <= main_stage_0_11;
        main_stage_0_13 <= main_stage_0_12;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_sva_duc <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
      ELSIF ( (COMP_LOOP_asn_itm_12 AND main_stage_0_13 AND ccs_ccore_en AND (NOT(CONV_SL_1_1(rem_12cyc_st_12_3_2=STD_LOGIC_VECTOR'("11")))))
          = '1' ) THEN
        result_sva_duc <= result_sva_duc_mx0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_12_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_12_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( COMP_LOOP_and_26_cse = '1' ) THEN
        rem_12cyc_st_12_3_2 <= rem_12cyc_st_11_3_2;
        rem_12cyc_st_12_1_0 <= rem_12cyc_st_11_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_cse = '1' ) THEN
        rem_12_cmp_1_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_3_2_63_0, mut_3_3_63_0,
            mut_3_4_63_0, mut_3_5_63_0, mut_3_6_63_0, mut_3_7_63_0, mut_3_8_63_0,
            mut_3_9_63_0, mut_3_10_63_0, mut_3_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_294
            & and_dcpl_300 & and_dcpl_306 & and_dcpl_312 & and_dcpl_318 & and_dcpl_324
            & and_dcpl_330 & and_dcpl_336 & and_dcpl_342 & and_dcpl_348 & and_tmp_35));
        rem_12_cmp_1_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_2_2_63_0, mut_2_3_63_0,
            mut_2_4_63_0, mut_2_5_63_0, mut_2_6_63_0, mut_2_7_63_0, mut_2_8_63_0,
            mut_2_9_63_0, mut_2_10_63_0, mut_2_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_294
            & and_dcpl_300 & and_dcpl_306 & and_dcpl_312 & and_dcpl_318 & and_dcpl_324
            & and_dcpl_330 & and_dcpl_336 & and_dcpl_342 & and_dcpl_348 & and_tmp_35));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_2_cse = '1' ) THEN
        rem_12_cmp_2_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_5_2_63_0, mut_5_3_63_0,
            mut_5_4_63_0, mut_5_5_63_0, mut_5_6_63_0, mut_5_7_63_0, mut_5_8_63_0,
            mut_5_9_63_0, mut_5_10_63_0, mut_5_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_356
            & and_dcpl_360 & and_dcpl_364 & and_dcpl_368 & and_dcpl_372 & and_dcpl_376
            & and_dcpl_379 & and_dcpl_382 & and_dcpl_385 & and_dcpl_388 & mux_tmp_76));
        rem_12_cmp_2_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_4_2_63_0, mut_4_3_63_0,
            mut_4_4_63_0, mut_4_5_63_0, mut_4_6_63_0, mut_4_7_63_0, mut_4_8_63_0,
            mut_4_9_63_0, mut_4_10_63_0, mut_4_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_356
            & and_dcpl_360 & and_dcpl_364 & and_dcpl_368 & and_dcpl_372 & and_dcpl_376
            & and_dcpl_379 & and_dcpl_382 & and_dcpl_385 & and_dcpl_388 & mux_tmp_76));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_4_cse = '1' ) THEN
        rem_12_cmp_3_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_7_2_63_0, mut_7_3_63_0,
            mut_7_4_63_0, mut_7_5_63_0, mut_7_6_63_0, mut_7_7_63_0, mut_7_8_63_0,
            mut_7_9_63_0, mut_7_10_63_0, mut_7_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_394
            & and_dcpl_397 & and_dcpl_400 & and_dcpl_403 & and_dcpl_406 & and_dcpl_409
            & and_dcpl_413 & and_dcpl_417 & and_dcpl_421 & and_dcpl_425 & and_tmp_80));
        rem_12_cmp_3_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_6_2_63_0, mut_6_3_63_0,
            mut_6_4_63_0, mut_6_5_63_0, mut_6_6_63_0, mut_6_7_63_0, mut_6_8_63_0,
            mut_6_9_63_0, mut_6_10_63_0, mut_6_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_394
            & and_dcpl_397 & and_dcpl_400 & and_dcpl_403 & and_dcpl_406 & and_dcpl_409
            & and_dcpl_413 & and_dcpl_417 & and_dcpl_421 & and_dcpl_425 & and_tmp_80));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_6_cse = '1' ) THEN
        rem_12_cmp_4_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_9_2_63_0, mut_9_3_63_0,
            mut_9_4_63_0, mut_9_5_63_0, mut_9_6_63_0, mut_9_7_63_0, mut_9_8_63_0,
            mut_9_9_63_0, mut_9_10_63_0, mut_9_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_431
            & and_dcpl_433 & and_dcpl_435 & and_dcpl_437 & and_dcpl_439 & and_dcpl_442
            & and_dcpl_445 & and_dcpl_448 & and_dcpl_451 & and_dcpl_454 & mux_tmp_141));
        rem_12_cmp_4_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_8_2_63_0, mut_8_3_63_0,
            mut_8_4_63_0, mut_8_5_63_0, mut_8_6_63_0, mut_8_7_63_0, mut_8_8_63_0,
            mut_8_9_63_0, mut_8_10_63_0, mut_8_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_431
            & and_dcpl_433 & and_dcpl_435 & and_dcpl_437 & and_dcpl_439 & and_dcpl_442
            & and_dcpl_445 & and_dcpl_448 & and_dcpl_451 & and_dcpl_454 & mux_tmp_141));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_8_cse = '1' ) THEN
        rem_12_cmp_5_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_11_2_63_0, mut_11_3_63_0,
            mut_11_4_63_0, mut_11_5_63_0, mut_11_6_63_0, mut_11_7_63_0, mut_11_8_63_0,
            mut_11_9_63_0, mut_11_10_63_0, mut_11_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_461
            & and_dcpl_465 & and_dcpl_469 & and_dcpl_473 & and_dcpl_477 & and_dcpl_480
            & and_dcpl_483 & and_dcpl_486 & and_dcpl_489 & and_dcpl_492 & and_tmp_125));
        rem_12_cmp_5_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_10_2_63_0, mut_10_3_63_0,
            mut_10_4_63_0, mut_10_5_63_0, mut_10_6_63_0, mut_10_7_63_0, mut_10_8_63_0,
            mut_10_9_63_0, mut_10_10_63_0, mut_10_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_461
            & and_dcpl_465 & and_dcpl_469 & and_dcpl_473 & and_dcpl_477 & and_dcpl_480
            & and_dcpl_483 & and_dcpl_486 & and_dcpl_489 & and_dcpl_492 & and_tmp_125));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_10_cse = '1' ) THEN
        rem_12_cmp_6_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_13_2_63_0, mut_13_3_63_0,
            mut_13_4_63_0, mut_13_5_63_0, mut_13_6_63_0, mut_13_7_63_0, mut_13_8_63_0,
            mut_13_9_63_0, mut_13_10_63_0, mut_13_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_498
            & and_dcpl_500 & and_dcpl_502 & and_dcpl_504 & and_dcpl_506 & and_dcpl_508
            & and_dcpl_510 & and_dcpl_512 & and_dcpl_514 & and_dcpl_516 & mux_tmp_206));
        rem_12_cmp_6_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_12_2_63_0, mut_12_3_63_0,
            mut_12_4_63_0, mut_12_5_63_0, mut_12_6_63_0, mut_12_7_63_0, mut_12_8_63_0,
            mut_12_9_63_0, mut_12_10_63_0, mut_12_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_498
            & and_dcpl_500 & and_dcpl_502 & and_dcpl_504 & and_dcpl_506 & and_dcpl_508
            & and_dcpl_510 & and_dcpl_512 & and_dcpl_514 & and_dcpl_516 & mux_tmp_206));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_12_cse = '1' ) THEN
        rem_12_cmp_7_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_15_2_63_0, mut_15_3_63_0,
            mut_15_4_63_0, mut_15_5_63_0, mut_15_6_63_0, mut_15_7_63_0, mut_15_8_63_0,
            mut_15_9_63_0, mut_15_10_63_0, mut_15_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_520
            & and_dcpl_523 & and_dcpl_526 & and_dcpl_529 & and_dcpl_532 & and_dcpl_534
            & and_dcpl_536 & and_dcpl_538 & and_dcpl_540 & and_dcpl_542 & and_tmp_170));
        rem_12_cmp_7_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_14_2_63_0, mut_14_3_63_0,
            mut_14_4_63_0, mut_14_5_63_0, mut_14_6_63_0, mut_14_7_63_0, mut_14_8_63_0,
            mut_14_9_63_0, mut_14_10_63_0, mut_14_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_520
            & and_dcpl_523 & and_dcpl_526 & and_dcpl_529 & and_dcpl_532 & and_dcpl_534
            & and_dcpl_536 & and_dcpl_538 & and_dcpl_540 & and_dcpl_542 & and_tmp_170));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_14_cse = '1' ) THEN
        rem_12_cmp_8_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_17_2_63_0, mut_17_3_63_0,
            mut_17_4_63_0, mut_17_5_63_0, mut_17_6_63_0, mut_17_7_63_0, mut_17_8_63_0,
            mut_17_9_63_0, mut_17_10_63_0, mut_17_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_546
            & and_dcpl_548 & and_dcpl_550 & and_dcpl_552 & and_dcpl_554 & and_dcpl_556
            & and_dcpl_558 & and_dcpl_560 & and_dcpl_562 & and_dcpl_564 & mux_tmp_271));
        rem_12_cmp_8_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_16_2_63_0, mut_16_3_63_0,
            mut_16_4_63_0, mut_16_5_63_0, mut_16_6_63_0, mut_16_7_63_0, mut_16_8_63_0,
            mut_16_9_63_0, mut_16_10_63_0, mut_16_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_546
            & and_dcpl_548 & and_dcpl_550 & and_dcpl_552 & and_dcpl_554 & and_dcpl_556
            & and_dcpl_558 & and_dcpl_560 & and_dcpl_562 & and_dcpl_564 & mux_tmp_271));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_16_cse = '1' ) THEN
        rem_12_cmp_9_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_19_2_63_0, mut_19_3_63_0,
            mut_19_4_63_0, mut_19_5_63_0, mut_19_6_63_0, mut_19_7_63_0, mut_19_8_63_0,
            mut_19_9_63_0, mut_19_10_63_0, mut_19_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_569
            & and_dcpl_573 & and_dcpl_577 & and_dcpl_581 & and_dcpl_585 & and_dcpl_589
            & and_dcpl_593 & and_dcpl_597 & and_dcpl_601 & and_dcpl_605 & and_tmp_206));
        rem_12_cmp_9_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_18_2_63_0, mut_18_3_63_0,
            mut_18_4_63_0, mut_18_5_63_0, mut_18_6_63_0, mut_18_7_63_0, mut_18_8_63_0,
            mut_18_9_63_0, mut_18_10_63_0, mut_18_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_569
            & and_dcpl_573 & and_dcpl_577 & and_dcpl_581 & and_dcpl_585 & and_dcpl_589
            & and_dcpl_593 & and_dcpl_597 & and_dcpl_601 & and_dcpl_605 & and_tmp_206));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_18_cse = '1' ) THEN
        rem_12_cmp_10_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_21_2_63_0, mut_21_3_63_0,
            mut_21_4_63_0, mut_21_5_63_0, mut_21_6_63_0, mut_21_7_63_0, mut_21_8_63_0,
            mut_21_9_63_0, mut_21_10_63_0, mut_21_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_610
            & and_dcpl_612 & and_dcpl_614 & and_dcpl_616 & and_dcpl_618 & and_dcpl_622
            & and_dcpl_625 & and_dcpl_628 & and_dcpl_631 & and_dcpl_634 & mux_tmp_354));
        rem_12_cmp_10_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_20_2_63_0,
            mut_20_3_63_0, mut_20_4_63_0, mut_20_5_63_0, mut_20_6_63_0, mut_20_7_63_0,
            mut_20_8_63_0, mut_20_9_63_0, mut_20_10_63_0, mut_20_11_63_0, STD_LOGIC_VECTOR'(
            and_dcpl_610 & and_dcpl_612 & and_dcpl_614 & and_dcpl_616 & and_dcpl_618
            & and_dcpl_622 & and_dcpl_625 & and_dcpl_628 & and_dcpl_631 & and_dcpl_634
            & mux_tmp_354));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_20_cse = '1' ) THEN
        rem_12_cmp_11_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_23_2_63_0, mut_23_3_63_0,
            mut_23_4_63_0, mut_23_5_63_0, mut_23_6_63_0, mut_23_7_63_0, mut_23_8_63_0,
            mut_23_9_63_0, mut_23_10_63_0, mut_23_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_638
            & and_dcpl_641 & and_dcpl_644 & and_dcpl_647 & and_dcpl_650 & and_dcpl_653
            & and_dcpl_657 & and_dcpl_661 & and_dcpl_665 & and_dcpl_669 & and_tmp_233));
        rem_12_cmp_11_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_22_2_63_0,
            mut_22_3_63_0, mut_22_4_63_0, mut_22_5_63_0, mut_22_6_63_0, mut_22_7_63_0,
            mut_22_8_63_0, mut_22_9_63_0, mut_22_10_63_0, mut_22_11_63_0, STD_LOGIC_VECTOR'(
            and_dcpl_638 & and_dcpl_641 & and_dcpl_644 & and_dcpl_647 & and_dcpl_650
            & and_dcpl_653 & and_dcpl_657 & and_dcpl_661 & and_dcpl_665 & and_dcpl_669
            & and_tmp_233));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_22_cse = '1' ) THEN
        rem_12_cmp_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_1_2_63_0, mut_1_3_63_0,
            mut_1_4_63_0, mut_1_5_63_0, mut_1_6_63_0, mut_1_7_63_0, mut_1_8_63_0,
            mut_1_9_63_0, mut_1_10_63_0, mut_1_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_673
            & and_dcpl_675 & and_dcpl_677 & and_dcpl_679 & and_dcpl_681 & and_dcpl_684
            & and_dcpl_687 & and_dcpl_690 & and_dcpl_693 & and_dcpl_696 & mux_tmp_437));
        rem_12_cmp_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_2_63_0, mut_3_63_0,
            mut_4_63_0, mut_5_63_0, mut_6_63_0, mut_7_63_0, mut_8_63_0, mut_9_63_0,
            mut_10_63_0, mut_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_673 & and_dcpl_675
            & and_dcpl_677 & and_dcpl_679 & and_dcpl_681 & and_dcpl_684 & and_dcpl_687
            & and_dcpl_690 & and_dcpl_693 & and_dcpl_696 & mux_tmp_437));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_28_cse = '1' ) THEN
        mut_3_11_63_0 <= mut_3_10_63_0;
        mut_2_11_63_0 <= mut_2_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_30_cse = '1' ) THEN
        mut_5_11_63_0 <= mut_5_10_63_0;
        mut_4_11_63_0 <= mut_4_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_32_cse = '1' ) THEN
        mut_7_11_63_0 <= mut_7_10_63_0;
        mut_6_11_63_0 <= mut_6_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_34_cse = '1' ) THEN
        mut_9_11_63_0 <= mut_9_10_63_0;
        mut_8_11_63_0 <= mut_8_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_36_cse = '1' ) THEN
        mut_11_11_63_0 <= mut_11_10_63_0;
        mut_10_11_63_0 <= mut_10_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_38_cse = '1' ) THEN
        mut_13_11_63_0 <= mut_13_10_63_0;
        mut_12_11_63_0 <= mut_12_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_40_cse = '1' ) THEN
        mut_15_11_63_0 <= mut_15_10_63_0;
        mut_14_11_63_0 <= mut_14_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_42_cse = '1' ) THEN
        mut_17_11_63_0 <= mut_17_10_63_0;
        mut_16_11_63_0 <= mut_16_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_44_cse = '1' ) THEN
        mut_19_11_63_0 <= mut_19_10_63_0;
        mut_18_11_63_0 <= mut_18_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_46_cse = '1' ) THEN
        mut_21_11_63_0 <= mut_21_10_63_0;
        mut_20_11_63_0 <= mut_20_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_48_cse = '1' ) THEN
        mut_23_11_63_0 <= mut_23_10_63_0;
        mut_22_11_63_0 <= mut_22_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_50_cse = '1' ) THEN
        mut_1_11_63_0 <= mut_1_10_63_0;
        mut_11_63_0 <= mut_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_11_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_11_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( COMP_LOOP_and_52_cse = '1' ) THEN
        rem_12cyc_st_11_3_2 <= rem_12cyc_st_10_3_2;
        rem_12cyc_st_11_1_0 <= rem_12cyc_st_10_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_54_cse = '1' ) THEN
        mut_3_10_63_0 <= mut_3_9_63_0;
        mut_2_10_63_0 <= mut_2_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_56_cse = '1' ) THEN
        mut_5_10_63_0 <= mut_5_9_63_0;
        mut_4_10_63_0 <= mut_4_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_58_cse = '1' ) THEN
        mut_7_10_63_0 <= mut_7_9_63_0;
        mut_6_10_63_0 <= mut_6_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_60_cse = '1' ) THEN
        mut_9_10_63_0 <= mut_9_9_63_0;
        mut_8_10_63_0 <= mut_8_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_62_cse = '1' ) THEN
        mut_11_10_63_0 <= mut_11_9_63_0;
        mut_10_10_63_0 <= mut_10_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_64_cse = '1' ) THEN
        mut_13_10_63_0 <= mut_13_9_63_0;
        mut_12_10_63_0 <= mut_12_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_66_cse = '1' ) THEN
        mut_15_10_63_0 <= mut_15_9_63_0;
        mut_14_10_63_0 <= mut_14_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_68_cse = '1' ) THEN
        mut_17_10_63_0 <= mut_17_9_63_0;
        mut_16_10_63_0 <= mut_16_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_70_cse = '1' ) THEN
        mut_19_10_63_0 <= mut_19_9_63_0;
        mut_18_10_63_0 <= mut_18_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_72_cse = '1' ) THEN
        mut_21_10_63_0 <= mut_21_9_63_0;
        mut_20_10_63_0 <= mut_20_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_74_cse = '1' ) THEN
        mut_23_10_63_0 <= mut_23_9_63_0;
        mut_22_10_63_0 <= mut_22_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_76_cse = '1' ) THEN
        mut_1_10_63_0 <= mut_1_9_63_0;
        mut_10_63_0 <= mut_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_10_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_10_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( COMP_LOOP_and_78_cse = '1' ) THEN
        rem_12cyc_st_10_3_2 <= rem_12cyc_st_9_3_2;
        rem_12cyc_st_10_1_0 <= rem_12cyc_st_9_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_80_cse = '1' ) THEN
        mut_3_9_63_0 <= mut_3_8_63_0;
        mut_2_9_63_0 <= mut_2_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_82_cse = '1' ) THEN
        mut_5_9_63_0 <= mut_5_8_63_0;
        mut_4_9_63_0 <= mut_4_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_84_cse = '1' ) THEN
        mut_7_9_63_0 <= mut_7_8_63_0;
        mut_6_9_63_0 <= mut_6_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_86_cse = '1' ) THEN
        mut_9_9_63_0 <= mut_9_8_63_0;
        mut_8_9_63_0 <= mut_8_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_88_cse = '1' ) THEN
        mut_11_9_63_0 <= mut_11_8_63_0;
        mut_10_9_63_0 <= mut_10_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_90_cse = '1' ) THEN
        mut_13_9_63_0 <= mut_13_8_63_0;
        mut_12_9_63_0 <= mut_12_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_92_cse = '1' ) THEN
        mut_15_9_63_0 <= mut_15_8_63_0;
        mut_14_9_63_0 <= mut_14_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_94_cse = '1' ) THEN
        mut_17_9_63_0 <= mut_17_8_63_0;
        mut_16_9_63_0 <= mut_16_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_96_cse = '1' ) THEN
        mut_19_9_63_0 <= mut_19_8_63_0;
        mut_18_9_63_0 <= mut_18_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_98_cse = '1' ) THEN
        mut_21_9_63_0 <= mut_21_8_63_0;
        mut_20_9_63_0 <= mut_20_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_100_cse = '1' ) THEN
        mut_23_9_63_0 <= mut_23_8_63_0;
        mut_22_9_63_0 <= mut_22_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_102_cse = '1' ) THEN
        mut_1_9_63_0 <= mut_1_8_63_0;
        mut_9_63_0 <= mut_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_9_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_9_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( COMP_LOOP_and_104_cse = '1' ) THEN
        rem_12cyc_st_9_3_2 <= rem_12cyc_st_8_3_2;
        rem_12cyc_st_9_1_0 <= rem_12cyc_st_8_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_106_cse = '1' ) THEN
        mut_3_8_63_0 <= mut_3_7_63_0;
        mut_2_8_63_0 <= mut_2_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_108_cse = '1' ) THEN
        mut_5_8_63_0 <= mut_5_7_63_0;
        mut_4_8_63_0 <= mut_4_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_110_cse = '1' ) THEN
        mut_7_8_63_0 <= mut_7_7_63_0;
        mut_6_8_63_0 <= mut_6_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_112_cse = '1' ) THEN
        mut_9_8_63_0 <= mut_9_7_63_0;
        mut_8_8_63_0 <= mut_8_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_114_cse = '1' ) THEN
        mut_11_8_63_0 <= mut_11_7_63_0;
        mut_10_8_63_0 <= mut_10_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_116_cse = '1' ) THEN
        mut_13_8_63_0 <= mut_13_7_63_0;
        mut_12_8_63_0 <= mut_12_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_118_cse = '1' ) THEN
        mut_15_8_63_0 <= mut_15_7_63_0;
        mut_14_8_63_0 <= mut_14_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_120_cse = '1' ) THEN
        mut_17_8_63_0 <= mut_17_7_63_0;
        mut_16_8_63_0 <= mut_16_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_122_cse = '1' ) THEN
        mut_19_8_63_0 <= mut_19_7_63_0;
        mut_18_8_63_0 <= mut_18_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_124_cse = '1' ) THEN
        mut_21_8_63_0 <= mut_21_7_63_0;
        mut_20_8_63_0 <= mut_20_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_126_cse = '1' ) THEN
        mut_23_8_63_0 <= mut_23_7_63_0;
        mut_22_8_63_0 <= mut_22_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_128_cse = '1' ) THEN
        mut_1_8_63_0 <= mut_1_7_63_0;
        mut_8_63_0 <= mut_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_8_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_8_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( COMP_LOOP_and_130_cse = '1' ) THEN
        rem_12cyc_st_8_3_2 <= rem_12cyc_st_7_3_2;
        rem_12cyc_st_8_1_0 <= rem_12cyc_st_7_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_132_cse = '1' ) THEN
        mut_3_7_63_0 <= mut_3_6_63_0;
        mut_2_7_63_0 <= mut_2_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_134_cse = '1' ) THEN
        mut_5_7_63_0 <= mut_5_6_63_0;
        mut_4_7_63_0 <= mut_4_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_136_cse = '1' ) THEN
        mut_7_7_63_0 <= mut_7_6_63_0;
        mut_6_7_63_0 <= mut_6_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_138_cse = '1' ) THEN
        mut_9_7_63_0 <= mut_9_6_63_0;
        mut_8_7_63_0 <= mut_8_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_140_cse = '1' ) THEN
        mut_11_7_63_0 <= mut_11_6_63_0;
        mut_10_7_63_0 <= mut_10_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_142_cse = '1' ) THEN
        mut_13_7_63_0 <= mut_13_6_63_0;
        mut_12_7_63_0 <= mut_12_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_144_cse = '1' ) THEN
        mut_15_7_63_0 <= mut_15_6_63_0;
        mut_14_7_63_0 <= mut_14_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_146_cse = '1' ) THEN
        mut_17_7_63_0 <= mut_17_6_63_0;
        mut_16_7_63_0 <= mut_16_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_148_cse = '1' ) THEN
        mut_19_7_63_0 <= mut_19_6_63_0;
        mut_18_7_63_0 <= mut_18_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_150_cse = '1' ) THEN
        mut_21_7_63_0 <= mut_21_6_63_0;
        mut_20_7_63_0 <= mut_20_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_152_cse = '1' ) THEN
        mut_23_7_63_0 <= mut_23_6_63_0;
        mut_22_7_63_0 <= mut_22_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_154_cse = '1' ) THEN
        mut_1_7_63_0 <= mut_1_6_63_0;
        mut_7_63_0 <= mut_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_7_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_7_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( COMP_LOOP_and_156_cse = '1' ) THEN
        rem_12cyc_st_7_3_2 <= rem_12cyc_st_6_3_2;
        rem_12cyc_st_7_1_0 <= rem_12cyc_st_6_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_158_cse = '1' ) THEN
        mut_3_6_63_0 <= mut_3_5_63_0;
        mut_2_6_63_0 <= mut_2_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_160_cse = '1' ) THEN
        mut_5_6_63_0 <= mut_5_5_63_0;
        mut_4_6_63_0 <= mut_4_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_162_cse = '1' ) THEN
        mut_7_6_63_0 <= mut_7_5_63_0;
        mut_6_6_63_0 <= mut_6_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_164_cse = '1' ) THEN
        mut_9_6_63_0 <= mut_9_5_63_0;
        mut_8_6_63_0 <= mut_8_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_166_cse = '1' ) THEN
        mut_11_6_63_0 <= mut_11_5_63_0;
        mut_10_6_63_0 <= mut_10_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_168_cse = '1' ) THEN
        mut_13_6_63_0 <= mut_13_5_63_0;
        mut_12_6_63_0 <= mut_12_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_170_cse = '1' ) THEN
        mut_15_6_63_0 <= mut_15_5_63_0;
        mut_14_6_63_0 <= mut_14_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_172_cse = '1' ) THEN
        mut_17_6_63_0 <= mut_17_5_63_0;
        mut_16_6_63_0 <= mut_16_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_174_cse = '1' ) THEN
        mut_19_6_63_0 <= mut_19_5_63_0;
        mut_18_6_63_0 <= mut_18_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_176_cse = '1' ) THEN
        mut_21_6_63_0 <= mut_21_5_63_0;
        mut_20_6_63_0 <= mut_20_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_178_cse = '1' ) THEN
        mut_23_6_63_0 <= mut_23_5_63_0;
        mut_22_6_63_0 <= mut_22_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_180_cse = '1' ) THEN
        mut_1_6_63_0 <= mut_1_5_63_0;
        mut_6_63_0 <= mut_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_182_cse = '1' ) THEN
        m_buf_sva_6 <= m_buf_sva_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_6_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_6_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( COMP_LOOP_and_182_cse = '1' ) THEN
        rem_12cyc_st_6_3_2 <= rem_12cyc_st_5_3_2;
        rem_12cyc_st_6_1_0 <= rem_12cyc_st_5_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_184_cse = '1' ) THEN
        mut_3_5_63_0 <= mut_3_4_63_0;
        mut_2_5_63_0 <= mut_2_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_186_cse = '1' ) THEN
        mut_5_5_63_0 <= mut_5_4_63_0;
        mut_4_5_63_0 <= mut_4_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_188_cse = '1' ) THEN
        mut_7_5_63_0 <= mut_7_4_63_0;
        mut_6_5_63_0 <= mut_6_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_190_cse = '1' ) THEN
        mut_9_5_63_0 <= mut_9_4_63_0;
        mut_8_5_63_0 <= mut_8_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_192_cse = '1' ) THEN
        mut_11_5_63_0 <= mut_11_4_63_0;
        mut_10_5_63_0 <= mut_10_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_194_cse = '1' ) THEN
        mut_13_5_63_0 <= mut_13_4_63_0;
        mut_12_5_63_0 <= mut_12_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_196_cse = '1' ) THEN
        mut_15_5_63_0 <= mut_15_4_63_0;
        mut_14_5_63_0 <= mut_14_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_198_cse = '1' ) THEN
        mut_17_5_63_0 <= mut_17_4_63_0;
        mut_16_5_63_0 <= mut_16_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_200_cse = '1' ) THEN
        mut_19_5_63_0 <= mut_19_4_63_0;
        mut_18_5_63_0 <= mut_18_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_202_cse = '1' ) THEN
        mut_21_5_63_0 <= mut_21_4_63_0;
        mut_20_5_63_0 <= mut_20_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_204_cse = '1' ) THEN
        mut_23_5_63_0 <= mut_23_4_63_0;
        mut_22_5_63_0 <= mut_22_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_206_cse = '1' ) THEN
        mut_1_5_63_0 <= mut_1_4_63_0;
        mut_5_63_0 <= mut_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_208_cse = '1' ) THEN
        m_buf_sva_5 <= m_buf_sva_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_5_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_5_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( COMP_LOOP_and_208_cse = '1' ) THEN
        rem_12cyc_st_5_3_2 <= rem_12cyc_st_4_3_2;
        rem_12cyc_st_5_1_0 <= rem_12cyc_st_4_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_210_cse = '1' ) THEN
        mut_3_4_63_0 <= mut_3_3_63_0;
        mut_2_4_63_0 <= mut_2_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_212_cse = '1' ) THEN
        mut_5_4_63_0 <= mut_5_3_63_0;
        mut_4_4_63_0 <= mut_4_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_214_cse = '1' ) THEN
        mut_7_4_63_0 <= mut_7_3_63_0;
        mut_6_4_63_0 <= mut_6_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_216_cse = '1' ) THEN
        mut_9_4_63_0 <= mut_9_3_63_0;
        mut_8_4_63_0 <= mut_8_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_218_cse = '1' ) THEN
        mut_11_4_63_0 <= mut_11_3_63_0;
        mut_10_4_63_0 <= mut_10_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_220_cse = '1' ) THEN
        mut_13_4_63_0 <= mut_13_3_63_0;
        mut_12_4_63_0 <= mut_12_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_222_cse = '1' ) THEN
        mut_15_4_63_0 <= mut_15_3_63_0;
        mut_14_4_63_0 <= mut_14_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_224_cse = '1' ) THEN
        mut_17_4_63_0 <= mut_17_3_63_0;
        mut_16_4_63_0 <= mut_16_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_226_cse = '1' ) THEN
        mut_19_4_63_0 <= mut_19_3_63_0;
        mut_18_4_63_0 <= mut_18_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_228_cse = '1' ) THEN
        mut_21_4_63_0 <= mut_21_3_63_0;
        mut_20_4_63_0 <= mut_20_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_230_cse = '1' ) THEN
        mut_23_4_63_0 <= mut_23_3_63_0;
        mut_22_4_63_0 <= mut_22_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_232_cse = '1' ) THEN
        mut_1_4_63_0 <= mut_1_3_63_0;
        mut_4_63_0 <= mut_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_234_cse = '1' ) THEN
        m_buf_sva_4 <= m_buf_sva_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_4_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_4_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( COMP_LOOP_and_234_cse = '1' ) THEN
        rem_12cyc_st_4_3_2 <= rem_12cyc_st_3_3_2;
        rem_12cyc_st_4_1_0 <= rem_12cyc_st_3_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_236_cse = '1' ) THEN
        mut_3_3_63_0 <= mut_3_2_63_0;
        mut_2_3_63_0 <= mut_2_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_238_cse = '1' ) THEN
        mut_5_3_63_0 <= mut_5_2_63_0;
        mut_4_3_63_0 <= mut_4_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_240_cse = '1' ) THEN
        mut_7_3_63_0 <= mut_7_2_63_0;
        mut_6_3_63_0 <= mut_6_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_242_cse = '1' ) THEN
        mut_9_3_63_0 <= mut_9_2_63_0;
        mut_8_3_63_0 <= mut_8_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_244_cse = '1' ) THEN
        mut_11_3_63_0 <= mut_11_2_63_0;
        mut_10_3_63_0 <= mut_10_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_246_cse = '1' ) THEN
        mut_13_3_63_0 <= mut_13_2_63_0;
        mut_12_3_63_0 <= mut_12_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_248_cse = '1' ) THEN
        mut_15_3_63_0 <= mut_15_2_63_0;
        mut_14_3_63_0 <= mut_14_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_250_cse = '1' ) THEN
        mut_17_3_63_0 <= mut_17_2_63_0;
        mut_16_3_63_0 <= mut_16_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_252_cse = '1' ) THEN
        mut_19_3_63_0 <= mut_19_2_63_0;
        mut_18_3_63_0 <= mut_18_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_254_cse = '1' ) THEN
        mut_21_3_63_0 <= mut_21_2_63_0;
        mut_20_3_63_0 <= mut_20_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_256_cse = '1' ) THEN
        mut_23_3_63_0 <= mut_23_2_63_0;
        mut_22_3_63_0 <= mut_22_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_258_cse = '1' ) THEN
        mut_1_3_63_0 <= mut_1_2_63_0;
        mut_3_63_0 <= mut_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_260_cse = '1' ) THEN
        m_buf_sva_3 <= m_buf_sva_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_3_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_3_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( COMP_LOOP_and_260_cse = '1' ) THEN
        rem_12cyc_st_3_3_2 <= rem_12cyc_st_2_3_2;
        rem_12cyc_st_3_1_0 <= rem_12cyc_st_2_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_262_cse = '1' ) THEN
        mut_3_2_63_0 <= rem_12_cmp_1_b_63_0;
        mut_2_2_63_0 <= rem_12_cmp_1_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_264_cse = '1' ) THEN
        mut_5_2_63_0 <= rem_12_cmp_2_b_63_0;
        mut_4_2_63_0 <= rem_12_cmp_2_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_266_cse = '1' ) THEN
        mut_7_2_63_0 <= rem_12_cmp_3_b_63_0;
        mut_6_2_63_0 <= rem_12_cmp_3_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_268_cse = '1' ) THEN
        mut_9_2_63_0 <= rem_12_cmp_4_b_63_0;
        mut_8_2_63_0 <= rem_12_cmp_4_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_270_cse = '1' ) THEN
        mut_11_2_63_0 <= rem_12_cmp_5_b_63_0;
        mut_10_2_63_0 <= rem_12_cmp_5_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_272_cse = '1' ) THEN
        mut_13_2_63_0 <= rem_12_cmp_6_b_63_0;
        mut_12_2_63_0 <= rem_12_cmp_6_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_274_cse = '1' ) THEN
        mut_15_2_63_0 <= rem_12_cmp_7_b_63_0;
        mut_14_2_63_0 <= rem_12_cmp_7_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_276_cse = '1' ) THEN
        mut_17_2_63_0 <= rem_12_cmp_8_b_63_0;
        mut_16_2_63_0 <= rem_12_cmp_8_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_278_cse = '1' ) THEN
        mut_19_2_63_0 <= rem_12_cmp_9_b_63_0;
        mut_18_2_63_0 <= rem_12_cmp_9_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_280_cse = '1' ) THEN
        mut_21_2_63_0 <= rem_12_cmp_10_b_63_0;
        mut_20_2_63_0 <= rem_12_cmp_10_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_282_cse = '1' ) THEN
        mut_23_2_63_0 <= rem_12_cmp_11_b_63_0;
        mut_22_2_63_0 <= rem_12_cmp_11_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_284_cse = '1' ) THEN
        mut_1_2_63_0 <= rem_12_cmp_b_63_0;
        mut_2_63_0 <= rem_12_cmp_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_286_cse = '1' ) THEN
        m_buf_sva_2 <= m_buf_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_2_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_2_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( COMP_LOOP_and_286_cse = '1' ) THEN
        rem_12cyc_st_2_3_2 <= rem_12cyc_3_2;
        rem_12cyc_st_2_1_0 <= rem_12cyc_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( COMP_LOOP_and_24_cse = '1' ) THEN
        m_buf_sva_1 <= m_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( COMP_LOOP_and_24_cse = '1' ) THEN
        rem_12cyc_3_2 <= COMP_LOOP_acc_tmp;
        rem_12cyc_1_0 <= COMP_LOOP_acc_1_tmp(1 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  qelse_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(result_sva_duc_mx0) + UNSIGNED(m_buf_sva_12),
      64));
  mux_8_nl <= MUX_s_1_2_2((rem_12_cmp_1_z(63)), (rem_12_cmp_3_z(63)), rem_12cyc_st_12_1_0(1));
  mux_7_nl <= MUX_s_1_2_2((rem_12_cmp_2_z(63)), (rem_12_cmp_4_z(63)), rem_12cyc_st_12_1_0(1));
  mux_9_nl <= MUX_s_1_2_2(mux_8_nl, mux_7_nl, rem_12cyc_st_12_1_0(0));
  mux_5_nl <= MUX_s_1_2_2((rem_12_cmp_9_z(63)), (rem_12_cmp_11_z(63)), rem_12cyc_st_12_1_0(1));
  mux_4_nl <= MUX_s_1_2_2((rem_12_cmp_10_z(63)), (rem_12_cmp_z(63)), rem_12cyc_st_12_1_0(1));
  mux_6_nl <= MUX_s_1_2_2(mux_5_nl, mux_4_nl, rem_12cyc_st_12_1_0(0));
  mux_10_nl <= MUX_s_1_2_2(mux_9_nl, mux_6_nl, rem_12cyc_st_12_3_2(1));
  mux_1_nl <= MUX_s_1_2_2((rem_12_cmp_5_z(63)), (rem_12_cmp_7_z(63)), rem_12cyc_st_12_1_0(1));
  mux_nl <= MUX_s_1_2_2((rem_12_cmp_6_z(63)), (rem_12_cmp_8_z(63)), rem_12cyc_st_12_1_0(1));
  mux_2_nl <= MUX_s_1_2_2(mux_1_nl, mux_nl, rem_12cyc_st_12_1_0(0));
  mux_3_nl <= MUX_s_1_2_2(mux_2_nl, (result_sva_duc(63)), rem_12cyc_st_12_3_2(1));
  mux_11_nl <= MUX_s_1_2_2(mux_10_nl, mux_3_nl, rem_12cyc_st_12_3_2(0));
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    modulo
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;
USE work.mgc_comps.ALL;


ENTITY modulo IS
  PORT(
    base_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    m_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    return_rsc_z : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    ccs_ccore_start_rsc_dat : IN STD_LOGIC;
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_srst : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC
  );
END modulo;

ARCHITECTURE v1 OF modulo IS
  -- Default Constants

  COMPONENT modulo_core
    PORT(
      base_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      m_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      return_rsc_z : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      ccs_ccore_start_rsc_dat : IN STD_LOGIC;
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_srst : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL modulo_core_inst_base_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_core_inst_m_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_core_inst_return_rsc_z : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  modulo_core_inst : modulo_core
    PORT MAP(
      base_rsc_dat => modulo_core_inst_base_rsc_dat,
      m_rsc_dat => modulo_core_inst_m_rsc_dat,
      return_rsc_z => modulo_core_inst_return_rsc_z,
      ccs_ccore_start_rsc_dat => ccs_ccore_start_rsc_dat,
      ccs_ccore_clk => ccs_ccore_clk,
      ccs_ccore_srst => ccs_ccore_srst,
      ccs_ccore_en => ccs_ccore_en
    );
  modulo_core_inst_base_rsc_dat <= base_rsc_dat;
  modulo_core_inst_m_rsc_dat <= m_rsc_dat;
  return_rsc_z <= modulo_core_inst_return_rsc_z;

END v1;




--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_comps_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_shift_comps_v5 IS

COMPONENT mgc_shift_l_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_shift_comps_v5;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_shift_l_v5 IS
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_shift_l_v5;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_shift_l_v5 IS

  FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1 > arg2) THEN
      RETURN(arg1) ;
    ELSE
      RETURN(arg2) ;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(SIGNED(result), arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE)
  RETURN UNSIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, '0', olen);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE)
  RETURN SIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen);
  END;

BEGIN
UNSGNED:  IF signd_a = 0 GENERATE
    z <= std_logic_vector(fshl_stdar(unsigned(a), unsigned(s), width_z));
  END GENERATE;
SGNED:  IF signd_a /= 0 GENERATE
    z <= std_logic_vector(fshl_stdar(  signed(a), unsigned(s), width_z));
  END GENERATE;
END beh;

--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Mon Aug  2 20:57:22 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_40_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_40_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_40_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_40_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_39_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_39_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_39_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_39_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_38_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_38_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_38_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_38_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_37_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_37_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_37_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_37_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_36_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_36_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_36_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_36_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_35_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_35_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_35_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_35_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_34_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_34_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_34_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_34_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_33_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_33_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_33_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_33_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_32_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_32_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_32_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_32_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_31_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_31_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_31_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_31_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_30_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_30_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_30_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_30_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_29_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_29_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_29_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_29_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_28_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_28_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_28_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_28_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_27_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_27_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_27_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_27_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_26_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_26_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_26_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_26_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_25_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_25_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_25_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_25_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen;

ARCHITECTURE v7 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
    COMP_LOOP_C_31_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_62_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_93_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_124_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_155_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_186_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_217_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_248_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_279_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_310_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_341_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_372_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_403_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_434_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_465_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_496_tr0 : IN STD_LOGIC;
    VEC_LOOP_C_0_tr0 : IN STD_LOGIC;
    STAGE_LOOP_C_1_tr0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_core_core_fsm;

ARCHITECTURE v7 OF inPlaceNTT_DIF_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for inPlaceNTT_DIF_core_core_fsm_1
  TYPE inPlaceNTT_DIF_core_core_fsm_1_ST IS (main_C_0, STAGE_LOOP_C_0, COMP_LOOP_C_0,
      COMP_LOOP_C_1, COMP_LOOP_C_2, COMP_LOOP_C_3, COMP_LOOP_C_4, COMP_LOOP_C_5,
      COMP_LOOP_C_6, COMP_LOOP_C_7, COMP_LOOP_C_8, COMP_LOOP_C_9, COMP_LOOP_C_10,
      COMP_LOOP_C_11, COMP_LOOP_C_12, COMP_LOOP_C_13, COMP_LOOP_C_14, COMP_LOOP_C_15,
      COMP_LOOP_C_16, COMP_LOOP_C_17, COMP_LOOP_C_18, COMP_LOOP_C_19, COMP_LOOP_C_20,
      COMP_LOOP_C_21, COMP_LOOP_C_22, COMP_LOOP_C_23, COMP_LOOP_C_24, COMP_LOOP_C_25,
      COMP_LOOP_C_26, COMP_LOOP_C_27, COMP_LOOP_C_28, COMP_LOOP_C_29, COMP_LOOP_C_30,
      COMP_LOOP_C_31, COMP_LOOP_C_32, COMP_LOOP_C_33, COMP_LOOP_C_34, COMP_LOOP_C_35,
      COMP_LOOP_C_36, COMP_LOOP_C_37, COMP_LOOP_C_38, COMP_LOOP_C_39, COMP_LOOP_C_40,
      COMP_LOOP_C_41, COMP_LOOP_C_42, COMP_LOOP_C_43, COMP_LOOP_C_44, COMP_LOOP_C_45,
      COMP_LOOP_C_46, COMP_LOOP_C_47, COMP_LOOP_C_48, COMP_LOOP_C_49, COMP_LOOP_C_50,
      COMP_LOOP_C_51, COMP_LOOP_C_52, COMP_LOOP_C_53, COMP_LOOP_C_54, COMP_LOOP_C_55,
      COMP_LOOP_C_56, COMP_LOOP_C_57, COMP_LOOP_C_58, COMP_LOOP_C_59, COMP_LOOP_C_60,
      COMP_LOOP_C_61, COMP_LOOP_C_62, COMP_LOOP_C_63, COMP_LOOP_C_64, COMP_LOOP_C_65,
      COMP_LOOP_C_66, COMP_LOOP_C_67, COMP_LOOP_C_68, COMP_LOOP_C_69, COMP_LOOP_C_70,
      COMP_LOOP_C_71, COMP_LOOP_C_72, COMP_LOOP_C_73, COMP_LOOP_C_74, COMP_LOOP_C_75,
      COMP_LOOP_C_76, COMP_LOOP_C_77, COMP_LOOP_C_78, COMP_LOOP_C_79, COMP_LOOP_C_80,
      COMP_LOOP_C_81, COMP_LOOP_C_82, COMP_LOOP_C_83, COMP_LOOP_C_84, COMP_LOOP_C_85,
      COMP_LOOP_C_86, COMP_LOOP_C_87, COMP_LOOP_C_88, COMP_LOOP_C_89, COMP_LOOP_C_90,
      COMP_LOOP_C_91, COMP_LOOP_C_92, COMP_LOOP_C_93, COMP_LOOP_C_94, COMP_LOOP_C_95,
      COMP_LOOP_C_96, COMP_LOOP_C_97, COMP_LOOP_C_98, COMP_LOOP_C_99, COMP_LOOP_C_100,
      COMP_LOOP_C_101, COMP_LOOP_C_102, COMP_LOOP_C_103, COMP_LOOP_C_104, COMP_LOOP_C_105,
      COMP_LOOP_C_106, COMP_LOOP_C_107, COMP_LOOP_C_108, COMP_LOOP_C_109, COMP_LOOP_C_110,
      COMP_LOOP_C_111, COMP_LOOP_C_112, COMP_LOOP_C_113, COMP_LOOP_C_114, COMP_LOOP_C_115,
      COMP_LOOP_C_116, COMP_LOOP_C_117, COMP_LOOP_C_118, COMP_LOOP_C_119, COMP_LOOP_C_120,
      COMP_LOOP_C_121, COMP_LOOP_C_122, COMP_LOOP_C_123, COMP_LOOP_C_124, COMP_LOOP_C_125,
      COMP_LOOP_C_126, COMP_LOOP_C_127, COMP_LOOP_C_128, COMP_LOOP_C_129, COMP_LOOP_C_130,
      COMP_LOOP_C_131, COMP_LOOP_C_132, COMP_LOOP_C_133, COMP_LOOP_C_134, COMP_LOOP_C_135,
      COMP_LOOP_C_136, COMP_LOOP_C_137, COMP_LOOP_C_138, COMP_LOOP_C_139, COMP_LOOP_C_140,
      COMP_LOOP_C_141, COMP_LOOP_C_142, COMP_LOOP_C_143, COMP_LOOP_C_144, COMP_LOOP_C_145,
      COMP_LOOP_C_146, COMP_LOOP_C_147, COMP_LOOP_C_148, COMP_LOOP_C_149, COMP_LOOP_C_150,
      COMP_LOOP_C_151, COMP_LOOP_C_152, COMP_LOOP_C_153, COMP_LOOP_C_154, COMP_LOOP_C_155,
      COMP_LOOP_C_156, COMP_LOOP_C_157, COMP_LOOP_C_158, COMP_LOOP_C_159, COMP_LOOP_C_160,
      COMP_LOOP_C_161, COMP_LOOP_C_162, COMP_LOOP_C_163, COMP_LOOP_C_164, COMP_LOOP_C_165,
      COMP_LOOP_C_166, COMP_LOOP_C_167, COMP_LOOP_C_168, COMP_LOOP_C_169, COMP_LOOP_C_170,
      COMP_LOOP_C_171, COMP_LOOP_C_172, COMP_LOOP_C_173, COMP_LOOP_C_174, COMP_LOOP_C_175,
      COMP_LOOP_C_176, COMP_LOOP_C_177, COMP_LOOP_C_178, COMP_LOOP_C_179, COMP_LOOP_C_180,
      COMP_LOOP_C_181, COMP_LOOP_C_182, COMP_LOOP_C_183, COMP_LOOP_C_184, COMP_LOOP_C_185,
      COMP_LOOP_C_186, COMP_LOOP_C_187, COMP_LOOP_C_188, COMP_LOOP_C_189, COMP_LOOP_C_190,
      COMP_LOOP_C_191, COMP_LOOP_C_192, COMP_LOOP_C_193, COMP_LOOP_C_194, COMP_LOOP_C_195,
      COMP_LOOP_C_196, COMP_LOOP_C_197, COMP_LOOP_C_198, COMP_LOOP_C_199, COMP_LOOP_C_200,
      COMP_LOOP_C_201, COMP_LOOP_C_202, COMP_LOOP_C_203, COMP_LOOP_C_204, COMP_LOOP_C_205,
      COMP_LOOP_C_206, COMP_LOOP_C_207, COMP_LOOP_C_208, COMP_LOOP_C_209, COMP_LOOP_C_210,
      COMP_LOOP_C_211, COMP_LOOP_C_212, COMP_LOOP_C_213, COMP_LOOP_C_214, COMP_LOOP_C_215,
      COMP_LOOP_C_216, COMP_LOOP_C_217, COMP_LOOP_C_218, COMP_LOOP_C_219, COMP_LOOP_C_220,
      COMP_LOOP_C_221, COMP_LOOP_C_222, COMP_LOOP_C_223, COMP_LOOP_C_224, COMP_LOOP_C_225,
      COMP_LOOP_C_226, COMP_LOOP_C_227, COMP_LOOP_C_228, COMP_LOOP_C_229, COMP_LOOP_C_230,
      COMP_LOOP_C_231, COMP_LOOP_C_232, COMP_LOOP_C_233, COMP_LOOP_C_234, COMP_LOOP_C_235,
      COMP_LOOP_C_236, COMP_LOOP_C_237, COMP_LOOP_C_238, COMP_LOOP_C_239, COMP_LOOP_C_240,
      COMP_LOOP_C_241, COMP_LOOP_C_242, COMP_LOOP_C_243, COMP_LOOP_C_244, COMP_LOOP_C_245,
      COMP_LOOP_C_246, COMP_LOOP_C_247, COMP_LOOP_C_248, COMP_LOOP_C_249, COMP_LOOP_C_250,
      COMP_LOOP_C_251, COMP_LOOP_C_252, COMP_LOOP_C_253, COMP_LOOP_C_254, COMP_LOOP_C_255,
      COMP_LOOP_C_256, COMP_LOOP_C_257, COMP_LOOP_C_258, COMP_LOOP_C_259, COMP_LOOP_C_260,
      COMP_LOOP_C_261, COMP_LOOP_C_262, COMP_LOOP_C_263, COMP_LOOP_C_264, COMP_LOOP_C_265,
      COMP_LOOP_C_266, COMP_LOOP_C_267, COMP_LOOP_C_268, COMP_LOOP_C_269, COMP_LOOP_C_270,
      COMP_LOOP_C_271, COMP_LOOP_C_272, COMP_LOOP_C_273, COMP_LOOP_C_274, COMP_LOOP_C_275,
      COMP_LOOP_C_276, COMP_LOOP_C_277, COMP_LOOP_C_278, COMP_LOOP_C_279, COMP_LOOP_C_280,
      COMP_LOOP_C_281, COMP_LOOP_C_282, COMP_LOOP_C_283, COMP_LOOP_C_284, COMP_LOOP_C_285,
      COMP_LOOP_C_286, COMP_LOOP_C_287, COMP_LOOP_C_288, COMP_LOOP_C_289, COMP_LOOP_C_290,
      COMP_LOOP_C_291, COMP_LOOP_C_292, COMP_LOOP_C_293, COMP_LOOP_C_294, COMP_LOOP_C_295,
      COMP_LOOP_C_296, COMP_LOOP_C_297, COMP_LOOP_C_298, COMP_LOOP_C_299, COMP_LOOP_C_300,
      COMP_LOOP_C_301, COMP_LOOP_C_302, COMP_LOOP_C_303, COMP_LOOP_C_304, COMP_LOOP_C_305,
      COMP_LOOP_C_306, COMP_LOOP_C_307, COMP_LOOP_C_308, COMP_LOOP_C_309, COMP_LOOP_C_310,
      COMP_LOOP_C_311, COMP_LOOP_C_312, COMP_LOOP_C_313, COMP_LOOP_C_314, COMP_LOOP_C_315,
      COMP_LOOP_C_316, COMP_LOOP_C_317, COMP_LOOP_C_318, COMP_LOOP_C_319, COMP_LOOP_C_320,
      COMP_LOOP_C_321, COMP_LOOP_C_322, COMP_LOOP_C_323, COMP_LOOP_C_324, COMP_LOOP_C_325,
      COMP_LOOP_C_326, COMP_LOOP_C_327, COMP_LOOP_C_328, COMP_LOOP_C_329, COMP_LOOP_C_330,
      COMP_LOOP_C_331, COMP_LOOP_C_332, COMP_LOOP_C_333, COMP_LOOP_C_334, COMP_LOOP_C_335,
      COMP_LOOP_C_336, COMP_LOOP_C_337, COMP_LOOP_C_338, COMP_LOOP_C_339, COMP_LOOP_C_340,
      COMP_LOOP_C_341, COMP_LOOP_C_342, COMP_LOOP_C_343, COMP_LOOP_C_344, COMP_LOOP_C_345,
      COMP_LOOP_C_346, COMP_LOOP_C_347, COMP_LOOP_C_348, COMP_LOOP_C_349, COMP_LOOP_C_350,
      COMP_LOOP_C_351, COMP_LOOP_C_352, COMP_LOOP_C_353, COMP_LOOP_C_354, COMP_LOOP_C_355,
      COMP_LOOP_C_356, COMP_LOOP_C_357, COMP_LOOP_C_358, COMP_LOOP_C_359, COMP_LOOP_C_360,
      COMP_LOOP_C_361, COMP_LOOP_C_362, COMP_LOOP_C_363, COMP_LOOP_C_364, COMP_LOOP_C_365,
      COMP_LOOP_C_366, COMP_LOOP_C_367, COMP_LOOP_C_368, COMP_LOOP_C_369, COMP_LOOP_C_370,
      COMP_LOOP_C_371, COMP_LOOP_C_372, COMP_LOOP_C_373, COMP_LOOP_C_374, COMP_LOOP_C_375,
      COMP_LOOP_C_376, COMP_LOOP_C_377, COMP_LOOP_C_378, COMP_LOOP_C_379, COMP_LOOP_C_380,
      COMP_LOOP_C_381, COMP_LOOP_C_382, COMP_LOOP_C_383, COMP_LOOP_C_384, COMP_LOOP_C_385,
      COMP_LOOP_C_386, COMP_LOOP_C_387, COMP_LOOP_C_388, COMP_LOOP_C_389, COMP_LOOP_C_390,
      COMP_LOOP_C_391, COMP_LOOP_C_392, COMP_LOOP_C_393, COMP_LOOP_C_394, COMP_LOOP_C_395,
      COMP_LOOP_C_396, COMP_LOOP_C_397, COMP_LOOP_C_398, COMP_LOOP_C_399, COMP_LOOP_C_400,
      COMP_LOOP_C_401, COMP_LOOP_C_402, COMP_LOOP_C_403, COMP_LOOP_C_404, COMP_LOOP_C_405,
      COMP_LOOP_C_406, COMP_LOOP_C_407, COMP_LOOP_C_408, COMP_LOOP_C_409, COMP_LOOP_C_410,
      COMP_LOOP_C_411, COMP_LOOP_C_412, COMP_LOOP_C_413, COMP_LOOP_C_414, COMP_LOOP_C_415,
      COMP_LOOP_C_416, COMP_LOOP_C_417, COMP_LOOP_C_418, COMP_LOOP_C_419, COMP_LOOP_C_420,
      COMP_LOOP_C_421, COMP_LOOP_C_422, COMP_LOOP_C_423, COMP_LOOP_C_424, COMP_LOOP_C_425,
      COMP_LOOP_C_426, COMP_LOOP_C_427, COMP_LOOP_C_428, COMP_LOOP_C_429, COMP_LOOP_C_430,
      COMP_LOOP_C_431, COMP_LOOP_C_432, COMP_LOOP_C_433, COMP_LOOP_C_434, COMP_LOOP_C_435,
      COMP_LOOP_C_436, COMP_LOOP_C_437, COMP_LOOP_C_438, COMP_LOOP_C_439, COMP_LOOP_C_440,
      COMP_LOOP_C_441, COMP_LOOP_C_442, COMP_LOOP_C_443, COMP_LOOP_C_444, COMP_LOOP_C_445,
      COMP_LOOP_C_446, COMP_LOOP_C_447, COMP_LOOP_C_448, COMP_LOOP_C_449, COMP_LOOP_C_450,
      COMP_LOOP_C_451, COMP_LOOP_C_452, COMP_LOOP_C_453, COMP_LOOP_C_454, COMP_LOOP_C_455,
      COMP_LOOP_C_456, COMP_LOOP_C_457, COMP_LOOP_C_458, COMP_LOOP_C_459, COMP_LOOP_C_460,
      COMP_LOOP_C_461, COMP_LOOP_C_462, COMP_LOOP_C_463, COMP_LOOP_C_464, COMP_LOOP_C_465,
      COMP_LOOP_C_466, COMP_LOOP_C_467, COMP_LOOP_C_468, COMP_LOOP_C_469, COMP_LOOP_C_470,
      COMP_LOOP_C_471, COMP_LOOP_C_472, COMP_LOOP_C_473, COMP_LOOP_C_474, COMP_LOOP_C_475,
      COMP_LOOP_C_476, COMP_LOOP_C_477, COMP_LOOP_C_478, COMP_LOOP_C_479, COMP_LOOP_C_480,
      COMP_LOOP_C_481, COMP_LOOP_C_482, COMP_LOOP_C_483, COMP_LOOP_C_484, COMP_LOOP_C_485,
      COMP_LOOP_C_486, COMP_LOOP_C_487, COMP_LOOP_C_488, COMP_LOOP_C_489, COMP_LOOP_C_490,
      COMP_LOOP_C_491, COMP_LOOP_C_492, COMP_LOOP_C_493, COMP_LOOP_C_494, COMP_LOOP_C_495,
      COMP_LOOP_C_496, VEC_LOOP_C_0, STAGE_LOOP_C_1, main_C_1);

  SIGNAL state_var : inPlaceNTT_DIF_core_core_fsm_1_ST;
  SIGNAL state_var_NS : inPlaceNTT_DIF_core_core_fsm_1_ST;

BEGIN
  inPlaceNTT_DIF_core_core_fsm_1 : PROCESS (COMP_LOOP_C_31_tr0, COMP_LOOP_C_62_tr0,
      COMP_LOOP_C_93_tr0, COMP_LOOP_C_124_tr0, COMP_LOOP_C_155_tr0, COMP_LOOP_C_186_tr0,
      COMP_LOOP_C_217_tr0, COMP_LOOP_C_248_tr0, COMP_LOOP_C_279_tr0, COMP_LOOP_C_310_tr0,
      COMP_LOOP_C_341_tr0, COMP_LOOP_C_372_tr0, COMP_LOOP_C_403_tr0, COMP_LOOP_C_434_tr0,
      COMP_LOOP_C_465_tr0, COMP_LOOP_C_496_tr0, VEC_LOOP_C_0_tr0, STAGE_LOOP_C_1_tr0,
      state_var)
  BEGIN
    CASE state_var IS
      WHEN STAGE_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000000001");
        state_var_NS <= COMP_LOOP_C_0;
      WHEN COMP_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000000010");
        state_var_NS <= COMP_LOOP_C_1;
      WHEN COMP_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000000011");
        state_var_NS <= COMP_LOOP_C_2;
      WHEN COMP_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000000100");
        state_var_NS <= COMP_LOOP_C_3;
      WHEN COMP_LOOP_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000000101");
        state_var_NS <= COMP_LOOP_C_4;
      WHEN COMP_LOOP_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000000110");
        state_var_NS <= COMP_LOOP_C_5;
      WHEN COMP_LOOP_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000000111");
        state_var_NS <= COMP_LOOP_C_6;
      WHEN COMP_LOOP_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000001000");
        state_var_NS <= COMP_LOOP_C_7;
      WHEN COMP_LOOP_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000001001");
        state_var_NS <= COMP_LOOP_C_8;
      WHEN COMP_LOOP_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000001010");
        state_var_NS <= COMP_LOOP_C_9;
      WHEN COMP_LOOP_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000001011");
        state_var_NS <= COMP_LOOP_C_10;
      WHEN COMP_LOOP_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000001100");
        state_var_NS <= COMP_LOOP_C_11;
      WHEN COMP_LOOP_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000001101");
        state_var_NS <= COMP_LOOP_C_12;
      WHEN COMP_LOOP_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000001110");
        state_var_NS <= COMP_LOOP_C_13;
      WHEN COMP_LOOP_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000001111");
        state_var_NS <= COMP_LOOP_C_14;
      WHEN COMP_LOOP_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000010000");
        state_var_NS <= COMP_LOOP_C_15;
      WHEN COMP_LOOP_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000010001");
        state_var_NS <= COMP_LOOP_C_16;
      WHEN COMP_LOOP_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000010010");
        state_var_NS <= COMP_LOOP_C_17;
      WHEN COMP_LOOP_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000010011");
        state_var_NS <= COMP_LOOP_C_18;
      WHEN COMP_LOOP_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000010100");
        state_var_NS <= COMP_LOOP_C_19;
      WHEN COMP_LOOP_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000010101");
        state_var_NS <= COMP_LOOP_C_20;
      WHEN COMP_LOOP_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000010110");
        state_var_NS <= COMP_LOOP_C_21;
      WHEN COMP_LOOP_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000010111");
        state_var_NS <= COMP_LOOP_C_22;
      WHEN COMP_LOOP_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000011000");
        state_var_NS <= COMP_LOOP_C_23;
      WHEN COMP_LOOP_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000011001");
        state_var_NS <= COMP_LOOP_C_24;
      WHEN COMP_LOOP_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000011010");
        state_var_NS <= COMP_LOOP_C_25;
      WHEN COMP_LOOP_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000011011");
        state_var_NS <= COMP_LOOP_C_26;
      WHEN COMP_LOOP_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000011100");
        state_var_NS <= COMP_LOOP_C_27;
      WHEN COMP_LOOP_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000011101");
        state_var_NS <= COMP_LOOP_C_28;
      WHEN COMP_LOOP_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000011110");
        state_var_NS <= COMP_LOOP_C_29;
      WHEN COMP_LOOP_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000011111");
        state_var_NS <= COMP_LOOP_C_30;
      WHEN COMP_LOOP_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000100000");
        state_var_NS <= COMP_LOOP_C_31;
      WHEN COMP_LOOP_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000100001");
        IF ( COMP_LOOP_C_31_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_32;
        END IF;
      WHEN COMP_LOOP_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000100010");
        state_var_NS <= COMP_LOOP_C_33;
      WHEN COMP_LOOP_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000100011");
        state_var_NS <= COMP_LOOP_C_34;
      WHEN COMP_LOOP_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000100100");
        state_var_NS <= COMP_LOOP_C_35;
      WHEN COMP_LOOP_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000100101");
        state_var_NS <= COMP_LOOP_C_36;
      WHEN COMP_LOOP_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000100110");
        state_var_NS <= COMP_LOOP_C_37;
      WHEN COMP_LOOP_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000100111");
        state_var_NS <= COMP_LOOP_C_38;
      WHEN COMP_LOOP_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000101000");
        state_var_NS <= COMP_LOOP_C_39;
      WHEN COMP_LOOP_C_39 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000101001");
        state_var_NS <= COMP_LOOP_C_40;
      WHEN COMP_LOOP_C_40 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000101010");
        state_var_NS <= COMP_LOOP_C_41;
      WHEN COMP_LOOP_C_41 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000101011");
        state_var_NS <= COMP_LOOP_C_42;
      WHEN COMP_LOOP_C_42 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000101100");
        state_var_NS <= COMP_LOOP_C_43;
      WHEN COMP_LOOP_C_43 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000101101");
        state_var_NS <= COMP_LOOP_C_44;
      WHEN COMP_LOOP_C_44 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000101110");
        state_var_NS <= COMP_LOOP_C_45;
      WHEN COMP_LOOP_C_45 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000101111");
        state_var_NS <= COMP_LOOP_C_46;
      WHEN COMP_LOOP_C_46 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000110000");
        state_var_NS <= COMP_LOOP_C_47;
      WHEN COMP_LOOP_C_47 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000110001");
        state_var_NS <= COMP_LOOP_C_48;
      WHEN COMP_LOOP_C_48 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000110010");
        state_var_NS <= COMP_LOOP_C_49;
      WHEN COMP_LOOP_C_49 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000110011");
        state_var_NS <= COMP_LOOP_C_50;
      WHEN COMP_LOOP_C_50 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000110100");
        state_var_NS <= COMP_LOOP_C_51;
      WHEN COMP_LOOP_C_51 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000110101");
        state_var_NS <= COMP_LOOP_C_52;
      WHEN COMP_LOOP_C_52 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000110110");
        state_var_NS <= COMP_LOOP_C_53;
      WHEN COMP_LOOP_C_53 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000110111");
        state_var_NS <= COMP_LOOP_C_54;
      WHEN COMP_LOOP_C_54 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000111000");
        state_var_NS <= COMP_LOOP_C_55;
      WHEN COMP_LOOP_C_55 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000111001");
        state_var_NS <= COMP_LOOP_C_56;
      WHEN COMP_LOOP_C_56 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000111010");
        state_var_NS <= COMP_LOOP_C_57;
      WHEN COMP_LOOP_C_57 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000111011");
        state_var_NS <= COMP_LOOP_C_58;
      WHEN COMP_LOOP_C_58 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000111100");
        state_var_NS <= COMP_LOOP_C_59;
      WHEN COMP_LOOP_C_59 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000111101");
        state_var_NS <= COMP_LOOP_C_60;
      WHEN COMP_LOOP_C_60 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000111110");
        state_var_NS <= COMP_LOOP_C_61;
      WHEN COMP_LOOP_C_61 =>
        fsm_output <= STD_LOGIC_VECTOR'( "000111111");
        state_var_NS <= COMP_LOOP_C_62;
      WHEN COMP_LOOP_C_62 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001000000");
        IF ( COMP_LOOP_C_62_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_63;
        END IF;
      WHEN COMP_LOOP_C_63 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001000001");
        state_var_NS <= COMP_LOOP_C_64;
      WHEN COMP_LOOP_C_64 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001000010");
        state_var_NS <= COMP_LOOP_C_65;
      WHEN COMP_LOOP_C_65 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001000011");
        state_var_NS <= COMP_LOOP_C_66;
      WHEN COMP_LOOP_C_66 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001000100");
        state_var_NS <= COMP_LOOP_C_67;
      WHEN COMP_LOOP_C_67 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001000101");
        state_var_NS <= COMP_LOOP_C_68;
      WHEN COMP_LOOP_C_68 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001000110");
        state_var_NS <= COMP_LOOP_C_69;
      WHEN COMP_LOOP_C_69 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001000111");
        state_var_NS <= COMP_LOOP_C_70;
      WHEN COMP_LOOP_C_70 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001001000");
        state_var_NS <= COMP_LOOP_C_71;
      WHEN COMP_LOOP_C_71 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001001001");
        state_var_NS <= COMP_LOOP_C_72;
      WHEN COMP_LOOP_C_72 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001001010");
        state_var_NS <= COMP_LOOP_C_73;
      WHEN COMP_LOOP_C_73 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001001011");
        state_var_NS <= COMP_LOOP_C_74;
      WHEN COMP_LOOP_C_74 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001001100");
        state_var_NS <= COMP_LOOP_C_75;
      WHEN COMP_LOOP_C_75 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001001101");
        state_var_NS <= COMP_LOOP_C_76;
      WHEN COMP_LOOP_C_76 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001001110");
        state_var_NS <= COMP_LOOP_C_77;
      WHEN COMP_LOOP_C_77 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001001111");
        state_var_NS <= COMP_LOOP_C_78;
      WHEN COMP_LOOP_C_78 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001010000");
        state_var_NS <= COMP_LOOP_C_79;
      WHEN COMP_LOOP_C_79 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001010001");
        state_var_NS <= COMP_LOOP_C_80;
      WHEN COMP_LOOP_C_80 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001010010");
        state_var_NS <= COMP_LOOP_C_81;
      WHEN COMP_LOOP_C_81 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001010011");
        state_var_NS <= COMP_LOOP_C_82;
      WHEN COMP_LOOP_C_82 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001010100");
        state_var_NS <= COMP_LOOP_C_83;
      WHEN COMP_LOOP_C_83 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001010101");
        state_var_NS <= COMP_LOOP_C_84;
      WHEN COMP_LOOP_C_84 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001010110");
        state_var_NS <= COMP_LOOP_C_85;
      WHEN COMP_LOOP_C_85 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001010111");
        state_var_NS <= COMP_LOOP_C_86;
      WHEN COMP_LOOP_C_86 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001011000");
        state_var_NS <= COMP_LOOP_C_87;
      WHEN COMP_LOOP_C_87 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001011001");
        state_var_NS <= COMP_LOOP_C_88;
      WHEN COMP_LOOP_C_88 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001011010");
        state_var_NS <= COMP_LOOP_C_89;
      WHEN COMP_LOOP_C_89 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001011011");
        state_var_NS <= COMP_LOOP_C_90;
      WHEN COMP_LOOP_C_90 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001011100");
        state_var_NS <= COMP_LOOP_C_91;
      WHEN COMP_LOOP_C_91 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001011101");
        state_var_NS <= COMP_LOOP_C_92;
      WHEN COMP_LOOP_C_92 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001011110");
        state_var_NS <= COMP_LOOP_C_93;
      WHEN COMP_LOOP_C_93 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001011111");
        IF ( COMP_LOOP_C_93_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_94;
        END IF;
      WHEN COMP_LOOP_C_94 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001100000");
        state_var_NS <= COMP_LOOP_C_95;
      WHEN COMP_LOOP_C_95 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001100001");
        state_var_NS <= COMP_LOOP_C_96;
      WHEN COMP_LOOP_C_96 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001100010");
        state_var_NS <= COMP_LOOP_C_97;
      WHEN COMP_LOOP_C_97 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001100011");
        state_var_NS <= COMP_LOOP_C_98;
      WHEN COMP_LOOP_C_98 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001100100");
        state_var_NS <= COMP_LOOP_C_99;
      WHEN COMP_LOOP_C_99 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001100101");
        state_var_NS <= COMP_LOOP_C_100;
      WHEN COMP_LOOP_C_100 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001100110");
        state_var_NS <= COMP_LOOP_C_101;
      WHEN COMP_LOOP_C_101 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001100111");
        state_var_NS <= COMP_LOOP_C_102;
      WHEN COMP_LOOP_C_102 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001101000");
        state_var_NS <= COMP_LOOP_C_103;
      WHEN COMP_LOOP_C_103 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001101001");
        state_var_NS <= COMP_LOOP_C_104;
      WHEN COMP_LOOP_C_104 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001101010");
        state_var_NS <= COMP_LOOP_C_105;
      WHEN COMP_LOOP_C_105 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001101011");
        state_var_NS <= COMP_LOOP_C_106;
      WHEN COMP_LOOP_C_106 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001101100");
        state_var_NS <= COMP_LOOP_C_107;
      WHEN COMP_LOOP_C_107 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001101101");
        state_var_NS <= COMP_LOOP_C_108;
      WHEN COMP_LOOP_C_108 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001101110");
        state_var_NS <= COMP_LOOP_C_109;
      WHEN COMP_LOOP_C_109 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001101111");
        state_var_NS <= COMP_LOOP_C_110;
      WHEN COMP_LOOP_C_110 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001110000");
        state_var_NS <= COMP_LOOP_C_111;
      WHEN COMP_LOOP_C_111 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001110001");
        state_var_NS <= COMP_LOOP_C_112;
      WHEN COMP_LOOP_C_112 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001110010");
        state_var_NS <= COMP_LOOP_C_113;
      WHEN COMP_LOOP_C_113 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001110011");
        state_var_NS <= COMP_LOOP_C_114;
      WHEN COMP_LOOP_C_114 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001110100");
        state_var_NS <= COMP_LOOP_C_115;
      WHEN COMP_LOOP_C_115 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001110101");
        state_var_NS <= COMP_LOOP_C_116;
      WHEN COMP_LOOP_C_116 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001110110");
        state_var_NS <= COMP_LOOP_C_117;
      WHEN COMP_LOOP_C_117 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001110111");
        state_var_NS <= COMP_LOOP_C_118;
      WHEN COMP_LOOP_C_118 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001111000");
        state_var_NS <= COMP_LOOP_C_119;
      WHEN COMP_LOOP_C_119 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001111001");
        state_var_NS <= COMP_LOOP_C_120;
      WHEN COMP_LOOP_C_120 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001111010");
        state_var_NS <= COMP_LOOP_C_121;
      WHEN COMP_LOOP_C_121 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001111011");
        state_var_NS <= COMP_LOOP_C_122;
      WHEN COMP_LOOP_C_122 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001111100");
        state_var_NS <= COMP_LOOP_C_123;
      WHEN COMP_LOOP_C_123 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001111101");
        state_var_NS <= COMP_LOOP_C_124;
      WHEN COMP_LOOP_C_124 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001111110");
        IF ( COMP_LOOP_C_124_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_125;
        END IF;
      WHEN COMP_LOOP_C_125 =>
        fsm_output <= STD_LOGIC_VECTOR'( "001111111");
        state_var_NS <= COMP_LOOP_C_126;
      WHEN COMP_LOOP_C_126 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010000000");
        state_var_NS <= COMP_LOOP_C_127;
      WHEN COMP_LOOP_C_127 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010000001");
        state_var_NS <= COMP_LOOP_C_128;
      WHEN COMP_LOOP_C_128 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010000010");
        state_var_NS <= COMP_LOOP_C_129;
      WHEN COMP_LOOP_C_129 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010000011");
        state_var_NS <= COMP_LOOP_C_130;
      WHEN COMP_LOOP_C_130 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010000100");
        state_var_NS <= COMP_LOOP_C_131;
      WHEN COMP_LOOP_C_131 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010000101");
        state_var_NS <= COMP_LOOP_C_132;
      WHEN COMP_LOOP_C_132 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010000110");
        state_var_NS <= COMP_LOOP_C_133;
      WHEN COMP_LOOP_C_133 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010000111");
        state_var_NS <= COMP_LOOP_C_134;
      WHEN COMP_LOOP_C_134 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010001000");
        state_var_NS <= COMP_LOOP_C_135;
      WHEN COMP_LOOP_C_135 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010001001");
        state_var_NS <= COMP_LOOP_C_136;
      WHEN COMP_LOOP_C_136 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010001010");
        state_var_NS <= COMP_LOOP_C_137;
      WHEN COMP_LOOP_C_137 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010001011");
        state_var_NS <= COMP_LOOP_C_138;
      WHEN COMP_LOOP_C_138 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010001100");
        state_var_NS <= COMP_LOOP_C_139;
      WHEN COMP_LOOP_C_139 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010001101");
        state_var_NS <= COMP_LOOP_C_140;
      WHEN COMP_LOOP_C_140 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010001110");
        state_var_NS <= COMP_LOOP_C_141;
      WHEN COMP_LOOP_C_141 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010001111");
        state_var_NS <= COMP_LOOP_C_142;
      WHEN COMP_LOOP_C_142 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010010000");
        state_var_NS <= COMP_LOOP_C_143;
      WHEN COMP_LOOP_C_143 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010010001");
        state_var_NS <= COMP_LOOP_C_144;
      WHEN COMP_LOOP_C_144 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010010010");
        state_var_NS <= COMP_LOOP_C_145;
      WHEN COMP_LOOP_C_145 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010010011");
        state_var_NS <= COMP_LOOP_C_146;
      WHEN COMP_LOOP_C_146 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010010100");
        state_var_NS <= COMP_LOOP_C_147;
      WHEN COMP_LOOP_C_147 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010010101");
        state_var_NS <= COMP_LOOP_C_148;
      WHEN COMP_LOOP_C_148 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010010110");
        state_var_NS <= COMP_LOOP_C_149;
      WHEN COMP_LOOP_C_149 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010010111");
        state_var_NS <= COMP_LOOP_C_150;
      WHEN COMP_LOOP_C_150 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010011000");
        state_var_NS <= COMP_LOOP_C_151;
      WHEN COMP_LOOP_C_151 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010011001");
        state_var_NS <= COMP_LOOP_C_152;
      WHEN COMP_LOOP_C_152 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010011010");
        state_var_NS <= COMP_LOOP_C_153;
      WHEN COMP_LOOP_C_153 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010011011");
        state_var_NS <= COMP_LOOP_C_154;
      WHEN COMP_LOOP_C_154 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010011100");
        state_var_NS <= COMP_LOOP_C_155;
      WHEN COMP_LOOP_C_155 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010011101");
        IF ( COMP_LOOP_C_155_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_156;
        END IF;
      WHEN COMP_LOOP_C_156 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010011110");
        state_var_NS <= COMP_LOOP_C_157;
      WHEN COMP_LOOP_C_157 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010011111");
        state_var_NS <= COMP_LOOP_C_158;
      WHEN COMP_LOOP_C_158 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010100000");
        state_var_NS <= COMP_LOOP_C_159;
      WHEN COMP_LOOP_C_159 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010100001");
        state_var_NS <= COMP_LOOP_C_160;
      WHEN COMP_LOOP_C_160 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010100010");
        state_var_NS <= COMP_LOOP_C_161;
      WHEN COMP_LOOP_C_161 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010100011");
        state_var_NS <= COMP_LOOP_C_162;
      WHEN COMP_LOOP_C_162 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010100100");
        state_var_NS <= COMP_LOOP_C_163;
      WHEN COMP_LOOP_C_163 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010100101");
        state_var_NS <= COMP_LOOP_C_164;
      WHEN COMP_LOOP_C_164 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010100110");
        state_var_NS <= COMP_LOOP_C_165;
      WHEN COMP_LOOP_C_165 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010100111");
        state_var_NS <= COMP_LOOP_C_166;
      WHEN COMP_LOOP_C_166 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010101000");
        state_var_NS <= COMP_LOOP_C_167;
      WHEN COMP_LOOP_C_167 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010101001");
        state_var_NS <= COMP_LOOP_C_168;
      WHEN COMP_LOOP_C_168 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010101010");
        state_var_NS <= COMP_LOOP_C_169;
      WHEN COMP_LOOP_C_169 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010101011");
        state_var_NS <= COMP_LOOP_C_170;
      WHEN COMP_LOOP_C_170 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010101100");
        state_var_NS <= COMP_LOOP_C_171;
      WHEN COMP_LOOP_C_171 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010101101");
        state_var_NS <= COMP_LOOP_C_172;
      WHEN COMP_LOOP_C_172 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010101110");
        state_var_NS <= COMP_LOOP_C_173;
      WHEN COMP_LOOP_C_173 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010101111");
        state_var_NS <= COMP_LOOP_C_174;
      WHEN COMP_LOOP_C_174 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010110000");
        state_var_NS <= COMP_LOOP_C_175;
      WHEN COMP_LOOP_C_175 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010110001");
        state_var_NS <= COMP_LOOP_C_176;
      WHEN COMP_LOOP_C_176 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010110010");
        state_var_NS <= COMP_LOOP_C_177;
      WHEN COMP_LOOP_C_177 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010110011");
        state_var_NS <= COMP_LOOP_C_178;
      WHEN COMP_LOOP_C_178 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010110100");
        state_var_NS <= COMP_LOOP_C_179;
      WHEN COMP_LOOP_C_179 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010110101");
        state_var_NS <= COMP_LOOP_C_180;
      WHEN COMP_LOOP_C_180 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010110110");
        state_var_NS <= COMP_LOOP_C_181;
      WHEN COMP_LOOP_C_181 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010110111");
        state_var_NS <= COMP_LOOP_C_182;
      WHEN COMP_LOOP_C_182 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010111000");
        state_var_NS <= COMP_LOOP_C_183;
      WHEN COMP_LOOP_C_183 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010111001");
        state_var_NS <= COMP_LOOP_C_184;
      WHEN COMP_LOOP_C_184 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010111010");
        state_var_NS <= COMP_LOOP_C_185;
      WHEN COMP_LOOP_C_185 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010111011");
        state_var_NS <= COMP_LOOP_C_186;
      WHEN COMP_LOOP_C_186 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010111100");
        IF ( COMP_LOOP_C_186_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_187;
        END IF;
      WHEN COMP_LOOP_C_187 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010111101");
        state_var_NS <= COMP_LOOP_C_188;
      WHEN COMP_LOOP_C_188 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010111110");
        state_var_NS <= COMP_LOOP_C_189;
      WHEN COMP_LOOP_C_189 =>
        fsm_output <= STD_LOGIC_VECTOR'( "010111111");
        state_var_NS <= COMP_LOOP_C_190;
      WHEN COMP_LOOP_C_190 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011000000");
        state_var_NS <= COMP_LOOP_C_191;
      WHEN COMP_LOOP_C_191 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011000001");
        state_var_NS <= COMP_LOOP_C_192;
      WHEN COMP_LOOP_C_192 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011000010");
        state_var_NS <= COMP_LOOP_C_193;
      WHEN COMP_LOOP_C_193 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011000011");
        state_var_NS <= COMP_LOOP_C_194;
      WHEN COMP_LOOP_C_194 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011000100");
        state_var_NS <= COMP_LOOP_C_195;
      WHEN COMP_LOOP_C_195 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011000101");
        state_var_NS <= COMP_LOOP_C_196;
      WHEN COMP_LOOP_C_196 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011000110");
        state_var_NS <= COMP_LOOP_C_197;
      WHEN COMP_LOOP_C_197 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011000111");
        state_var_NS <= COMP_LOOP_C_198;
      WHEN COMP_LOOP_C_198 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011001000");
        state_var_NS <= COMP_LOOP_C_199;
      WHEN COMP_LOOP_C_199 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011001001");
        state_var_NS <= COMP_LOOP_C_200;
      WHEN COMP_LOOP_C_200 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011001010");
        state_var_NS <= COMP_LOOP_C_201;
      WHEN COMP_LOOP_C_201 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011001011");
        state_var_NS <= COMP_LOOP_C_202;
      WHEN COMP_LOOP_C_202 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011001100");
        state_var_NS <= COMP_LOOP_C_203;
      WHEN COMP_LOOP_C_203 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011001101");
        state_var_NS <= COMP_LOOP_C_204;
      WHEN COMP_LOOP_C_204 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011001110");
        state_var_NS <= COMP_LOOP_C_205;
      WHEN COMP_LOOP_C_205 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011001111");
        state_var_NS <= COMP_LOOP_C_206;
      WHEN COMP_LOOP_C_206 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011010000");
        state_var_NS <= COMP_LOOP_C_207;
      WHEN COMP_LOOP_C_207 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011010001");
        state_var_NS <= COMP_LOOP_C_208;
      WHEN COMP_LOOP_C_208 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011010010");
        state_var_NS <= COMP_LOOP_C_209;
      WHEN COMP_LOOP_C_209 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011010011");
        state_var_NS <= COMP_LOOP_C_210;
      WHEN COMP_LOOP_C_210 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011010100");
        state_var_NS <= COMP_LOOP_C_211;
      WHEN COMP_LOOP_C_211 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011010101");
        state_var_NS <= COMP_LOOP_C_212;
      WHEN COMP_LOOP_C_212 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011010110");
        state_var_NS <= COMP_LOOP_C_213;
      WHEN COMP_LOOP_C_213 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011010111");
        state_var_NS <= COMP_LOOP_C_214;
      WHEN COMP_LOOP_C_214 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011011000");
        state_var_NS <= COMP_LOOP_C_215;
      WHEN COMP_LOOP_C_215 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011011001");
        state_var_NS <= COMP_LOOP_C_216;
      WHEN COMP_LOOP_C_216 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011011010");
        state_var_NS <= COMP_LOOP_C_217;
      WHEN COMP_LOOP_C_217 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011011011");
        IF ( COMP_LOOP_C_217_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_218;
        END IF;
      WHEN COMP_LOOP_C_218 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011011100");
        state_var_NS <= COMP_LOOP_C_219;
      WHEN COMP_LOOP_C_219 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011011101");
        state_var_NS <= COMP_LOOP_C_220;
      WHEN COMP_LOOP_C_220 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011011110");
        state_var_NS <= COMP_LOOP_C_221;
      WHEN COMP_LOOP_C_221 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011011111");
        state_var_NS <= COMP_LOOP_C_222;
      WHEN COMP_LOOP_C_222 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011100000");
        state_var_NS <= COMP_LOOP_C_223;
      WHEN COMP_LOOP_C_223 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011100001");
        state_var_NS <= COMP_LOOP_C_224;
      WHEN COMP_LOOP_C_224 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011100010");
        state_var_NS <= COMP_LOOP_C_225;
      WHEN COMP_LOOP_C_225 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011100011");
        state_var_NS <= COMP_LOOP_C_226;
      WHEN COMP_LOOP_C_226 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011100100");
        state_var_NS <= COMP_LOOP_C_227;
      WHEN COMP_LOOP_C_227 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011100101");
        state_var_NS <= COMP_LOOP_C_228;
      WHEN COMP_LOOP_C_228 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011100110");
        state_var_NS <= COMP_LOOP_C_229;
      WHEN COMP_LOOP_C_229 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011100111");
        state_var_NS <= COMP_LOOP_C_230;
      WHEN COMP_LOOP_C_230 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011101000");
        state_var_NS <= COMP_LOOP_C_231;
      WHEN COMP_LOOP_C_231 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011101001");
        state_var_NS <= COMP_LOOP_C_232;
      WHEN COMP_LOOP_C_232 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011101010");
        state_var_NS <= COMP_LOOP_C_233;
      WHEN COMP_LOOP_C_233 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011101011");
        state_var_NS <= COMP_LOOP_C_234;
      WHEN COMP_LOOP_C_234 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011101100");
        state_var_NS <= COMP_LOOP_C_235;
      WHEN COMP_LOOP_C_235 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011101101");
        state_var_NS <= COMP_LOOP_C_236;
      WHEN COMP_LOOP_C_236 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011101110");
        state_var_NS <= COMP_LOOP_C_237;
      WHEN COMP_LOOP_C_237 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011101111");
        state_var_NS <= COMP_LOOP_C_238;
      WHEN COMP_LOOP_C_238 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011110000");
        state_var_NS <= COMP_LOOP_C_239;
      WHEN COMP_LOOP_C_239 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011110001");
        state_var_NS <= COMP_LOOP_C_240;
      WHEN COMP_LOOP_C_240 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011110010");
        state_var_NS <= COMP_LOOP_C_241;
      WHEN COMP_LOOP_C_241 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011110011");
        state_var_NS <= COMP_LOOP_C_242;
      WHEN COMP_LOOP_C_242 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011110100");
        state_var_NS <= COMP_LOOP_C_243;
      WHEN COMP_LOOP_C_243 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011110101");
        state_var_NS <= COMP_LOOP_C_244;
      WHEN COMP_LOOP_C_244 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011110110");
        state_var_NS <= COMP_LOOP_C_245;
      WHEN COMP_LOOP_C_245 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011110111");
        state_var_NS <= COMP_LOOP_C_246;
      WHEN COMP_LOOP_C_246 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011111000");
        state_var_NS <= COMP_LOOP_C_247;
      WHEN COMP_LOOP_C_247 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011111001");
        state_var_NS <= COMP_LOOP_C_248;
      WHEN COMP_LOOP_C_248 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011111010");
        IF ( COMP_LOOP_C_248_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_249;
        END IF;
      WHEN COMP_LOOP_C_249 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011111011");
        state_var_NS <= COMP_LOOP_C_250;
      WHEN COMP_LOOP_C_250 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011111100");
        state_var_NS <= COMP_LOOP_C_251;
      WHEN COMP_LOOP_C_251 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011111101");
        state_var_NS <= COMP_LOOP_C_252;
      WHEN COMP_LOOP_C_252 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011111110");
        state_var_NS <= COMP_LOOP_C_253;
      WHEN COMP_LOOP_C_253 =>
        fsm_output <= STD_LOGIC_VECTOR'( "011111111");
        state_var_NS <= COMP_LOOP_C_254;
      WHEN COMP_LOOP_C_254 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100000000");
        state_var_NS <= COMP_LOOP_C_255;
      WHEN COMP_LOOP_C_255 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100000001");
        state_var_NS <= COMP_LOOP_C_256;
      WHEN COMP_LOOP_C_256 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100000010");
        state_var_NS <= COMP_LOOP_C_257;
      WHEN COMP_LOOP_C_257 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100000011");
        state_var_NS <= COMP_LOOP_C_258;
      WHEN COMP_LOOP_C_258 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100000100");
        state_var_NS <= COMP_LOOP_C_259;
      WHEN COMP_LOOP_C_259 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100000101");
        state_var_NS <= COMP_LOOP_C_260;
      WHEN COMP_LOOP_C_260 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100000110");
        state_var_NS <= COMP_LOOP_C_261;
      WHEN COMP_LOOP_C_261 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100000111");
        state_var_NS <= COMP_LOOP_C_262;
      WHEN COMP_LOOP_C_262 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100001000");
        state_var_NS <= COMP_LOOP_C_263;
      WHEN COMP_LOOP_C_263 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100001001");
        state_var_NS <= COMP_LOOP_C_264;
      WHEN COMP_LOOP_C_264 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100001010");
        state_var_NS <= COMP_LOOP_C_265;
      WHEN COMP_LOOP_C_265 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100001011");
        state_var_NS <= COMP_LOOP_C_266;
      WHEN COMP_LOOP_C_266 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100001100");
        state_var_NS <= COMP_LOOP_C_267;
      WHEN COMP_LOOP_C_267 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100001101");
        state_var_NS <= COMP_LOOP_C_268;
      WHEN COMP_LOOP_C_268 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100001110");
        state_var_NS <= COMP_LOOP_C_269;
      WHEN COMP_LOOP_C_269 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100001111");
        state_var_NS <= COMP_LOOP_C_270;
      WHEN COMP_LOOP_C_270 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100010000");
        state_var_NS <= COMP_LOOP_C_271;
      WHEN COMP_LOOP_C_271 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100010001");
        state_var_NS <= COMP_LOOP_C_272;
      WHEN COMP_LOOP_C_272 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100010010");
        state_var_NS <= COMP_LOOP_C_273;
      WHEN COMP_LOOP_C_273 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100010011");
        state_var_NS <= COMP_LOOP_C_274;
      WHEN COMP_LOOP_C_274 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100010100");
        state_var_NS <= COMP_LOOP_C_275;
      WHEN COMP_LOOP_C_275 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100010101");
        state_var_NS <= COMP_LOOP_C_276;
      WHEN COMP_LOOP_C_276 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100010110");
        state_var_NS <= COMP_LOOP_C_277;
      WHEN COMP_LOOP_C_277 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100010111");
        state_var_NS <= COMP_LOOP_C_278;
      WHEN COMP_LOOP_C_278 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100011000");
        state_var_NS <= COMP_LOOP_C_279;
      WHEN COMP_LOOP_C_279 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100011001");
        IF ( COMP_LOOP_C_279_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_280;
        END IF;
      WHEN COMP_LOOP_C_280 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100011010");
        state_var_NS <= COMP_LOOP_C_281;
      WHEN COMP_LOOP_C_281 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100011011");
        state_var_NS <= COMP_LOOP_C_282;
      WHEN COMP_LOOP_C_282 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100011100");
        state_var_NS <= COMP_LOOP_C_283;
      WHEN COMP_LOOP_C_283 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100011101");
        state_var_NS <= COMP_LOOP_C_284;
      WHEN COMP_LOOP_C_284 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100011110");
        state_var_NS <= COMP_LOOP_C_285;
      WHEN COMP_LOOP_C_285 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100011111");
        state_var_NS <= COMP_LOOP_C_286;
      WHEN COMP_LOOP_C_286 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100100000");
        state_var_NS <= COMP_LOOP_C_287;
      WHEN COMP_LOOP_C_287 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100100001");
        state_var_NS <= COMP_LOOP_C_288;
      WHEN COMP_LOOP_C_288 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100100010");
        state_var_NS <= COMP_LOOP_C_289;
      WHEN COMP_LOOP_C_289 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100100011");
        state_var_NS <= COMP_LOOP_C_290;
      WHEN COMP_LOOP_C_290 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100100100");
        state_var_NS <= COMP_LOOP_C_291;
      WHEN COMP_LOOP_C_291 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100100101");
        state_var_NS <= COMP_LOOP_C_292;
      WHEN COMP_LOOP_C_292 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100100110");
        state_var_NS <= COMP_LOOP_C_293;
      WHEN COMP_LOOP_C_293 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100100111");
        state_var_NS <= COMP_LOOP_C_294;
      WHEN COMP_LOOP_C_294 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100101000");
        state_var_NS <= COMP_LOOP_C_295;
      WHEN COMP_LOOP_C_295 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100101001");
        state_var_NS <= COMP_LOOP_C_296;
      WHEN COMP_LOOP_C_296 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100101010");
        state_var_NS <= COMP_LOOP_C_297;
      WHEN COMP_LOOP_C_297 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100101011");
        state_var_NS <= COMP_LOOP_C_298;
      WHEN COMP_LOOP_C_298 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100101100");
        state_var_NS <= COMP_LOOP_C_299;
      WHEN COMP_LOOP_C_299 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100101101");
        state_var_NS <= COMP_LOOP_C_300;
      WHEN COMP_LOOP_C_300 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100101110");
        state_var_NS <= COMP_LOOP_C_301;
      WHEN COMP_LOOP_C_301 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100101111");
        state_var_NS <= COMP_LOOP_C_302;
      WHEN COMP_LOOP_C_302 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100110000");
        state_var_NS <= COMP_LOOP_C_303;
      WHEN COMP_LOOP_C_303 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100110001");
        state_var_NS <= COMP_LOOP_C_304;
      WHEN COMP_LOOP_C_304 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100110010");
        state_var_NS <= COMP_LOOP_C_305;
      WHEN COMP_LOOP_C_305 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100110011");
        state_var_NS <= COMP_LOOP_C_306;
      WHEN COMP_LOOP_C_306 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100110100");
        state_var_NS <= COMP_LOOP_C_307;
      WHEN COMP_LOOP_C_307 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100110101");
        state_var_NS <= COMP_LOOP_C_308;
      WHEN COMP_LOOP_C_308 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100110110");
        state_var_NS <= COMP_LOOP_C_309;
      WHEN COMP_LOOP_C_309 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100110111");
        state_var_NS <= COMP_LOOP_C_310;
      WHEN COMP_LOOP_C_310 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100111000");
        IF ( COMP_LOOP_C_310_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_311;
        END IF;
      WHEN COMP_LOOP_C_311 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100111001");
        state_var_NS <= COMP_LOOP_C_312;
      WHEN COMP_LOOP_C_312 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100111010");
        state_var_NS <= COMP_LOOP_C_313;
      WHEN COMP_LOOP_C_313 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100111011");
        state_var_NS <= COMP_LOOP_C_314;
      WHEN COMP_LOOP_C_314 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100111100");
        state_var_NS <= COMP_LOOP_C_315;
      WHEN COMP_LOOP_C_315 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100111101");
        state_var_NS <= COMP_LOOP_C_316;
      WHEN COMP_LOOP_C_316 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100111110");
        state_var_NS <= COMP_LOOP_C_317;
      WHEN COMP_LOOP_C_317 =>
        fsm_output <= STD_LOGIC_VECTOR'( "100111111");
        state_var_NS <= COMP_LOOP_C_318;
      WHEN COMP_LOOP_C_318 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101000000");
        state_var_NS <= COMP_LOOP_C_319;
      WHEN COMP_LOOP_C_319 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101000001");
        state_var_NS <= COMP_LOOP_C_320;
      WHEN COMP_LOOP_C_320 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101000010");
        state_var_NS <= COMP_LOOP_C_321;
      WHEN COMP_LOOP_C_321 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101000011");
        state_var_NS <= COMP_LOOP_C_322;
      WHEN COMP_LOOP_C_322 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101000100");
        state_var_NS <= COMP_LOOP_C_323;
      WHEN COMP_LOOP_C_323 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101000101");
        state_var_NS <= COMP_LOOP_C_324;
      WHEN COMP_LOOP_C_324 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101000110");
        state_var_NS <= COMP_LOOP_C_325;
      WHEN COMP_LOOP_C_325 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101000111");
        state_var_NS <= COMP_LOOP_C_326;
      WHEN COMP_LOOP_C_326 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101001000");
        state_var_NS <= COMP_LOOP_C_327;
      WHEN COMP_LOOP_C_327 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101001001");
        state_var_NS <= COMP_LOOP_C_328;
      WHEN COMP_LOOP_C_328 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101001010");
        state_var_NS <= COMP_LOOP_C_329;
      WHEN COMP_LOOP_C_329 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101001011");
        state_var_NS <= COMP_LOOP_C_330;
      WHEN COMP_LOOP_C_330 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101001100");
        state_var_NS <= COMP_LOOP_C_331;
      WHEN COMP_LOOP_C_331 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101001101");
        state_var_NS <= COMP_LOOP_C_332;
      WHEN COMP_LOOP_C_332 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101001110");
        state_var_NS <= COMP_LOOP_C_333;
      WHEN COMP_LOOP_C_333 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101001111");
        state_var_NS <= COMP_LOOP_C_334;
      WHEN COMP_LOOP_C_334 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101010000");
        state_var_NS <= COMP_LOOP_C_335;
      WHEN COMP_LOOP_C_335 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101010001");
        state_var_NS <= COMP_LOOP_C_336;
      WHEN COMP_LOOP_C_336 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101010010");
        state_var_NS <= COMP_LOOP_C_337;
      WHEN COMP_LOOP_C_337 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101010011");
        state_var_NS <= COMP_LOOP_C_338;
      WHEN COMP_LOOP_C_338 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101010100");
        state_var_NS <= COMP_LOOP_C_339;
      WHEN COMP_LOOP_C_339 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101010101");
        state_var_NS <= COMP_LOOP_C_340;
      WHEN COMP_LOOP_C_340 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101010110");
        state_var_NS <= COMP_LOOP_C_341;
      WHEN COMP_LOOP_C_341 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101010111");
        IF ( COMP_LOOP_C_341_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_342;
        END IF;
      WHEN COMP_LOOP_C_342 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101011000");
        state_var_NS <= COMP_LOOP_C_343;
      WHEN COMP_LOOP_C_343 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101011001");
        state_var_NS <= COMP_LOOP_C_344;
      WHEN COMP_LOOP_C_344 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101011010");
        state_var_NS <= COMP_LOOP_C_345;
      WHEN COMP_LOOP_C_345 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101011011");
        state_var_NS <= COMP_LOOP_C_346;
      WHEN COMP_LOOP_C_346 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101011100");
        state_var_NS <= COMP_LOOP_C_347;
      WHEN COMP_LOOP_C_347 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101011101");
        state_var_NS <= COMP_LOOP_C_348;
      WHEN COMP_LOOP_C_348 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101011110");
        state_var_NS <= COMP_LOOP_C_349;
      WHEN COMP_LOOP_C_349 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101011111");
        state_var_NS <= COMP_LOOP_C_350;
      WHEN COMP_LOOP_C_350 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101100000");
        state_var_NS <= COMP_LOOP_C_351;
      WHEN COMP_LOOP_C_351 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101100001");
        state_var_NS <= COMP_LOOP_C_352;
      WHEN COMP_LOOP_C_352 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101100010");
        state_var_NS <= COMP_LOOP_C_353;
      WHEN COMP_LOOP_C_353 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101100011");
        state_var_NS <= COMP_LOOP_C_354;
      WHEN COMP_LOOP_C_354 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101100100");
        state_var_NS <= COMP_LOOP_C_355;
      WHEN COMP_LOOP_C_355 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101100101");
        state_var_NS <= COMP_LOOP_C_356;
      WHEN COMP_LOOP_C_356 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101100110");
        state_var_NS <= COMP_LOOP_C_357;
      WHEN COMP_LOOP_C_357 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101100111");
        state_var_NS <= COMP_LOOP_C_358;
      WHEN COMP_LOOP_C_358 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101101000");
        state_var_NS <= COMP_LOOP_C_359;
      WHEN COMP_LOOP_C_359 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101101001");
        state_var_NS <= COMP_LOOP_C_360;
      WHEN COMP_LOOP_C_360 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101101010");
        state_var_NS <= COMP_LOOP_C_361;
      WHEN COMP_LOOP_C_361 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101101011");
        state_var_NS <= COMP_LOOP_C_362;
      WHEN COMP_LOOP_C_362 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101101100");
        state_var_NS <= COMP_LOOP_C_363;
      WHEN COMP_LOOP_C_363 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101101101");
        state_var_NS <= COMP_LOOP_C_364;
      WHEN COMP_LOOP_C_364 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101101110");
        state_var_NS <= COMP_LOOP_C_365;
      WHEN COMP_LOOP_C_365 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101101111");
        state_var_NS <= COMP_LOOP_C_366;
      WHEN COMP_LOOP_C_366 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101110000");
        state_var_NS <= COMP_LOOP_C_367;
      WHEN COMP_LOOP_C_367 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101110001");
        state_var_NS <= COMP_LOOP_C_368;
      WHEN COMP_LOOP_C_368 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101110010");
        state_var_NS <= COMP_LOOP_C_369;
      WHEN COMP_LOOP_C_369 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101110011");
        state_var_NS <= COMP_LOOP_C_370;
      WHEN COMP_LOOP_C_370 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101110100");
        state_var_NS <= COMP_LOOP_C_371;
      WHEN COMP_LOOP_C_371 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101110101");
        state_var_NS <= COMP_LOOP_C_372;
      WHEN COMP_LOOP_C_372 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101110110");
        IF ( COMP_LOOP_C_372_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_373;
        END IF;
      WHEN COMP_LOOP_C_373 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101110111");
        state_var_NS <= COMP_LOOP_C_374;
      WHEN COMP_LOOP_C_374 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101111000");
        state_var_NS <= COMP_LOOP_C_375;
      WHEN COMP_LOOP_C_375 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101111001");
        state_var_NS <= COMP_LOOP_C_376;
      WHEN COMP_LOOP_C_376 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101111010");
        state_var_NS <= COMP_LOOP_C_377;
      WHEN COMP_LOOP_C_377 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101111011");
        state_var_NS <= COMP_LOOP_C_378;
      WHEN COMP_LOOP_C_378 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101111100");
        state_var_NS <= COMP_LOOP_C_379;
      WHEN COMP_LOOP_C_379 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101111101");
        state_var_NS <= COMP_LOOP_C_380;
      WHEN COMP_LOOP_C_380 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101111110");
        state_var_NS <= COMP_LOOP_C_381;
      WHEN COMP_LOOP_C_381 =>
        fsm_output <= STD_LOGIC_VECTOR'( "101111111");
        state_var_NS <= COMP_LOOP_C_382;
      WHEN COMP_LOOP_C_382 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110000000");
        state_var_NS <= COMP_LOOP_C_383;
      WHEN COMP_LOOP_C_383 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110000001");
        state_var_NS <= COMP_LOOP_C_384;
      WHEN COMP_LOOP_C_384 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110000010");
        state_var_NS <= COMP_LOOP_C_385;
      WHEN COMP_LOOP_C_385 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110000011");
        state_var_NS <= COMP_LOOP_C_386;
      WHEN COMP_LOOP_C_386 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110000100");
        state_var_NS <= COMP_LOOP_C_387;
      WHEN COMP_LOOP_C_387 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110000101");
        state_var_NS <= COMP_LOOP_C_388;
      WHEN COMP_LOOP_C_388 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110000110");
        state_var_NS <= COMP_LOOP_C_389;
      WHEN COMP_LOOP_C_389 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110000111");
        state_var_NS <= COMP_LOOP_C_390;
      WHEN COMP_LOOP_C_390 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110001000");
        state_var_NS <= COMP_LOOP_C_391;
      WHEN COMP_LOOP_C_391 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110001001");
        state_var_NS <= COMP_LOOP_C_392;
      WHEN COMP_LOOP_C_392 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110001010");
        state_var_NS <= COMP_LOOP_C_393;
      WHEN COMP_LOOP_C_393 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110001011");
        state_var_NS <= COMP_LOOP_C_394;
      WHEN COMP_LOOP_C_394 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110001100");
        state_var_NS <= COMP_LOOP_C_395;
      WHEN COMP_LOOP_C_395 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110001101");
        state_var_NS <= COMP_LOOP_C_396;
      WHEN COMP_LOOP_C_396 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110001110");
        state_var_NS <= COMP_LOOP_C_397;
      WHEN COMP_LOOP_C_397 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110001111");
        state_var_NS <= COMP_LOOP_C_398;
      WHEN COMP_LOOP_C_398 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110010000");
        state_var_NS <= COMP_LOOP_C_399;
      WHEN COMP_LOOP_C_399 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110010001");
        state_var_NS <= COMP_LOOP_C_400;
      WHEN COMP_LOOP_C_400 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110010010");
        state_var_NS <= COMP_LOOP_C_401;
      WHEN COMP_LOOP_C_401 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110010011");
        state_var_NS <= COMP_LOOP_C_402;
      WHEN COMP_LOOP_C_402 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110010100");
        state_var_NS <= COMP_LOOP_C_403;
      WHEN COMP_LOOP_C_403 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110010101");
        IF ( COMP_LOOP_C_403_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_404;
        END IF;
      WHEN COMP_LOOP_C_404 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110010110");
        state_var_NS <= COMP_LOOP_C_405;
      WHEN COMP_LOOP_C_405 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110010111");
        state_var_NS <= COMP_LOOP_C_406;
      WHEN COMP_LOOP_C_406 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110011000");
        state_var_NS <= COMP_LOOP_C_407;
      WHEN COMP_LOOP_C_407 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110011001");
        state_var_NS <= COMP_LOOP_C_408;
      WHEN COMP_LOOP_C_408 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110011010");
        state_var_NS <= COMP_LOOP_C_409;
      WHEN COMP_LOOP_C_409 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110011011");
        state_var_NS <= COMP_LOOP_C_410;
      WHEN COMP_LOOP_C_410 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110011100");
        state_var_NS <= COMP_LOOP_C_411;
      WHEN COMP_LOOP_C_411 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110011101");
        state_var_NS <= COMP_LOOP_C_412;
      WHEN COMP_LOOP_C_412 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110011110");
        state_var_NS <= COMP_LOOP_C_413;
      WHEN COMP_LOOP_C_413 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110011111");
        state_var_NS <= COMP_LOOP_C_414;
      WHEN COMP_LOOP_C_414 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110100000");
        state_var_NS <= COMP_LOOP_C_415;
      WHEN COMP_LOOP_C_415 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110100001");
        state_var_NS <= COMP_LOOP_C_416;
      WHEN COMP_LOOP_C_416 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110100010");
        state_var_NS <= COMP_LOOP_C_417;
      WHEN COMP_LOOP_C_417 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110100011");
        state_var_NS <= COMP_LOOP_C_418;
      WHEN COMP_LOOP_C_418 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110100100");
        state_var_NS <= COMP_LOOP_C_419;
      WHEN COMP_LOOP_C_419 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110100101");
        state_var_NS <= COMP_LOOP_C_420;
      WHEN COMP_LOOP_C_420 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110100110");
        state_var_NS <= COMP_LOOP_C_421;
      WHEN COMP_LOOP_C_421 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110100111");
        state_var_NS <= COMP_LOOP_C_422;
      WHEN COMP_LOOP_C_422 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110101000");
        state_var_NS <= COMP_LOOP_C_423;
      WHEN COMP_LOOP_C_423 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110101001");
        state_var_NS <= COMP_LOOP_C_424;
      WHEN COMP_LOOP_C_424 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110101010");
        state_var_NS <= COMP_LOOP_C_425;
      WHEN COMP_LOOP_C_425 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110101011");
        state_var_NS <= COMP_LOOP_C_426;
      WHEN COMP_LOOP_C_426 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110101100");
        state_var_NS <= COMP_LOOP_C_427;
      WHEN COMP_LOOP_C_427 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110101101");
        state_var_NS <= COMP_LOOP_C_428;
      WHEN COMP_LOOP_C_428 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110101110");
        state_var_NS <= COMP_LOOP_C_429;
      WHEN COMP_LOOP_C_429 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110101111");
        state_var_NS <= COMP_LOOP_C_430;
      WHEN COMP_LOOP_C_430 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110110000");
        state_var_NS <= COMP_LOOP_C_431;
      WHEN COMP_LOOP_C_431 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110110001");
        state_var_NS <= COMP_LOOP_C_432;
      WHEN COMP_LOOP_C_432 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110110010");
        state_var_NS <= COMP_LOOP_C_433;
      WHEN COMP_LOOP_C_433 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110110011");
        state_var_NS <= COMP_LOOP_C_434;
      WHEN COMP_LOOP_C_434 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110110100");
        IF ( COMP_LOOP_C_434_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_435;
        END IF;
      WHEN COMP_LOOP_C_435 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110110101");
        state_var_NS <= COMP_LOOP_C_436;
      WHEN COMP_LOOP_C_436 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110110110");
        state_var_NS <= COMP_LOOP_C_437;
      WHEN COMP_LOOP_C_437 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110110111");
        state_var_NS <= COMP_LOOP_C_438;
      WHEN COMP_LOOP_C_438 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110111000");
        state_var_NS <= COMP_LOOP_C_439;
      WHEN COMP_LOOP_C_439 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110111001");
        state_var_NS <= COMP_LOOP_C_440;
      WHEN COMP_LOOP_C_440 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110111010");
        state_var_NS <= COMP_LOOP_C_441;
      WHEN COMP_LOOP_C_441 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110111011");
        state_var_NS <= COMP_LOOP_C_442;
      WHEN COMP_LOOP_C_442 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110111100");
        state_var_NS <= COMP_LOOP_C_443;
      WHEN COMP_LOOP_C_443 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110111101");
        state_var_NS <= COMP_LOOP_C_444;
      WHEN COMP_LOOP_C_444 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110111110");
        state_var_NS <= COMP_LOOP_C_445;
      WHEN COMP_LOOP_C_445 =>
        fsm_output <= STD_LOGIC_VECTOR'( "110111111");
        state_var_NS <= COMP_LOOP_C_446;
      WHEN COMP_LOOP_C_446 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111000000");
        state_var_NS <= COMP_LOOP_C_447;
      WHEN COMP_LOOP_C_447 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111000001");
        state_var_NS <= COMP_LOOP_C_448;
      WHEN COMP_LOOP_C_448 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111000010");
        state_var_NS <= COMP_LOOP_C_449;
      WHEN COMP_LOOP_C_449 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111000011");
        state_var_NS <= COMP_LOOP_C_450;
      WHEN COMP_LOOP_C_450 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111000100");
        state_var_NS <= COMP_LOOP_C_451;
      WHEN COMP_LOOP_C_451 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111000101");
        state_var_NS <= COMP_LOOP_C_452;
      WHEN COMP_LOOP_C_452 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111000110");
        state_var_NS <= COMP_LOOP_C_453;
      WHEN COMP_LOOP_C_453 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111000111");
        state_var_NS <= COMP_LOOP_C_454;
      WHEN COMP_LOOP_C_454 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111001000");
        state_var_NS <= COMP_LOOP_C_455;
      WHEN COMP_LOOP_C_455 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111001001");
        state_var_NS <= COMP_LOOP_C_456;
      WHEN COMP_LOOP_C_456 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111001010");
        state_var_NS <= COMP_LOOP_C_457;
      WHEN COMP_LOOP_C_457 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111001011");
        state_var_NS <= COMP_LOOP_C_458;
      WHEN COMP_LOOP_C_458 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111001100");
        state_var_NS <= COMP_LOOP_C_459;
      WHEN COMP_LOOP_C_459 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111001101");
        state_var_NS <= COMP_LOOP_C_460;
      WHEN COMP_LOOP_C_460 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111001110");
        state_var_NS <= COMP_LOOP_C_461;
      WHEN COMP_LOOP_C_461 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111001111");
        state_var_NS <= COMP_LOOP_C_462;
      WHEN COMP_LOOP_C_462 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111010000");
        state_var_NS <= COMP_LOOP_C_463;
      WHEN COMP_LOOP_C_463 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111010001");
        state_var_NS <= COMP_LOOP_C_464;
      WHEN COMP_LOOP_C_464 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111010010");
        state_var_NS <= COMP_LOOP_C_465;
      WHEN COMP_LOOP_C_465 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111010011");
        IF ( COMP_LOOP_C_465_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_466;
        END IF;
      WHEN COMP_LOOP_C_466 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111010100");
        state_var_NS <= COMP_LOOP_C_467;
      WHEN COMP_LOOP_C_467 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111010101");
        state_var_NS <= COMP_LOOP_C_468;
      WHEN COMP_LOOP_C_468 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111010110");
        state_var_NS <= COMP_LOOP_C_469;
      WHEN COMP_LOOP_C_469 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111010111");
        state_var_NS <= COMP_LOOP_C_470;
      WHEN COMP_LOOP_C_470 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111011000");
        state_var_NS <= COMP_LOOP_C_471;
      WHEN COMP_LOOP_C_471 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111011001");
        state_var_NS <= COMP_LOOP_C_472;
      WHEN COMP_LOOP_C_472 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111011010");
        state_var_NS <= COMP_LOOP_C_473;
      WHEN COMP_LOOP_C_473 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111011011");
        state_var_NS <= COMP_LOOP_C_474;
      WHEN COMP_LOOP_C_474 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111011100");
        state_var_NS <= COMP_LOOP_C_475;
      WHEN COMP_LOOP_C_475 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111011101");
        state_var_NS <= COMP_LOOP_C_476;
      WHEN COMP_LOOP_C_476 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111011110");
        state_var_NS <= COMP_LOOP_C_477;
      WHEN COMP_LOOP_C_477 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111011111");
        state_var_NS <= COMP_LOOP_C_478;
      WHEN COMP_LOOP_C_478 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111100000");
        state_var_NS <= COMP_LOOP_C_479;
      WHEN COMP_LOOP_C_479 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111100001");
        state_var_NS <= COMP_LOOP_C_480;
      WHEN COMP_LOOP_C_480 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111100010");
        state_var_NS <= COMP_LOOP_C_481;
      WHEN COMP_LOOP_C_481 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111100011");
        state_var_NS <= COMP_LOOP_C_482;
      WHEN COMP_LOOP_C_482 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111100100");
        state_var_NS <= COMP_LOOP_C_483;
      WHEN COMP_LOOP_C_483 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111100101");
        state_var_NS <= COMP_LOOP_C_484;
      WHEN COMP_LOOP_C_484 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111100110");
        state_var_NS <= COMP_LOOP_C_485;
      WHEN COMP_LOOP_C_485 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111100111");
        state_var_NS <= COMP_LOOP_C_486;
      WHEN COMP_LOOP_C_486 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111101000");
        state_var_NS <= COMP_LOOP_C_487;
      WHEN COMP_LOOP_C_487 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111101001");
        state_var_NS <= COMP_LOOP_C_488;
      WHEN COMP_LOOP_C_488 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111101010");
        state_var_NS <= COMP_LOOP_C_489;
      WHEN COMP_LOOP_C_489 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111101011");
        state_var_NS <= COMP_LOOP_C_490;
      WHEN COMP_LOOP_C_490 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111101100");
        state_var_NS <= COMP_LOOP_C_491;
      WHEN COMP_LOOP_C_491 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111101101");
        state_var_NS <= COMP_LOOP_C_492;
      WHEN COMP_LOOP_C_492 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111101110");
        state_var_NS <= COMP_LOOP_C_493;
      WHEN COMP_LOOP_C_493 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111101111");
        state_var_NS <= COMP_LOOP_C_494;
      WHEN COMP_LOOP_C_494 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111110000");
        state_var_NS <= COMP_LOOP_C_495;
      WHEN COMP_LOOP_C_495 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111110001");
        state_var_NS <= COMP_LOOP_C_496;
      WHEN COMP_LOOP_C_496 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111110010");
        IF ( COMP_LOOP_C_496_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN VEC_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111110011");
        IF ( VEC_LOOP_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN STAGE_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111110100");
        IF ( STAGE_LOOP_C_1_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSE
          state_var_NS <= STAGE_LOOP_C_0;
        END IF;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "111110101");
        state_var_NS <= main_C_0;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "000000000");
        state_var_NS <= STAGE_LOOP_C_0;
    END CASE;
  END PROCESS inPlaceNTT_DIF_core_core_fsm_1;

  inPlaceNTT_DIF_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        state_var <= state_var_NS;
      END IF;
    END IF;
  END PROCESS inPlaceNTT_DIF_core_core_fsm_1_REG;

END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_core_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_core_wait_dp IS
  PORT(
    ensig_cgo_iro : IN STD_LOGIC;
    ensig_cgo : IN STD_LOGIC;
    COMP_LOOP_1_modulo_cmp_ccs_ccore_en : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_core_wait_dp;

ARCHITECTURE v7 OF inPlaceNTT_DIF_core_wait_dp IS
  -- Default Constants

BEGIN
  COMP_LOOP_1_modulo_cmp_ccs_ccore_en <= ensig_cgo OR ensig_cgo_iro;
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    vec_rsc_0_0_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_1_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_2_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_3_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_4_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_5_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_6_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_7_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_8_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_9_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_10_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_11_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_12_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_13_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_14_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_15_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_0_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_0_i_radr_d : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_1_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_2_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_3_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_4_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_5_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_6_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_7_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_8_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_8_i_radr_d : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_9_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_10_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_11_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_12_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_13_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_14_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_15_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_0_i_d_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_radr_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_0_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_0_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_1_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_2_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_3_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_4_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_5_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_6_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_7_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_8_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_9_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_10_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_11_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_12_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_13_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_14_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_15_i_we_d_pff : OUT STD_LOGIC;
    twiddle_rsc_0_1_i_radr_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_2_i_radr_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_4_i_radr_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0)
  );
END inPlaceNTT_DIF_core;

ARCHITECTURE v7 OF inPlaceNTT_DIF_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL p_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_cmp_return_rsc_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_cmp_ccs_ccore_en : STD_LOGIC;
  SIGNAL fsm_output : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL or_dcpl_5 : STD_LOGIC;
  SIGNAL and_dcpl_5 : STD_LOGIC;
  SIGNAL nor_tmp_10 : STD_LOGIC;
  SIGNAL or_tmp_29 : STD_LOGIC;
  SIGNAL nor_tmp_47 : STD_LOGIC;
  SIGNAL nor_tmp_115 : STD_LOGIC;
  SIGNAL mux_tmp_439 : STD_LOGIC;
  SIGNAL mux_tmp_538 : STD_LOGIC;
  SIGNAL mux_tmp_929 : STD_LOGIC;
  SIGNAL nand_tmp_13 : STD_LOGIC;
  SIGNAL and_dcpl_45 : STD_LOGIC;
  SIGNAL and_dcpl_46 : STD_LOGIC;
  SIGNAL and_dcpl_47 : STD_LOGIC;
  SIGNAL and_dcpl_48 : STD_LOGIC;
  SIGNAL and_dcpl_51 : STD_LOGIC;
  SIGNAL and_dcpl_53 : STD_LOGIC;
  SIGNAL and_dcpl_54 : STD_LOGIC;
  SIGNAL and_dcpl_55 : STD_LOGIC;
  SIGNAL and_dcpl_57 : STD_LOGIC;
  SIGNAL and_dcpl_58 : STD_LOGIC;
  SIGNAL nor_tmp_339 : STD_LOGIC;
  SIGNAL mux_tmp_1062 : STD_LOGIC;
  SIGNAL mux_tmp_1065 : STD_LOGIC;
  SIGNAL mux_tmp_1067 : STD_LOGIC;
  SIGNAL and_dcpl_60 : STD_LOGIC;
  SIGNAL and_dcpl_61 : STD_LOGIC;
  SIGNAL and_dcpl_62 : STD_LOGIC;
  SIGNAL and_dcpl_63 : STD_LOGIC;
  SIGNAL and_dcpl_64 : STD_LOGIC;
  SIGNAL and_dcpl_65 : STD_LOGIC;
  SIGNAL and_dcpl_66 : STD_LOGIC;
  SIGNAL and_dcpl_67 : STD_LOGIC;
  SIGNAL and_dcpl_69 : STD_LOGIC;
  SIGNAL and_dcpl_70 : STD_LOGIC;
  SIGNAL and_dcpl_71 : STD_LOGIC;
  SIGNAL and_dcpl_72 : STD_LOGIC;
  SIGNAL and_dcpl_74 : STD_LOGIC;
  SIGNAL and_dcpl_75 : STD_LOGIC;
  SIGNAL and_dcpl_77 : STD_LOGIC;
  SIGNAL and_dcpl_79 : STD_LOGIC;
  SIGNAL and_dcpl_81 : STD_LOGIC;
  SIGNAL and_dcpl_82 : STD_LOGIC;
  SIGNAL and_dcpl_83 : STD_LOGIC;
  SIGNAL and_dcpl_85 : STD_LOGIC;
  SIGNAL and_dcpl_86 : STD_LOGIC;
  SIGNAL and_dcpl_87 : STD_LOGIC;
  SIGNAL and_dcpl_88 : STD_LOGIC;
  SIGNAL and_dcpl_89 : STD_LOGIC;
  SIGNAL and_dcpl_91 : STD_LOGIC;
  SIGNAL and_dcpl_92 : STD_LOGIC;
  SIGNAL and_dcpl_93 : STD_LOGIC;
  SIGNAL and_dcpl_95 : STD_LOGIC;
  SIGNAL and_dcpl_96 : STD_LOGIC;
  SIGNAL and_dcpl_97 : STD_LOGIC;
  SIGNAL and_dcpl_99 : STD_LOGIC;
  SIGNAL and_dcpl_100 : STD_LOGIC;
  SIGNAL and_dcpl_102 : STD_LOGIC;
  SIGNAL and_dcpl_103 : STD_LOGIC;
  SIGNAL and_dcpl_104 : STD_LOGIC;
  SIGNAL and_dcpl_105 : STD_LOGIC;
  SIGNAL and_dcpl_107 : STD_LOGIC;
  SIGNAL and_dcpl_108 : STD_LOGIC;
  SIGNAL and_dcpl_110 : STD_LOGIC;
  SIGNAL and_dcpl_111 : STD_LOGIC;
  SIGNAL and_dcpl_112 : STD_LOGIC;
  SIGNAL and_dcpl_113 : STD_LOGIC;
  SIGNAL and_dcpl_115 : STD_LOGIC;
  SIGNAL and_dcpl_116 : STD_LOGIC;
  SIGNAL and_dcpl_118 : STD_LOGIC;
  SIGNAL and_dcpl_119 : STD_LOGIC;
  SIGNAL and_dcpl_120 : STD_LOGIC;
  SIGNAL and_dcpl_121 : STD_LOGIC;
  SIGNAL and_dcpl_123 : STD_LOGIC;
  SIGNAL and_dcpl_124 : STD_LOGIC;
  SIGNAL and_dcpl_125 : STD_LOGIC;
  SIGNAL and_dcpl_127 : STD_LOGIC;
  SIGNAL and_dcpl_128 : STD_LOGIC;
  SIGNAL and_dcpl_130 : STD_LOGIC;
  SIGNAL and_dcpl_131 : STD_LOGIC;
  SIGNAL and_dcpl_136 : STD_LOGIC;
  SIGNAL and_dcpl_141 : STD_LOGIC;
  SIGNAL and_dcpl_146 : STD_LOGIC;
  SIGNAL and_dcpl_151 : STD_LOGIC;
  SIGNAL and_dcpl_156 : STD_LOGIC;
  SIGNAL and_dcpl_161 : STD_LOGIC;
  SIGNAL and_dcpl_166 : STD_LOGIC;
  SIGNAL not_tmp_395 : STD_LOGIC;
  SIGNAL not_tmp_399 : STD_LOGIC;
  SIGNAL and_dcpl_171 : STD_LOGIC;
  SIGNAL and_dcpl_175 : STD_LOGIC;
  SIGNAL and_dcpl_180 : STD_LOGIC;
  SIGNAL and_dcpl_181 : STD_LOGIC;
  SIGNAL and_dcpl_182 : STD_LOGIC;
  SIGNAL and_dcpl_183 : STD_LOGIC;
  SIGNAL and_dcpl_184 : STD_LOGIC;
  SIGNAL and_dcpl_186 : STD_LOGIC;
  SIGNAL or_tmp_2077 : STD_LOGIC;
  SIGNAL and_dcpl_188 : STD_LOGIC;
  SIGNAL and_dcpl_189 : STD_LOGIC;
  SIGNAL and_dcpl_190 : STD_LOGIC;
  SIGNAL and_dcpl_191 : STD_LOGIC;
  SIGNAL and_dcpl_192 : STD_LOGIC;
  SIGNAL and_dcpl_193 : STD_LOGIC;
  SIGNAL and_dcpl_195 : STD_LOGIC;
  SIGNAL and_dcpl_196 : STD_LOGIC;
  SIGNAL and_dcpl_197 : STD_LOGIC;
  SIGNAL and_dcpl_198 : STD_LOGIC;
  SIGNAL and_dcpl_202 : STD_LOGIC;
  SIGNAL and_dcpl_207 : STD_LOGIC;
  SIGNAL mux_tmp_2224 : STD_LOGIC;
  SIGNAL mux_tmp_2225 : STD_LOGIC;
  SIGNAL mux_tmp_2229 : STD_LOGIC;
  SIGNAL or_tmp_2258 : STD_LOGIC;
  SIGNAL mux_tmp_2237 : STD_LOGIC;
  SIGNAL not_tmp_676 : STD_LOGIC;
  SIGNAL nor_tmp_480 : STD_LOGIC;
  SIGNAL mux_tmp_2238 : STD_LOGIC;
  SIGNAL or_tmp_2266 : STD_LOGIC;
  SIGNAL mux_tmp_2245 : STD_LOGIC;
  SIGNAL mux_tmp_2246 : STD_LOGIC;
  SIGNAL mux_tmp_2249 : STD_LOGIC;
  SIGNAL and_dcpl_220 : STD_LOGIC;
  SIGNAL and_dcpl_222 : STD_LOGIC;
  SIGNAL and_dcpl_223 : STD_LOGIC;
  SIGNAL and_dcpl_225 : STD_LOGIC;
  SIGNAL and_dcpl_226 : STD_LOGIC;
  SIGNAL and_dcpl_227 : STD_LOGIC;
  SIGNAL and_dcpl_228 : STD_LOGIC;
  SIGNAL and_dcpl_229 : STD_LOGIC;
  SIGNAL and_dcpl_230 : STD_LOGIC;
  SIGNAL and_dcpl_231 : STD_LOGIC;
  SIGNAL and_dcpl_232 : STD_LOGIC;
  SIGNAL and_dcpl_233 : STD_LOGIC;
  SIGNAL and_dcpl_234 : STD_LOGIC;
  SIGNAL and_dcpl_235 : STD_LOGIC;
  SIGNAL and_dcpl_236 : STD_LOGIC;
  SIGNAL or_tmp_2274 : STD_LOGIC;
  SIGNAL mux_tmp_2256 : STD_LOGIC;
  SIGNAL mux_tmp_2257 : STD_LOGIC;
  SIGNAL mux_tmp_2258 : STD_LOGIC;
  SIGNAL mux_tmp_2259 : STD_LOGIC;
  SIGNAL or_tmp_2277 : STD_LOGIC;
  SIGNAL or_tmp_2279 : STD_LOGIC;
  SIGNAL mux_tmp_2264 : STD_LOGIC;
  SIGNAL or_dcpl_182 : STD_LOGIC;
  SIGNAL or_dcpl_183 : STD_LOGIC;
  SIGNAL or_dcpl_184 : STD_LOGIC;
  SIGNAL mux_tmp_2282 : STD_LOGIC;
  SIGNAL nor_tmp_489 : STD_LOGIC;
  SIGNAL mux_tmp_2288 : STD_LOGIC;
  SIGNAL mux_tmp_2291 : STD_LOGIC;
  SIGNAL mux_tmp_2292 : STD_LOGIC;
  SIGNAL not_tmp_703 : STD_LOGIC;
  SIGNAL or_tmp_2300 : STD_LOGIC;
  SIGNAL or_dcpl_190 : STD_LOGIC;
  SIGNAL and_dcpl_248 : STD_LOGIC;
  SIGNAL and_dcpl_252 : STD_LOGIC;
  SIGNAL and_dcpl_255 : STD_LOGIC;
  SIGNAL nor_tmp_499 : STD_LOGIC;
  SIGNAL mux_tmp_2311 : STD_LOGIC;
  SIGNAL and_dcpl_258 : STD_LOGIC;
  SIGNAL mux_tmp_2318 : STD_LOGIC;
  SIGNAL and_dcpl_262 : STD_LOGIC;
  SIGNAL nor_tmp_507 : STD_LOGIC;
  SIGNAL and_tmp_28 : STD_LOGIC;
  SIGNAL mux_tmp_2325 : STD_LOGIC;
  SIGNAL mux_tmp_2328 : STD_LOGIC;
  SIGNAL nor_tmp_509 : STD_LOGIC;
  SIGNAL and_dcpl_266 : STD_LOGIC;
  SIGNAL not_tmp_727 : STD_LOGIC;
  SIGNAL and_dcpl_270 : STD_LOGIC;
  SIGNAL nor_tmp_515 : STD_LOGIC;
  SIGNAL mux_tmp_2344 : STD_LOGIC;
  SIGNAL mux_tmp_2347 : STD_LOGIC;
  SIGNAL mux_tmp_2348 : STD_LOGIC;
  SIGNAL mux_tmp_2351 : STD_LOGIC;
  SIGNAL and_dcpl_271 : STD_LOGIC;
  SIGNAL mux_tmp_2357 : STD_LOGIC;
  SIGNAL mux_tmp_2365 : STD_LOGIC;
  SIGNAL mux_tmp_2369 : STD_LOGIC;
  SIGNAL nor_tmp_528 : STD_LOGIC;
  SIGNAL nor_tmp_530 : STD_LOGIC;
  SIGNAL mux_tmp_2384 : STD_LOGIC;
  SIGNAL nor_tmp_537 : STD_LOGIC;
  SIGNAL mux_tmp_2392 : STD_LOGIC;
  SIGNAL mux_tmp_2395 : STD_LOGIC;
  SIGNAL nor_tmp_538 : STD_LOGIC;
  SIGNAL mux_tmp_2401 : STD_LOGIC;
  SIGNAL nor_tmp_544 : STD_LOGIC;
  SIGNAL mux_tmp_2410 : STD_LOGIC;
  SIGNAL nor_tmp_547 : STD_LOGIC;
  SIGNAL nor_tmp_548 : STD_LOGIC;
  SIGNAL not_tmp_762 : STD_LOGIC;
  SIGNAL or_dcpl_207 : STD_LOGIC;
  SIGNAL and_dcpl_277 : STD_LOGIC;
  SIGNAL or_tmp_2358 : STD_LOGIC;
  SIGNAL mux_tmp_2447 : STD_LOGIC;
  SIGNAL nand_tmp_100 : STD_LOGIC;
  SIGNAL mux_tmp_2450 : STD_LOGIC;
  SIGNAL or_tmp_2362 : STD_LOGIC;
  SIGNAL and_dcpl_286 : STD_LOGIC;
  SIGNAL or_tmp_2384 : STD_LOGIC;
  SIGNAL COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_13_psp_sva_1 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_4_sva_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL VEC_LOOP_j_10_0_sva_9_0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_10_tmp_mul_idiv_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_nor_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_13_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_1_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_14_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_3_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_16_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_9_tmp_lshift_itm : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_nor_6_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_19_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_11_tmp_mul_idiv_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_2_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_6_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_10_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_14_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_4_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_8_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_12_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_2_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_6_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_10_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_14_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_4_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_8_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_12_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_1_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_5_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_9_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_13_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_3_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_7_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_11_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_15_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_11_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_14_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_17_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_20_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_13_psp_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_16_psp_sva : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_19_psp_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_13_tmp_mul_idiv_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_5_tmp_mul_idiv_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_psp_sva : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_k_10_4_sva_5_0 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_2_sva_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL nor_1796_tmp : STD_LOGIC;
  SIGNAL nor_1798_tmp : STD_LOGIC;
  SIGNAL and_342_tmp : STD_LOGIC;
  SIGNAL and_341_tmp : STD_LOGIC;
  SIGNAL and_332_tmp : STD_LOGIC;
  SIGNAL and_314_m1c : STD_LOGIC;
  SIGNAL reg_COMP_LOOP_k_10_4_ftd : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL mux_1128_cse : STD_LOGIC;
  SIGNAL nand_271_cse : STD_LOGIC;
  SIGNAL nand_272_cse : STD_LOGIC;
  SIGNAL mux_1191_cse : STD_LOGIC;
  SIGNAL nor_346_cse : STD_LOGIC;
  SIGNAL nor_351_cse : STD_LOGIC;
  SIGNAL nor_1528_cse : STD_LOGIC;
  SIGNAL nand_265_cse : STD_LOGIC;
  SIGNAL mux_1378_cse : STD_LOGIC;
  SIGNAL nand_219_cse : STD_LOGIC;
  SIGNAL mux_1628_cse : STD_LOGIC;
  SIGNAL nand_211_cse : STD_LOGIC;
  SIGNAL nand_212_cse : STD_LOGIC;
  SIGNAL mux_1691_cse : STD_LOGIC;
  SIGNAL and_523_cse : STD_LOGIC;
  SIGNAL mux_1878_cse : STD_LOGIC;
  SIGNAL nand_122_cse : STD_LOGIC;
  SIGNAL nand_121_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_triosy_0_15_obj_ld_cse : STD_LOGIC;
  SIGNAL reg_ensig_cgo_cse : STD_LOGIC;
  SIGNAL and_421_cse : STD_LOGIC;
  SIGNAL and_831_cse : STD_LOGIC;
  SIGNAL and_407_cse : STD_LOGIC;
  SIGNAL and_733_cse : STD_LOGIC;
  SIGNAL or_432_cse : STD_LOGIC;
  SIGNAL and_674_cse : STD_LOGIC;
  SIGNAL and_675_cse : STD_LOGIC;
  SIGNAL nand_301_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_2_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_1_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_21_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_29_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_14_cse : STD_LOGIC;
  SIGNAL and_570_cse : STD_LOGIC;
  SIGNAL or_2729_cse : STD_LOGIC;
  SIGNAL and_712_cse : STD_LOGIC;
  SIGNAL nor_1792_cse : STD_LOGIC;
  SIGNAL nor_1630_cse : STD_LOGIC;
  SIGNAL nor_1624_cse : STD_LOGIC;
  SIGNAL or_36_cse : STD_LOGIC;
  SIGNAL mux_228_cse : STD_LOGIC;
  SIGNAL nor_572_cse : STD_LOGIC;
  SIGNAL or_2732_cse : STD_LOGIC;
  SIGNAL or_455_cse : STD_LOGIC;
  SIGNAL or_454_cse : STD_LOGIC;
  SIGNAL mux_464_cse : STD_LOGIC;
  SIGNAL or_610_cse : STD_LOGIC;
  SIGNAL mux_1116_cse : STD_LOGIC;
  SIGNAL nor_1523_cse : STD_LOGIC;
  SIGNAL nor_1526_cse : STD_LOGIC;
  SIGNAL nor_1527_cse : STD_LOGIC;
  SIGNAL mux_1241_cse : STD_LOGIC;
  SIGNAL nor_1402_cse : STD_LOGIC;
  SIGNAL nor_1405_cse : STD_LOGIC;
  SIGNAL nor_1406_cse : STD_LOGIC;
  SIGNAL mux_1366_cse : STD_LOGIC;
  SIGNAL nor_1286_cse : STD_LOGIC;
  SIGNAL nor_1289_cse : STD_LOGIC;
  SIGNAL nor_1290_cse : STD_LOGIC;
  SIGNAL nand_268_cse : STD_LOGIC;
  SIGNAL mux_1491_cse : STD_LOGIC;
  SIGNAL nand_261_cse : STD_LOGIC;
  SIGNAL nand_226_cse : STD_LOGIC;
  SIGNAL and_529_cse : STD_LOGIC;
  SIGNAL nor_1173_cse : STD_LOGIC;
  SIGNAL nor_1174_cse : STD_LOGIC;
  SIGNAL mux_1616_cse : STD_LOGIC;
  SIGNAL nand_222_cse : STD_LOGIC;
  SIGNAL nand_223_cse : STD_LOGIC;
  SIGNAL nor_1056_cse : STD_LOGIC;
  SIGNAL nor_1059_cse : STD_LOGIC;
  SIGNAL nor_1060_cse : STD_LOGIC;
  SIGNAL mux_1741_cse : STD_LOGIC;
  SIGNAL and_506_cse : STD_LOGIC;
  SIGNAL nor_944_cse : STD_LOGIC;
  SIGNAL nor_945_cse : STD_LOGIC;
  SIGNAL mux_1866_cse : STD_LOGIC;
  SIGNAL nand_184_cse : STD_LOGIC;
  SIGNAL nand_185_cse : STD_LOGIC;
  SIGNAL and_490_cse : STD_LOGIC;
  SIGNAL nor_837_cse : STD_LOGIC;
  SIGNAL nor_838_cse : STD_LOGIC;
  SIGNAL nand_170_cse : STD_LOGIC;
  SIGNAL mux_1991_cse : STD_LOGIC;
  SIGNAL nand_157_cse : STD_LOGIC;
  SIGNAL and_450_cse : STD_LOGIC;
  SIGNAL and_836_cse : STD_LOGIC;
  SIGNAL and_453_cse : STD_LOGIC;
  SIGNAL nor_1767_cse : STD_LOGIC;
  SIGNAL or_2589_cse : STD_LOGIC;
  SIGNAL or_2697_cse : STD_LOGIC;
  SIGNAL or_2487_cse : STD_LOGIC;
  SIGNAL or_2486_cse : STD_LOGIC;
  SIGNAL or_2612_cse : STD_LOGIC;
  SIGNAL or_2635_cse : STD_LOGIC;
  SIGNAL nor_1554_cse : STD_LOGIC;
  SIGNAL nor_1435_cse : STD_LOGIC;
  SIGNAL nor_1317_cse : STD_LOGIC;
  SIGNAL nor_1200_cse : STD_LOGIC;
  SIGNAL mux_1441_cse : STD_LOGIC;
  SIGNAL nor_1086_cse : STD_LOGIC;
  SIGNAL nor_970_cse : STD_LOGIC;
  SIGNAL nor_860_cse : STD_LOGIC;
  SIGNAL nor_761_cse : STD_LOGIC;
  SIGNAL mux_1941_cse : STD_LOGIC;
  SIGNAL mux_955_cse : STD_LOGIC;
  SIGNAL and_728_cse : STD_LOGIC;
  SIGNAL mux_559_cse : STD_LOGIC;
  SIGNAL or_2626_cse : STD_LOGIC;
  SIGNAL or_2621_cse : STD_LOGIC;
  SIGNAL and_655_cse : STD_LOGIC;
  SIGNAL or_611_cse : STD_LOGIC;
  SIGNAL mux_952_cse : STD_LOGIC;
  SIGNAL mux_949_cse : STD_LOGIC;
  SIGNAL mux_965_cse : STD_LOGIC;
  SIGNAL mux_2255_rmff : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL p_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_psp_sva : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL mux_2303_itm : STD_LOGIC;
  SIGNAL mux_2383_itm : STD_LOGIC;
  SIGNAL mux_2398_itm : STD_LOGIC;
  SIGNAL mux_2410_itm : STD_LOGIC;
  SIGNAL mux_2424_itm : STD_LOGIC;
  SIGNAL mux_2435_itm : STD_LOGIC;
  SIGNAL mux_2442_itm : STD_LOGIC;
  SIGNAL mux_2444_itm : STD_LOGIC;
  SIGNAL mux_2449_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_1_tmp_lshift_itm : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL z_out : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL z_out_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL and_dcpl_356 : STD_LOGIC;
  SIGNAL z_out_2 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL and_dcpl_360 : STD_LOGIC;
  SIGNAL and_dcpl_362 : STD_LOGIC;
  SIGNAL and_dcpl_366 : STD_LOGIC;
  SIGNAL and_dcpl_367 : STD_LOGIC;
  SIGNAL and_dcpl_370 : STD_LOGIC;
  SIGNAL and_dcpl_373 : STD_LOGIC;
  SIGNAL and_dcpl_374 : STD_LOGIC;
  SIGNAL and_dcpl_376 : STD_LOGIC;
  SIGNAL and_dcpl_377 : STD_LOGIC;
  SIGNAL and_dcpl_378 : STD_LOGIC;
  SIGNAL and_dcpl_380 : STD_LOGIC;
  SIGNAL and_dcpl_383 : STD_LOGIC;
  SIGNAL and_dcpl_384 : STD_LOGIC;
  SIGNAL and_dcpl_385 : STD_LOGIC;
  SIGNAL and_dcpl_386 : STD_LOGIC;
  SIGNAL and_dcpl_387 : STD_LOGIC;
  SIGNAL and_dcpl_389 : STD_LOGIC;
  SIGNAL and_dcpl_390 : STD_LOGIC;
  SIGNAL and_dcpl_391 : STD_LOGIC;
  SIGNAL and_dcpl_394 : STD_LOGIC;
  SIGNAL and_dcpl_395 : STD_LOGIC;
  SIGNAL and_dcpl_396 : STD_LOGIC;
  SIGNAL and_dcpl_397 : STD_LOGIC;
  SIGNAL and_dcpl_399 : STD_LOGIC;
  SIGNAL and_dcpl_400 : STD_LOGIC;
  SIGNAL and_dcpl_401 : STD_LOGIC;
  SIGNAL and_dcpl_404 : STD_LOGIC;
  SIGNAL and_dcpl_405 : STD_LOGIC;
  SIGNAL and_dcpl_406 : STD_LOGIC;
  SIGNAL and_dcpl_409 : STD_LOGIC;
  SIGNAL and_dcpl_410 : STD_LOGIC;
  SIGNAL and_dcpl_411 : STD_LOGIC;
  SIGNAL and_dcpl_412 : STD_LOGIC;
  SIGNAL and_dcpl_413 : STD_LOGIC;
  SIGNAL and_dcpl_414 : STD_LOGIC;
  SIGNAL and_dcpl_415 : STD_LOGIC;
  SIGNAL and_dcpl_416 : STD_LOGIC;
  SIGNAL and_dcpl_417 : STD_LOGIC;
  SIGNAL and_dcpl_418 : STD_LOGIC;
  SIGNAL and_dcpl_419 : STD_LOGIC;
  SIGNAL and_dcpl_420 : STD_LOGIC;
  SIGNAL and_dcpl_421 : STD_LOGIC;
  SIGNAL and_dcpl_422 : STD_LOGIC;
  SIGNAL and_dcpl_425 : STD_LOGIC;
  SIGNAL and_dcpl_426 : STD_LOGIC;
  SIGNAL and_dcpl_427 : STD_LOGIC;
  SIGNAL and_dcpl_428 : STD_LOGIC;
  SIGNAL and_dcpl_429 : STD_LOGIC;
  SIGNAL and_dcpl_430 : STD_LOGIC;
  SIGNAL and_dcpl_431 : STD_LOGIC;
  SIGNAL z_out_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL and_dcpl_447 : STD_LOGIC;
  SIGNAL z_out_4 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL and_dcpl_465 : STD_LOGIC;
  SIGNAL and_dcpl_467 : STD_LOGIC;
  SIGNAL and_dcpl_475 : STD_LOGIC;
  SIGNAL and_dcpl_477 : STD_LOGIC;
  SIGNAL and_dcpl_480 : STD_LOGIC;
  SIGNAL and_dcpl_482 : STD_LOGIC;
  SIGNAL and_dcpl_484 : STD_LOGIC;
  SIGNAL and_dcpl_486 : STD_LOGIC;
  SIGNAL and_dcpl_495 : STD_LOGIC;
  SIGNAL and_dcpl_571 : STD_LOGIC;
  SIGNAL and_dcpl_577 : STD_LOGIC;
  SIGNAL and_dcpl_589 : STD_LOGIC;
  SIGNAL z_out_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_LOOP_i_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_1_tmp_acc_cse_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_2_tmp_lshift_ncse_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL tmp_33_sva_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_33_sva_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_33_sva_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_33_sva_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_33_sva_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_33_sva_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_33_sva_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_33_sva_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_33_sva_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_33_sva_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_33_sva_11 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_33_sva_12 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_33_sva_13 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_33_sva_14 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_33_sva_15 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_3_tmp_lshift_ncse_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL tmp_36_sva_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_36_sva_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_6_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_12_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_13_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_14_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_62_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_64_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_65_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_66_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_68_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_69_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_70_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_72_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_5_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_51_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_52_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_77_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_54_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_79_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_80_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_81_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_57_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_83_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_84_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_85_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_86_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_87_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_88_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_89_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_9_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_91_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_92_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_137_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_94_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_139_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_140_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_141_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_97_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_143_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_144_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_145_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_146_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_147_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_148_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_149_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_1_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_and_185_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_13_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_131_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_132_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_197_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_134_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_199_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_200_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_201_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_137_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_203_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_204_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_205_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_206_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_207_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_208_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_209_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_2_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_and_244_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_17_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_171_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_172_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_257_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_174_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_259_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_260_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_261_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_177_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_263_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_264_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_265_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_266_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_267_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_268_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_269_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_3_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_21_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_211_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_212_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_317_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_214_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_319_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_320_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_321_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_217_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_323_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_324_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_325_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_326_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_327_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_328_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_329_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_4_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_25_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_251_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_252_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_377_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_254_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_379_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_380_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_381_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_257_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_383_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_384_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_385_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_386_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_387_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_388_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_389_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_5_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_29_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_291_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_292_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_437_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_294_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_439_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_440_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_441_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_297_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_443_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_444_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_445_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_446_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_447_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_448_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_449_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_6_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_33_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_331_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_332_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_497_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_334_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_499_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_500_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_501_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_337_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_503_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_504_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_505_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_506_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_507_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_508_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_509_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_37_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_371_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_372_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_557_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_374_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_559_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_560_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_561_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_377_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_563_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_564_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_565_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_566_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_567_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_568_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_569_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_7_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_41_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_411_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_412_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_617_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_414_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_619_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_620_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_621_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_417_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_623_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_624_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_625_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_626_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_627_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_628_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_629_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_8_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_45_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_451_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_452_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_677_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_454_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_679_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_680_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_681_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_457_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_683_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_684_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_685_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_686_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_687_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_688_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_689_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_9_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_49_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_491_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_492_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_737_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_494_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_739_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_740_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_741_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_497_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_743_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_744_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_745_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_746_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_747_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_748_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_749_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_53_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_531_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_532_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_797_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_534_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_799_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_800_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_801_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_537_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_803_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_804_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_805_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_806_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_807_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_808_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_809_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_57_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_571_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_572_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_857_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_574_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_859_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_860_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_861_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_577_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_863_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_864_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_865_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_866_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_867_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_868_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_869_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_12_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_12_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_61_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_611_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_612_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_917_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_614_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_919_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_920_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_921_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_617_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_923_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_924_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_925_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_926_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_927_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_928_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_929_itm : STD_LOGIC;
  SIGNAL STAGE_LOOP_i_3_0_sva_mx0c1 : STD_LOGIC;
  SIGNAL VEC_LOOP_j_10_0_sva_9_0_mx0c0 : STD_LOGIC;
  SIGNAL COMP_LOOP_k_10_4_sva_2 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_mux1h_4_itm_mx0w3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_33_sva_13_mx0w1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_10_acc_8_itm_mx0c2 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm_mx0c3 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm_mx0c6 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm_mx0c9 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm_mx0c12 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm_mx0c15 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm_mx0c18 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm_mx0c21 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm_mx0c24 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm_mx0c27 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm_mx0c30 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm_mx0c33 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm_mx0c36 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm_mx0c39 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm_mx0c42 : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm_mx0c47 : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_155 : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_157 : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_159 : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_161 : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_167 : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_16_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_14_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_15_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_16_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_or_17_ssc : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_27_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_17_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_1_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_23_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_3_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_6_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_19_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_31_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_20_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_21_cse : STD_LOGIC;
  SIGNAL nor_724_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_19_cse : STD_LOGIC;
  SIGNAL nor_712_cse : STD_LOGIC;
  SIGNAL nor_704_cse : STD_LOGIC;
  SIGNAL mux_2131_cse : STD_LOGIC;
  SIGNAL nor_691_cse : STD_LOGIC;
  SIGNAL nor_682_cse : STD_LOGIC;
  SIGNAL nor_670_cse : STD_LOGIC;
  SIGNAL nor_662_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_46_cse : STD_LOGIC;
  SIGNAL nor_647_cse : STD_LOGIC;
  SIGNAL nor_639_cse : STD_LOGIC;
  SIGNAL nor_627_cse : STD_LOGIC;
  SIGNAL nor_619_cse : STD_LOGIC;
  SIGNAL mux_2208_cse : STD_LOGIC;
  SIGNAL nor_606_cse : STD_LOGIC;
  SIGNAL nor_597_cse : STD_LOGIC;
  SIGNAL nor_589_cse : STD_LOGIC;
  SIGNAL and_427_cse : STD_LOGIC;
  SIGNAL mux_2465_cse : STD_LOGIC;
  SIGNAL mux_2169_cse : STD_LOGIC;
  SIGNAL and_1025_cse : STD_LOGIC;
  SIGNAL and_1028_cse : STD_LOGIC;
  SIGNAL and_1044_cse : STD_LOGIC;
  SIGNAL and_1046_cse : STD_LOGIC;
  SIGNAL and_1051_cse : STD_LOGIC;
  SIGNAL and_1052_cse : STD_LOGIC;
  SIGNAL and_1055_cse : STD_LOGIC;
  SIGNAL and_1056_cse : STD_LOGIC;
  SIGNAL and_1060_cse : STD_LOGIC;
  SIGNAL and_1061_cse : STD_LOGIC;
  SIGNAL and_1064_cse : STD_LOGIC;
  SIGNAL and_1037_cse : STD_LOGIC;
  SIGNAL and_1040_cse : STD_LOGIC;
  SIGNAL or_tmp_2410 : STD_LOGIC;
  SIGNAL or_2259_cse_1 : STD_LOGIC;
  SIGNAL and_1189_cse : STD_LOGIC;
  SIGNAL and_1191_cse : STD_LOGIC;
  SIGNAL and_1190_cse : STD_LOGIC;
  SIGNAL nand_324_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_or_40_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_621_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_or_41_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_or_43_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_622_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_or_47_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_or_52_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_or_54_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_or_18_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_2_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_3_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_4_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_5_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_6_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_7_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_8_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_9_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_10_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_11_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_12_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_13_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_14_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_15_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_16_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL STAGE_LOOP_acc_itm_4_1 : STD_LOGIC;
  SIGNAL COMP_LOOP_mux_361_cse : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL nor_1871_nl : STD_LOGIC;
  SIGNAL and_1183_nl : STD_LOGIC;
  SIGNAL nor_1589_nl : STD_LOGIC;
  SIGNAL nor_1590_nl : STD_LOGIC;
  SIGNAL mux_1190_nl : STD_LOGIC;
  SIGNAL nor_1529_nl : STD_LOGIC;
  SIGNAL nor_1530_nl : STD_LOGIC;
  SIGNAL nor_1352_nl : STD_LOGIC;
  SIGNAL nor_1353_nl : STD_LOGIC;
  SIGNAL nor_1291_nl : STD_LOGIC;
  SIGNAL mux_1440_nl : STD_LOGIC;
  SIGNAL nor_1293_nl : STD_LOGIC;
  SIGNAL nor_1121_nl : STD_LOGIC;
  SIGNAL nor_1122_nl : STD_LOGIC;
  SIGNAL mux_1690_nl : STD_LOGIC;
  SIGNAL nor_1061_nl : STD_LOGIC;
  SIGNAL nor_1062_nl : STD_LOGIC;
  SIGNAL and_503_nl : STD_LOGIC;
  SIGNAL nor_893_nl : STD_LOGIC;
  SIGNAL and_493_nl : STD_LOGIC;
  SIGNAL mux_1940_nl : STD_LOGIC;
  SIGNAL nor_839_nl : STD_LOGIC;
  SIGNAL mux_2254_nl : STD_LOGIC;
  SIGNAL mux_2253_nl : STD_LOGIC;
  SIGNAL mux_2252_nl : STD_LOGIC;
  SIGNAL mux_2251_nl : STD_LOGIC;
  SIGNAL mux_2250_nl : STD_LOGIC;
  SIGNAL mux_2249_nl : STD_LOGIC;
  SIGNAL mux_2245_nl : STD_LOGIC;
  SIGNAL mux_2242_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_j_not_1_nl : STD_LOGIC;
  SIGNAL nor_1870_nl : STD_LOGIC;
  SIGNAL and_nl : STD_LOGIC;
  SIGNAL nand_nl : STD_LOGIC;
  SIGNAL mux_1074_nl : STD_LOGIC;
  SIGNAL nor_1622_nl : STD_LOGIC;
  SIGNAL and_568_nl : STD_LOGIC;
  SIGNAL mux_2558_nl : STD_LOGIC;
  SIGNAL or_nl : STD_LOGIC;
  SIGNAL mux_nl : STD_LOGIC;
  SIGNAL nand_325_nl : STD_LOGIC;
  SIGNAL nand_323_nl : STD_LOGIC;
  SIGNAL mux_2309_nl : STD_LOGIC;
  SIGNAL mux_2308_nl : STD_LOGIC;
  SIGNAL mux_2312_nl : STD_LOGIC;
  SIGNAL and_270_nl : STD_LOGIC;
  SIGNAL mux_2314_nl : STD_LOGIC;
  SIGNAL nand_320_nl : STD_LOGIC;
  SIGNAL mux_2315_nl : STD_LOGIC;
  SIGNAL nand_111_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_3_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_2317_nl : STD_LOGIC;
  SIGNAL mux_2316_nl : STD_LOGIC;
  SIGNAL mux_2319_nl : STD_LOGIC;
  SIGNAL mux_2318_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_12_nl : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL mux_2321_nl : STD_LOGIC;
  SIGNAL mux_2320_nl : STD_LOGIC;
  SIGNAL nand_110_nl : STD_LOGIC;
  SIGNAL mux_2326_nl : STD_LOGIC;
  SIGNAL and_823_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_5_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_2327_nl : STD_LOGIC;
  SIGNAL and_412_nl : STD_LOGIC;
  SIGNAL mux_2332_nl : STD_LOGIC;
  SIGNAL mux_2331_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_6_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_2335_nl : STD_LOGIC;
  SIGNAL mux_2334_nl : STD_LOGIC;
  SIGNAL mux_2333_nl : STD_LOGIC;
  SIGNAL and_408_nl : STD_LOGIC;
  SIGNAL mux_2338_nl : STD_LOGIC;
  SIGNAL mux_2336_nl : STD_LOGIC;
  SIGNAL mux_2340_nl : STD_LOGIC;
  SIGNAL mux_2339_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_7_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_2341_nl : STD_LOGIC;
  SIGNAL and_405_nl : STD_LOGIC;
  SIGNAL mux_2346_nl : STD_LOGIC;
  SIGNAL mux_2345_nl : STD_LOGIC;
  SIGNAL mux_2349_nl : STD_LOGIC;
  SIGNAL mux_2348_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_15_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL mux_2352_nl : STD_LOGIC;
  SIGNAL mux_2351_nl : STD_LOGIC;
  SIGNAL mux_2350_nl : STD_LOGIC;
  SIGNAL mux_2354_nl : STD_LOGIC;
  SIGNAL and_296_nl : STD_LOGIC;
  SIGNAL mux_2355_nl : STD_LOGIC;
  SIGNAL and_397_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_9_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_2356_nl : STD_LOGIC;
  SIGNAL and_299_nl : STD_LOGIC;
  SIGNAL mux_2364_nl : STD_LOGIC;
  SIGNAL mux_2368_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_2372_nl : STD_LOGIC;
  SIGNAL mux_2371_nl : STD_LOGIC;
  SIGNAL mux_2375_nl : STD_LOGIC;
  SIGNAL mux_2378_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_11_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL and_390_nl : STD_LOGIC;
  SIGNAL mux_2389_nl : STD_LOGIC;
  SIGNAL mux_2392_nl : STD_LOGIC;
  SIGNAL mux_2391_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_18_nl : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL mux_2395_nl : STD_LOGIC;
  SIGNAL mux_2394_nl : STD_LOGIC;
  SIGNAL mux_2400_nl : STD_LOGIC;
  SIGNAL mux_2399_nl : STD_LOGIC;
  SIGNAL nor_581_nl : STD_LOGIC;
  SIGNAL and_379_nl : STD_LOGIC;
  SIGNAL and_380_nl : STD_LOGIC;
  SIGNAL mux_2402_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_13_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_2405_nl : STD_LOGIC;
  SIGNAL mux_2415_nl : STD_LOGIC;
  SIGNAL mux_2418_nl : STD_LOGIC;
  SIGNAL mux_2417_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_14_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_2422_nl : STD_LOGIC;
  SIGNAL mux_2421_nl : STD_LOGIC;
  SIGNAL mux_2426_nl : STD_LOGIC;
  SIGNAL mux_2425_nl : STD_LOGIC;
  SIGNAL nor_580_nl : STD_LOGIC;
  SIGNAL mux_2428_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_15_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_2431_nl : STD_LOGIC;
  SIGNAL mux_2436_nl : STD_LOGIC;
  SIGNAL mux_2438_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_21_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL nor_298_nl : STD_LOGIC;
  SIGNAL or_614_nl : STD_LOGIC;
  SIGNAL mux_951_nl : STD_LOGIC;
  SIGNAL nor_1642_nl : STD_LOGIC;
  SIGNAL and_303_nl : STD_LOGIC;
  SIGNAL and_363_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL and_304_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_17_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_19_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_20_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_21_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_23_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_24_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_25_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_26_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_27_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_28_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_29_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_11_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_12_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_14_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_17_nl : STD_LOGIC;
  SIGNAL and_311_nl : STD_LOGIC;
  SIGNAL mux_2565_nl : STD_LOGIC;
  SIGNAL mux_2564_nl : STD_LOGIC;
  SIGNAL or_2758_nl : STD_LOGIC;
  SIGNAL mux_2563_nl : STD_LOGIC;
  SIGNAL mux_2562_nl : STD_LOGIC;
  SIGNAL mux_2561_nl : STD_LOGIC;
  SIGNAL mux_2560_nl : STD_LOGIC;
  SIGNAL or_2756_nl : STD_LOGIC;
  SIGNAL or_2754_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_33_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_55_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_56_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_57_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_58_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_59_nl : STD_LOGIC;
  SIGNAL mux_2463_nl : STD_LOGIC;
  SIGNAL mux_2462_nl : STD_LOGIC;
  SIGNAL mux_2461_nl : STD_LOGIC;
  SIGNAL mux_2460_nl : STD_LOGIC;
  SIGNAL mux_2459_nl : STD_LOGIC;
  SIGNAL mux_2458_nl : STD_LOGIC;
  SIGNAL or_2563_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_23_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_mux_9_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_or_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_2_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_3_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_4_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_5_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_6_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_7_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_8_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_9_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_11_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_12_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_13_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_14_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_15_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_21_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_22_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_42_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_43_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_44_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_45_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_46_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_7_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_47_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_48_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_49_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_50_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_51_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_52_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_53_nl : STD_LOGIC;
  SIGNAL and_336_nl : STD_LOGIC;
  SIGNAL and_340_nl : STD_LOGIC;
  SIGNAL mux_2504_nl : STD_LOGIC;
  SIGNAL mux_2503_nl : STD_LOGIC;
  SIGNAL mux_2502_nl : STD_LOGIC;
  SIGNAL mux_2501_nl : STD_LOGIC;
  SIGNAL or_2595_nl : STD_LOGIC;
  SIGNAL mux_2500_nl : STD_LOGIC;
  SIGNAL mux_2499_nl : STD_LOGIC;
  SIGNAL or_2593_nl : STD_LOGIC;
  SIGNAL or_2591_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_36_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_37_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_38_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_39_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_40_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_41_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_20_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_21_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_22_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_23_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_24_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_25_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_26_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_27_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_28_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_29_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_30_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_31_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_32_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_33_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_34_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_35_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_17_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_18_nl : STD_LOGIC;
  SIGNAL mux_2518_nl : STD_LOGIC;
  SIGNAL mux_2517_nl : STD_LOGIC;
  SIGNAL mux_2516_nl : STD_LOGIC;
  SIGNAL mux_2515_nl : STD_LOGIC;
  SIGNAL mux_2514_nl : STD_LOGIC;
  SIGNAL mux_2520_nl : STD_LOGIC;
  SIGNAL mux_2519_nl : STD_LOGIC;
  SIGNAL and_357_nl : STD_LOGIC;
  SIGNAL mux_2532_nl : STD_LOGIC;
  SIGNAL mux_2531_nl : STD_LOGIC;
  SIGNAL mux_2530_nl : STD_LOGIC;
  SIGNAL mux_2529_nl : STD_LOGIC;
  SIGNAL mux_2528_nl : STD_LOGIC;
  SIGNAL mux_2527_nl : STD_LOGIC;
  SIGNAL mux_2526_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_7_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_8_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_9_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_11_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_12_nl : STD_LOGIC;
  SIGNAL mux_2542_nl : STD_LOGIC;
  SIGNAL nor_568_nl : STD_LOGIC;
  SIGNAL mux_2541_nl : STD_LOGIC;
  SIGNAL mux_2540_nl : STD_LOGIC;
  SIGNAL mux_2539_nl : STD_LOGIC;
  SIGNAL mux_2546_nl : STD_LOGIC;
  SIGNAL mux_2545_nl : STD_LOGIC;
  SIGNAL mux_2544_nl : STD_LOGIC;
  SIGNAL mux_2543_nl : STD_LOGIC;
  SIGNAL and_352_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_2_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_3_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_4_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_5_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_6_nl : STD_LOGIC;
  SIGNAL mux_2553_nl : STD_LOGIC;
  SIGNAL mux_2552_nl : STD_LOGIC;
  SIGNAL mux_2551_nl : STD_LOGIC;
  SIGNAL mux_561_nl : STD_LOGIC;
  SIGNAL mux_560_nl : STD_LOGIC;
  SIGNAL mux_2556_nl : STD_LOGIC;
  SIGNAL mux_2555_nl : STD_LOGIC;
  SIGNAL mux_2554_nl : STD_LOGIC;
  SIGNAL or_2625_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_2_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_3_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_4_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_5_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_6_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_7_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_8_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_9_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_10_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_11_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_12_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_13_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_14_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_15_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_16_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL and_313_nl : STD_LOGIC;
  SIGNAL mux_1080_nl : STD_LOGIC;
  SIGNAL and_565_nl : STD_LOGIC;
  SIGNAL or_714_nl : STD_LOGIC;
  SIGNAL nand_22_nl : STD_LOGIC;
  SIGNAL mux_1083_nl : STD_LOGIC;
  SIGNAL nand_23_nl : STD_LOGIC;
  SIGNAL mux_1085_nl : STD_LOGIC;
  SIGNAL or_712_nl : STD_LOGIC;
  SIGNAL or_762_nl : STD_LOGIC;
  SIGNAL mux_1115_nl : STD_LOGIC;
  SIGNAL or_760_nl : STD_LOGIC;
  SIGNAL or_758_nl : STD_LOGIC;
  SIGNAL nor_1479_nl : STD_LOGIC;
  SIGNAL mux_1240_nl : STD_LOGIC;
  SIGNAL nor_1480_nl : STD_LOGIC;
  SIGNAL nor_1481_nl : STD_LOGIC;
  SIGNAL or_1150_nl : STD_LOGIC;
  SIGNAL mux_1365_nl : STD_LOGIC;
  SIGNAL or_1148_nl : STD_LOGIC;
  SIGNAL or_1146_nl : STD_LOGIC;
  SIGNAL nor_1242_nl : STD_LOGIC;
  SIGNAL mux_1490_nl : STD_LOGIC;
  SIGNAL nor_1243_nl : STD_LOGIC;
  SIGNAL nor_1244_nl : STD_LOGIC;
  SIGNAL or_1538_nl : STD_LOGIC;
  SIGNAL mux_1615_nl : STD_LOGIC;
  SIGNAL or_1536_nl : STD_LOGIC;
  SIGNAL or_1534_nl : STD_LOGIC;
  SIGNAL nor_1012_nl : STD_LOGIC;
  SIGNAL mux_1740_nl : STD_LOGIC;
  SIGNAL nor_1013_nl : STD_LOGIC;
  SIGNAL nor_1014_nl : STD_LOGIC;
  SIGNAL nand_322_nl : STD_LOGIC;
  SIGNAL mux_1865_nl : STD_LOGIC;
  SIGNAL or_1922_nl : STD_LOGIC;
  SIGNAL or_1920_nl : STD_LOGIC;
  SIGNAL and_835_nl : STD_LOGIC;
  SIGNAL mux_1990_nl : STD_LOGIC;
  SIGNAL nor_795_nl : STD_LOGIC;
  SIGNAL nor_796_nl : STD_LOGIC;
  SIGNAL or_2430_nl : STD_LOGIC;
  SIGNAL or_2434_nl : STD_LOGIC;
  SIGNAL or_2435_nl : STD_LOGIC;
  SIGNAL or_2443_nl : STD_LOGIC;
  SIGNAL mux_2263_nl : STD_LOGIC;
  SIGNAL or_2444_nl : STD_LOGIC;
  SIGNAL or_2440_nl : STD_LOGIC;
  SIGNAL mux_2267_nl : STD_LOGIC;
  SIGNAL nand_114_nl : STD_LOGIC;
  SIGNAL nand_113_nl : STD_LOGIC;
  SIGNAL or_2455_nl : STD_LOGIC;
  SIGNAL or_2482_nl : STD_LOGIC;
  SIGNAL or_2481_nl : STD_LOGIC;
  SIGNAL mux_2302_nl : STD_LOGIC;
  SIGNAL mux_2306_nl : STD_LOGIC;
  SIGNAL mux_2305_nl : STD_LOGIC;
  SIGNAL and_416_nl : STD_LOGIC;
  SIGNAL mux_22_nl : STD_LOGIC;
  SIGNAL mux_2325_nl : STD_LOGIC;
  SIGNAL mux_2324_nl : STD_LOGIC;
  SIGNAL mux_2323_nl : STD_LOGIC;
  SIGNAL or_2497_nl : STD_LOGIC;
  SIGNAL mux_61_nl : STD_LOGIC;
  SIGNAL mux_2328_nl : STD_LOGIC;
  SIGNAL and_411_nl : STD_LOGIC;
  SIGNAL mux_2329_nl : STD_LOGIC;
  SIGNAL mux_2343_nl : STD_LOGIC;
  SIGNAL mux_2342_nl : STD_LOGIC;
  SIGNAL and_403_nl : STD_LOGIC;
  SIGNAL or_2507_nl : STD_LOGIC;
  SIGNAL or_2506_nl : STD_LOGIC;
  SIGNAL and_401_nl : STD_LOGIC;
  SIGNAL mux_2353_nl : STD_LOGIC;
  SIGNAL and_398_nl : STD_LOGIC;
  SIGNAL mux_2359_nl : STD_LOGIC;
  SIGNAL mux_2358_nl : STD_LOGIC;
  SIGNAL mux_2357_nl : STD_LOGIC;
  SIGNAL and_396_nl : STD_LOGIC;
  SIGNAL mux_2362_nl : STD_LOGIC;
  SIGNAL mux_2361_nl : STD_LOGIC;
  SIGNAL and_566_nl : STD_LOGIC;
  SIGNAL mux_2374_nl : STD_LOGIC;
  SIGNAL and_392_nl : STD_LOGIC;
  SIGNAL mux_2382_nl : STD_LOGIC;
  SIGNAL mux_2381_nl : STD_LOGIC;
  SIGNAL and_388_nl : STD_LOGIC;
  SIGNAL mux_2387_nl : STD_LOGIC;
  SIGNAL mux_2386_nl : STD_LOGIC;
  SIGNAL mux_2397_nl : STD_LOGIC;
  SIGNAL mux_2409_nl : STD_LOGIC;
  SIGNAL mux_2408_nl : STD_LOGIC;
  SIGNAL mux_2407_nl : STD_LOGIC;
  SIGNAL and_376_nl : STD_LOGIC;
  SIGNAL mux_2413_nl : STD_LOGIC;
  SIGNAL mux_2412_nl : STD_LOGIC;
  SIGNAL and_372_nl : STD_LOGIC;
  SIGNAL and_370_nl : STD_LOGIC;
  SIGNAL mux_2434_nl : STD_LOGIC;
  SIGNAL mux_2433_nl : STD_LOGIC;
  SIGNAL and_366_nl : STD_LOGIC;
  SIGNAL mux_2441_nl : STD_LOGIC;
  SIGNAL mux_2440_nl : STD_LOGIC;
  SIGNAL mux_2443_nl : STD_LOGIC;
  SIGNAL mux_2448_nl : STD_LOGIC;
  SIGNAL or_427_nl : STD_LOGIC;
  SIGNAL or_2571_nl : STD_LOGIC;
  SIGNAL mux_2468_nl : STD_LOGIC;
  SIGNAL and_361_nl : STD_LOGIC;
  SIGNAL nor_577_nl : STD_LOGIC;
  SIGNAL nor_576_nl : STD_LOGIC;
  SIGNAL mux_2471_nl : STD_LOGIC;
  SIGNAL nand_103_nl : STD_LOGIC;
  SIGNAL and_360_nl : STD_LOGIC;
  SIGNAL mux_2470_nl : STD_LOGIC;
  SIGNAL nand_101_nl : STD_LOGIC;
  SIGNAL mux_2467_nl : STD_LOGIC;
  SIGNAL or_2569_nl : STD_LOGIC;
  SIGNAL STAGE_LOOP_acc_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL mux_2498_nl : STD_LOGIC;
  SIGNAL nor_575_nl : STD_LOGIC;
  SIGNAL mux_27_nl : STD_LOGIC;
  SIGNAL or_44_nl : STD_LOGIC;
  SIGNAL mux_2509_nl : STD_LOGIC;
  SIGNAL mux_2508_nl : STD_LOGIC;
  SIGNAL mux_2507_nl : STD_LOGIC;
  SIGNAL nand_107_nl : STD_LOGIC;
  SIGNAL mux_2512_nl : STD_LOGIC;
  SIGNAL nor_570_nl : STD_LOGIC;
  SIGNAL mux_2511_nl : STD_LOGIC;
  SIGNAL mux_2510_nl : STD_LOGIC;
  SIGNAL mux_2525_nl : STD_LOGIC;
  SIGNAL mux_2524_nl : STD_LOGIC;
  SIGNAL mux_2523_nl : STD_LOGIC;
  SIGNAL and_354_nl : STD_LOGIC;
  SIGNAL mux_2522_nl : STD_LOGIC;
  SIGNAL and_356_nl : STD_LOGIC;
  SIGNAL mux_2538_nl : STD_LOGIC;
  SIGNAL mux_2537_nl : STD_LOGIC;
  SIGNAL mux_2536_nl : STD_LOGIC;
  SIGNAL mux_234_nl : STD_LOGIC;
  SIGNAL nor_1750_nl : STD_LOGIC;
  SIGNAL mux_233_nl : STD_LOGIC;
  SIGNAL mux_232_nl : STD_LOGIC;
  SIGNAL mux_1089_nl : STD_LOGIC;
  SIGNAL mux_1088_nl : STD_LOGIC;
  SIGNAL or_715_nl : STD_LOGIC;
  SIGNAL mux_1087_nl : STD_LOGIC;
  SIGNAL or_711_nl : STD_LOGIC;
  SIGNAL and_94_nl : STD_LOGIC;
  SIGNAL and_99_nl : STD_LOGIC;
  SIGNAL and_106_nl : STD_LOGIC;
  SIGNAL and_110_nl : STD_LOGIC;
  SIGNAL and_116_nl : STD_LOGIC;
  SIGNAL and_120_nl : STD_LOGIC;
  SIGNAL and_124_nl : STD_LOGIC;
  SIGNAL and_127_nl : STD_LOGIC;
  SIGNAL and_132_nl : STD_LOGIC;
  SIGNAL and_135_nl : STD_LOGIC;
  SIGNAL and_140_nl : STD_LOGIC;
  SIGNAL and_143_nl : STD_LOGIC;
  SIGNAL and_148_nl : STD_LOGIC;
  SIGNAL and_152_nl : STD_LOGIC;
  SIGNAL and_155_nl : STD_LOGIC;
  SIGNAL and_158_nl : STD_LOGIC;
  SIGNAL and_159_nl : STD_LOGIC;
  SIGNAL and_160_nl : STD_LOGIC;
  SIGNAL and_161_nl : STD_LOGIC;
  SIGNAL and_163_nl : STD_LOGIC;
  SIGNAL and_164_nl : STD_LOGIC;
  SIGNAL and_165_nl : STD_LOGIC;
  SIGNAL and_166_nl : STD_LOGIC;
  SIGNAL and_168_nl : STD_LOGIC;
  SIGNAL and_169_nl : STD_LOGIC;
  SIGNAL and_170_nl : STD_LOGIC;
  SIGNAL and_171_nl : STD_LOGIC;
  SIGNAL and_173_nl : STD_LOGIC;
  SIGNAL and_174_nl : STD_LOGIC;
  SIGNAL and_175_nl : STD_LOGIC;
  SIGNAL and_176_nl : STD_LOGIC;
  SIGNAL and_178_nl : STD_LOGIC;
  SIGNAL and_179_nl : STD_LOGIC;
  SIGNAL and_180_nl : STD_LOGIC;
  SIGNAL and_181_nl : STD_LOGIC;
  SIGNAL and_183_nl : STD_LOGIC;
  SIGNAL and_184_nl : STD_LOGIC;
  SIGNAL and_185_nl : STD_LOGIC;
  SIGNAL and_186_nl : STD_LOGIC;
  SIGNAL and_188_nl : STD_LOGIC;
  SIGNAL and_189_nl : STD_LOGIC;
  SIGNAL and_190_nl : STD_LOGIC;
  SIGNAL and_191_nl : STD_LOGIC;
  SIGNAL and_193_nl : STD_LOGIC;
  SIGNAL and_194_nl : STD_LOGIC;
  SIGNAL and_195_nl : STD_LOGIC;
  SIGNAL and_196_nl : STD_LOGIC;
  SIGNAL nor_1596_nl : STD_LOGIC;
  SIGNAL mux_1119_nl : STD_LOGIC;
  SIGNAL mux_1118_nl : STD_LOGIC;
  SIGNAL nor_1597_nl : STD_LOGIC;
  SIGNAL mux_1117_nl : STD_LOGIC;
  SIGNAL or_763_nl : STD_LOGIC;
  SIGNAL mux_1114_nl : STD_LOGIC;
  SIGNAL mux_1113_nl : STD_LOGIC;
  SIGNAL or_757_nl : STD_LOGIC;
  SIGNAL or_755_nl : STD_LOGIC;
  SIGNAL mux_1112_nl : STD_LOGIC;
  SIGNAL or_753_nl : STD_LOGIC;
  SIGNAL or_752_nl : STD_LOGIC;
  SIGNAL mux_1111_nl : STD_LOGIC;
  SIGNAL mux_1110_nl : STD_LOGIC;
  SIGNAL mux_1109_nl : STD_LOGIC;
  SIGNAL nor_1598_nl : STD_LOGIC;
  SIGNAL nor_1599_nl : STD_LOGIC;
  SIGNAL mux_1108_nl : STD_LOGIC;
  SIGNAL nor_1600_nl : STD_LOGIC;
  SIGNAL nor_1601_nl : STD_LOGIC;
  SIGNAL mux_1107_nl : STD_LOGIC;
  SIGNAL mux_1106_nl : STD_LOGIC;
  SIGNAL nor_1602_nl : STD_LOGIC;
  SIGNAL nor_1603_nl : STD_LOGIC;
  SIGNAL mux_1105_nl : STD_LOGIC;
  SIGNAL nor_1604_nl : STD_LOGIC;
  SIGNAL nor_1605_nl : STD_LOGIC;
  SIGNAL mux_1104_nl : STD_LOGIC;
  SIGNAL mux_1103_nl : STD_LOGIC;
  SIGNAL mux_1102_nl : STD_LOGIC;
  SIGNAL mux_1101_nl : STD_LOGIC;
  SIGNAL nor_1606_nl : STD_LOGIC;
  SIGNAL nor_1607_nl : STD_LOGIC;
  SIGNAL mux_1100_nl : STD_LOGIC;
  SIGNAL nor_1608_nl : STD_LOGIC;
  SIGNAL nor_1609_nl : STD_LOGIC;
  SIGNAL mux_1099_nl : STD_LOGIC;
  SIGNAL mux_1098_nl : STD_LOGIC;
  SIGNAL nor_1610_nl : STD_LOGIC;
  SIGNAL nor_1611_nl : STD_LOGIC;
  SIGNAL mux_1097_nl : STD_LOGIC;
  SIGNAL nor_1612_nl : STD_LOGIC;
  SIGNAL nor_1613_nl : STD_LOGIC;
  SIGNAL mux_1096_nl : STD_LOGIC;
  SIGNAL mux_1095_nl : STD_LOGIC;
  SIGNAL mux_1094_nl : STD_LOGIC;
  SIGNAL nor_1614_nl : STD_LOGIC;
  SIGNAL nor_1615_nl : STD_LOGIC;
  SIGNAL mux_1093_nl : STD_LOGIC;
  SIGNAL nor_1616_nl : STD_LOGIC;
  SIGNAL nor_1617_nl : STD_LOGIC;
  SIGNAL mux_1092_nl : STD_LOGIC;
  SIGNAL mux_1091_nl : STD_LOGIC;
  SIGNAL nor_1618_nl : STD_LOGIC;
  SIGNAL nor_1619_nl : STD_LOGIC;
  SIGNAL mux_1090_nl : STD_LOGIC;
  SIGNAL nor_1620_nl : STD_LOGIC;
  SIGNAL nor_1621_nl : STD_LOGIC;
  SIGNAL mux_1150_nl : STD_LOGIC;
  SIGNAL mux_1149_nl : STD_LOGIC;
  SIGNAL mux_1148_nl : STD_LOGIC;
  SIGNAL nor_1569_nl : STD_LOGIC;
  SIGNAL mux_1147_nl : STD_LOGIC;
  SIGNAL mux_1146_nl : STD_LOGIC;
  SIGNAL nor_1570_nl : STD_LOGIC;
  SIGNAL nor_1571_nl : STD_LOGIC;
  SIGNAL nor_1572_nl : STD_LOGIC;
  SIGNAL mux_1145_nl : STD_LOGIC;
  SIGNAL mux_1144_nl : STD_LOGIC;
  SIGNAL mux_1143_nl : STD_LOGIC;
  SIGNAL nor_1573_nl : STD_LOGIC;
  SIGNAL nor_1574_nl : STD_LOGIC;
  SIGNAL nor_1575_nl : STD_LOGIC;
  SIGNAL nor_1576_nl : STD_LOGIC;
  SIGNAL mux_1142_nl : STD_LOGIC;
  SIGNAL mux_1141_nl : STD_LOGIC;
  SIGNAL mux_1140_nl : STD_LOGIC;
  SIGNAL nor_1577_nl : STD_LOGIC;
  SIGNAL mux_1139_nl : STD_LOGIC;
  SIGNAL nor_1578_nl : STD_LOGIC;
  SIGNAL nor_1579_nl : STD_LOGIC;
  SIGNAL nor_1580_nl : STD_LOGIC;
  SIGNAL mux_1138_nl : STD_LOGIC;
  SIGNAL nor_1581_nl : STD_LOGIC;
  SIGNAL mux_1137_nl : STD_LOGIC;
  SIGNAL mux_1136_nl : STD_LOGIC;
  SIGNAL nor_1582_nl : STD_LOGIC;
  SIGNAL nor_1583_nl : STD_LOGIC;
  SIGNAL nor_1584_nl : STD_LOGIC;
  SIGNAL mux_1135_nl : STD_LOGIC;
  SIGNAL mux_1134_nl : STD_LOGIC;
  SIGNAL mux_1133_nl : STD_LOGIC;
  SIGNAL and_561_nl : STD_LOGIC;
  SIGNAL mux_1132_nl : STD_LOGIC;
  SIGNAL nor_1585_nl : STD_LOGIC;
  SIGNAL nor_1586_nl : STD_LOGIC;
  SIGNAL nor_1587_nl : STD_LOGIC;
  SIGNAL mux_1131_nl : STD_LOGIC;
  SIGNAL or_785_nl : STD_LOGIC;
  SIGNAL or_783_nl : STD_LOGIC;
  SIGNAL mux_1130_nl : STD_LOGIC;
  SIGNAL nor_1588_nl : STD_LOGIC;
  SIGNAL mux_1129_nl : STD_LOGIC;
  SIGNAL or_781_nl : STD_LOGIC;
  SIGNAL or_779_nl : STD_LOGIC;
  SIGNAL and_562_nl : STD_LOGIC;
  SIGNAL mux_1127_nl : STD_LOGIC;
  SIGNAL nor_1591_nl : STD_LOGIC;
  SIGNAL mux_1126_nl : STD_LOGIC;
  SIGNAL mux_1125_nl : STD_LOGIC;
  SIGNAL or_775_nl : STD_LOGIC;
  SIGNAL or_773_nl : STD_LOGIC;
  SIGNAL mux_1124_nl : STD_LOGIC;
  SIGNAL or_772_nl : STD_LOGIC;
  SIGNAL or_770_nl : STD_LOGIC;
  SIGNAL and_563_nl : STD_LOGIC;
  SIGNAL mux_1123_nl : STD_LOGIC;
  SIGNAL mux_1122_nl : STD_LOGIC;
  SIGNAL nor_1592_nl : STD_LOGIC;
  SIGNAL nor_1593_nl : STD_LOGIC;
  SIGNAL mux_1121_nl : STD_LOGIC;
  SIGNAL nor_1594_nl : STD_LOGIC;
  SIGNAL nor_1595_nl : STD_LOGIC;
  SIGNAL nor_1539_nl : STD_LOGIC;
  SIGNAL mux_1181_nl : STD_LOGIC;
  SIGNAL mux_1180_nl : STD_LOGIC;
  SIGNAL and_560_nl : STD_LOGIC;
  SIGNAL mux_1179_nl : STD_LOGIC;
  SIGNAL nor_1540_nl : STD_LOGIC;
  SIGNAL mux_1176_nl : STD_LOGIC;
  SIGNAL mux_1175_nl : STD_LOGIC;
  SIGNAL nor_1541_nl : STD_LOGIC;
  SIGNAL nor_1542_nl : STD_LOGIC;
  SIGNAL mux_1174_nl : STD_LOGIC;
  SIGNAL nor_1543_nl : STD_LOGIC;
  SIGNAL nor_1544_nl : STD_LOGIC;
  SIGNAL mux_1173_nl : STD_LOGIC;
  SIGNAL mux_1172_nl : STD_LOGIC;
  SIGNAL mux_1171_nl : STD_LOGIC;
  SIGNAL nor_1545_nl : STD_LOGIC;
  SIGNAL nor_1546_nl : STD_LOGIC;
  SIGNAL mux_1170_nl : STD_LOGIC;
  SIGNAL nor_1547_nl : STD_LOGIC;
  SIGNAL nor_1548_nl : STD_LOGIC;
  SIGNAL mux_1169_nl : STD_LOGIC;
  SIGNAL mux_1168_nl : STD_LOGIC;
  SIGNAL nor_1549_nl : STD_LOGIC;
  SIGNAL nor_1550_nl : STD_LOGIC;
  SIGNAL mux_1167_nl : STD_LOGIC;
  SIGNAL nor_1551_nl : STD_LOGIC;
  SIGNAL nor_1552_nl : STD_LOGIC;
  SIGNAL mux_1166_nl : STD_LOGIC;
  SIGNAL mux_1165_nl : STD_LOGIC;
  SIGNAL mux_1164_nl : STD_LOGIC;
  SIGNAL mux_1163_nl : STD_LOGIC;
  SIGNAL nor_1553_nl : STD_LOGIC;
  SIGNAL mux_1162_nl : STD_LOGIC;
  SIGNAL nor_1556_nl : STD_LOGIC;
  SIGNAL mux_1161_nl : STD_LOGIC;
  SIGNAL mux_1160_nl : STD_LOGIC;
  SIGNAL nor_1557_nl : STD_LOGIC;
  SIGNAL mux_1159_nl : STD_LOGIC;
  SIGNAL nor_1560_nl : STD_LOGIC;
  SIGNAL mux_1158_nl : STD_LOGIC;
  SIGNAL mux_1157_nl : STD_LOGIC;
  SIGNAL mux_1156_nl : STD_LOGIC;
  SIGNAL nor_1561_nl : STD_LOGIC;
  SIGNAL nor_1562_nl : STD_LOGIC;
  SIGNAL mux_1155_nl : STD_LOGIC;
  SIGNAL nor_1563_nl : STD_LOGIC;
  SIGNAL nor_1564_nl : STD_LOGIC;
  SIGNAL mux_1154_nl : STD_LOGIC;
  SIGNAL mux_1153_nl : STD_LOGIC;
  SIGNAL nor_1565_nl : STD_LOGIC;
  SIGNAL nor_1566_nl : STD_LOGIC;
  SIGNAL mux_1152_nl : STD_LOGIC;
  SIGNAL nor_1567_nl : STD_LOGIC;
  SIGNAL nor_1568_nl : STD_LOGIC;
  SIGNAL mux_1213_nl : STD_LOGIC;
  SIGNAL mux_1212_nl : STD_LOGIC;
  SIGNAL mux_1211_nl : STD_LOGIC;
  SIGNAL mux_1210_nl : STD_LOGIC;
  SIGNAL nor_1506_nl : STD_LOGIC;
  SIGNAL nor_1507_nl : STD_LOGIC;
  SIGNAL mux_1209_nl : STD_LOGIC;
  SIGNAL nor_1508_nl : STD_LOGIC;
  SIGNAL nor_1509_nl : STD_LOGIC;
  SIGNAL mux_1208_nl : STD_LOGIC;
  SIGNAL mux_1207_nl : STD_LOGIC;
  SIGNAL nor_1510_nl : STD_LOGIC;
  SIGNAL nor_1511_nl : STD_LOGIC;
  SIGNAL nor_1512_nl : STD_LOGIC;
  SIGNAL mux_1206_nl : STD_LOGIC;
  SIGNAL mux_1205_nl : STD_LOGIC;
  SIGNAL mux_1204_nl : STD_LOGIC;
  SIGNAL nor_1513_nl : STD_LOGIC;
  SIGNAL nor_1514_nl : STD_LOGIC;
  SIGNAL mux_1203_nl : STD_LOGIC;
  SIGNAL nor_1515_nl : STD_LOGIC;
  SIGNAL nor_1516_nl : STD_LOGIC;
  SIGNAL mux_1202_nl : STD_LOGIC;
  SIGNAL mux_1201_nl : STD_LOGIC;
  SIGNAL nor_1517_nl : STD_LOGIC;
  SIGNAL nor_1518_nl : STD_LOGIC;
  SIGNAL mux_1200_nl : STD_LOGIC;
  SIGNAL mux_1199_nl : STD_LOGIC;
  SIGNAL nor_1519_nl : STD_LOGIC;
  SIGNAL nor_1520_nl : STD_LOGIC;
  SIGNAL nor_1521_nl : STD_LOGIC;
  SIGNAL and_557_nl : STD_LOGIC;
  SIGNAL mux_1198_nl : STD_LOGIC;
  SIGNAL mux_1197_nl : STD_LOGIC;
  SIGNAL mux_1196_nl : STD_LOGIC;
  SIGNAL mux_1195_nl : STD_LOGIC;
  SIGNAL and_558_nl : STD_LOGIC;
  SIGNAL mux_1194_nl : STD_LOGIC;
  SIGNAL nor_1524_nl : STD_LOGIC;
  SIGNAL nor_1525_nl : STD_LOGIC;
  SIGNAL mux_1193_nl : STD_LOGIC;
  SIGNAL mux_1192_nl : STD_LOGIC;
  SIGNAL and_559_nl : STD_LOGIC;
  SIGNAL mux_1189_nl : STD_LOGIC;
  SIGNAL mux_1188_nl : STD_LOGIC;
  SIGNAL mux_1187_nl : STD_LOGIC;
  SIGNAL nor_1531_nl : STD_LOGIC;
  SIGNAL nor_1532_nl : STD_LOGIC;
  SIGNAL mux_1186_nl : STD_LOGIC;
  SIGNAL nor_1533_nl : STD_LOGIC;
  SIGNAL nor_1534_nl : STD_LOGIC;
  SIGNAL mux_1185_nl : STD_LOGIC;
  SIGNAL mux_1184_nl : STD_LOGIC;
  SIGNAL nor_1535_nl : STD_LOGIC;
  SIGNAL nor_1536_nl : STD_LOGIC;
  SIGNAL mux_1183_nl : STD_LOGIC;
  SIGNAL nor_1537_nl : STD_LOGIC;
  SIGNAL nor_1538_nl : STD_LOGIC;
  SIGNAL nor_1477_nl : STD_LOGIC;
  SIGNAL mux_1244_nl : STD_LOGIC;
  SIGNAL mux_1243_nl : STD_LOGIC;
  SIGNAL nor_1478_nl : STD_LOGIC;
  SIGNAL mux_1242_nl : STD_LOGIC;
  SIGNAL nand_31_nl : STD_LOGIC;
  SIGNAL mux_1239_nl : STD_LOGIC;
  SIGNAL mux_1238_nl : STD_LOGIC;
  SIGNAL or_952_nl : STD_LOGIC;
  SIGNAL or_950_nl : STD_LOGIC;
  SIGNAL mux_1237_nl : STD_LOGIC;
  SIGNAL or_948_nl : STD_LOGIC;
  SIGNAL or_947_nl : STD_LOGIC;
  SIGNAL mux_1236_nl : STD_LOGIC;
  SIGNAL mux_1235_nl : STD_LOGIC;
  SIGNAL mux_1234_nl : STD_LOGIC;
  SIGNAL nor_1482_nl : STD_LOGIC;
  SIGNAL nor_1483_nl : STD_LOGIC;
  SIGNAL mux_1233_nl : STD_LOGIC;
  SIGNAL nor_1484_nl : STD_LOGIC;
  SIGNAL nor_1485_nl : STD_LOGIC;
  SIGNAL mux_1232_nl : STD_LOGIC;
  SIGNAL mux_1231_nl : STD_LOGIC;
  SIGNAL nor_1486_nl : STD_LOGIC;
  SIGNAL nor_1487_nl : STD_LOGIC;
  SIGNAL mux_1230_nl : STD_LOGIC;
  SIGNAL nor_1488_nl : STD_LOGIC;
  SIGNAL nor_1489_nl : STD_LOGIC;
  SIGNAL mux_1229_nl : STD_LOGIC;
  SIGNAL mux_1228_nl : STD_LOGIC;
  SIGNAL mux_1227_nl : STD_LOGIC;
  SIGNAL mux_1226_nl : STD_LOGIC;
  SIGNAL nor_1490_nl : STD_LOGIC;
  SIGNAL nor_1491_nl : STD_LOGIC;
  SIGNAL mux_1225_nl : STD_LOGIC;
  SIGNAL nor_1492_nl : STD_LOGIC;
  SIGNAL nor_1493_nl : STD_LOGIC;
  SIGNAL mux_1224_nl : STD_LOGIC;
  SIGNAL mux_1223_nl : STD_LOGIC;
  SIGNAL nor_1494_nl : STD_LOGIC;
  SIGNAL nor_1495_nl : STD_LOGIC;
  SIGNAL mux_1222_nl : STD_LOGIC;
  SIGNAL nor_1496_nl : STD_LOGIC;
  SIGNAL nor_1497_nl : STD_LOGIC;
  SIGNAL mux_1221_nl : STD_LOGIC;
  SIGNAL mux_1220_nl : STD_LOGIC;
  SIGNAL mux_1219_nl : STD_LOGIC;
  SIGNAL nor_1498_nl : STD_LOGIC;
  SIGNAL nor_1499_nl : STD_LOGIC;
  SIGNAL mux_1218_nl : STD_LOGIC;
  SIGNAL nor_1500_nl : STD_LOGIC;
  SIGNAL nor_1501_nl : STD_LOGIC;
  SIGNAL mux_1217_nl : STD_LOGIC;
  SIGNAL mux_1216_nl : STD_LOGIC;
  SIGNAL nor_1502_nl : STD_LOGIC;
  SIGNAL nor_1503_nl : STD_LOGIC;
  SIGNAL mux_1215_nl : STD_LOGIC;
  SIGNAL nor_1504_nl : STD_LOGIC;
  SIGNAL nor_1505_nl : STD_LOGIC;
  SIGNAL mux_1275_nl : STD_LOGIC;
  SIGNAL mux_1274_nl : STD_LOGIC;
  SIGNAL mux_1273_nl : STD_LOGIC;
  SIGNAL nor_1450_nl : STD_LOGIC;
  SIGNAL mux_1272_nl : STD_LOGIC;
  SIGNAL mux_1271_nl : STD_LOGIC;
  SIGNAL nor_1451_nl : STD_LOGIC;
  SIGNAL nor_1452_nl : STD_LOGIC;
  SIGNAL nor_1453_nl : STD_LOGIC;
  SIGNAL mux_1270_nl : STD_LOGIC;
  SIGNAL mux_1269_nl : STD_LOGIC;
  SIGNAL mux_1268_nl : STD_LOGIC;
  SIGNAL nor_1454_nl : STD_LOGIC;
  SIGNAL nor_1455_nl : STD_LOGIC;
  SIGNAL nor_1456_nl : STD_LOGIC;
  SIGNAL nor_1457_nl : STD_LOGIC;
  SIGNAL mux_1267_nl : STD_LOGIC;
  SIGNAL mux_1266_nl : STD_LOGIC;
  SIGNAL mux_1265_nl : STD_LOGIC;
  SIGNAL nor_1458_nl : STD_LOGIC;
  SIGNAL mux_1264_nl : STD_LOGIC;
  SIGNAL nor_1459_nl : STD_LOGIC;
  SIGNAL nor_1460_nl : STD_LOGIC;
  SIGNAL nor_1461_nl : STD_LOGIC;
  SIGNAL mux_1263_nl : STD_LOGIC;
  SIGNAL nor_1462_nl : STD_LOGIC;
  SIGNAL mux_1262_nl : STD_LOGIC;
  SIGNAL mux_1261_nl : STD_LOGIC;
  SIGNAL nor_1463_nl : STD_LOGIC;
  SIGNAL nor_1464_nl : STD_LOGIC;
  SIGNAL nor_1465_nl : STD_LOGIC;
  SIGNAL mux_1260_nl : STD_LOGIC;
  SIGNAL mux_1259_nl : STD_LOGIC;
  SIGNAL mux_1258_nl : STD_LOGIC;
  SIGNAL and_554_nl : STD_LOGIC;
  SIGNAL mux_1257_nl : STD_LOGIC;
  SIGNAL nor_1466_nl : STD_LOGIC;
  SIGNAL nor_1467_nl : STD_LOGIC;
  SIGNAL nor_1468_nl : STD_LOGIC;
  SIGNAL mux_1256_nl : STD_LOGIC;
  SIGNAL or_979_nl : STD_LOGIC;
  SIGNAL or_977_nl : STD_LOGIC;
  SIGNAL mux_1255_nl : STD_LOGIC;
  SIGNAL nor_1469_nl : STD_LOGIC;
  SIGNAL mux_1254_nl : STD_LOGIC;
  SIGNAL or_975_nl : STD_LOGIC;
  SIGNAL or_973_nl : STD_LOGIC;
  SIGNAL and_555_nl : STD_LOGIC;
  SIGNAL mux_1252_nl : STD_LOGIC;
  SIGNAL nor_1472_nl : STD_LOGIC;
  SIGNAL mux_1251_nl : STD_LOGIC;
  SIGNAL mux_1250_nl : STD_LOGIC;
  SIGNAL or_969_nl : STD_LOGIC;
  SIGNAL or_967_nl : STD_LOGIC;
  SIGNAL mux_1249_nl : STD_LOGIC;
  SIGNAL or_966_nl : STD_LOGIC;
  SIGNAL or_964_nl : STD_LOGIC;
  SIGNAL and_556_nl : STD_LOGIC;
  SIGNAL mux_1248_nl : STD_LOGIC;
  SIGNAL mux_1247_nl : STD_LOGIC;
  SIGNAL nor_1473_nl : STD_LOGIC;
  SIGNAL nor_1474_nl : STD_LOGIC;
  SIGNAL mux_1246_nl : STD_LOGIC;
  SIGNAL nor_1475_nl : STD_LOGIC;
  SIGNAL nor_1476_nl : STD_LOGIC;
  SIGNAL nor_1418_nl : STD_LOGIC;
  SIGNAL mux_1306_nl : STD_LOGIC;
  SIGNAL mux_1305_nl : STD_LOGIC;
  SIGNAL and_552_nl : STD_LOGIC;
  SIGNAL mux_1304_nl : STD_LOGIC;
  SIGNAL and_553_nl : STD_LOGIC;
  SIGNAL mux_1301_nl : STD_LOGIC;
  SIGNAL mux_1300_nl : STD_LOGIC;
  SIGNAL nor_1422_nl : STD_LOGIC;
  SIGNAL nor_1423_nl : STD_LOGIC;
  SIGNAL mux_1299_nl : STD_LOGIC;
  SIGNAL nor_1424_nl : STD_LOGIC;
  SIGNAL nor_1425_nl : STD_LOGIC;
  SIGNAL mux_1298_nl : STD_LOGIC;
  SIGNAL mux_1297_nl : STD_LOGIC;
  SIGNAL mux_1296_nl : STD_LOGIC;
  SIGNAL nor_1426_nl : STD_LOGIC;
  SIGNAL nor_1427_nl : STD_LOGIC;
  SIGNAL mux_1295_nl : STD_LOGIC;
  SIGNAL nor_1428_nl : STD_LOGIC;
  SIGNAL nor_1429_nl : STD_LOGIC;
  SIGNAL mux_1294_nl : STD_LOGIC;
  SIGNAL mux_1293_nl : STD_LOGIC;
  SIGNAL nor_1430_nl : STD_LOGIC;
  SIGNAL nor_1431_nl : STD_LOGIC;
  SIGNAL mux_1292_nl : STD_LOGIC;
  SIGNAL nor_1432_nl : STD_LOGIC;
  SIGNAL nor_1433_nl : STD_LOGIC;
  SIGNAL mux_1291_nl : STD_LOGIC;
  SIGNAL mux_1290_nl : STD_LOGIC;
  SIGNAL mux_1289_nl : STD_LOGIC;
  SIGNAL mux_1288_nl : STD_LOGIC;
  SIGNAL nor_1434_nl : STD_LOGIC;
  SIGNAL mux_1287_nl : STD_LOGIC;
  SIGNAL nor_1437_nl : STD_LOGIC;
  SIGNAL mux_1286_nl : STD_LOGIC;
  SIGNAL mux_1285_nl : STD_LOGIC;
  SIGNAL nor_1438_nl : STD_LOGIC;
  SIGNAL mux_1284_nl : STD_LOGIC;
  SIGNAL nor_1441_nl : STD_LOGIC;
  SIGNAL mux_1283_nl : STD_LOGIC;
  SIGNAL mux_1282_nl : STD_LOGIC;
  SIGNAL mux_1281_nl : STD_LOGIC;
  SIGNAL nor_1442_nl : STD_LOGIC;
  SIGNAL nor_1443_nl : STD_LOGIC;
  SIGNAL mux_1280_nl : STD_LOGIC;
  SIGNAL nor_1444_nl : STD_LOGIC;
  SIGNAL nor_1445_nl : STD_LOGIC;
  SIGNAL mux_1279_nl : STD_LOGIC;
  SIGNAL mux_1278_nl : STD_LOGIC;
  SIGNAL nor_1446_nl : STD_LOGIC;
  SIGNAL nor_1447_nl : STD_LOGIC;
  SIGNAL mux_1277_nl : STD_LOGIC;
  SIGNAL nor_1448_nl : STD_LOGIC;
  SIGNAL nor_1449_nl : STD_LOGIC;
  SIGNAL mux_1338_nl : STD_LOGIC;
  SIGNAL mux_1337_nl : STD_LOGIC;
  SIGNAL mux_1336_nl : STD_LOGIC;
  SIGNAL mux_1335_nl : STD_LOGIC;
  SIGNAL nor_1385_nl : STD_LOGIC;
  SIGNAL nor_1386_nl : STD_LOGIC;
  SIGNAL mux_1334_nl : STD_LOGIC;
  SIGNAL nor_1387_nl : STD_LOGIC;
  SIGNAL nor_1388_nl : STD_LOGIC;
  SIGNAL mux_1333_nl : STD_LOGIC;
  SIGNAL mux_1332_nl : STD_LOGIC;
  SIGNAL nor_1389_nl : STD_LOGIC;
  SIGNAL nor_1390_nl : STD_LOGIC;
  SIGNAL nor_1391_nl : STD_LOGIC;
  SIGNAL mux_1331_nl : STD_LOGIC;
  SIGNAL mux_1330_nl : STD_LOGIC;
  SIGNAL mux_1329_nl : STD_LOGIC;
  SIGNAL nor_1392_nl : STD_LOGIC;
  SIGNAL nor_1393_nl : STD_LOGIC;
  SIGNAL mux_1328_nl : STD_LOGIC;
  SIGNAL nor_1394_nl : STD_LOGIC;
  SIGNAL nor_1395_nl : STD_LOGIC;
  SIGNAL mux_1327_nl : STD_LOGIC;
  SIGNAL mux_1326_nl : STD_LOGIC;
  SIGNAL nor_1396_nl : STD_LOGIC;
  SIGNAL nor_1397_nl : STD_LOGIC;
  SIGNAL mux_1325_nl : STD_LOGIC;
  SIGNAL mux_1324_nl : STD_LOGIC;
  SIGNAL nor_1398_nl : STD_LOGIC;
  SIGNAL nor_1399_nl : STD_LOGIC;
  SIGNAL nor_1400_nl : STD_LOGIC;
  SIGNAL and_549_nl : STD_LOGIC;
  SIGNAL mux_1323_nl : STD_LOGIC;
  SIGNAL mux_1322_nl : STD_LOGIC;
  SIGNAL mux_1321_nl : STD_LOGIC;
  SIGNAL mux_1320_nl : STD_LOGIC;
  SIGNAL and_550_nl : STD_LOGIC;
  SIGNAL mux_1319_nl : STD_LOGIC;
  SIGNAL nor_1403_nl : STD_LOGIC;
  SIGNAL nor_1404_nl : STD_LOGIC;
  SIGNAL mux_1318_nl : STD_LOGIC;
  SIGNAL mux_1317_nl : STD_LOGIC;
  SIGNAL and_551_nl : STD_LOGIC;
  SIGNAL mux_1314_nl : STD_LOGIC;
  SIGNAL mux_1313_nl : STD_LOGIC;
  SIGNAL mux_1312_nl : STD_LOGIC;
  SIGNAL nor_1410_nl : STD_LOGIC;
  SIGNAL nor_1411_nl : STD_LOGIC;
  SIGNAL mux_1311_nl : STD_LOGIC;
  SIGNAL nor_1412_nl : STD_LOGIC;
  SIGNAL nor_1413_nl : STD_LOGIC;
  SIGNAL mux_1310_nl : STD_LOGIC;
  SIGNAL mux_1309_nl : STD_LOGIC;
  SIGNAL nor_1414_nl : STD_LOGIC;
  SIGNAL nor_1415_nl : STD_LOGIC;
  SIGNAL mux_1308_nl : STD_LOGIC;
  SIGNAL nor_1416_nl : STD_LOGIC;
  SIGNAL nor_1417_nl : STD_LOGIC;
  SIGNAL nor_1359_nl : STD_LOGIC;
  SIGNAL mux_1369_nl : STD_LOGIC;
  SIGNAL mux_1368_nl : STD_LOGIC;
  SIGNAL nor_1360_nl : STD_LOGIC;
  SIGNAL mux_1367_nl : STD_LOGIC;
  SIGNAL or_1151_nl : STD_LOGIC;
  SIGNAL mux_1364_nl : STD_LOGIC;
  SIGNAL mux_1363_nl : STD_LOGIC;
  SIGNAL or_1145_nl : STD_LOGIC;
  SIGNAL or_1143_nl : STD_LOGIC;
  SIGNAL mux_1362_nl : STD_LOGIC;
  SIGNAL or_1141_nl : STD_LOGIC;
  SIGNAL or_1140_nl : STD_LOGIC;
  SIGNAL mux_1361_nl : STD_LOGIC;
  SIGNAL mux_1360_nl : STD_LOGIC;
  SIGNAL mux_1359_nl : STD_LOGIC;
  SIGNAL nor_1361_nl : STD_LOGIC;
  SIGNAL nor_1362_nl : STD_LOGIC;
  SIGNAL mux_1358_nl : STD_LOGIC;
  SIGNAL nor_1363_nl : STD_LOGIC;
  SIGNAL nor_1364_nl : STD_LOGIC;
  SIGNAL mux_1357_nl : STD_LOGIC;
  SIGNAL mux_1356_nl : STD_LOGIC;
  SIGNAL nor_1365_nl : STD_LOGIC;
  SIGNAL nor_1366_nl : STD_LOGIC;
  SIGNAL mux_1355_nl : STD_LOGIC;
  SIGNAL nor_1367_nl : STD_LOGIC;
  SIGNAL nor_1368_nl : STD_LOGIC;
  SIGNAL mux_1354_nl : STD_LOGIC;
  SIGNAL mux_1353_nl : STD_LOGIC;
  SIGNAL mux_1352_nl : STD_LOGIC;
  SIGNAL mux_1351_nl : STD_LOGIC;
  SIGNAL nor_1369_nl : STD_LOGIC;
  SIGNAL nor_1370_nl : STD_LOGIC;
  SIGNAL mux_1350_nl : STD_LOGIC;
  SIGNAL nor_1371_nl : STD_LOGIC;
  SIGNAL nor_1372_nl : STD_LOGIC;
  SIGNAL mux_1349_nl : STD_LOGIC;
  SIGNAL mux_1348_nl : STD_LOGIC;
  SIGNAL nor_1373_nl : STD_LOGIC;
  SIGNAL nor_1374_nl : STD_LOGIC;
  SIGNAL mux_1347_nl : STD_LOGIC;
  SIGNAL nor_1375_nl : STD_LOGIC;
  SIGNAL nor_1376_nl : STD_LOGIC;
  SIGNAL mux_1346_nl : STD_LOGIC;
  SIGNAL mux_1345_nl : STD_LOGIC;
  SIGNAL mux_1344_nl : STD_LOGIC;
  SIGNAL nor_1377_nl : STD_LOGIC;
  SIGNAL nor_1378_nl : STD_LOGIC;
  SIGNAL mux_1343_nl : STD_LOGIC;
  SIGNAL nor_1379_nl : STD_LOGIC;
  SIGNAL nor_1380_nl : STD_LOGIC;
  SIGNAL mux_1342_nl : STD_LOGIC;
  SIGNAL mux_1341_nl : STD_LOGIC;
  SIGNAL nor_1381_nl : STD_LOGIC;
  SIGNAL nor_1382_nl : STD_LOGIC;
  SIGNAL mux_1340_nl : STD_LOGIC;
  SIGNAL nor_1383_nl : STD_LOGIC;
  SIGNAL nor_1384_nl : STD_LOGIC;
  SIGNAL mux_1400_nl : STD_LOGIC;
  SIGNAL mux_1399_nl : STD_LOGIC;
  SIGNAL mux_1398_nl : STD_LOGIC;
  SIGNAL nor_1332_nl : STD_LOGIC;
  SIGNAL mux_1397_nl : STD_LOGIC;
  SIGNAL mux_1396_nl : STD_LOGIC;
  SIGNAL nor_1333_nl : STD_LOGIC;
  SIGNAL nor_1334_nl : STD_LOGIC;
  SIGNAL nor_1335_nl : STD_LOGIC;
  SIGNAL mux_1395_nl : STD_LOGIC;
  SIGNAL mux_1394_nl : STD_LOGIC;
  SIGNAL mux_1393_nl : STD_LOGIC;
  SIGNAL nor_1336_nl : STD_LOGIC;
  SIGNAL nor_1337_nl : STD_LOGIC;
  SIGNAL nor_1338_nl : STD_LOGIC;
  SIGNAL nor_1339_nl : STD_LOGIC;
  SIGNAL mux_1392_nl : STD_LOGIC;
  SIGNAL mux_1391_nl : STD_LOGIC;
  SIGNAL mux_1390_nl : STD_LOGIC;
  SIGNAL nor_1340_nl : STD_LOGIC;
  SIGNAL mux_1389_nl : STD_LOGIC;
  SIGNAL nor_1341_nl : STD_LOGIC;
  SIGNAL nor_1342_nl : STD_LOGIC;
  SIGNAL nor_1343_nl : STD_LOGIC;
  SIGNAL mux_1388_nl : STD_LOGIC;
  SIGNAL nor_1344_nl : STD_LOGIC;
  SIGNAL mux_1387_nl : STD_LOGIC;
  SIGNAL mux_1386_nl : STD_LOGIC;
  SIGNAL nor_1345_nl : STD_LOGIC;
  SIGNAL nor_1346_nl : STD_LOGIC;
  SIGNAL nor_1347_nl : STD_LOGIC;
  SIGNAL mux_1385_nl : STD_LOGIC;
  SIGNAL mux_1384_nl : STD_LOGIC;
  SIGNAL mux_1383_nl : STD_LOGIC;
  SIGNAL and_546_nl : STD_LOGIC;
  SIGNAL mux_1382_nl : STD_LOGIC;
  SIGNAL nor_1348_nl : STD_LOGIC;
  SIGNAL nor_1349_nl : STD_LOGIC;
  SIGNAL nor_1350_nl : STD_LOGIC;
  SIGNAL mux_1381_nl : STD_LOGIC;
  SIGNAL or_1173_nl : STD_LOGIC;
  SIGNAL or_1171_nl : STD_LOGIC;
  SIGNAL mux_1380_nl : STD_LOGIC;
  SIGNAL nor_1351_nl : STD_LOGIC;
  SIGNAL mux_1379_nl : STD_LOGIC;
  SIGNAL or_1169_nl : STD_LOGIC;
  SIGNAL or_1167_nl : STD_LOGIC;
  SIGNAL and_547_nl : STD_LOGIC;
  SIGNAL mux_1377_nl : STD_LOGIC;
  SIGNAL nor_1354_nl : STD_LOGIC;
  SIGNAL mux_1376_nl : STD_LOGIC;
  SIGNAL mux_1375_nl : STD_LOGIC;
  SIGNAL or_1163_nl : STD_LOGIC;
  SIGNAL or_1161_nl : STD_LOGIC;
  SIGNAL mux_1374_nl : STD_LOGIC;
  SIGNAL or_1160_nl : STD_LOGIC;
  SIGNAL or_1158_nl : STD_LOGIC;
  SIGNAL and_548_nl : STD_LOGIC;
  SIGNAL mux_1373_nl : STD_LOGIC;
  SIGNAL mux_1372_nl : STD_LOGIC;
  SIGNAL nor_1355_nl : STD_LOGIC;
  SIGNAL nor_1356_nl : STD_LOGIC;
  SIGNAL mux_1371_nl : STD_LOGIC;
  SIGNAL nor_1357_nl : STD_LOGIC;
  SIGNAL nor_1358_nl : STD_LOGIC;
  SIGNAL nor_1302_nl : STD_LOGIC;
  SIGNAL mux_1431_nl : STD_LOGIC;
  SIGNAL mux_1430_nl : STD_LOGIC;
  SIGNAL and_545_nl : STD_LOGIC;
  SIGNAL mux_1429_nl : STD_LOGIC;
  SIGNAL nor_1303_nl : STD_LOGIC;
  SIGNAL mux_1426_nl : STD_LOGIC;
  SIGNAL mux_1425_nl : STD_LOGIC;
  SIGNAL nor_1304_nl : STD_LOGIC;
  SIGNAL nor_1305_nl : STD_LOGIC;
  SIGNAL mux_1424_nl : STD_LOGIC;
  SIGNAL nor_1306_nl : STD_LOGIC;
  SIGNAL nor_1307_nl : STD_LOGIC;
  SIGNAL mux_1423_nl : STD_LOGIC;
  SIGNAL mux_1422_nl : STD_LOGIC;
  SIGNAL mux_1421_nl : STD_LOGIC;
  SIGNAL nor_1308_nl : STD_LOGIC;
  SIGNAL nor_1309_nl : STD_LOGIC;
  SIGNAL mux_1420_nl : STD_LOGIC;
  SIGNAL nor_1310_nl : STD_LOGIC;
  SIGNAL nor_1311_nl : STD_LOGIC;
  SIGNAL mux_1419_nl : STD_LOGIC;
  SIGNAL mux_1418_nl : STD_LOGIC;
  SIGNAL nor_1312_nl : STD_LOGIC;
  SIGNAL nor_1313_nl : STD_LOGIC;
  SIGNAL mux_1417_nl : STD_LOGIC;
  SIGNAL nor_1314_nl : STD_LOGIC;
  SIGNAL nor_1315_nl : STD_LOGIC;
  SIGNAL mux_1416_nl : STD_LOGIC;
  SIGNAL mux_1415_nl : STD_LOGIC;
  SIGNAL mux_1414_nl : STD_LOGIC;
  SIGNAL mux_1413_nl : STD_LOGIC;
  SIGNAL nor_1316_nl : STD_LOGIC;
  SIGNAL mux_1412_nl : STD_LOGIC;
  SIGNAL nor_1319_nl : STD_LOGIC;
  SIGNAL mux_1411_nl : STD_LOGIC;
  SIGNAL mux_1410_nl : STD_LOGIC;
  SIGNAL nor_1320_nl : STD_LOGIC;
  SIGNAL mux_1409_nl : STD_LOGIC;
  SIGNAL nor_1323_nl : STD_LOGIC;
  SIGNAL mux_1408_nl : STD_LOGIC;
  SIGNAL mux_1407_nl : STD_LOGIC;
  SIGNAL mux_1406_nl : STD_LOGIC;
  SIGNAL nor_1324_nl : STD_LOGIC;
  SIGNAL nor_1325_nl : STD_LOGIC;
  SIGNAL mux_1405_nl : STD_LOGIC;
  SIGNAL nor_1326_nl : STD_LOGIC;
  SIGNAL nor_1327_nl : STD_LOGIC;
  SIGNAL mux_1404_nl : STD_LOGIC;
  SIGNAL mux_1403_nl : STD_LOGIC;
  SIGNAL nor_1328_nl : STD_LOGIC;
  SIGNAL nor_1329_nl : STD_LOGIC;
  SIGNAL mux_1402_nl : STD_LOGIC;
  SIGNAL nor_1330_nl : STD_LOGIC;
  SIGNAL nor_1331_nl : STD_LOGIC;
  SIGNAL mux_1463_nl : STD_LOGIC;
  SIGNAL mux_1462_nl : STD_LOGIC;
  SIGNAL mux_1461_nl : STD_LOGIC;
  SIGNAL mux_1460_nl : STD_LOGIC;
  SIGNAL nor_1269_nl : STD_LOGIC;
  SIGNAL nor_1270_nl : STD_LOGIC;
  SIGNAL mux_1459_nl : STD_LOGIC;
  SIGNAL nor_1271_nl : STD_LOGIC;
  SIGNAL nor_1272_nl : STD_LOGIC;
  SIGNAL mux_1458_nl : STD_LOGIC;
  SIGNAL mux_1457_nl : STD_LOGIC;
  SIGNAL nor_1273_nl : STD_LOGIC;
  SIGNAL nor_1274_nl : STD_LOGIC;
  SIGNAL nor_1275_nl : STD_LOGIC;
  SIGNAL mux_1456_nl : STD_LOGIC;
  SIGNAL mux_1455_nl : STD_LOGIC;
  SIGNAL mux_1454_nl : STD_LOGIC;
  SIGNAL nor_1276_nl : STD_LOGIC;
  SIGNAL nor_1277_nl : STD_LOGIC;
  SIGNAL mux_1453_nl : STD_LOGIC;
  SIGNAL nor_1278_nl : STD_LOGIC;
  SIGNAL nor_1279_nl : STD_LOGIC;
  SIGNAL mux_1452_nl : STD_LOGIC;
  SIGNAL mux_1451_nl : STD_LOGIC;
  SIGNAL nor_1280_nl : STD_LOGIC;
  SIGNAL nor_1281_nl : STD_LOGIC;
  SIGNAL mux_1450_nl : STD_LOGIC;
  SIGNAL mux_1449_nl : STD_LOGIC;
  SIGNAL nor_1282_nl : STD_LOGIC;
  SIGNAL nor_1283_nl : STD_LOGIC;
  SIGNAL nor_1284_nl : STD_LOGIC;
  SIGNAL and_542_nl : STD_LOGIC;
  SIGNAL mux_1448_nl : STD_LOGIC;
  SIGNAL mux_1447_nl : STD_LOGIC;
  SIGNAL mux_1446_nl : STD_LOGIC;
  SIGNAL mux_1445_nl : STD_LOGIC;
  SIGNAL and_543_nl : STD_LOGIC;
  SIGNAL mux_1444_nl : STD_LOGIC;
  SIGNAL nor_1287_nl : STD_LOGIC;
  SIGNAL nor_1288_nl : STD_LOGIC;
  SIGNAL mux_1443_nl : STD_LOGIC;
  SIGNAL mux_1442_nl : STD_LOGIC;
  SIGNAL and_544_nl : STD_LOGIC;
  SIGNAL mux_1439_nl : STD_LOGIC;
  SIGNAL mux_1438_nl : STD_LOGIC;
  SIGNAL mux_1437_nl : STD_LOGIC;
  SIGNAL nor_1294_nl : STD_LOGIC;
  SIGNAL nor_1295_nl : STD_LOGIC;
  SIGNAL mux_1436_nl : STD_LOGIC;
  SIGNAL nor_1296_nl : STD_LOGIC;
  SIGNAL nor_1297_nl : STD_LOGIC;
  SIGNAL mux_1435_nl : STD_LOGIC;
  SIGNAL mux_1434_nl : STD_LOGIC;
  SIGNAL nor_1298_nl : STD_LOGIC;
  SIGNAL nor_1299_nl : STD_LOGIC;
  SIGNAL mux_1433_nl : STD_LOGIC;
  SIGNAL nor_1300_nl : STD_LOGIC;
  SIGNAL nor_1301_nl : STD_LOGIC;
  SIGNAL nor_1240_nl : STD_LOGIC;
  SIGNAL mux_1494_nl : STD_LOGIC;
  SIGNAL mux_1493_nl : STD_LOGIC;
  SIGNAL nor_1241_nl : STD_LOGIC;
  SIGNAL mux_1492_nl : STD_LOGIC;
  SIGNAL nand_47_nl : STD_LOGIC;
  SIGNAL mux_1489_nl : STD_LOGIC;
  SIGNAL mux_1488_nl : STD_LOGIC;
  SIGNAL or_1340_nl : STD_LOGIC;
  SIGNAL or_1338_nl : STD_LOGIC;
  SIGNAL mux_1487_nl : STD_LOGIC;
  SIGNAL or_1336_nl : STD_LOGIC;
  SIGNAL or_1335_nl : STD_LOGIC;
  SIGNAL mux_1486_nl : STD_LOGIC;
  SIGNAL mux_1485_nl : STD_LOGIC;
  SIGNAL mux_1484_nl : STD_LOGIC;
  SIGNAL nor_1245_nl : STD_LOGIC;
  SIGNAL nor_1246_nl : STD_LOGIC;
  SIGNAL mux_1483_nl : STD_LOGIC;
  SIGNAL nor_1247_nl : STD_LOGIC;
  SIGNAL nor_1248_nl : STD_LOGIC;
  SIGNAL mux_1482_nl : STD_LOGIC;
  SIGNAL mux_1481_nl : STD_LOGIC;
  SIGNAL nor_1249_nl : STD_LOGIC;
  SIGNAL nor_1250_nl : STD_LOGIC;
  SIGNAL mux_1480_nl : STD_LOGIC;
  SIGNAL nor_1251_nl : STD_LOGIC;
  SIGNAL nor_1252_nl : STD_LOGIC;
  SIGNAL mux_1479_nl : STD_LOGIC;
  SIGNAL mux_1478_nl : STD_LOGIC;
  SIGNAL mux_1477_nl : STD_LOGIC;
  SIGNAL mux_1476_nl : STD_LOGIC;
  SIGNAL nor_1253_nl : STD_LOGIC;
  SIGNAL nor_1254_nl : STD_LOGIC;
  SIGNAL mux_1475_nl : STD_LOGIC;
  SIGNAL nor_1255_nl : STD_LOGIC;
  SIGNAL nor_1256_nl : STD_LOGIC;
  SIGNAL mux_1474_nl : STD_LOGIC;
  SIGNAL mux_1473_nl : STD_LOGIC;
  SIGNAL nor_1257_nl : STD_LOGIC;
  SIGNAL nor_1258_nl : STD_LOGIC;
  SIGNAL mux_1472_nl : STD_LOGIC;
  SIGNAL nor_1259_nl : STD_LOGIC;
  SIGNAL nor_1260_nl : STD_LOGIC;
  SIGNAL mux_1471_nl : STD_LOGIC;
  SIGNAL mux_1470_nl : STD_LOGIC;
  SIGNAL mux_1469_nl : STD_LOGIC;
  SIGNAL nor_1261_nl : STD_LOGIC;
  SIGNAL nor_1262_nl : STD_LOGIC;
  SIGNAL mux_1468_nl : STD_LOGIC;
  SIGNAL nor_1263_nl : STD_LOGIC;
  SIGNAL nor_1264_nl : STD_LOGIC;
  SIGNAL mux_1467_nl : STD_LOGIC;
  SIGNAL mux_1466_nl : STD_LOGIC;
  SIGNAL nor_1265_nl : STD_LOGIC;
  SIGNAL nor_1266_nl : STD_LOGIC;
  SIGNAL mux_1465_nl : STD_LOGIC;
  SIGNAL nor_1267_nl : STD_LOGIC;
  SIGNAL nor_1268_nl : STD_LOGIC;
  SIGNAL mux_1525_nl : STD_LOGIC;
  SIGNAL mux_1524_nl : STD_LOGIC;
  SIGNAL mux_1523_nl : STD_LOGIC;
  SIGNAL nor_1213_nl : STD_LOGIC;
  SIGNAL mux_1522_nl : STD_LOGIC;
  SIGNAL mux_1521_nl : STD_LOGIC;
  SIGNAL nor_1214_nl : STD_LOGIC;
  SIGNAL nor_1215_nl : STD_LOGIC;
  SIGNAL nor_1216_nl : STD_LOGIC;
  SIGNAL mux_1520_nl : STD_LOGIC;
  SIGNAL mux_1519_nl : STD_LOGIC;
  SIGNAL mux_1518_nl : STD_LOGIC;
  SIGNAL nor_1217_nl : STD_LOGIC;
  SIGNAL nor_1218_nl : STD_LOGIC;
  SIGNAL nor_1219_nl : STD_LOGIC;
  SIGNAL nor_1220_nl : STD_LOGIC;
  SIGNAL mux_1517_nl : STD_LOGIC;
  SIGNAL mux_1516_nl : STD_LOGIC;
  SIGNAL mux_1515_nl : STD_LOGIC;
  SIGNAL nor_1221_nl : STD_LOGIC;
  SIGNAL mux_1514_nl : STD_LOGIC;
  SIGNAL nor_1222_nl : STD_LOGIC;
  SIGNAL nor_1223_nl : STD_LOGIC;
  SIGNAL nor_1224_nl : STD_LOGIC;
  SIGNAL mux_1513_nl : STD_LOGIC;
  SIGNAL nor_1225_nl : STD_LOGIC;
  SIGNAL mux_1512_nl : STD_LOGIC;
  SIGNAL mux_1511_nl : STD_LOGIC;
  SIGNAL nor_1226_nl : STD_LOGIC;
  SIGNAL nor_1227_nl : STD_LOGIC;
  SIGNAL nor_1228_nl : STD_LOGIC;
  SIGNAL mux_1510_nl : STD_LOGIC;
  SIGNAL mux_1509_nl : STD_LOGIC;
  SIGNAL mux_1508_nl : STD_LOGIC;
  SIGNAL and_539_nl : STD_LOGIC;
  SIGNAL mux_1507_nl : STD_LOGIC;
  SIGNAL nor_1229_nl : STD_LOGIC;
  SIGNAL nor_1230_nl : STD_LOGIC;
  SIGNAL nor_1231_nl : STD_LOGIC;
  SIGNAL mux_1506_nl : STD_LOGIC;
  SIGNAL or_1367_nl : STD_LOGIC;
  SIGNAL or_1365_nl : STD_LOGIC;
  SIGNAL mux_1505_nl : STD_LOGIC;
  SIGNAL nor_1232_nl : STD_LOGIC;
  SIGNAL mux_1504_nl : STD_LOGIC;
  SIGNAL or_1363_nl : STD_LOGIC;
  SIGNAL or_1361_nl : STD_LOGIC;
  SIGNAL and_540_nl : STD_LOGIC;
  SIGNAL mux_1502_nl : STD_LOGIC;
  SIGNAL nor_1235_nl : STD_LOGIC;
  SIGNAL mux_1501_nl : STD_LOGIC;
  SIGNAL mux_1500_nl : STD_LOGIC;
  SIGNAL or_1357_nl : STD_LOGIC;
  SIGNAL or_1355_nl : STD_LOGIC;
  SIGNAL mux_1499_nl : STD_LOGIC;
  SIGNAL or_1354_nl : STD_LOGIC;
  SIGNAL or_1352_nl : STD_LOGIC;
  SIGNAL and_541_nl : STD_LOGIC;
  SIGNAL mux_1498_nl : STD_LOGIC;
  SIGNAL mux_1497_nl : STD_LOGIC;
  SIGNAL nor_1236_nl : STD_LOGIC;
  SIGNAL nor_1237_nl : STD_LOGIC;
  SIGNAL mux_1496_nl : STD_LOGIC;
  SIGNAL nor_1238_nl : STD_LOGIC;
  SIGNAL nor_1239_nl : STD_LOGIC;
  SIGNAL nor_1184_nl : STD_LOGIC;
  SIGNAL mux_1556_nl : STD_LOGIC;
  SIGNAL mux_1555_nl : STD_LOGIC;
  SIGNAL and_534_nl : STD_LOGIC;
  SIGNAL mux_1554_nl : STD_LOGIC;
  SIGNAL and_535_nl : STD_LOGIC;
  SIGNAL mux_1551_nl : STD_LOGIC;
  SIGNAL mux_1550_nl : STD_LOGIC;
  SIGNAL nor_1188_nl : STD_LOGIC;
  SIGNAL nor_1189_nl : STD_LOGIC;
  SIGNAL mux_1549_nl : STD_LOGIC;
  SIGNAL nor_1190_nl : STD_LOGIC;
  SIGNAL nor_1191_nl : STD_LOGIC;
  SIGNAL mux_1548_nl : STD_LOGIC;
  SIGNAL mux_1547_nl : STD_LOGIC;
  SIGNAL mux_1546_nl : STD_LOGIC;
  SIGNAL nor_1192_nl : STD_LOGIC;
  SIGNAL nor_1193_nl : STD_LOGIC;
  SIGNAL mux_1545_nl : STD_LOGIC;
  SIGNAL and_536_nl : STD_LOGIC;
  SIGNAL nor_1194_nl : STD_LOGIC;
  SIGNAL mux_1544_nl : STD_LOGIC;
  SIGNAL mux_1543_nl : STD_LOGIC;
  SIGNAL and_842_nl : STD_LOGIC;
  SIGNAL nor_1196_nl : STD_LOGIC;
  SIGNAL mux_1542_nl : STD_LOGIC;
  SIGNAL nor_1197_nl : STD_LOGIC;
  SIGNAL nor_1198_nl : STD_LOGIC;
  SIGNAL mux_1541_nl : STD_LOGIC;
  SIGNAL mux_1540_nl : STD_LOGIC;
  SIGNAL mux_1539_nl : STD_LOGIC;
  SIGNAL mux_1538_nl : STD_LOGIC;
  SIGNAL nor_1199_nl : STD_LOGIC;
  SIGNAL mux_1537_nl : STD_LOGIC;
  SIGNAL nor_1201_nl : STD_LOGIC;
  SIGNAL mux_1536_nl : STD_LOGIC;
  SIGNAL mux_1535_nl : STD_LOGIC;
  SIGNAL and_853_nl : STD_LOGIC;
  SIGNAL mux_1534_nl : STD_LOGIC;
  SIGNAL nor_1205_nl : STD_LOGIC;
  SIGNAL mux_1533_nl : STD_LOGIC;
  SIGNAL mux_1532_nl : STD_LOGIC;
  SIGNAL mux_1531_nl : STD_LOGIC;
  SIGNAL nor_1206_nl : STD_LOGIC;
  SIGNAL nor_1207_nl : STD_LOGIC;
  SIGNAL mux_1530_nl : STD_LOGIC;
  SIGNAL and_538_nl : STD_LOGIC;
  SIGNAL nor_1208_nl : STD_LOGIC;
  SIGNAL mux_1529_nl : STD_LOGIC;
  SIGNAL mux_1528_nl : STD_LOGIC;
  SIGNAL and_872_nl : STD_LOGIC;
  SIGNAL nor_1210_nl : STD_LOGIC;
  SIGNAL mux_1527_nl : STD_LOGIC;
  SIGNAL nor_1211_nl : STD_LOGIC;
  SIGNAL nor_1212_nl : STD_LOGIC;
  SIGNAL mux_1588_nl : STD_LOGIC;
  SIGNAL mux_1587_nl : STD_LOGIC;
  SIGNAL mux_1586_nl : STD_LOGIC;
  SIGNAL mux_1585_nl : STD_LOGIC;
  SIGNAL nor_1154_nl : STD_LOGIC;
  SIGNAL nor_1155_nl : STD_LOGIC;
  SIGNAL mux_1584_nl : STD_LOGIC;
  SIGNAL nor_1156_nl : STD_LOGIC;
  SIGNAL nor_1157_nl : STD_LOGIC;
  SIGNAL mux_1583_nl : STD_LOGIC;
  SIGNAL mux_1582_nl : STD_LOGIC;
  SIGNAL nor_1158_nl : STD_LOGIC;
  SIGNAL nor_1159_nl : STD_LOGIC;
  SIGNAL nor_1160_nl : STD_LOGIC;
  SIGNAL mux_1581_nl : STD_LOGIC;
  SIGNAL mux_1580_nl : STD_LOGIC;
  SIGNAL mux_1579_nl : STD_LOGIC;
  SIGNAL nor_1161_nl : STD_LOGIC;
  SIGNAL and_852_nl : STD_LOGIC;
  SIGNAL mux_1578_nl : STD_LOGIC;
  SIGNAL and_858_nl : STD_LOGIC;
  SIGNAL nor_1164_nl : STD_LOGIC;
  SIGNAL mux_1577_nl : STD_LOGIC;
  SIGNAL mux_1576_nl : STD_LOGIC;
  SIGNAL and_870_nl : STD_LOGIC;
  SIGNAL and_871_nl : STD_LOGIC;
  SIGNAL mux_1575_nl : STD_LOGIC;
  SIGNAL mux_1574_nl : STD_LOGIC;
  SIGNAL nor_1167_nl : STD_LOGIC;
  SIGNAL nor_1168_nl : STD_LOGIC;
  SIGNAL nor_1169_nl : STD_LOGIC;
  SIGNAL and_528_nl : STD_LOGIC;
  SIGNAL mux_1573_nl : STD_LOGIC;
  SIGNAL mux_1572_nl : STD_LOGIC;
  SIGNAL mux_1571_nl : STD_LOGIC;
  SIGNAL mux_1570_nl : STD_LOGIC;
  SIGNAL and_530_nl : STD_LOGIC;
  SIGNAL mux_1569_nl : STD_LOGIC;
  SIGNAL nor_1171_nl : STD_LOGIC;
  SIGNAL nor_1172_nl : STD_LOGIC;
  SIGNAL mux_1568_nl : STD_LOGIC;
  SIGNAL mux_1567_nl : STD_LOGIC;
  SIGNAL and_531_nl : STD_LOGIC;
  SIGNAL mux_1564_nl : STD_LOGIC;
  SIGNAL mux_1563_nl : STD_LOGIC;
  SIGNAL mux_1562_nl : STD_LOGIC;
  SIGNAL nor_1178_nl : STD_LOGIC;
  SIGNAL nor_1179_nl : STD_LOGIC;
  SIGNAL mux_1561_nl : STD_LOGIC;
  SIGNAL nor_1180_nl : STD_LOGIC;
  SIGNAL nor_1181_nl : STD_LOGIC;
  SIGNAL mux_1560_nl : STD_LOGIC;
  SIGNAL mux_1559_nl : STD_LOGIC;
  SIGNAL and_532_nl : STD_LOGIC;
  SIGNAL nor_1182_nl : STD_LOGIC;
  SIGNAL mux_1558_nl : STD_LOGIC;
  SIGNAL and_533_nl : STD_LOGIC;
  SIGNAL nor_1183_nl : STD_LOGIC;
  SIGNAL nor_1128_nl : STD_LOGIC;
  SIGNAL mux_1619_nl : STD_LOGIC;
  SIGNAL mux_1618_nl : STD_LOGIC;
  SIGNAL nor_1129_nl : STD_LOGIC;
  SIGNAL mux_1617_nl : STD_LOGIC;
  SIGNAL or_1539_nl : STD_LOGIC;
  SIGNAL mux_1614_nl : STD_LOGIC;
  SIGNAL mux_1613_nl : STD_LOGIC;
  SIGNAL or_1533_nl : STD_LOGIC;
  SIGNAL or_1531_nl : STD_LOGIC;
  SIGNAL mux_1612_nl : STD_LOGIC;
  SIGNAL or_1529_nl : STD_LOGIC;
  SIGNAL or_1528_nl : STD_LOGIC;
  SIGNAL mux_1611_nl : STD_LOGIC;
  SIGNAL mux_1610_nl : STD_LOGIC;
  SIGNAL mux_1609_nl : STD_LOGIC;
  SIGNAL nor_1130_nl : STD_LOGIC;
  SIGNAL nor_1131_nl : STD_LOGIC;
  SIGNAL mux_1608_nl : STD_LOGIC;
  SIGNAL nor_1132_nl : STD_LOGIC;
  SIGNAL nor_1133_nl : STD_LOGIC;
  SIGNAL mux_1607_nl : STD_LOGIC;
  SIGNAL mux_1606_nl : STD_LOGIC;
  SIGNAL nor_1134_nl : STD_LOGIC;
  SIGNAL nor_1135_nl : STD_LOGIC;
  SIGNAL mux_1605_nl : STD_LOGIC;
  SIGNAL nor_1136_nl : STD_LOGIC;
  SIGNAL nor_1137_nl : STD_LOGIC;
  SIGNAL mux_1604_nl : STD_LOGIC;
  SIGNAL mux_1603_nl : STD_LOGIC;
  SIGNAL mux_1602_nl : STD_LOGIC;
  SIGNAL mux_1601_nl : STD_LOGIC;
  SIGNAL nor_1138_nl : STD_LOGIC;
  SIGNAL nor_1139_nl : STD_LOGIC;
  SIGNAL mux_1600_nl : STD_LOGIC;
  SIGNAL nor_1140_nl : STD_LOGIC;
  SIGNAL nor_1141_nl : STD_LOGIC;
  SIGNAL mux_1599_nl : STD_LOGIC;
  SIGNAL mux_1598_nl : STD_LOGIC;
  SIGNAL nor_1142_nl : STD_LOGIC;
  SIGNAL nor_1143_nl : STD_LOGIC;
  SIGNAL mux_1597_nl : STD_LOGIC;
  SIGNAL nor_1144_nl : STD_LOGIC;
  SIGNAL nor_1145_nl : STD_LOGIC;
  SIGNAL mux_1596_nl : STD_LOGIC;
  SIGNAL mux_1595_nl : STD_LOGIC;
  SIGNAL mux_1594_nl : STD_LOGIC;
  SIGNAL nor_1146_nl : STD_LOGIC;
  SIGNAL nor_1147_nl : STD_LOGIC;
  SIGNAL mux_1593_nl : STD_LOGIC;
  SIGNAL nor_1148_nl : STD_LOGIC;
  SIGNAL nor_1149_nl : STD_LOGIC;
  SIGNAL mux_1592_nl : STD_LOGIC;
  SIGNAL mux_1591_nl : STD_LOGIC;
  SIGNAL nor_1150_nl : STD_LOGIC;
  SIGNAL nor_1151_nl : STD_LOGIC;
  SIGNAL mux_1590_nl : STD_LOGIC;
  SIGNAL nor_1152_nl : STD_LOGIC;
  SIGNAL nor_1153_nl : STD_LOGIC;
  SIGNAL mux_1650_nl : STD_LOGIC;
  SIGNAL mux_1649_nl : STD_LOGIC;
  SIGNAL mux_1648_nl : STD_LOGIC;
  SIGNAL nor_1101_nl : STD_LOGIC;
  SIGNAL mux_1647_nl : STD_LOGIC;
  SIGNAL mux_1646_nl : STD_LOGIC;
  SIGNAL nor_1102_nl : STD_LOGIC;
  SIGNAL nor_1103_nl : STD_LOGIC;
  SIGNAL nor_1104_nl : STD_LOGIC;
  SIGNAL mux_1645_nl : STD_LOGIC;
  SIGNAL mux_1644_nl : STD_LOGIC;
  SIGNAL mux_1643_nl : STD_LOGIC;
  SIGNAL nor_1105_nl : STD_LOGIC;
  SIGNAL nor_1106_nl : STD_LOGIC;
  SIGNAL nor_1107_nl : STD_LOGIC;
  SIGNAL nor_1108_nl : STD_LOGIC;
  SIGNAL mux_1642_nl : STD_LOGIC;
  SIGNAL mux_1641_nl : STD_LOGIC;
  SIGNAL mux_1640_nl : STD_LOGIC;
  SIGNAL nor_1109_nl : STD_LOGIC;
  SIGNAL mux_1639_nl : STD_LOGIC;
  SIGNAL nor_1110_nl : STD_LOGIC;
  SIGNAL nor_1111_nl : STD_LOGIC;
  SIGNAL nor_1112_nl : STD_LOGIC;
  SIGNAL mux_1638_nl : STD_LOGIC;
  SIGNAL nor_1113_nl : STD_LOGIC;
  SIGNAL mux_1637_nl : STD_LOGIC;
  SIGNAL mux_1636_nl : STD_LOGIC;
  SIGNAL nor_1114_nl : STD_LOGIC;
  SIGNAL nor_1115_nl : STD_LOGIC;
  SIGNAL nor_1116_nl : STD_LOGIC;
  SIGNAL mux_1635_nl : STD_LOGIC;
  SIGNAL mux_1634_nl : STD_LOGIC;
  SIGNAL mux_1633_nl : STD_LOGIC;
  SIGNAL and_525_nl : STD_LOGIC;
  SIGNAL mux_1632_nl : STD_LOGIC;
  SIGNAL nor_1117_nl : STD_LOGIC;
  SIGNAL nor_1118_nl : STD_LOGIC;
  SIGNAL nor_1119_nl : STD_LOGIC;
  SIGNAL mux_1631_nl : STD_LOGIC;
  SIGNAL or_1561_nl : STD_LOGIC;
  SIGNAL or_1559_nl : STD_LOGIC;
  SIGNAL mux_1630_nl : STD_LOGIC;
  SIGNAL nor_1120_nl : STD_LOGIC;
  SIGNAL mux_1629_nl : STD_LOGIC;
  SIGNAL or_1557_nl : STD_LOGIC;
  SIGNAL or_1555_nl : STD_LOGIC;
  SIGNAL and_526_nl : STD_LOGIC;
  SIGNAL mux_1627_nl : STD_LOGIC;
  SIGNAL nor_1123_nl : STD_LOGIC;
  SIGNAL mux_1626_nl : STD_LOGIC;
  SIGNAL mux_1625_nl : STD_LOGIC;
  SIGNAL or_1551_nl : STD_LOGIC;
  SIGNAL or_1549_nl : STD_LOGIC;
  SIGNAL mux_1624_nl : STD_LOGIC;
  SIGNAL or_1548_nl : STD_LOGIC;
  SIGNAL or_1546_nl : STD_LOGIC;
  SIGNAL and_527_nl : STD_LOGIC;
  SIGNAL mux_1623_nl : STD_LOGIC;
  SIGNAL mux_1622_nl : STD_LOGIC;
  SIGNAL nor_1124_nl : STD_LOGIC;
  SIGNAL nor_1125_nl : STD_LOGIC;
  SIGNAL mux_1621_nl : STD_LOGIC;
  SIGNAL nor_1126_nl : STD_LOGIC;
  SIGNAL nor_1127_nl : STD_LOGIC;
  SIGNAL nor_1071_nl : STD_LOGIC;
  SIGNAL mux_1681_nl : STD_LOGIC;
  SIGNAL mux_1680_nl : STD_LOGIC;
  SIGNAL and_524_nl : STD_LOGIC;
  SIGNAL mux_1679_nl : STD_LOGIC;
  SIGNAL nor_1072_nl : STD_LOGIC;
  SIGNAL mux_1676_nl : STD_LOGIC;
  SIGNAL mux_1675_nl : STD_LOGIC;
  SIGNAL nor_1073_nl : STD_LOGIC;
  SIGNAL nor_1074_nl : STD_LOGIC;
  SIGNAL mux_1674_nl : STD_LOGIC;
  SIGNAL nor_1075_nl : STD_LOGIC;
  SIGNAL nor_1076_nl : STD_LOGIC;
  SIGNAL mux_1673_nl : STD_LOGIC;
  SIGNAL mux_1672_nl : STD_LOGIC;
  SIGNAL mux_1671_nl : STD_LOGIC;
  SIGNAL nor_1077_nl : STD_LOGIC;
  SIGNAL nor_1078_nl : STD_LOGIC;
  SIGNAL mux_1670_nl : STD_LOGIC;
  SIGNAL nor_1079_nl : STD_LOGIC;
  SIGNAL nor_1080_nl : STD_LOGIC;
  SIGNAL mux_1669_nl : STD_LOGIC;
  SIGNAL mux_1668_nl : STD_LOGIC;
  SIGNAL nor_1081_nl : STD_LOGIC;
  SIGNAL nor_1082_nl : STD_LOGIC;
  SIGNAL mux_1667_nl : STD_LOGIC;
  SIGNAL nor_1083_nl : STD_LOGIC;
  SIGNAL nor_1084_nl : STD_LOGIC;
  SIGNAL mux_1666_nl : STD_LOGIC;
  SIGNAL mux_1665_nl : STD_LOGIC;
  SIGNAL mux_1664_nl : STD_LOGIC;
  SIGNAL mux_1663_nl : STD_LOGIC;
  SIGNAL nor_1085_nl : STD_LOGIC;
  SIGNAL mux_1662_nl : STD_LOGIC;
  SIGNAL nor_1088_nl : STD_LOGIC;
  SIGNAL mux_1661_nl : STD_LOGIC;
  SIGNAL mux_1660_nl : STD_LOGIC;
  SIGNAL nor_1089_nl : STD_LOGIC;
  SIGNAL mux_1659_nl : STD_LOGIC;
  SIGNAL nor_1092_nl : STD_LOGIC;
  SIGNAL mux_1658_nl : STD_LOGIC;
  SIGNAL mux_1657_nl : STD_LOGIC;
  SIGNAL mux_1656_nl : STD_LOGIC;
  SIGNAL nor_1093_nl : STD_LOGIC;
  SIGNAL nor_1094_nl : STD_LOGIC;
  SIGNAL mux_1655_nl : STD_LOGIC;
  SIGNAL nor_1095_nl : STD_LOGIC;
  SIGNAL nor_1096_nl : STD_LOGIC;
  SIGNAL mux_1654_nl : STD_LOGIC;
  SIGNAL mux_1653_nl : STD_LOGIC;
  SIGNAL nor_1097_nl : STD_LOGIC;
  SIGNAL nor_1098_nl : STD_LOGIC;
  SIGNAL mux_1652_nl : STD_LOGIC;
  SIGNAL nor_1099_nl : STD_LOGIC;
  SIGNAL nor_1100_nl : STD_LOGIC;
  SIGNAL mux_1713_nl : STD_LOGIC;
  SIGNAL mux_1712_nl : STD_LOGIC;
  SIGNAL mux_1711_nl : STD_LOGIC;
  SIGNAL mux_1710_nl : STD_LOGIC;
  SIGNAL nor_1039_nl : STD_LOGIC;
  SIGNAL nor_1040_nl : STD_LOGIC;
  SIGNAL mux_1709_nl : STD_LOGIC;
  SIGNAL nor_1041_nl : STD_LOGIC;
  SIGNAL nor_1042_nl : STD_LOGIC;
  SIGNAL mux_1708_nl : STD_LOGIC;
  SIGNAL mux_1707_nl : STD_LOGIC;
  SIGNAL nor_1043_nl : STD_LOGIC;
  SIGNAL nor_1044_nl : STD_LOGIC;
  SIGNAL nor_1045_nl : STD_LOGIC;
  SIGNAL mux_1706_nl : STD_LOGIC;
  SIGNAL mux_1705_nl : STD_LOGIC;
  SIGNAL mux_1704_nl : STD_LOGIC;
  SIGNAL nor_1046_nl : STD_LOGIC;
  SIGNAL nor_1047_nl : STD_LOGIC;
  SIGNAL mux_1703_nl : STD_LOGIC;
  SIGNAL nor_1048_nl : STD_LOGIC;
  SIGNAL nor_1049_nl : STD_LOGIC;
  SIGNAL mux_1702_nl : STD_LOGIC;
  SIGNAL mux_1701_nl : STD_LOGIC;
  SIGNAL nor_1050_nl : STD_LOGIC;
  SIGNAL nor_1051_nl : STD_LOGIC;
  SIGNAL mux_1700_nl : STD_LOGIC;
  SIGNAL mux_1699_nl : STD_LOGIC;
  SIGNAL nor_1052_nl : STD_LOGIC;
  SIGNAL nor_1053_nl : STD_LOGIC;
  SIGNAL nor_1054_nl : STD_LOGIC;
  SIGNAL and_520_nl : STD_LOGIC;
  SIGNAL mux_1698_nl : STD_LOGIC;
  SIGNAL mux_1697_nl : STD_LOGIC;
  SIGNAL mux_1696_nl : STD_LOGIC;
  SIGNAL mux_1695_nl : STD_LOGIC;
  SIGNAL and_521_nl : STD_LOGIC;
  SIGNAL mux_1694_nl : STD_LOGIC;
  SIGNAL nor_1057_nl : STD_LOGIC;
  SIGNAL nor_1058_nl : STD_LOGIC;
  SIGNAL mux_1693_nl : STD_LOGIC;
  SIGNAL mux_1692_nl : STD_LOGIC;
  SIGNAL and_522_nl : STD_LOGIC;
  SIGNAL mux_1689_nl : STD_LOGIC;
  SIGNAL mux_1688_nl : STD_LOGIC;
  SIGNAL mux_1687_nl : STD_LOGIC;
  SIGNAL nor_1063_nl : STD_LOGIC;
  SIGNAL nor_1064_nl : STD_LOGIC;
  SIGNAL mux_1686_nl : STD_LOGIC;
  SIGNAL nor_1065_nl : STD_LOGIC;
  SIGNAL nor_1066_nl : STD_LOGIC;
  SIGNAL mux_1685_nl : STD_LOGIC;
  SIGNAL mux_1684_nl : STD_LOGIC;
  SIGNAL nor_1067_nl : STD_LOGIC;
  SIGNAL nor_1068_nl : STD_LOGIC;
  SIGNAL mux_1683_nl : STD_LOGIC;
  SIGNAL nor_1069_nl : STD_LOGIC;
  SIGNAL nor_1070_nl : STD_LOGIC;
  SIGNAL nor_1010_nl : STD_LOGIC;
  SIGNAL mux_1744_nl : STD_LOGIC;
  SIGNAL mux_1743_nl : STD_LOGIC;
  SIGNAL nor_1011_nl : STD_LOGIC;
  SIGNAL mux_1742_nl : STD_LOGIC;
  SIGNAL nand_63_nl : STD_LOGIC;
  SIGNAL mux_1739_nl : STD_LOGIC;
  SIGNAL mux_1738_nl : STD_LOGIC;
  SIGNAL or_1728_nl : STD_LOGIC;
  SIGNAL or_1726_nl : STD_LOGIC;
  SIGNAL mux_1737_nl : STD_LOGIC;
  SIGNAL or_1724_nl : STD_LOGIC;
  SIGNAL or_1723_nl : STD_LOGIC;
  SIGNAL mux_1736_nl : STD_LOGIC;
  SIGNAL mux_1735_nl : STD_LOGIC;
  SIGNAL mux_1734_nl : STD_LOGIC;
  SIGNAL nor_1015_nl : STD_LOGIC;
  SIGNAL nor_1016_nl : STD_LOGIC;
  SIGNAL mux_1733_nl : STD_LOGIC;
  SIGNAL nor_1017_nl : STD_LOGIC;
  SIGNAL nor_1018_nl : STD_LOGIC;
  SIGNAL mux_1732_nl : STD_LOGIC;
  SIGNAL mux_1731_nl : STD_LOGIC;
  SIGNAL nor_1019_nl : STD_LOGIC;
  SIGNAL nor_1020_nl : STD_LOGIC;
  SIGNAL mux_1730_nl : STD_LOGIC;
  SIGNAL nor_1021_nl : STD_LOGIC;
  SIGNAL nor_1022_nl : STD_LOGIC;
  SIGNAL mux_1729_nl : STD_LOGIC;
  SIGNAL mux_1728_nl : STD_LOGIC;
  SIGNAL mux_1727_nl : STD_LOGIC;
  SIGNAL mux_1726_nl : STD_LOGIC;
  SIGNAL nor_1023_nl : STD_LOGIC;
  SIGNAL nor_1024_nl : STD_LOGIC;
  SIGNAL mux_1725_nl : STD_LOGIC;
  SIGNAL nor_1025_nl : STD_LOGIC;
  SIGNAL nor_1026_nl : STD_LOGIC;
  SIGNAL mux_1724_nl : STD_LOGIC;
  SIGNAL mux_1723_nl : STD_LOGIC;
  SIGNAL nor_1027_nl : STD_LOGIC;
  SIGNAL nor_1028_nl : STD_LOGIC;
  SIGNAL mux_1722_nl : STD_LOGIC;
  SIGNAL nor_1029_nl : STD_LOGIC;
  SIGNAL nor_1030_nl : STD_LOGIC;
  SIGNAL mux_1721_nl : STD_LOGIC;
  SIGNAL mux_1720_nl : STD_LOGIC;
  SIGNAL mux_1719_nl : STD_LOGIC;
  SIGNAL nor_1031_nl : STD_LOGIC;
  SIGNAL nor_1032_nl : STD_LOGIC;
  SIGNAL mux_1718_nl : STD_LOGIC;
  SIGNAL nor_1033_nl : STD_LOGIC;
  SIGNAL nor_1034_nl : STD_LOGIC;
  SIGNAL mux_1717_nl : STD_LOGIC;
  SIGNAL mux_1716_nl : STD_LOGIC;
  SIGNAL nor_1035_nl : STD_LOGIC;
  SIGNAL nor_1036_nl : STD_LOGIC;
  SIGNAL mux_1715_nl : STD_LOGIC;
  SIGNAL nor_1037_nl : STD_LOGIC;
  SIGNAL nor_1038_nl : STD_LOGIC;
  SIGNAL mux_1775_nl : STD_LOGIC;
  SIGNAL mux_1774_nl : STD_LOGIC;
  SIGNAL mux_1773_nl : STD_LOGIC;
  SIGNAL nor_983_nl : STD_LOGIC;
  SIGNAL mux_1772_nl : STD_LOGIC;
  SIGNAL mux_1771_nl : STD_LOGIC;
  SIGNAL nor_984_nl : STD_LOGIC;
  SIGNAL nor_985_nl : STD_LOGIC;
  SIGNAL nor_986_nl : STD_LOGIC;
  SIGNAL mux_1770_nl : STD_LOGIC;
  SIGNAL mux_1769_nl : STD_LOGIC;
  SIGNAL mux_1768_nl : STD_LOGIC;
  SIGNAL nor_987_nl : STD_LOGIC;
  SIGNAL nor_988_nl : STD_LOGIC;
  SIGNAL nor_989_nl : STD_LOGIC;
  SIGNAL nor_990_nl : STD_LOGIC;
  SIGNAL mux_1767_nl : STD_LOGIC;
  SIGNAL mux_1766_nl : STD_LOGIC;
  SIGNAL mux_1765_nl : STD_LOGIC;
  SIGNAL nor_991_nl : STD_LOGIC;
  SIGNAL mux_1764_nl : STD_LOGIC;
  SIGNAL nor_992_nl : STD_LOGIC;
  SIGNAL nor_993_nl : STD_LOGIC;
  SIGNAL nor_994_nl : STD_LOGIC;
  SIGNAL mux_1763_nl : STD_LOGIC;
  SIGNAL nor_995_nl : STD_LOGIC;
  SIGNAL mux_1762_nl : STD_LOGIC;
  SIGNAL mux_1761_nl : STD_LOGIC;
  SIGNAL nor_996_nl : STD_LOGIC;
  SIGNAL nor_997_nl : STD_LOGIC;
  SIGNAL nor_998_nl : STD_LOGIC;
  SIGNAL mux_1760_nl : STD_LOGIC;
  SIGNAL mux_1759_nl : STD_LOGIC;
  SIGNAL mux_1758_nl : STD_LOGIC;
  SIGNAL and_517_nl : STD_LOGIC;
  SIGNAL mux_1757_nl : STD_LOGIC;
  SIGNAL nor_999_nl : STD_LOGIC;
  SIGNAL nor_1000_nl : STD_LOGIC;
  SIGNAL nor_1001_nl : STD_LOGIC;
  SIGNAL mux_1756_nl : STD_LOGIC;
  SIGNAL or_1755_nl : STD_LOGIC;
  SIGNAL or_1753_nl : STD_LOGIC;
  SIGNAL mux_1755_nl : STD_LOGIC;
  SIGNAL nor_1002_nl : STD_LOGIC;
  SIGNAL mux_1754_nl : STD_LOGIC;
  SIGNAL or_1751_nl : STD_LOGIC;
  SIGNAL or_1749_nl : STD_LOGIC;
  SIGNAL and_518_nl : STD_LOGIC;
  SIGNAL mux_1752_nl : STD_LOGIC;
  SIGNAL nor_1005_nl : STD_LOGIC;
  SIGNAL mux_1751_nl : STD_LOGIC;
  SIGNAL mux_1750_nl : STD_LOGIC;
  SIGNAL or_1745_nl : STD_LOGIC;
  SIGNAL or_1743_nl : STD_LOGIC;
  SIGNAL mux_1749_nl : STD_LOGIC;
  SIGNAL or_1742_nl : STD_LOGIC;
  SIGNAL or_1740_nl : STD_LOGIC;
  SIGNAL and_519_nl : STD_LOGIC;
  SIGNAL mux_1748_nl : STD_LOGIC;
  SIGNAL mux_1747_nl : STD_LOGIC;
  SIGNAL nor_1006_nl : STD_LOGIC;
  SIGNAL nor_1007_nl : STD_LOGIC;
  SIGNAL mux_1746_nl : STD_LOGIC;
  SIGNAL nor_1008_nl : STD_LOGIC;
  SIGNAL nor_1009_nl : STD_LOGIC;
  SIGNAL nor_954_nl : STD_LOGIC;
  SIGNAL mux_1806_nl : STD_LOGIC;
  SIGNAL mux_1805_nl : STD_LOGIC;
  SIGNAL and_512_nl : STD_LOGIC;
  SIGNAL mux_1804_nl : STD_LOGIC;
  SIGNAL and_513_nl : STD_LOGIC;
  SIGNAL mux_1801_nl : STD_LOGIC;
  SIGNAL mux_1800_nl : STD_LOGIC;
  SIGNAL nor_958_nl : STD_LOGIC;
  SIGNAL nor_959_nl : STD_LOGIC;
  SIGNAL mux_1799_nl : STD_LOGIC;
  SIGNAL nor_960_nl : STD_LOGIC;
  SIGNAL nor_961_nl : STD_LOGIC;
  SIGNAL mux_1798_nl : STD_LOGIC;
  SIGNAL mux_1797_nl : STD_LOGIC;
  SIGNAL mux_1796_nl : STD_LOGIC;
  SIGNAL nor_962_nl : STD_LOGIC;
  SIGNAL nor_963_nl : STD_LOGIC;
  SIGNAL mux_1795_nl : STD_LOGIC;
  SIGNAL and_514_nl : STD_LOGIC;
  SIGNAL nor_964_nl : STD_LOGIC;
  SIGNAL mux_1794_nl : STD_LOGIC;
  SIGNAL mux_1793_nl : STD_LOGIC;
  SIGNAL and_841_nl : STD_LOGIC;
  SIGNAL nor_966_nl : STD_LOGIC;
  SIGNAL mux_1792_nl : STD_LOGIC;
  SIGNAL nor_967_nl : STD_LOGIC;
  SIGNAL nor_968_nl : STD_LOGIC;
  SIGNAL mux_1791_nl : STD_LOGIC;
  SIGNAL mux_1790_nl : STD_LOGIC;
  SIGNAL mux_1789_nl : STD_LOGIC;
  SIGNAL mux_1788_nl : STD_LOGIC;
  SIGNAL nor_969_nl : STD_LOGIC;
  SIGNAL mux_1787_nl : STD_LOGIC;
  SIGNAL nor_971_nl : STD_LOGIC;
  SIGNAL mux_1786_nl : STD_LOGIC;
  SIGNAL mux_1785_nl : STD_LOGIC;
  SIGNAL and_851_nl : STD_LOGIC;
  SIGNAL mux_1784_nl : STD_LOGIC;
  SIGNAL nor_975_nl : STD_LOGIC;
  SIGNAL mux_1783_nl : STD_LOGIC;
  SIGNAL mux_1782_nl : STD_LOGIC;
  SIGNAL mux_1781_nl : STD_LOGIC;
  SIGNAL nor_976_nl : STD_LOGIC;
  SIGNAL nor_977_nl : STD_LOGIC;
  SIGNAL mux_1780_nl : STD_LOGIC;
  SIGNAL and_516_nl : STD_LOGIC;
  SIGNAL nor_978_nl : STD_LOGIC;
  SIGNAL mux_1779_nl : STD_LOGIC;
  SIGNAL mux_1778_nl : STD_LOGIC;
  SIGNAL and_869_nl : STD_LOGIC;
  SIGNAL nor_980_nl : STD_LOGIC;
  SIGNAL mux_1777_nl : STD_LOGIC;
  SIGNAL nor_981_nl : STD_LOGIC;
  SIGNAL nor_982_nl : STD_LOGIC;
  SIGNAL mux_1838_nl : STD_LOGIC;
  SIGNAL mux_1837_nl : STD_LOGIC;
  SIGNAL mux_1836_nl : STD_LOGIC;
  SIGNAL mux_1835_nl : STD_LOGIC;
  SIGNAL nor_925_nl : STD_LOGIC;
  SIGNAL nor_926_nl : STD_LOGIC;
  SIGNAL mux_1834_nl : STD_LOGIC;
  SIGNAL nor_927_nl : STD_LOGIC;
  SIGNAL nor_928_nl : STD_LOGIC;
  SIGNAL mux_1833_nl : STD_LOGIC;
  SIGNAL mux_1832_nl : STD_LOGIC;
  SIGNAL nor_929_nl : STD_LOGIC;
  SIGNAL nor_930_nl : STD_LOGIC;
  SIGNAL nor_931_nl : STD_LOGIC;
  SIGNAL mux_1831_nl : STD_LOGIC;
  SIGNAL mux_1830_nl : STD_LOGIC;
  SIGNAL mux_1829_nl : STD_LOGIC;
  SIGNAL nor_932_nl : STD_LOGIC;
  SIGNAL and_850_nl : STD_LOGIC;
  SIGNAL mux_1828_nl : STD_LOGIC;
  SIGNAL and_857_nl : STD_LOGIC;
  SIGNAL nor_935_nl : STD_LOGIC;
  SIGNAL mux_1827_nl : STD_LOGIC;
  SIGNAL mux_1826_nl : STD_LOGIC;
  SIGNAL and_867_nl : STD_LOGIC;
  SIGNAL and_868_nl : STD_LOGIC;
  SIGNAL mux_1825_nl : STD_LOGIC;
  SIGNAL mux_1824_nl : STD_LOGIC;
  SIGNAL nor_938_nl : STD_LOGIC;
  SIGNAL nor_939_nl : STD_LOGIC;
  SIGNAL nor_940_nl : STD_LOGIC;
  SIGNAL and_505_nl : STD_LOGIC;
  SIGNAL mux_1823_nl : STD_LOGIC;
  SIGNAL mux_1822_nl : STD_LOGIC;
  SIGNAL mux_1821_nl : STD_LOGIC;
  SIGNAL mux_1820_nl : STD_LOGIC;
  SIGNAL and_507_nl : STD_LOGIC;
  SIGNAL mux_1819_nl : STD_LOGIC;
  SIGNAL nor_942_nl : STD_LOGIC;
  SIGNAL nor_943_nl : STD_LOGIC;
  SIGNAL mux_1818_nl : STD_LOGIC;
  SIGNAL mux_1817_nl : STD_LOGIC;
  SIGNAL and_508_nl : STD_LOGIC;
  SIGNAL mux_1814_nl : STD_LOGIC;
  SIGNAL mux_1813_nl : STD_LOGIC;
  SIGNAL mux_1812_nl : STD_LOGIC;
  SIGNAL nor_948_nl : STD_LOGIC;
  SIGNAL nor_949_nl : STD_LOGIC;
  SIGNAL mux_1811_nl : STD_LOGIC;
  SIGNAL nor_950_nl : STD_LOGIC;
  SIGNAL nor_951_nl : STD_LOGIC;
  SIGNAL mux_1810_nl : STD_LOGIC;
  SIGNAL mux_1809_nl : STD_LOGIC;
  SIGNAL and_510_nl : STD_LOGIC;
  SIGNAL nor_952_nl : STD_LOGIC;
  SIGNAL mux_1808_nl : STD_LOGIC;
  SIGNAL and_511_nl : STD_LOGIC;
  SIGNAL nor_953_nl : STD_LOGIC;
  SIGNAL nor_899_nl : STD_LOGIC;
  SIGNAL mux_1869_nl : STD_LOGIC;
  SIGNAL mux_1868_nl : STD_LOGIC;
  SIGNAL nor_900_nl : STD_LOGIC;
  SIGNAL mux_1867_nl : STD_LOGIC;
  SIGNAL or_1925_nl : STD_LOGIC;
  SIGNAL mux_1864_nl : STD_LOGIC;
  SIGNAL mux_1863_nl : STD_LOGIC;
  SIGNAL or_1919_nl : STD_LOGIC;
  SIGNAL or_1918_nl : STD_LOGIC;
  SIGNAL mux_1862_nl : STD_LOGIC;
  SIGNAL or_1916_nl : STD_LOGIC;
  SIGNAL or_1915_nl : STD_LOGIC;
  SIGNAL mux_1861_nl : STD_LOGIC;
  SIGNAL mux_1860_nl : STD_LOGIC;
  SIGNAL mux_1859_nl : STD_LOGIC;
  SIGNAL nor_901_nl : STD_LOGIC;
  SIGNAL nor_902_nl : STD_LOGIC;
  SIGNAL mux_1858_nl : STD_LOGIC;
  SIGNAL nor_903_nl : STD_LOGIC;
  SIGNAL nor_904_nl : STD_LOGIC;
  SIGNAL mux_1857_nl : STD_LOGIC;
  SIGNAL mux_1856_nl : STD_LOGIC;
  SIGNAL nor_905_nl : STD_LOGIC;
  SIGNAL nor_906_nl : STD_LOGIC;
  SIGNAL mux_1855_nl : STD_LOGIC;
  SIGNAL nor_907_nl : STD_LOGIC;
  SIGNAL nor_908_nl : STD_LOGIC;
  SIGNAL mux_1854_nl : STD_LOGIC;
  SIGNAL mux_1853_nl : STD_LOGIC;
  SIGNAL mux_1852_nl : STD_LOGIC;
  SIGNAL mux_1851_nl : STD_LOGIC;
  SIGNAL nor_909_nl : STD_LOGIC;
  SIGNAL nor_910_nl : STD_LOGIC;
  SIGNAL mux_1850_nl : STD_LOGIC;
  SIGNAL nor_911_nl : STD_LOGIC;
  SIGNAL nor_912_nl : STD_LOGIC;
  SIGNAL mux_1849_nl : STD_LOGIC;
  SIGNAL mux_1848_nl : STD_LOGIC;
  SIGNAL nor_913_nl : STD_LOGIC;
  SIGNAL nor_914_nl : STD_LOGIC;
  SIGNAL mux_1847_nl : STD_LOGIC;
  SIGNAL nor_915_nl : STD_LOGIC;
  SIGNAL nor_916_nl : STD_LOGIC;
  SIGNAL mux_1846_nl : STD_LOGIC;
  SIGNAL mux_1845_nl : STD_LOGIC;
  SIGNAL mux_1844_nl : STD_LOGIC;
  SIGNAL nor_917_nl : STD_LOGIC;
  SIGNAL nor_918_nl : STD_LOGIC;
  SIGNAL mux_1843_nl : STD_LOGIC;
  SIGNAL nor_919_nl : STD_LOGIC;
  SIGNAL nor_920_nl : STD_LOGIC;
  SIGNAL mux_1842_nl : STD_LOGIC;
  SIGNAL mux_1841_nl : STD_LOGIC;
  SIGNAL nor_921_nl : STD_LOGIC;
  SIGNAL nor_922_nl : STD_LOGIC;
  SIGNAL mux_1840_nl : STD_LOGIC;
  SIGNAL nor_923_nl : STD_LOGIC;
  SIGNAL nor_924_nl : STD_LOGIC;
  SIGNAL mux_1900_nl : STD_LOGIC;
  SIGNAL mux_1899_nl : STD_LOGIC;
  SIGNAL mux_1898_nl : STD_LOGIC;
  SIGNAL nor_873_nl : STD_LOGIC;
  SIGNAL mux_1897_nl : STD_LOGIC;
  SIGNAL mux_1896_nl : STD_LOGIC;
  SIGNAL nor_874_nl : STD_LOGIC;
  SIGNAL nor_875_nl : STD_LOGIC;
  SIGNAL nor_876_nl : STD_LOGIC;
  SIGNAL mux_1895_nl : STD_LOGIC;
  SIGNAL mux_1894_nl : STD_LOGIC;
  SIGNAL mux_1893_nl : STD_LOGIC;
  SIGNAL nor_877_nl : STD_LOGIC;
  SIGNAL nor_878_nl : STD_LOGIC;
  SIGNAL nor_879_nl : STD_LOGIC;
  SIGNAL nor_880_nl : STD_LOGIC;
  SIGNAL mux_1892_nl : STD_LOGIC;
  SIGNAL mux_1891_nl : STD_LOGIC;
  SIGNAL mux_1890_nl : STD_LOGIC;
  SIGNAL nor_881_nl : STD_LOGIC;
  SIGNAL mux_1889_nl : STD_LOGIC;
  SIGNAL nor_882_nl : STD_LOGIC;
  SIGNAL nor_883_nl : STD_LOGIC;
  SIGNAL nor_884_nl : STD_LOGIC;
  SIGNAL mux_1888_nl : STD_LOGIC;
  SIGNAL nor_885_nl : STD_LOGIC;
  SIGNAL mux_1887_nl : STD_LOGIC;
  SIGNAL mux_1886_nl : STD_LOGIC;
  SIGNAL nor_886_nl : STD_LOGIC;
  SIGNAL nor_887_nl : STD_LOGIC;
  SIGNAL nor_888_nl : STD_LOGIC;
  SIGNAL mux_1885_nl : STD_LOGIC;
  SIGNAL mux_1884_nl : STD_LOGIC;
  SIGNAL mux_1883_nl : STD_LOGIC;
  SIGNAL and_501_nl : STD_LOGIC;
  SIGNAL mux_1882_nl : STD_LOGIC;
  SIGNAL nor_889_nl : STD_LOGIC;
  SIGNAL nor_890_nl : STD_LOGIC;
  SIGNAL nor_891_nl : STD_LOGIC;
  SIGNAL mux_1881_nl : STD_LOGIC;
  SIGNAL or_1947_nl : STD_LOGIC;
  SIGNAL or_1945_nl : STD_LOGIC;
  SIGNAL mux_1880_nl : STD_LOGIC;
  SIGNAL nor_892_nl : STD_LOGIC;
  SIGNAL mux_1879_nl : STD_LOGIC;
  SIGNAL or_1943_nl : STD_LOGIC;
  SIGNAL or_1941_nl : STD_LOGIC;
  SIGNAL and_502_nl : STD_LOGIC;
  SIGNAL mux_1877_nl : STD_LOGIC;
  SIGNAL nor_894_nl : STD_LOGIC;
  SIGNAL mux_1876_nl : STD_LOGIC;
  SIGNAL mux_1875_nl : STD_LOGIC;
  SIGNAL or_1937_nl : STD_LOGIC;
  SIGNAL or_1935_nl : STD_LOGIC;
  SIGNAL mux_1874_nl : STD_LOGIC;
  SIGNAL or_1934_nl : STD_LOGIC;
  SIGNAL or_1932_nl : STD_LOGIC;
  SIGNAL and_504_nl : STD_LOGIC;
  SIGNAL mux_1873_nl : STD_LOGIC;
  SIGNAL mux_1872_nl : STD_LOGIC;
  SIGNAL nor_895_nl : STD_LOGIC;
  SIGNAL nor_896_nl : STD_LOGIC;
  SIGNAL mux_1871_nl : STD_LOGIC;
  SIGNAL nor_897_nl : STD_LOGIC;
  SIGNAL nor_898_nl : STD_LOGIC;
  SIGNAL nor_846_nl : STD_LOGIC;
  SIGNAL mux_1931_nl : STD_LOGIC;
  SIGNAL mux_1930_nl : STD_LOGIC;
  SIGNAL and_497_nl : STD_LOGIC;
  SIGNAL mux_1929_nl : STD_LOGIC;
  SIGNAL nor_847_nl : STD_LOGIC;
  SIGNAL mux_1926_nl : STD_LOGIC;
  SIGNAL mux_1925_nl : STD_LOGIC;
  SIGNAL nor_848_nl : STD_LOGIC;
  SIGNAL nor_849_nl : STD_LOGIC;
  SIGNAL mux_1924_nl : STD_LOGIC;
  SIGNAL nor_850_nl : STD_LOGIC;
  SIGNAL nor_851_nl : STD_LOGIC;
  SIGNAL mux_1923_nl : STD_LOGIC;
  SIGNAL mux_1922_nl : STD_LOGIC;
  SIGNAL mux_1921_nl : STD_LOGIC;
  SIGNAL nor_852_nl : STD_LOGIC;
  SIGNAL nor_853_nl : STD_LOGIC;
  SIGNAL mux_1920_nl : STD_LOGIC;
  SIGNAL and_498_nl : STD_LOGIC;
  SIGNAL nor_854_nl : STD_LOGIC;
  SIGNAL mux_1919_nl : STD_LOGIC;
  SIGNAL mux_1918_nl : STD_LOGIC;
  SIGNAL and_840_nl : STD_LOGIC;
  SIGNAL nor_856_nl : STD_LOGIC;
  SIGNAL mux_1917_nl : STD_LOGIC;
  SIGNAL nor_857_nl : STD_LOGIC;
  SIGNAL nor_858_nl : STD_LOGIC;
  SIGNAL mux_1916_nl : STD_LOGIC;
  SIGNAL mux_1915_nl : STD_LOGIC;
  SIGNAL mux_1914_nl : STD_LOGIC;
  SIGNAL mux_1913_nl : STD_LOGIC;
  SIGNAL nor_859_nl : STD_LOGIC;
  SIGNAL mux_1912_nl : STD_LOGIC;
  SIGNAL nor_861_nl : STD_LOGIC;
  SIGNAL mux_1911_nl : STD_LOGIC;
  SIGNAL mux_1910_nl : STD_LOGIC;
  SIGNAL and_849_nl : STD_LOGIC;
  SIGNAL mux_1909_nl : STD_LOGIC;
  SIGNAL nor_865_nl : STD_LOGIC;
  SIGNAL mux_1908_nl : STD_LOGIC;
  SIGNAL mux_1907_nl : STD_LOGIC;
  SIGNAL mux_1906_nl : STD_LOGIC;
  SIGNAL nor_866_nl : STD_LOGIC;
  SIGNAL nor_867_nl : STD_LOGIC;
  SIGNAL mux_1905_nl : STD_LOGIC;
  SIGNAL and_500_nl : STD_LOGIC;
  SIGNAL nor_868_nl : STD_LOGIC;
  SIGNAL mux_1904_nl : STD_LOGIC;
  SIGNAL mux_1903_nl : STD_LOGIC;
  SIGNAL and_866_nl : STD_LOGIC;
  SIGNAL nor_870_nl : STD_LOGIC;
  SIGNAL mux_1902_nl : STD_LOGIC;
  SIGNAL nor_871_nl : STD_LOGIC;
  SIGNAL nor_872_nl : STD_LOGIC;
  SIGNAL mux_1963_nl : STD_LOGIC;
  SIGNAL mux_1962_nl : STD_LOGIC;
  SIGNAL mux_1961_nl : STD_LOGIC;
  SIGNAL mux_1960_nl : STD_LOGIC;
  SIGNAL nor_818_nl : STD_LOGIC;
  SIGNAL nor_819_nl : STD_LOGIC;
  SIGNAL mux_1959_nl : STD_LOGIC;
  SIGNAL nor_820_nl : STD_LOGIC;
  SIGNAL nor_821_nl : STD_LOGIC;
  SIGNAL mux_1958_nl : STD_LOGIC;
  SIGNAL mux_1957_nl : STD_LOGIC;
  SIGNAL nor_822_nl : STD_LOGIC;
  SIGNAL nor_823_nl : STD_LOGIC;
  SIGNAL nor_824_nl : STD_LOGIC;
  SIGNAL mux_1956_nl : STD_LOGIC;
  SIGNAL mux_1955_nl : STD_LOGIC;
  SIGNAL mux_1954_nl : STD_LOGIC;
  SIGNAL nor_825_nl : STD_LOGIC;
  SIGNAL and_848_nl : STD_LOGIC;
  SIGNAL mux_1953_nl : STD_LOGIC;
  SIGNAL and_856_nl : STD_LOGIC;
  SIGNAL nor_828_nl : STD_LOGIC;
  SIGNAL mux_1952_nl : STD_LOGIC;
  SIGNAL mux_1951_nl : STD_LOGIC;
  SIGNAL and_864_nl : STD_LOGIC;
  SIGNAL and_865_nl : STD_LOGIC;
  SIGNAL mux_1950_nl : STD_LOGIC;
  SIGNAL mux_1949_nl : STD_LOGIC;
  SIGNAL nor_831_nl : STD_LOGIC;
  SIGNAL nor_832_nl : STD_LOGIC;
  SIGNAL nor_833_nl : STD_LOGIC;
  SIGNAL and_489_nl : STD_LOGIC;
  SIGNAL mux_1948_nl : STD_LOGIC;
  SIGNAL mux_1947_nl : STD_LOGIC;
  SIGNAL mux_1946_nl : STD_LOGIC;
  SIGNAL mux_1945_nl : STD_LOGIC;
  SIGNAL and_491_nl : STD_LOGIC;
  SIGNAL mux_1944_nl : STD_LOGIC;
  SIGNAL nor_835_nl : STD_LOGIC;
  SIGNAL nor_836_nl : STD_LOGIC;
  SIGNAL mux_1943_nl : STD_LOGIC;
  SIGNAL mux_1942_nl : STD_LOGIC;
  SIGNAL and_492_nl : STD_LOGIC;
  SIGNAL mux_1939_nl : STD_LOGIC;
  SIGNAL mux_1938_nl : STD_LOGIC;
  SIGNAL mux_1937_nl : STD_LOGIC;
  SIGNAL nor_840_nl : STD_LOGIC;
  SIGNAL nor_841_nl : STD_LOGIC;
  SIGNAL mux_1936_nl : STD_LOGIC;
  SIGNAL nor_842_nl : STD_LOGIC;
  SIGNAL nor_843_nl : STD_LOGIC;
  SIGNAL mux_1935_nl : STD_LOGIC;
  SIGNAL mux_1934_nl : STD_LOGIC;
  SIGNAL and_495_nl : STD_LOGIC;
  SIGNAL nor_844_nl : STD_LOGIC;
  SIGNAL mux_1933_nl : STD_LOGIC;
  SIGNAL and_496_nl : STD_LOGIC;
  SIGNAL nor_845_nl : STD_LOGIC;
  SIGNAL nor_792_nl : STD_LOGIC;
  SIGNAL mux_1994_nl : STD_LOGIC;
  SIGNAL mux_1993_nl : STD_LOGIC;
  SIGNAL nor_793_nl : STD_LOGIC;
  SIGNAL mux_1992_nl : STD_LOGIC;
  SIGNAL nand_79_nl : STD_LOGIC;
  SIGNAL mux_1989_nl : STD_LOGIC;
  SIGNAL mux_1988_nl : STD_LOGIC;
  SIGNAL nand_156_nl : STD_LOGIC;
  SIGNAL or_2109_nl : STD_LOGIC;
  SIGNAL mux_1987_nl : STD_LOGIC;
  SIGNAL nand_158_nl : STD_LOGIC;
  SIGNAL or_2106_nl : STD_LOGIC;
  SIGNAL mux_1986_nl : STD_LOGIC;
  SIGNAL mux_1985_nl : STD_LOGIC;
  SIGNAL mux_1984_nl : STD_LOGIC;
  SIGNAL nor_797_nl : STD_LOGIC;
  SIGNAL nor_798_nl : STD_LOGIC;
  SIGNAL mux_1983_nl : STD_LOGIC;
  SIGNAL and_486_nl : STD_LOGIC;
  SIGNAL nor_799_nl : STD_LOGIC;
  SIGNAL mux_1982_nl : STD_LOGIC;
  SIGNAL mux_1981_nl : STD_LOGIC;
  SIGNAL and_839_nl : STD_LOGIC;
  SIGNAL nor_801_nl : STD_LOGIC;
  SIGNAL mux_1980_nl : STD_LOGIC;
  SIGNAL nor_802_nl : STD_LOGIC;
  SIGNAL nor_803_nl : STD_LOGIC;
  SIGNAL mux_1979_nl : STD_LOGIC;
  SIGNAL mux_1978_nl : STD_LOGIC;
  SIGNAL mux_1977_nl : STD_LOGIC;
  SIGNAL mux_1976_nl : STD_LOGIC;
  SIGNAL nor_804_nl : STD_LOGIC;
  SIGNAL nor_805_nl : STD_LOGIC;
  SIGNAL mux_1975_nl : STD_LOGIC;
  SIGNAL and_487_nl : STD_LOGIC;
  SIGNAL nor_806_nl : STD_LOGIC;
  SIGNAL mux_1974_nl : STD_LOGIC;
  SIGNAL mux_1973_nl : STD_LOGIC;
  SIGNAL and_847_nl : STD_LOGIC;
  SIGNAL nor_808_nl : STD_LOGIC;
  SIGNAL mux_1972_nl : STD_LOGIC;
  SIGNAL nor_809_nl : STD_LOGIC;
  SIGNAL nor_810_nl : STD_LOGIC;
  SIGNAL mux_1971_nl : STD_LOGIC;
  SIGNAL mux_1970_nl : STD_LOGIC;
  SIGNAL mux_1969_nl : STD_LOGIC;
  SIGNAL nor_811_nl : STD_LOGIC;
  SIGNAL nor_812_nl : STD_LOGIC;
  SIGNAL mux_1968_nl : STD_LOGIC;
  SIGNAL and_488_nl : STD_LOGIC;
  SIGNAL nor_813_nl : STD_LOGIC;
  SIGNAL mux_1967_nl : STD_LOGIC;
  SIGNAL mux_1966_nl : STD_LOGIC;
  SIGNAL and_863_nl : STD_LOGIC;
  SIGNAL nor_815_nl : STD_LOGIC;
  SIGNAL mux_1965_nl : STD_LOGIC;
  SIGNAL nor_816_nl : STD_LOGIC;
  SIGNAL nor_817_nl : STD_LOGIC;
  SIGNAL mux_2025_nl : STD_LOGIC;
  SIGNAL mux_2024_nl : STD_LOGIC;
  SIGNAL mux_2023_nl : STD_LOGIC;
  SIGNAL nor_769_nl : STD_LOGIC;
  SIGNAL mux_2022_nl : STD_LOGIC;
  SIGNAL mux_2021_nl : STD_LOGIC;
  SIGNAL nor_770_nl : STD_LOGIC;
  SIGNAL nor_771_nl : STD_LOGIC;
  SIGNAL nor_772_nl : STD_LOGIC;
  SIGNAL mux_2020_nl : STD_LOGIC;
  SIGNAL mux_2019_nl : STD_LOGIC;
  SIGNAL mux_2018_nl : STD_LOGIC;
  SIGNAL nor_773_nl : STD_LOGIC;
  SIGNAL nor_774_nl : STD_LOGIC;
  SIGNAL nor_775_nl : STD_LOGIC;
  SIGNAL nor_776_nl : STD_LOGIC;
  SIGNAL mux_2017_nl : STD_LOGIC;
  SIGNAL mux_2016_nl : STD_LOGIC;
  SIGNAL mux_2015_nl : STD_LOGIC;
  SIGNAL nor_777_nl : STD_LOGIC;
  SIGNAL mux_2014_nl : STD_LOGIC;
  SIGNAL nor_778_nl : STD_LOGIC;
  SIGNAL nor_779_nl : STD_LOGIC;
  SIGNAL nor_780_nl : STD_LOGIC;
  SIGNAL mux_2013_nl : STD_LOGIC;
  SIGNAL nor_781_nl : STD_LOGIC;
  SIGNAL mux_2012_nl : STD_LOGIC;
  SIGNAL mux_2011_nl : STD_LOGIC;
  SIGNAL nor_782_nl : STD_LOGIC;
  SIGNAL nor_783_nl : STD_LOGIC;
  SIGNAL nor_784_nl : STD_LOGIC;
  SIGNAL mux_2010_nl : STD_LOGIC;
  SIGNAL mux_2009_nl : STD_LOGIC;
  SIGNAL mux_2008_nl : STD_LOGIC;
  SIGNAL and_479_nl : STD_LOGIC;
  SIGNAL mux_2007_nl : STD_LOGIC;
  SIGNAL nor_785_nl : STD_LOGIC;
  SIGNAL and_480_nl : STD_LOGIC;
  SIGNAL nor_786_nl : STD_LOGIC;
  SIGNAL mux_2006_nl : STD_LOGIC;
  SIGNAL or_2136_nl : STD_LOGIC;
  SIGNAL nand_149_nl : STD_LOGIC;
  SIGNAL mux_2005_nl : STD_LOGIC;
  SIGNAL nor_787_nl : STD_LOGIC;
  SIGNAL mux_2004_nl : STD_LOGIC;
  SIGNAL or_2132_nl : STD_LOGIC;
  SIGNAL nand_150_nl : STD_LOGIC;
  SIGNAL and_481_nl : STD_LOGIC;
  SIGNAL mux_2002_nl : STD_LOGIC;
  SIGNAL nor_789_nl : STD_LOGIC;
  SIGNAL mux_2001_nl : STD_LOGIC;
  SIGNAL mux_2000_nl : STD_LOGIC;
  SIGNAL or_2126_nl : STD_LOGIC;
  SIGNAL nand_151_nl : STD_LOGIC;
  SIGNAL mux_1999_nl : STD_LOGIC;
  SIGNAL or_2123_nl : STD_LOGIC;
  SIGNAL nand_152_nl : STD_LOGIC;
  SIGNAL and_483_nl : STD_LOGIC;
  SIGNAL mux_1998_nl : STD_LOGIC;
  SIGNAL mux_1997_nl : STD_LOGIC;
  SIGNAL and_484_nl : STD_LOGIC;
  SIGNAL nor_790_nl : STD_LOGIC;
  SIGNAL mux_1996_nl : STD_LOGIC;
  SIGNAL and_485_nl : STD_LOGIC;
  SIGNAL nor_791_nl : STD_LOGIC;
  SIGNAL nor_751_nl : STD_LOGIC;
  SIGNAL mux_2056_nl : STD_LOGIC;
  SIGNAL mux_2055_nl : STD_LOGIC;
  SIGNAL and_463_nl : STD_LOGIC;
  SIGNAL mux_2054_nl : STD_LOGIC;
  SIGNAL and_464_nl : STD_LOGIC;
  SIGNAL mux_2051_nl : STD_LOGIC;
  SIGNAL mux_2050_nl : STD_LOGIC;
  SIGNAL and_465_nl : STD_LOGIC;
  SIGNAL nor_755_nl : STD_LOGIC;
  SIGNAL mux_2049_nl : STD_LOGIC;
  SIGNAL and_466_nl : STD_LOGIC;
  SIGNAL nor_756_nl : STD_LOGIC;
  SIGNAL mux_2048_nl : STD_LOGIC;
  SIGNAL mux_2047_nl : STD_LOGIC;
  SIGNAL mux_2046_nl : STD_LOGIC;
  SIGNAL and_467_nl : STD_LOGIC;
  SIGNAL nor_757_nl : STD_LOGIC;
  SIGNAL mux_2045_nl : STD_LOGIC;
  SIGNAL and_468_nl : STD_LOGIC;
  SIGNAL and_469_nl : STD_LOGIC;
  SIGNAL mux_2044_nl : STD_LOGIC;
  SIGNAL mux_2043_nl : STD_LOGIC;
  SIGNAL and_838_nl : STD_LOGIC;
  SIGNAL and_844_nl : STD_LOGIC;
  SIGNAL mux_2042_nl : STD_LOGIC;
  SIGNAL and_470_nl : STD_LOGIC;
  SIGNAL nor_760_nl : STD_LOGIC;
  SIGNAL mux_2041_nl : STD_LOGIC;
  SIGNAL mux_2040_nl : STD_LOGIC;
  SIGNAL mux_2039_nl : STD_LOGIC;
  SIGNAL mux_2038_nl : STD_LOGIC;
  SIGNAL and_471_nl : STD_LOGIC;
  SIGNAL mux_2037_nl : STD_LOGIC;
  SIGNAL and_473_nl : STD_LOGIC;
  SIGNAL mux_2036_nl : STD_LOGIC;
  SIGNAL mux_2035_nl : STD_LOGIC;
  SIGNAL and_846_nl : STD_LOGIC;
  SIGNAL mux_2034_nl : STD_LOGIC;
  SIGNAL nor_764_nl : STD_LOGIC;
  SIGNAL mux_2033_nl : STD_LOGIC;
  SIGNAL mux_2032_nl : STD_LOGIC;
  SIGNAL mux_2031_nl : STD_LOGIC;
  SIGNAL and_475_nl : STD_LOGIC;
  SIGNAL nor_765_nl : STD_LOGIC;
  SIGNAL mux_2030_nl : STD_LOGIC;
  SIGNAL and_476_nl : STD_LOGIC;
  SIGNAL and_477_nl : STD_LOGIC;
  SIGNAL mux_2029_nl : STD_LOGIC;
  SIGNAL mux_2028_nl : STD_LOGIC;
  SIGNAL and_861_nl : STD_LOGIC;
  SIGNAL and_862_nl : STD_LOGIC;
  SIGNAL mux_2027_nl : STD_LOGIC;
  SIGNAL and_478_nl : STD_LOGIC;
  SIGNAL nor_768_nl : STD_LOGIC;
  SIGNAL mux_2088_nl : STD_LOGIC;
  SIGNAL mux_2087_nl : STD_LOGIC;
  SIGNAL mux_2086_nl : STD_LOGIC;
  SIGNAL mux_2085_nl : STD_LOGIC;
  SIGNAL nor_731_nl : STD_LOGIC;
  SIGNAL nor_732_nl : STD_LOGIC;
  SIGNAL mux_2084_nl : STD_LOGIC;
  SIGNAL nor_733_nl : STD_LOGIC;
  SIGNAL nor_734_nl : STD_LOGIC;
  SIGNAL mux_2083_nl : STD_LOGIC;
  SIGNAL mux_2082_nl : STD_LOGIC;
  SIGNAL nor_735_nl : STD_LOGIC;
  SIGNAL nor_736_nl : STD_LOGIC;
  SIGNAL nor_737_nl : STD_LOGIC;
  SIGNAL mux_2081_nl : STD_LOGIC;
  SIGNAL mux_2080_nl : STD_LOGIC;
  SIGNAL mux_2079_nl : STD_LOGIC;
  SIGNAL and_447_nl : STD_LOGIC;
  SIGNAL and_845_nl : STD_LOGIC;
  SIGNAL mux_2078_nl : STD_LOGIC;
  SIGNAL and_854_nl : STD_LOGIC;
  SIGNAL nor_740_nl : STD_LOGIC;
  SIGNAL mux_2077_nl : STD_LOGIC;
  SIGNAL mux_2076_nl : STD_LOGIC;
  SIGNAL and_859_nl : STD_LOGIC;
  SIGNAL and_860_nl : STD_LOGIC;
  SIGNAL mux_2075_nl : STD_LOGIC;
  SIGNAL mux_2074_nl : STD_LOGIC;
  SIGNAL and_448_nl : STD_LOGIC;
  SIGNAL nor_743_nl : STD_LOGIC;
  SIGNAL nor_744_nl : STD_LOGIC;
  SIGNAL and_449_nl : STD_LOGIC;
  SIGNAL mux_2073_nl : STD_LOGIC;
  SIGNAL mux_2072_nl : STD_LOGIC;
  SIGNAL mux_2071_nl : STD_LOGIC;
  SIGNAL mux_2070_nl : STD_LOGIC;
  SIGNAL and_451_nl : STD_LOGIC;
  SIGNAL mux_2069_nl : STD_LOGIC;
  SIGNAL and_833_nl : STD_LOGIC;
  SIGNAL and_452_nl : STD_LOGIC;
  SIGNAL mux_2068_nl : STD_LOGIC;
  SIGNAL mux_2067_nl : STD_LOGIC;
  SIGNAL and_454_nl : STD_LOGIC;
  SIGNAL mux_2064_nl : STD_LOGIC;
  SIGNAL mux_2063_nl : STD_LOGIC;
  SIGNAL mux_2062_nl : STD_LOGIC;
  SIGNAL and_837_nl : STD_LOGIC;
  SIGNAL and_457_nl : STD_LOGIC;
  SIGNAL mux_2061_nl : STD_LOGIC;
  SIGNAL and_843_nl : STD_LOGIC;
  SIGNAL and_458_nl : STD_LOGIC;
  SIGNAL mux_2060_nl : STD_LOGIC;
  SIGNAL mux_2059_nl : STD_LOGIC;
  SIGNAL and_459_nl : STD_LOGIC;
  SIGNAL and_460_nl : STD_LOGIC;
  SIGNAL mux_2058_nl : STD_LOGIC;
  SIGNAL and_461_nl : STD_LOGIC;
  SIGNAL and_462_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_1_tmp_mul_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL mux_2097_nl : STD_LOGIC;
  SIGNAL mux_2096_nl : STD_LOGIC;
  SIGNAL or_2260_nl : STD_LOGIC;
  SIGNAL mux_2095_nl : STD_LOGIC;
  SIGNAL mux_2094_nl : STD_LOGIC;
  SIGNAL or_2257_nl : STD_LOGIC;
  SIGNAL mux_2093_nl : STD_LOGIC;
  SIGNAL mux_2092_nl : STD_LOGIC;
  SIGNAL mux_2091_nl : STD_LOGIC;
  SIGNAL or_2255_nl : STD_LOGIC;
  SIGNAL mux_2090_nl : STD_LOGIC;
  SIGNAL or_2254_nl : STD_LOGIC;
  SIGNAL or_2253_nl : STD_LOGIC;
  SIGNAL mux_2104_nl : STD_LOGIC;
  SIGNAL mux_2103_nl : STD_LOGIC;
  SIGNAL mux_2102_nl : STD_LOGIC;
  SIGNAL nor_723_nl : STD_LOGIC;
  SIGNAL mux_2115_nl : STD_LOGIC;
  SIGNAL mux_2114_nl : STD_LOGIC;
  SIGNAL mux_2113_nl : STD_LOGIC;
  SIGNAL mux_2112_nl : STD_LOGIC;
  SIGNAL nor_711_nl : STD_LOGIC;
  SIGNAL and_445_nl : STD_LOGIC;
  SIGNAL mux_2122_nl : STD_LOGIC;
  SIGNAL mux_2121_nl : STD_LOGIC;
  SIGNAL mux_2120_nl : STD_LOGIC;
  SIGNAL nor_703_nl : STD_LOGIC;
  SIGNAL nor_692_nl : STD_LOGIC;
  SIGNAL mux_2135_nl : STD_LOGIC;
  SIGNAL mux_2134_nl : STD_LOGIC;
  SIGNAL mux_2133_nl : STD_LOGIC;
  SIGNAL nor_689_nl : STD_LOGIC;
  SIGNAL nor_690_nl : STD_LOGIC;
  SIGNAL mux_2129_nl : STD_LOGIC;
  SIGNAL mux_2127_nl : STD_LOGIC;
  SIGNAL nor_696_nl : STD_LOGIC;
  SIGNAL mux_2142_nl : STD_LOGIC;
  SIGNAL mux_2141_nl : STD_LOGIC;
  SIGNAL mux_2140_nl : STD_LOGIC;
  SIGNAL nor_681_nl : STD_LOGIC;
  SIGNAL mux_2153_nl : STD_LOGIC;
  SIGNAL mux_2152_nl : STD_LOGIC;
  SIGNAL mux_2151_nl : STD_LOGIC;
  SIGNAL mux_2150_nl : STD_LOGIC;
  SIGNAL nor_669_nl : STD_LOGIC;
  SIGNAL and_443_nl : STD_LOGIC;
  SIGNAL mux_2160_nl : STD_LOGIC;
  SIGNAL mux_2159_nl : STD_LOGIC;
  SIGNAL mux_2158_nl : STD_LOGIC;
  SIGNAL nor_661_nl : STD_LOGIC;
  SIGNAL nor_650_nl : STD_LOGIC;
  SIGNAL mux_2174_nl : STD_LOGIC;
  SIGNAL mux_2173_nl : STD_LOGIC;
  SIGNAL mux_2172_nl : STD_LOGIC;
  SIGNAL nor_646_nl : STD_LOGIC;
  SIGNAL mux_2171_nl : STD_LOGIC;
  SIGNAL nor_648_nl : STD_LOGIC;
  SIGNAL mux_2167_nl : STD_LOGIC;
  SIGNAL mux_2165_nl : STD_LOGIC;
  SIGNAL nor_654_nl : STD_LOGIC;
  SIGNAL mux_2181_nl : STD_LOGIC;
  SIGNAL mux_2180_nl : STD_LOGIC;
  SIGNAL mux_2179_nl : STD_LOGIC;
  SIGNAL nor_638_nl : STD_LOGIC;
  SIGNAL mux_2192_nl : STD_LOGIC;
  SIGNAL mux_2191_nl : STD_LOGIC;
  SIGNAL mux_2190_nl : STD_LOGIC;
  SIGNAL mux_2189_nl : STD_LOGIC;
  SIGNAL nor_626_nl : STD_LOGIC;
  SIGNAL and_441_nl : STD_LOGIC;
  SIGNAL mux_2199_nl : STD_LOGIC;
  SIGNAL mux_2198_nl : STD_LOGIC;
  SIGNAL mux_2197_nl : STD_LOGIC;
  SIGNAL nor_618_nl : STD_LOGIC;
  SIGNAL nor_607_nl : STD_LOGIC;
  SIGNAL mux_2212_nl : STD_LOGIC;
  SIGNAL mux_2211_nl : STD_LOGIC;
  SIGNAL mux_2210_nl : STD_LOGIC;
  SIGNAL nor_604_nl : STD_LOGIC;
  SIGNAL nor_605_nl : STD_LOGIC;
  SIGNAL mux_2206_nl : STD_LOGIC;
  SIGNAL mux_2204_nl : STD_LOGIC;
  SIGNAL nor_611_nl : STD_LOGIC;
  SIGNAL mux_2219_nl : STD_LOGIC;
  SIGNAL mux_2218_nl : STD_LOGIC;
  SIGNAL mux_2217_nl : STD_LOGIC;
  SIGNAL nor_596_nl : STD_LOGIC;
  SIGNAL mux_2230_nl : STD_LOGIC;
  SIGNAL mux_2229_nl : STD_LOGIC;
  SIGNAL mux_2228_nl : STD_LOGIC;
  SIGNAL mux_2227_nl : STD_LOGIC;
  SIGNAL and_434_nl : STD_LOGIC;
  SIGNAL and_435_nl : STD_LOGIC;
  SIGNAL mux_2237_nl : STD_LOGIC;
  SIGNAL mux_2236_nl : STD_LOGIC;
  SIGNAL mux_2235_nl : STD_LOGIC;
  SIGNAL and_426_nl : STD_LOGIC;
  SIGNAL acc_nl : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_mux_358_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nand_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux_359_nl : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_and_260_nl : STD_LOGIC_VECTOR (53 DOWNTO 0);
  SIGNAL COMP_LOOP_mux1h_710_nl : STD_LOGIC_VECTOR (53 DOWNTO 0);
  SIGNAL COMP_LOOP_and_261_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_711_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_262_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_712_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_713_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_and_983_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_984_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_985_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_986_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_987_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_988_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_989_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_990_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_991_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_992_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_993_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_994_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_995_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_996_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_997_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_998_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_999_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1000_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1001_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1002_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1003_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1004_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1005_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1006_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1007_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1008_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1009_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1010_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1011_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1012_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1013_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1014_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1015_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1016_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1017_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1018_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1019_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1020_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1021_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1022_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1023_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1024_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1025_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1026_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1027_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1028_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1029_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1030_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1031_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1032_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1033_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1034_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1035_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1036_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_263_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_mux_8_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_264_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_714_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_715_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_or_61_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_716_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_62_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_717_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_2_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux_360_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_3_nl : STD_LOGIC;
  SIGNAL STAGE_LOOP_mux_4_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_mux1h_718_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_719_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1037_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1038_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1039_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1040_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1041_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1042_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1043_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1044_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1045_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1046_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1047_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1048_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1049_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1050_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1051_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_720_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1052_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1053_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1054_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1055_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1056_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1057_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1058_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1059_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1060_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1061_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1062_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1063_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1064_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1065_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1066_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_721_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_722_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1067_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1068_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1069_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1070_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1071_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1072_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1073_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1074_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1075_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1076_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1077_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1078_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1079_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1080_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1081_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_723_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_724_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_725_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_726_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1082_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1083_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1084_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1085_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1086_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1087_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1088_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1089_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1090_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1091_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1092_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1093_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1094_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1095_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1096_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_727_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_728_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_729_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_730_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_731_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_732_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_733_nl : STD_LOGIC;
  SIGNAL p_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL p_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT modulo
    PORT (
      base_rsc_dat : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      m_rsc_dat : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      return_rsc_z : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      ccs_ccore_start_rsc_dat : IN STD_LOGIC;
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_srst : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL COMP_LOOP_1_modulo_cmp_base_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_cmp_m_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_cmp_return_rsc_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_cmp_ccs_ccore_start_rsc_dat : STD_LOGIC;

  SIGNAL COMP_LOOP_1_tmp_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL COMP_LOOP_1_tmp_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_1_tmp_lshift_rg_z : STD_LOGIC_VECTOR (5 DOWNTO 0);

  SIGNAL COMP_LOOP_9_tmp_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL COMP_LOOP_9_tmp_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_9_tmp_lshift_rg_z : STD_LOGIC_VECTOR (10 DOWNTO 0);

  SIGNAL COMP_LOOP_2_tmp_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL COMP_LOOP_2_tmp_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_2_tmp_lshift_rg_z : STD_LOGIC_VECTOR (9 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_core_wait_dp
    PORT(
      ensig_cgo_iro : IN STD_LOGIC;
      ensig_cgo : IN STD_LOGIC;
      COMP_LOOP_1_modulo_cmp_ccs_ccore_en : OUT STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
      COMP_LOOP_C_31_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_62_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_93_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_124_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_155_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_186_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_217_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_248_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_279_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_310_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_341_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_372_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_403_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_434_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_465_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_496_tr0 : IN STD_LOGIC;
      VEC_LOOP_C_0_tr0 : IN STD_LOGIC;
      STAGE_LOOP_C_1_tr0 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (8 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_31_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_62_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_93_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_124_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_155_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_186_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_217_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_248_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_279_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_310_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_341_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_372_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_403_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_434_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_465_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_496_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_s_1_16_2(input_15 : STD_LOGIC;
  input_14 : STD_LOGIC;
  input_13 : STD_LOGIC;
  input_12 : STD_LOGIC;
  input_11 : STD_LOGIC;
  input_10 : STD_LOGIC;
  input_9 : STD_LOGIC;
  input_8 : STD_LOGIC;
  input_7 : STD_LOGIC;
  input_6 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(15 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
      tmp := sel(6);
      result := result or ( input_6 and tmp);
      tmp := sel(7);
      result := result or ( input_7 and tmp);
      tmp := sel(8);
      result := result or ( input_8 and tmp);
      tmp := sel(9);
      result := result or ( input_9 and tmp);
      tmp := sel(10);
      result := result or ( input_10 and tmp);
      tmp := sel(11);
      result := result or ( input_11 and tmp);
      tmp := sel(12);
      result := result or ( input_12 and tmp);
      tmp := sel(13);
      result := result or ( input_13 and tmp);
      tmp := sel(14);
      result := result or ( input_14 and tmp);
      tmp := sel(15);
      result := result or ( input_15 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_17_2(input_16 : STD_LOGIC;
  input_15 : STD_LOGIC;
  input_14 : STD_LOGIC;
  input_13 : STD_LOGIC;
  input_12 : STD_LOGIC;
  input_11 : STD_LOGIC;
  input_10 : STD_LOGIC;
  input_9 : STD_LOGIC;
  input_8 : STD_LOGIC;
  input_7 : STD_LOGIC;
  input_6 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(16 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
      tmp := sel(6);
      result := result or ( input_6 and tmp);
      tmp := sel(7);
      result := result or ( input_7 and tmp);
      tmp := sel(8);
      result := result or ( input_8 and tmp);
      tmp := sel(9);
      result := result or ( input_9 and tmp);
      tmp := sel(10);
      result := result or ( input_10 and tmp);
      tmp := sel(11);
      result := result or ( input_11 and tmp);
      tmp := sel(12);
      result := result or ( input_12 and tmp);
      tmp := sel(13);
      result := result or ( input_13 and tmp);
      tmp := sel(14);
      result := result or ( input_14 and tmp);
      tmp := sel(15);
      result := result or ( input_15 and tmp);
      tmp := sel(16);
      result := result or ( input_16 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_18_2(input_17 : STD_LOGIC;
  input_16 : STD_LOGIC;
  input_15 : STD_LOGIC;
  input_14 : STD_LOGIC;
  input_13 : STD_LOGIC;
  input_12 : STD_LOGIC;
  input_11 : STD_LOGIC;
  input_10 : STD_LOGIC;
  input_9 : STD_LOGIC;
  input_8 : STD_LOGIC;
  input_7 : STD_LOGIC;
  input_6 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(17 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
      tmp := sel(6);
      result := result or ( input_6 and tmp);
      tmp := sel(7);
      result := result or ( input_7 and tmp);
      tmp := sel(8);
      result := result or ( input_8 and tmp);
      tmp := sel(9);
      result := result or ( input_9 and tmp);
      tmp := sel(10);
      result := result or ( input_10 and tmp);
      tmp := sel(11);
      result := result or ( input_11 and tmp);
      tmp := sel(12);
      result := result or ( input_12 and tmp);
      tmp := sel(13);
      result := result or ( input_13 and tmp);
      tmp := sel(14);
      result := result or ( input_14 and tmp);
      tmp := sel(15);
      result := result or ( input_15 and tmp);
      tmp := sel(16);
      result := result or ( input_16 and tmp);
      tmp := sel(17);
      result := result or ( input_17 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_3_2(input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_4_2(input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_5_2(input_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_54_15_2(input_14 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(14 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(53 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(53 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_16_2(input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(15 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_19_2(input_18 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(18 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_3_2(input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_4_2(input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_6_2(input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_32_2(input_31 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_30 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_29 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_28 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_27 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_26 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_25 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_24 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_23 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_22 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_21 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_20 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(31 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
      tmp := (OTHERS=>sel( 20));
      result := result or ( input_20 and tmp);
      tmp := (OTHERS=>sel( 21));
      result := result or ( input_21 and tmp);
      tmp := (OTHERS=>sel( 22));
      result := result or ( input_22 and tmp);
      tmp := (OTHERS=>sel( 23));
      result := result or ( input_23 and tmp);
      tmp := (OTHERS=>sel( 24));
      result := result or ( input_24 and tmp);
      tmp := (OTHERS=>sel( 25));
      result := result or ( input_25 and tmp);
      tmp := (OTHERS=>sel( 26));
      result := result or ( input_26 and tmp);
      tmp := (OTHERS=>sel( 27));
      result := result or ( input_27 and tmp);
      tmp := (OTHERS=>sel( 28));
      result := result or ( input_28 and tmp);
      tmp := (OTHERS=>sel( 29));
      result := result or ( input_29 and tmp);
      tmp := (OTHERS=>sel( 30));
      result := result or ( input_30 and tmp);
      tmp := (OTHERS=>sel( 31));
      result := result or ( input_31 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_3_2(input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_4_2(input_3 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_6_2(input_5 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_8_20_2(input_19 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(19 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_10_2_2(input_0 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(9 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_11_2_2(input_0 : STD_LOGIC_VECTOR(10 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(10 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(10 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_4_2_2(input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_54_2_2(input_0 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(53 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(53 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_64_2_2(input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_6_2_2(input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_7_2_2(input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_8_2_2(input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION minimum(arg1,arg2:INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1<arg2)THEN
      RETURN arg1;
    ELSE
      RETURN arg2;
    END IF;
  END;

  FUNCTION maximum(arg1,arg2:INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1>arg2)THEN
      RETURN arg1;
    ELSE
      RETURN arg2;
    END IF;
  END;

  FUNCTION READSLICE_64_65(input_val:STD_LOGIC_VECTOR(64 DOWNTO 0);index:INTEGER)
  RETURN STD_LOGIC_VECTOR IS
    CONSTANT min_sat_index:INTEGER:= maximum( index, 0 );
    CONSTANT sat_index:INTEGER:= minimum( min_sat_index, 1);
  BEGIN
    RETURN input_val(sat_index+63 DOWNTO sat_index);
  END;

BEGIN
  p_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 5,
      width => 64
      )
    PORT MAP(
      dat => p_rsci_dat,
      idat => p_rsci_idat_1
    );
  p_rsci_dat <= p_rsc_dat;
  p_rsci_idat <= p_rsci_idat_1;

  vec_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_15_lz
    );
  vec_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_14_lz
    );
  vec_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_13_lz
    );
  vec_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_12_lz
    );
  vec_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_11_lz
    );
  vec_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_10_lz
    );
  vec_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_9_lz
    );
  vec_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_8_lz
    );
  vec_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_7_lz
    );
  vec_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_6_lz
    );
  vec_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_5_lz
    );
  vec_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_4_lz
    );
  vec_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_3_lz
    );
  vec_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_2_lz
    );
  vec_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_1_lz
    );
  vec_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_0_lz
    );
  p_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => p_rsc_triosy_lz
    );
  r_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => r_rsc_triosy_lz
    );
  twiddle_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_15_lz
    );
  twiddle_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_14_lz
    );
  twiddle_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_13_lz
    );
  twiddle_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_12_lz
    );
  twiddle_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_11_lz
    );
  twiddle_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_10_lz
    );
  twiddle_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_9_lz
    );
  twiddle_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_8_lz
    );
  twiddle_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_7_lz
    );
  twiddle_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_6_lz
    );
  twiddle_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_5_lz
    );
  twiddle_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_4_lz
    );
  twiddle_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_3_lz
    );
  twiddle_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_2_lz
    );
  twiddle_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_1_lz
    );
  twiddle_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_0_lz
    );
  COMP_LOOP_1_modulo_cmp : modulo
    PORT MAP(
      base_rsc_dat => COMP_LOOP_1_modulo_cmp_base_rsc_dat,
      m_rsc_dat => COMP_LOOP_1_modulo_cmp_m_rsc_dat,
      return_rsc_z => COMP_LOOP_1_modulo_cmp_return_rsc_z_1,
      ccs_ccore_start_rsc_dat => COMP_LOOP_1_modulo_cmp_ccs_ccore_start_rsc_dat,
      ccs_ccore_clk => clk,
      ccs_ccore_srst => rst,
      ccs_ccore_en => COMP_LOOP_1_modulo_cmp_ccs_ccore_en
    );
  COMP_LOOP_1_modulo_cmp_base_rsc_dat <= MUX_v_64_2_2(COMP_LOOP_10_acc_8_itm, (READSLICE_64_65(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_361_cse
      & '1') + UNSIGNED((MUX_v_64_2_2((NOT COMP_LOOP_10_acc_8_itm), (NOT z_out_7),
      COMP_LOOP_or_18_itm)) & '1'), 65)), 1)), MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2((NOT
      (MUX_s_1_2_2((MUX_s_1_2_2(((fsm_output(3)) AND (fsm_output(8)) AND (fsm_output(0))
      AND (fsm_output(5))), (NOT((fsm_output(3)) OR (fsm_output(8)) OR not_tmp_676)),
      fsm_output(4))), mux_tmp_2249, fsm_output(6)))), (MUX_s_1_2_2((NOT mux_tmp_2249),
      mux_tmp_2245, fsm_output(6))), fsm_output(1))), mux_tmp_2246, fsm_output(7))),
      (MUX_s_1_2_2(mux_tmp_2246, (MUX_s_1_2_2((MUX_s_1_2_2(((fsm_output(4)) OR mux_tmp_2238),
      (MUX_s_1_2_2(mux_tmp_2237, ((NOT (fsm_output(3))) OR (fsm_output(8)) OR not_tmp_676),
      fsm_output(4))), fsm_output(6))), (MUX_s_1_2_2((MUX_s_1_2_2(mux_tmp_2237, mux_tmp_2238,
      fsm_output(4))), (NOT((fsm_output(4)) AND (NOT mux_tmp_2237))), fsm_output(6))),
      fsm_output(1))), fsm_output(7))), fsm_output(2)));
  COMP_LOOP_1_modulo_cmp_m_rsc_dat <= p_sva;
  COMP_LOOP_1_modulo_cmp_return_rsc_z <= COMP_LOOP_1_modulo_cmp_return_rsc_z_1;
  COMP_LOOP_1_modulo_cmp_ccs_ccore_start_rsc_dat <= NOT (MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2(((fsm_output(3))
      OR mux_tmp_2258), mux_tmp_2257, and_421_cse)), (MUX_s_1_2_2(((fsm_output(0))
      OR (NOT (fsm_output(3))) OR mux_tmp_2259), or_tmp_2279, fsm_output(5))), fsm_output(4))),
      (MUX_s_1_2_2(mux_tmp_2264, (MUX_s_1_2_2((MUX_s_1_2_2(or_tmp_2277, mux_tmp_2257,
      fsm_output(0))), (NOT((fsm_output(3)) AND (NOT mux_tmp_2256))), fsm_output(5))),
      fsm_output(4))), fsm_output(6))), (MUX_s_1_2_2((MUX_s_1_2_2(mux_tmp_2264, (MUX_s_1_2_2(or_tmp_2277,
      mux_tmp_2257, (fsm_output(5)) OR (fsm_output(0)))), fsm_output(4))), (MUX_s_1_2_2((MUX_s_1_2_2(or_tmp_2277,
      (MUX_s_1_2_2(mux_tmp_2259, mux_tmp_2258, fsm_output(3))), and_421_cse)), ((fsm_output(5))
      OR (fsm_output(0)) OR mux_tmp_2257), fsm_output(4))), fsm_output(6))), fsm_output(1)));

  COMP_LOOP_1_tmp_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_l_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 0,
      width_s => 4,
      width_z => 6
      )
    PORT MAP(
      a => COMP_LOOP_1_tmp_lshift_rg_a,
      s => COMP_LOOP_1_tmp_lshift_rg_s,
      z => COMP_LOOP_1_tmp_lshift_rg_z
    );
  COMP_LOOP_1_tmp_lshift_rg_a(0) <= '1';
  COMP_LOOP_1_tmp_lshift_rg_s <= z_out_4;
  COMP_LOOP_1_tmp_lshift_itm <= COMP_LOOP_1_tmp_lshift_rg_z;

  COMP_LOOP_9_tmp_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_l_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 0,
      width_s => 4,
      width_z => 11
      )
    PORT MAP(
      a => COMP_LOOP_9_tmp_lshift_rg_a,
      s => COMP_LOOP_9_tmp_lshift_rg_s,
      z => COMP_LOOP_9_tmp_lshift_rg_z
    );
  COMP_LOOP_9_tmp_lshift_rg_a(0) <= '1';
  COMP_LOOP_9_tmp_lshift_rg_s <= MUX_v_4_2_2(STAGE_LOOP_i_3_0_sva, z_out_4, CONV_SL_1_1(fsm_output=STD_LOGIC_VECTOR'("000000010")));
  z_out <= COMP_LOOP_9_tmp_lshift_rg_z;

  COMP_LOOP_2_tmp_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_l_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 0,
      width_s => 4,
      width_z => 10
      )
    PORT MAP(
      a => COMP_LOOP_2_tmp_lshift_rg_a,
      s => COMP_LOOP_2_tmp_lshift_rg_s,
      z => COMP_LOOP_2_tmp_lshift_rg_z
    );
  COMP_LOOP_2_tmp_lshift_rg_a(0) <= '1';
  COMP_LOOP_2_tmp_lshift_rg_s <= MUX_v_4_2_2(COMP_LOOP_1_tmp_acc_cse_sva, z_out_4,
      CONV_SL_1_1(fsm_output=STD_LOGIC_VECTOR'("000000010")));
  z_out_1 <= COMP_LOOP_2_tmp_lshift_rg_z;

  inPlaceNTT_DIF_core_wait_dp_inst : inPlaceNTT_DIF_core_wait_dp
    PORT MAP(
      ensig_cgo_iro => mux_2255_rmff,
      ensig_cgo => reg_ensig_cgo_cse,
      COMP_LOOP_1_modulo_cmp_ccs_ccore_en => COMP_LOOP_1_modulo_cmp_ccs_ccore_en
    );
  inPlaceNTT_DIF_core_core_fsm_inst : inPlaceNTT_DIF_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      fsm_output => inPlaceNTT_DIF_core_core_fsm_inst_fsm_output,
      COMP_LOOP_C_31_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_31_tr0,
      COMP_LOOP_C_62_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_62_tr0,
      COMP_LOOP_C_93_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_93_tr0,
      COMP_LOOP_C_124_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_124_tr0,
      COMP_LOOP_C_155_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_155_tr0,
      COMP_LOOP_C_186_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_186_tr0,
      COMP_LOOP_C_217_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_217_tr0,
      COMP_LOOP_C_248_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_248_tr0,
      COMP_LOOP_C_279_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_279_tr0,
      COMP_LOOP_C_310_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_310_tr0,
      COMP_LOOP_C_341_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_341_tr0,
      COMP_LOOP_C_372_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_372_tr0,
      COMP_LOOP_C_403_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_403_tr0,
      COMP_LOOP_C_434_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_434_tr0,
      COMP_LOOP_C_465_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_465_tr0,
      COMP_LOOP_C_496_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_496_tr0,
      VEC_LOOP_C_0_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0,
      STAGE_LOOP_C_1_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0
    );
  fsm_output <= inPlaceNTT_DIF_core_core_fsm_inst_fsm_output;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_31_tr0 <= NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_62_tr0 <= NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_93_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_124_tr0 <= NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_155_tr0 <= NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_186_tr0 <= NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_217_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_248_tr0 <= NOT COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_279_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_310_tr0 <= NOT COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_341_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_372_tr0 <= NOT COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_403_tr0 <= NOT COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_434_tr0 <= NOT COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_465_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_496_tr0 <= NOT COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0 <= z_out_2(10);
  inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0 <= NOT STAGE_LOOP_acc_itm_4_1;

  nor_1589_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(2)) OR (COMP_LOOP_acc_16_psp_sva(0))
      OR (NOT COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  nor_1590_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      OR (fsm_output(7)) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1128_cse <= MUX_s_1_2_2(nor_1589_nl, nor_1590_nl, fsm_output(2));
  nor_346_cse <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) OR (NOT (fsm_output(5))));
  nor_1554_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(7)) OR not_tmp_395);
  nand_271_cse <= NOT((fsm_output(2)) AND (fsm_output(7)) AND (fsm_output(6)) AND
      (fsm_output(8)));
  nand_272_cse <= NOT((COMP_LOOP_acc_1_cse_sva(0)) AND CONV_SL_1_1(fsm_output(8 DOWNTO
      6)=STD_LOGIC_VECTOR'("111")));
  nor_1528_cse <= NOT((COMP_LOOP_acc_16_psp_sva(0)) OR (NOT COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm)
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1529_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("001")));
  mux_1190_nl <= MUX_s_1_2_2(nor_1528_cse, nor_1529_nl, fsm_output(2));
  nor_1530_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1191_cse <= MUX_s_1_2_2(mux_1190_nl, nor_1530_nl, VEC_LOOP_j_10_0_sva_9_0(2));
  nor_351_cse <= NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")));
  nor_1523_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1526_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1527_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nand_265_cse <= NOT((COMP_LOOP_acc_10_cse_10_1_15_sva(1)) AND (fsm_output(7)) AND
      (fsm_output(4)) AND (fsm_output(8)));
  nor_1435_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(7)) OR not_tmp_395);
  nor_1402_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1405_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1406_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1352_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(2))) OR (COMP_LOOP_acc_16_psp_sva(0))
      OR (NOT COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  nor_1353_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      OR (fsm_output(7)) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1378_cse <= MUX_s_1_2_2(nor_1352_nl, nor_1353_nl, fsm_output(2));
  nor_1317_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(7)) OR not_tmp_395);
  nor_1286_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1289_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1290_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1291_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  nor_1293_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("001")));
  mux_1440_nl <= MUX_s_1_2_2(nor_1528_cse, nor_1293_nl, fsm_output(2));
  mux_1441_cse <= MUX_s_1_2_2(nor_1291_nl, mux_1440_nl, VEC_LOOP_j_10_0_sva_9_0(2));
  nor_1200_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(7)) OR not_tmp_395);
  nand_226_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111")));
  and_529_cse <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_1173_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1174_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nand_219_cse <= NOT((COMP_LOOP_acc_10_cse_10_1_sva(3)) AND (fsm_output(7)) AND
      (fsm_output(4)) AND (fsm_output(8)));
  nor_1121_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(2)) OR (NOT (COMP_LOOP_acc_16_psp_sva(0)))
      OR (NOT COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  nor_1122_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      OR (fsm_output(7)) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1628_cse <= MUX_s_1_2_2(nor_1121_nl, nor_1122_nl, fsm_output(2));
  nor_1086_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(7)) OR not_tmp_395);
  nand_211_cse <= NOT((COMP_LOOP_acc_10_cse_10_1_sva(3)) AND (fsm_output(2)) AND
      (fsm_output(7)) AND (fsm_output(6)) AND (fsm_output(8)));
  nand_212_cse <= NOT((COMP_LOOP_acc_1_cse_sva(3)) AND (COMP_LOOP_acc_1_cse_sva(0))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111")));
  and_523_cse <= (COMP_LOOP_acc_16_psp_sva(0)) AND COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_1061_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("001")));
  mux_1690_nl <= MUX_s_1_2_2(and_523_cse, nor_1061_nl, fsm_output(2));
  nor_1062_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1691_cse <= MUX_s_1_2_2(mux_1690_nl, nor_1062_nl, VEC_LOOP_j_10_0_sva_9_0(2));
  nor_1056_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1059_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1060_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_970_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(7)) OR not_tmp_395);
  and_506_cse <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_944_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_945_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  and_503_nl <= (VEC_LOOP_j_10_0_sva_9_0(2)) AND (COMP_LOOP_acc_16_psp_sva(0)) AND
      COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm AND (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      AND (fsm_output(7)) AND (fsm_output(4)) AND (NOT (fsm_output(8)));
  nor_893_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      OR (fsm_output(7)) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1878_cse <= MUX_s_1_2_2(and_503_nl, nor_893_nl, fsm_output(2));
  nor_860_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(7)) OR not_tmp_395);
  and_490_cse <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_837_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_838_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nand_170_cse <= NOT((COMP_LOOP_acc_1_cse_sva(2)) AND (COMP_LOOP_acc_1_cse_sva(3))
      AND (COMP_LOOP_acc_1_cse_sva(0)) AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111")));
  and_493_nl <= (fsm_output(2)) AND CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO
      0)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(8
      DOWNTO 6)=STD_LOGIC_VECTOR'("001"));
  nor_839_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("001")));
  mux_1940_nl <= MUX_s_1_2_2(and_523_cse, nor_839_nl, fsm_output(2));
  mux_1941_cse <= MUX_s_1_2_2(and_493_nl, mux_1940_nl, VEC_LOOP_j_10_0_sva_9_0(2));
  nor_761_cse <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(7))))) OR not_tmp_395);
  and_450_cse <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  and_836_cse <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("100"));
  and_453_cse <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("010"));
  or_2259_cse_1 <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"));
  nand_122_cse <= NOT((z_out_3(0)) AND (fsm_output(4)));
  nand_121_cse <= NOT(CONV_SL_1_1(z_out_3(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      (fsm_output(4)));
  mux_2251_nl <= MUX_s_1_2_2((NOT mux_tmp_2224), mux_955_cse, fsm_output(7));
  mux_2252_nl <= MUX_s_1_2_2(mux_2251_nl, mux_965_cse, fsm_output(0));
  mux_2253_nl <= MUX_s_1_2_2(mux_tmp_2229, (NOT mux_2252_nl), fsm_output(5));
  mux_2254_nl <= MUX_s_1_2_2(mux_952_cse, mux_2253_nl, fsm_output(6));
  mux_2245_nl <= MUX_s_1_2_2(mux_tmp_2225, mux_949_cse, fsm_output(0));
  mux_2249_nl <= MUX_s_1_2_2(mux_tmp_2229, mux_2245_nl, fsm_output(5));
  mux_2242_nl <= MUX_s_1_2_2(mux_949_cse, (NOT mux_965_cse), fsm_output(5));
  mux_2250_nl <= MUX_s_1_2_2(mux_2249_nl, mux_2242_nl, fsm_output(6));
  mux_2255_rmff <= MUX_s_1_2_2(mux_2254_nl, mux_2250_nl, fsm_output(1));
  and_421_cse <= (fsm_output(5)) AND (fsm_output(0));
  nor_1624_cse <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")));
  and_1189_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  nand_324_cse <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111")));
  and_831_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_nor_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
  COMP_LOOP_tmp_nor_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
  COMP_LOOP_tmp_nor_1_cse <= NOT((z_out_3(3)) OR (z_out_3(2)) OR (z_out_3(0)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
  COMP_LOOP_tmp_nor_3_cse <= NOT((z_out_3(3)) OR (z_out_3(1)) OR (z_out_3(0)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
  COMP_LOOP_tmp_nor_6_cse <= NOT(CONV_SL_1_1(z_out_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
  nor_1767_cse <= NOT((fsm_output(5)) OR (fsm_output(0)));
  and_407_cse <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11"));
  and_733_cse <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11"));
  or_2729_cse <= (fsm_output(6)) OR (fsm_output(1)) OR (fsm_output(7)) OR (fsm_output(2));
  and_728_cse <= or_2729_cse AND (fsm_output(8));
  and_712_cse <= (fsm_output(0)) AND (fsm_output(3));
  or_432_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"));
  and_674_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"));
  and_675_cse <= (fsm_output(4)) AND (fsm_output(8));
  or_2697_cse <= (fsm_output(6)) OR (fsm_output(2));
  nand_301_cse <= NOT((fsm_output(7)) AND (fsm_output(4)) AND (fsm_output(8)));
  nor_298_nl <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10")));
  mux_955_cse <= MUX_s_1_2_2(and_675_cse, (fsm_output(4)), nor_298_nl);
  or_611_cse <= (fsm_output(2)) OR mux_tmp_929;
  nor_1642_nl <= NOT((fsm_output(4)) OR (fsm_output(8)));
  mux_951_nl <= MUX_s_1_2_2(nor_1642_nl, and_675_cse, fsm_output(3));
  or_614_nl <= (fsm_output(2)) OR (NOT mux_951_nl);
  mux_952_cse <= MUX_s_1_2_2(or_614_nl, nand_tmp_13, fsm_output(7));
  mux_949_cse <= MUX_s_1_2_2(nand_tmp_13, or_611_cse, fsm_output(7));
  mux_965_cse <= MUX_s_1_2_2((NOT nand_tmp_13), mux_955_cse, fsm_output(7));
  COMP_LOOP_tmp_or_1_cse <= and_dcpl_62 OR and_dcpl_189 OR and_dcpl_181 OR and_dcpl_190
      OR and_dcpl_183 OR and_dcpl_191 OR and_dcpl_184 OR and_dcpl_192;
  COMP_LOOP_tmp_or_2_cse <= and_dcpl_62 OR and_dcpl_65 OR and_dcpl_181 OR and_dcpl_190
      OR and_dcpl_183 OR and_dcpl_191 OR and_dcpl_184 OR and_dcpl_192;
  COMP_LOOP_or_27_cse <= and_dcpl_181 OR and_dcpl_190 OR and_dcpl_183 OR and_dcpl_191
      OR and_dcpl_184 OR and_dcpl_192;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_17_cse <= CONV_SL_1_1(z_out_3(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_19_cse <= CONV_SL_1_1(z_out_3(2 DOWNTO 0)=STD_LOGIC_VECTOR'("101"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_20_cse <= CONV_SL_1_1(z_out_3(2 DOWNTO 0)=STD_LOGIC_VECTOR'("110"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_21_cse <= CONV_SL_1_1(z_out_3(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"));
  COMP_LOOP_or_31_cse <= and_dcpl_195 OR and_dcpl_197 OR and_dcpl_198;
  COMP_LOOP_or_23_cse <= and_dcpl_189 OR and_dcpl_181 OR and_dcpl_190 OR and_dcpl_183
      OR and_dcpl_191 OR and_dcpl_184 OR and_dcpl_192;
  nor_1630_cse <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00")));
  and_1191_cse <= (COMP_LOOP_10_tmp_mul_idiv_sva(1)) AND COMP_LOOP_tmp_nor_14_itm;
  and_1190_cse <= (COMP_LOOP_10_tmp_mul_idiv_sva(2)) AND COMP_LOOP_tmp_nor_16_itm;
  and_314_m1c <= and_dcpl_51 AND and_dcpl_111;
  COMP_LOOP_tmp_or_29_cse <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_155 OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_157
      OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_159;
  COMP_LOOP_tmp_or_19_cse <= and_dcpl_65 OR and_dcpl_195 OR and_dcpl_197 OR and_dcpl_198;
  nor_572_cse <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  or_2589_cse <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00"));
  COMP_LOOP_tmp_or_21_cse <= and_dcpl_189 OR and_dcpl_195 OR and_dcpl_197 OR and_dcpl_198;
  COMP_LOOP_tmp_COMP_LOOP_tmp_nor_14_cse <= NOT(CONV_SL_1_1(COMP_LOOP_13_tmp_mul_idiv_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  and_570_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"));
  or_2612_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_nor_16_rgt <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR nor_1798_tmp);
  COMP_LOOP_tmp_and_14_rgt <= CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND (NOT nor_1798_tmp);
  COMP_LOOP_tmp_and_15_rgt <= CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND (NOT nor_1798_tmp);
  COMP_LOOP_tmp_and_16_rgt <= CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (NOT nor_1798_tmp);
  mux_228_cse <= MUX_s_1_2_2((NOT (fsm_output(7))), (fsm_output(7)), fsm_output(6));
  or_2621_cse <= and_570_cse OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_464_cse <= MUX_s_1_2_2((NOT (fsm_output(8))), (fsm_output(8)), fsm_output(7));
  mux_559_cse <= MUX_s_1_2_2(mux_464_cse, and_733_cse, fsm_output(6));
  or_455_cse <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  or_454_cse <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"));
  or_2626_cse <= (CONV_SL_1_1(fsm_output(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111")))
      OR (fsm_output(6));
  and_655_cse <= (((fsm_output(6)) AND (fsm_output(1)) AND (fsm_output(2))) OR (fsm_output(7)))
      AND (fsm_output(8));
  COMP_LOOP_1_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 &
      STD_LOGIC_VECTOR'( "0000")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_1_acc_10_itm_10_1_1 <= COMP_LOOP_1_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_acc_13_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0(9
      DOWNTO 2)) + UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 & STD_LOGIC_VECTOR'( "01")),
      8));
  COMP_LOOP_acc_1_cse_4_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0)
      + UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 & STD_LOGIC_VECTOR'( "0011")), 10));
  COMP_LOOP_acc_1_cse_2_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0)
      + UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 & STD_LOGIC_VECTOR'( "0001")), 10));
  COMP_LOOP_2_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 &
      STD_LOGIC_VECTOR'( "0001")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_2_acc_10_itm_10_1_1 <= COMP_LOOP_2_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_3_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 &
      STD_LOGIC_VECTOR'( "0010")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_3_acc_10_itm_10_1_1 <= COMP_LOOP_3_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_4_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 &
      STD_LOGIC_VECTOR'( "0011")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_4_acc_10_itm_10_1_1 <= COMP_LOOP_4_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_5_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 &
      STD_LOGIC_VECTOR'( "0100")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_5_acc_10_itm_10_1_1 <= COMP_LOOP_5_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_6_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 &
      STD_LOGIC_VECTOR'( "0101")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_6_acc_10_itm_10_1_1 <= COMP_LOOP_6_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_7_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 &
      STD_LOGIC_VECTOR'( "0110")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_7_acc_10_itm_10_1_1 <= COMP_LOOP_7_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_8_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 &
      STD_LOGIC_VECTOR'( "0111")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_8_acc_10_itm_10_1_1 <= COMP_LOOP_8_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_9_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 &
      STD_LOGIC_VECTOR'( "1000")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_9_acc_10_itm_10_1_1 <= COMP_LOOP_9_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_10_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 &
      STD_LOGIC_VECTOR'( "1001")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_10_acc_10_itm_10_1_1 <= COMP_LOOP_10_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_11_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 &
      STD_LOGIC_VECTOR'( "1010")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_11_acc_10_itm_10_1_1 <= COMP_LOOP_11_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_12_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 &
      STD_LOGIC_VECTOR'( "1011")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_12_acc_10_itm_10_1_1 <= COMP_LOOP_12_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_13_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 &
      STD_LOGIC_VECTOR'( "1100")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_13_acc_10_itm_10_1_1 <= COMP_LOOP_13_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_14_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 &
      STD_LOGIC_VECTOR'( "1101")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_14_acc_10_itm_10_1_1 <= COMP_LOOP_14_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_15_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 &
      STD_LOGIC_VECTOR'( "1110")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_15_acc_10_itm_10_1_1 <= COMP_LOOP_15_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_16_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 &
      STD_LOGIC_VECTOR'( "1111")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_16_acc_10_itm_10_1_1 <= COMP_LOOP_16_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_k_10_4_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0),
      6), 7) + UNSIGNED'( "0000001"), 7));
  COMP_LOOP_tmp_mux1h_4_itm_mx0w3 <= MUX1HOT_v_64_16_2(twiddle_rsc_0_0_i_q_d, tmp_33_sva_1,
      tmp_33_sva_2, tmp_33_sva_3, tmp_33_sva_4, tmp_33_sva_5, tmp_33_sva_6, tmp_33_sva_7,
      tmp_33_sva_8, tmp_33_sva_9, tmp_33_sva_10, tmp_33_sva_11, tmp_33_sva_12, tmp_33_sva_13,
      tmp_33_sva_14, tmp_33_sva_15, STD_LOGIC_VECTOR'( COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_itm
      & COMP_LOOP_tmp_COMP_LOOP_tmp_and_167 & and_1191_cse & COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm
      & and_1190_cse & COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm & COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm
      & COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm & COMP_LOOP_tmp_COMP_LOOP_tmp_and_161
      & COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm & COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm
      & COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm & COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm
      & COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm & COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm
      & COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm));
  nor_1792_cse <= NOT(CONV_SL_1_1(COMP_LOOP_11_tmp_mul_idiv_sva(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  and_313_nl <= CONV_SL_1_1(COMP_LOOP_11_tmp_mul_idiv_sva(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10"));
  tmp_33_sva_13_mx0w1 <= MUX1HOT_v_64_3_2(twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_4_i_q_d,
      twiddle_rsc_0_8_i_q_d, STD_LOGIC_VECTOR'( nor_1792_cse & (COMP_LOOP_11_tmp_mul_idiv_sva(1))
      & and_313_nl));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_155 <= (COMP_LOOP_11_tmp_mul_idiv_sva(0)) AND nor_1792_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_157 <= CONV_SL_1_1(COMP_LOOP_11_tmp_mul_idiv_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("010"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_159 <= CONV_SL_1_1(COMP_LOOP_11_tmp_mul_idiv_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("100"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_161 <= (COMP_LOOP_10_tmp_mul_idiv_sva(3)) AND COMP_LOOP_tmp_nor_19_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_167 <= (COMP_LOOP_10_tmp_mul_idiv_sva(0)) AND COMP_LOOP_tmp_nor_13_itm;
  or_dcpl_5 <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm;
  and_dcpl_5 <= nor_1630_cse AND (NOT (fsm_output(6)));
  or_36_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000"));
  nor_tmp_10 <= (fsm_output(3)) AND (fsm_output(2)) AND (fsm_output(1)) AND (fsm_output(6));
  or_tmp_29 <= and_674_cse OR (fsm_output(6));
  nor_tmp_47 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11"));
  or_2732_cse <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  nor_tmp_115 <= or_2732_cse AND (fsm_output(8));
  mux_tmp_439 <= MUX_s_1_2_2((NOT (fsm_output(8))), (fsm_output(8)), or_2732_cse);
  mux_tmp_538 <= MUX_s_1_2_2(mux_tmp_439, nor_tmp_115, and_674_cse);
  or_610_cse <= (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_tmp_929 <= MUX_s_1_2_2((NOT and_675_cse), or_610_cse, fsm_output(3));
  nand_tmp_13 <= NOT((fsm_output(2)) AND (NOT mux_tmp_929));
  and_dcpl_45 <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_46 <= NOT((fsm_output(3)) OR (fsm_output(0)));
  and_dcpl_47 <= and_dcpl_46 AND and_dcpl_45;
  and_dcpl_48 <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_51 <= and_dcpl_5 AND and_dcpl_48;
  and_dcpl_53 <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_54 <= and_dcpl_46 AND and_dcpl_53;
  and_dcpl_55 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_57 <= and_733_cse AND (fsm_output(6));
  and_dcpl_58 <= and_dcpl_57 AND and_dcpl_55;
  nor_tmp_339 <= or_2259_cse_1 AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111"));
  and_565_nl <= (fsm_output(2)) AND (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(7))
      AND (fsm_output(8));
  mux_1080_nl <= MUX_s_1_2_2(and_565_nl, and_dcpl_57, fsm_output(3));
  mux_tmp_1062 <= MUX_s_1_2_2(mux_1080_nl, nor_tmp_339, fsm_output(0));
  or_714_nl <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (NOT((fsm_output(1)) AND
      (fsm_output(6))));
  mux_1083_nl <= MUX_s_1_2_2((fsm_output(6)), (NOT (fsm_output(6))), fsm_output(1));
  nand_22_nl <= NOT((fsm_output(4)) AND (fsm_output(0)) AND mux_1083_nl);
  mux_tmp_1065 <= MUX_s_1_2_2(or_714_nl, nand_22_nl, fsm_output(5));
  nand_23_nl <= NOT((fsm_output(7)) AND (NOT mux_tmp_1065));
  or_712_nl <= (fsm_output(5)) OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(1))
      OR (fsm_output(6));
  mux_1085_nl <= MUX_s_1_2_2(mux_tmp_1065, or_712_nl, fsm_output(7));
  mux_tmp_1067 <= MUX_s_1_2_2(nand_23_nl, mux_1085_nl, fsm_output(2));
  and_dcpl_60 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_61 <= and_dcpl_5 AND and_dcpl_60;
  and_dcpl_62 <= and_dcpl_61 AND and_dcpl_47;
  and_dcpl_63 <= (NOT (fsm_output(3))) AND (fsm_output(0));
  and_dcpl_64 <= and_dcpl_63 AND and_dcpl_45;
  and_dcpl_65 <= and_dcpl_61 AND and_dcpl_64;
  and_dcpl_66 <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_67 <= and_dcpl_63 AND and_dcpl_66;
  and_dcpl_69 <= and_dcpl_46 AND and_dcpl_66;
  and_dcpl_70 <= and_dcpl_61 AND and_dcpl_69;
  and_dcpl_71 <= nor_1630_cse AND (fsm_output(6));
  and_dcpl_72 <= and_dcpl_71 AND and_dcpl_48;
  and_dcpl_74 <= and_dcpl_72 AND and_dcpl_64;
  and_dcpl_75 <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_77 <= and_712_cse AND and_dcpl_75;
  and_dcpl_79 <= and_dcpl_71 AND and_674_cse;
  and_dcpl_81 <= and_dcpl_72 AND and_dcpl_69;
  and_dcpl_82 <= (fsm_output(3)) AND (NOT (fsm_output(0)));
  and_dcpl_83 <= and_dcpl_82 AND and_dcpl_53;
  and_dcpl_85 <= and_712_cse AND and_dcpl_53;
  and_dcpl_86 <= and_dcpl_79 AND and_dcpl_85;
  and_dcpl_87 <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_88 <= and_dcpl_87 AND (NOT (fsm_output(6)));
  and_dcpl_89 <= and_dcpl_88 AND and_dcpl_55;
  and_dcpl_91 <= and_dcpl_82 AND and_dcpl_75;
  and_dcpl_92 <= and_dcpl_88 AND and_674_cse;
  and_dcpl_93 <= and_dcpl_92 AND and_dcpl_91;
  and_dcpl_95 <= and_dcpl_89 AND and_dcpl_85;
  and_dcpl_96 <= and_dcpl_87 AND (fsm_output(6));
  and_dcpl_97 <= and_dcpl_96 AND and_dcpl_60;
  and_dcpl_99 <= and_dcpl_96 AND and_dcpl_55;
  and_dcpl_100 <= and_dcpl_99 AND and_dcpl_91;
  and_dcpl_102 <= and_dcpl_97 AND and_dcpl_85;
  and_dcpl_103 <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_104 <= and_dcpl_103 AND (NOT (fsm_output(6)));
  and_dcpl_105 <= and_dcpl_104 AND and_dcpl_48;
  and_dcpl_107 <= and_dcpl_104 AND and_dcpl_60;
  and_dcpl_108 <= and_dcpl_107 AND and_dcpl_91;
  and_dcpl_110 <= and_dcpl_105 AND and_dcpl_85;
  and_dcpl_111 <= and_dcpl_63 AND and_dcpl_75;
  and_dcpl_112 <= and_dcpl_103 AND (fsm_output(6));
  and_dcpl_113 <= and_dcpl_112 AND and_674_cse;
  and_dcpl_115 <= and_dcpl_112 AND and_dcpl_48;
  and_dcpl_116 <= and_dcpl_115 AND and_dcpl_91;
  and_dcpl_118 <= and_dcpl_63 AND and_dcpl_53;
  and_dcpl_119 <= and_dcpl_113 AND and_dcpl_118;
  and_dcpl_120 <= and_733_cse AND (NOT (fsm_output(6)));
  and_dcpl_121 <= and_dcpl_120 AND and_dcpl_55;
  and_dcpl_123 <= and_dcpl_46 AND and_dcpl_75;
  and_dcpl_124 <= and_dcpl_120 AND and_674_cse;
  and_dcpl_125 <= and_dcpl_124 AND and_dcpl_123;
  and_dcpl_127 <= and_dcpl_121 AND and_dcpl_118;
  and_dcpl_128 <= and_dcpl_57 AND and_dcpl_60;
  and_dcpl_130 <= and_dcpl_58 AND and_dcpl_123;
  and_dcpl_131 <= and_dcpl_5 AND and_674_cse;
  and_dcpl_136 <= and_dcpl_71 AND and_dcpl_55;
  and_dcpl_141 <= and_dcpl_88 AND and_dcpl_60;
  and_dcpl_146 <= and_dcpl_96 AND and_dcpl_48;
  and_dcpl_151 <= and_dcpl_104 AND and_674_cse;
  and_dcpl_156 <= and_dcpl_112 AND and_dcpl_55;
  and_dcpl_161 <= and_dcpl_120 AND and_dcpl_60;
  and_dcpl_166 <= and_dcpl_57 AND and_dcpl_48;
  not_tmp_395 <= NOT((fsm_output(6)) AND (fsm_output(8)));
  or_762_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT
      (fsm_output(8)));
  or_760_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR (VEC_LOOP_j_10_0_sva_9_0(2)) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("100"));
  or_758_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010"));
  mux_1115_nl <= MUX_s_1_2_2(or_760_nl, or_758_nl, fsm_output(2));
  mux_1116_cse <= MUX_s_1_2_2(or_762_nl, mux_1115_nl, fsm_output(3));
  not_tmp_399 <= NOT((fsm_output(4)) AND (fsm_output(8)));
  nor_1479_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT
      (fsm_output(8))));
  nor_1480_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) OR (VEC_LOOP_j_10_0_sva_9_0(2))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1481_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  mux_1240_nl <= MUX_s_1_2_2(nor_1480_nl, nor_1481_nl, fsm_output(2));
  mux_1241_cse <= MUX_s_1_2_2(nor_1479_nl, mux_1240_nl, fsm_output(3));
  nand_268_cse <= NOT((COMP_LOOP_acc_10_cse_10_1_15_sva(1)) AND CONV_SL_1_1(fsm_output(8
      DOWNTO 6)=STD_LOGIC_VECTOR'("111")));
  nand_261_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111")));
  or_1150_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT
      (fsm_output(8)));
  or_1148_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100"));
  or_1146_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010"));
  mux_1365_nl <= MUX_s_1_2_2(or_1148_nl, or_1146_nl, fsm_output(2));
  mux_1366_cse <= MUX_s_1_2_2(or_1150_nl, mux_1365_nl, fsm_output(3));
  nor_1242_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT
      (fsm_output(8))));
  nor_1243_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1244_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  mux_1490_nl <= MUX_s_1_2_2(nor_1243_nl, nor_1244_nl, fsm_output(2));
  mux_1491_cse <= MUX_s_1_2_2(nor_1242_nl, mux_1490_nl, fsm_output(3));
  or_1538_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT
      (fsm_output(8)));
  or_1536_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR (VEC_LOOP_j_10_0_sva_9_0(2))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100"));
  or_1534_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010"));
  mux_1615_nl <= MUX_s_1_2_2(or_1536_nl, or_1534_nl, fsm_output(2));
  mux_1616_cse <= MUX_s_1_2_2(or_1538_nl, mux_1615_nl, fsm_output(3));
  nand_222_cse <= NOT((COMP_LOOP_acc_20_psp_sva(2)) AND CONV_SL_1_1(fsm_output(8
      DOWNTO 6)=STD_LOGIC_VECTOR'("111")));
  nand_223_cse <= NOT((COMP_LOOP_acc_10_cse_10_1_sva(3)) AND CONV_SL_1_1(fsm_output(8
      DOWNTO 6)=STD_LOGIC_VECTOR'("111")));
  nor_1012_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT
      (fsm_output(8))));
  nor_1013_nl <= NOT((NOT (COMP_LOOP_acc_16_psp_sva(0))) OR (VEC_LOOP_j_10_0_sva_9_0(2))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1014_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  mux_1740_nl <= MUX_s_1_2_2(nor_1013_nl, nor_1014_nl, fsm_output(2));
  mux_1741_cse <= MUX_s_1_2_2(nor_1012_nl, mux_1740_nl, fsm_output(3));
  nand_322_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (NOT (fsm_output(6))) AND (fsm_output(8)));
  or_1922_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100"));
  or_1920_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010"));
  mux_1865_nl <= MUX_s_1_2_2(or_1922_nl, or_1920_nl, fsm_output(2));
  mux_1866_cse <= MUX_s_1_2_2(nand_322_nl, mux_1865_nl, fsm_output(3));
  nand_184_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111")));
  nand_185_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111")));
  and_835_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (NOT (fsm_output(6))) AND (fsm_output(8));
  nor_795_nl <= NOT((NOT (COMP_LOOP_acc_16_psp_sva(0))) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_796_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  mux_1990_nl <= MUX_s_1_2_2(nor_795_nl, nor_796_nl, fsm_output(2));
  mux_1991_cse <= MUX_s_1_2_2(and_835_nl, mux_1990_nl, fsm_output(3));
  nand_157_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (NOT (fsm_output(7))));
  and_dcpl_171 <= (fsm_output(0)) AND (NOT (fsm_output(5)));
  and_dcpl_175 <= (or_36_cse XOR (fsm_output(4))) AND (NOT (fsm_output(8))) AND nor_572_cse
      AND and_dcpl_171;
  and_dcpl_180 <= (or_2259_cse_1 XOR (fsm_output(4))) AND nor_1630_cse AND (NOT (fsm_output(6)))
      AND (NOT (fsm_output(1))) AND nor_1767_cse;
  and_dcpl_181 <= and_dcpl_131 AND and_dcpl_47;
  and_dcpl_182 <= and_dcpl_82 AND and_dcpl_45;
  and_dcpl_183 <= and_dcpl_61 AND and_dcpl_182;
  and_dcpl_184 <= and_dcpl_131 AND and_dcpl_182;
  and_dcpl_186 <= nor_1630_cse AND CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("00"));
  or_tmp_2077 <= (fsm_output(4)) OR CONV_SL_1_1(COMP_LOOP_10_tmp_mul_idiv_sva(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0000"));
  and_dcpl_188 <= and_dcpl_5 AND and_dcpl_55;
  and_dcpl_189 <= and_dcpl_188 AND and_dcpl_47;
  and_dcpl_190 <= and_dcpl_51 AND and_dcpl_182;
  and_dcpl_191 <= and_dcpl_188 AND and_dcpl_182;
  and_dcpl_192 <= and_dcpl_51 AND and_dcpl_123;
  and_dcpl_193 <= and_dcpl_5 AND nor_1767_cse;
  and_dcpl_195 <= and_dcpl_131 AND and_dcpl_64;
  and_dcpl_196 <= and_712_cse AND and_dcpl_45;
  and_dcpl_197 <= and_dcpl_61 AND and_dcpl_196;
  and_dcpl_198 <= and_dcpl_131 AND and_dcpl_196;
  and_dcpl_202 <= and_dcpl_188 AND and_dcpl_196;
  and_dcpl_207 <= and_dcpl_51 AND and_dcpl_196;
  or_2430_nl <= (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(8));
  mux_tmp_2224 <= MUX_s_1_2_2(or_2430_nl, mux_tmp_929, fsm_output(2));
  mux_tmp_2225 <= MUX_s_1_2_2(mux_tmp_2224, or_611_cse, fsm_output(7));
  mux_tmp_2229 <= MUX_s_1_2_2(mux_952_cse, mux_tmp_2225, fsm_output(0));
  or_tmp_2258 <= (fsm_output(8)) OR (fsm_output(0)) OR (fsm_output(5));
  or_2434_nl <= (NOT (fsm_output(8))) OR (fsm_output(0)) OR (fsm_output(5));
  mux_tmp_2237 <= MUX_s_1_2_2(or_2434_nl, or_tmp_2258, fsm_output(3));
  not_tmp_676 <= NOT((fsm_output(0)) AND (fsm_output(5)));
  nor_tmp_480 <= (fsm_output(8)) AND (fsm_output(0)) AND (fsm_output(5));
  or_2435_nl <= (fsm_output(8)) OR not_tmp_676;
  mux_tmp_2238 <= MUX_s_1_2_2((NOT nor_tmp_480), or_2435_nl, fsm_output(3));
  or_tmp_2266 <= (NOT (fsm_output(3))) OR (NOT (fsm_output(8))) OR (fsm_output(0))
      OR (fsm_output(5));
  mux_2263_nl <= MUX_s_1_2_2((NOT (fsm_output(5))), (fsm_output(5)), fsm_output(0));
  or_2443_nl <= (fsm_output(3)) OR (fsm_output(8)) OR mux_2263_nl;
  mux_tmp_2245 <= MUX_s_1_2_2(or_2443_nl, or_tmp_2266, fsm_output(4));
  or_2444_nl <= (fsm_output(6)) OR mux_tmp_2245;
  or_2440_nl <= (NOT (fsm_output(6))) OR (fsm_output(4)) OR mux_tmp_2238;
  mux_tmp_2246 <= MUX_s_1_2_2(or_2444_nl, or_2440_nl, fsm_output(1));
  mux_2267_nl <= MUX_s_1_2_2((NOT or_tmp_2258), nor_tmp_480, fsm_output(3));
  mux_tmp_2249 <= MUX_s_1_2_2((NOT or_tmp_2266), mux_2267_nl, fsm_output(4));
  and_dcpl_220 <= and_dcpl_61 AND and_dcpl_67;
  and_dcpl_222 <= and_dcpl_71 AND and_dcpl_60 AND and_dcpl_47;
  and_dcpl_223 <= and_dcpl_72 AND and_dcpl_67;
  and_dcpl_225 <= and_dcpl_88 AND and_dcpl_48 AND and_dcpl_47;
  and_dcpl_226 <= and_dcpl_92 AND and_dcpl_77;
  and_dcpl_227 <= and_dcpl_92 AND and_dcpl_83;
  and_dcpl_228 <= and_dcpl_99 AND and_dcpl_77;
  and_dcpl_229 <= and_dcpl_99 AND and_dcpl_83;
  and_dcpl_230 <= and_dcpl_107 AND and_dcpl_77;
  and_dcpl_231 <= and_dcpl_107 AND and_dcpl_83;
  and_dcpl_232 <= and_dcpl_115 AND and_dcpl_77;
  and_dcpl_233 <= and_dcpl_115 AND and_dcpl_83;
  and_dcpl_234 <= and_dcpl_124 AND and_dcpl_111;
  and_dcpl_235 <= and_dcpl_124 AND and_dcpl_54;
  and_dcpl_236 <= and_dcpl_58 AND and_dcpl_111;
  or_tmp_2274 <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"));
  mux_tmp_2256 <= MUX_s_1_2_2(or_tmp_2274, or_454_cse, fsm_output(2));
  nand_114_nl <= NOT((fsm_output(2)) AND (fsm_output(7)) AND (fsm_output(8)));
  mux_tmp_2257 <= MUX_s_1_2_2(nand_114_nl, mux_tmp_2256, fsm_output(3));
  mux_tmp_2258 <= MUX_s_1_2_2(or_454_cse, or_455_cse, fsm_output(2));
  nand_113_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11")));
  mux_tmp_2259 <= MUX_s_1_2_2(nand_113_nl, or_tmp_2274, fsm_output(2));
  or_tmp_2277 <= (fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(8));
  or_tmp_2279 <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(8));
  or_2455_nl <= (fsm_output(0)) OR mux_tmp_2257;
  mux_tmp_2264 <= MUX_s_1_2_2(or_2455_nl, or_tmp_2279, fsm_output(5));
  or_dcpl_182 <= or_455_cse OR (fsm_output(6));
  or_dcpl_183 <= or_dcpl_182 OR CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01"));
  or_dcpl_184 <= or_dcpl_183 OR (fsm_output(3)) OR (fsm_output(0)) OR or_2589_cse;
  or_2482_nl <= (fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(7))
      OR (fsm_output(8));
  or_2481_nl <= (fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(6))
      OR (fsm_output(7)) OR (fsm_output(8));
  mux_tmp_2282 <= MUX_s_1_2_2(or_2482_nl, or_2481_nl, fsm_output(0));
  mux_2302_nl <= MUX_s_1_2_2((NOT mux_tmp_2282), nor_tmp_339, fsm_output(4));
  mux_2303_itm <= MUX_s_1_2_2(mux_2302_nl, and_dcpl_57, fsm_output(5));
  nor_tmp_489 <= (and_570_cse OR (fsm_output(6))) AND (fsm_output(7));
  mux_2306_nl <= MUX_s_1_2_2(mux_228_cse, nor_tmp_47, or_2259_cse_1);
  mux_2305_nl <= MUX_s_1_2_2(mux_228_cse, nor_tmp_47, or_36_cse);
  mux_tmp_2288 <= MUX_s_1_2_2(mux_2306_nl, mux_2305_nl, fsm_output(0));
  and_416_nl <= (fsm_output(3)) AND (fsm_output(2)) AND (fsm_output(6));
  mux_tmp_2291 <= MUX_s_1_2_2(nor_tmp_10, and_416_nl, fsm_output(0));
  or_2487_cse <= (fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(6));
  or_2486_cse <= (fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(6));
  mux_tmp_2292 <= MUX_s_1_2_2(or_2487_cse, or_2486_cse, fsm_output(0));
  not_tmp_703 <= NOT((fsm_output(4)) OR mux_tmp_2292);
  mux_22_nl <= MUX_s_1_2_2(or_2259_cse_1, or_36_cse, fsm_output(0));
  or_tmp_2300 <= (fsm_output(4)) OR mux_22_nl;
  or_dcpl_190 <= CONV_SL_1_1(fsm_output(5 DOWNTO 3)/=STD_LOGIC_VECTOR'("000"));
  and_dcpl_248 <= (or_tmp_2300 XOR (fsm_output(5))) AND and_dcpl_5;
  or_2497_nl <= (fsm_output(1)) OR (NOT (fsm_output(6)));
  mux_2323_nl <= MUX_s_1_2_2(or_2497_nl, (fsm_output(6)), or_2259_cse_1);
  mux_61_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), (fsm_output(6)), or_36_cse);
  mux_2324_nl <= MUX_s_1_2_2(mux_2323_nl, mux_61_nl, fsm_output(0));
  mux_2325_nl <= MUX_s_1_2_2(mux_2324_nl, (fsm_output(6)), or_2589_cse);
  and_dcpl_252 <= (NOT mux_2325_nl) AND nor_1630_cse;
  and_411_nl <= (CONV_SL_1_1(fsm_output(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")))
      AND (fsm_output(6));
  mux_2328_nl <= MUX_s_1_2_2(not_tmp_703, and_411_nl, fsm_output(5));
  and_dcpl_255 <= (NOT mux_2328_nl) AND nor_1630_cse;
  nor_tmp_499 <= ((fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(6))) AND (fsm_output(7));
  mux_2329_nl <= MUX_s_1_2_2(nor_tmp_47, nor_tmp_499, fsm_output(3));
  mux_tmp_2311 <= MUX_s_1_2_2(nor_tmp_489, mux_2329_nl, fsm_output(0));
  and_dcpl_258 <= (or_2697_cse OR and_1189_cse OR or_dcpl_190) AND nor_1630_cse;
  mux_tmp_2318 <= MUX_s_1_2_2(mux_tmp_2288, nor_tmp_47, fsm_output(4));
  and_403_nl <= or_2626_cse AND (fsm_output(7));
  mux_2342_nl <= MUX_s_1_2_2(mux_tmp_2288, and_403_nl, fsm_output(4));
  mux_2343_nl <= MUX_s_1_2_2(mux_2342_nl, (fsm_output(7)), fsm_output(5));
  and_dcpl_262 <= NOT(mux_2343_nl OR (fsm_output(8)));
  nor_tmp_507 <= or_432_cse AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11"));
  and_tmp_28 <= (fsm_output(3)) AND nor_tmp_507;
  or_2507_nl <= (fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(7));
  or_2506_nl <= (fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(6))
      OR (fsm_output(7));
  mux_tmp_2325 <= MUX_s_1_2_2(or_2507_nl, or_2506_nl, fsm_output(0));
  and_401_nl <= (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(7));
  mux_tmp_2328 <= MUX_s_1_2_2(and_tmp_28, and_401_nl, fsm_output(0));
  nor_tmp_509 <= (fsm_output(3)) AND (fsm_output(2)) AND (fsm_output(6)) AND (fsm_output(7));
  and_398_nl <= ((CONV_SL_1_1(fsm_output(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1111")))
      OR (fsm_output(6))) AND (fsm_output(7));
  mux_2353_nl <= MUX_s_1_2_2(mux_tmp_2318, and_398_nl, fsm_output(5));
  and_dcpl_266 <= NOT(mux_2353_nl OR (fsm_output(8)));
  not_tmp_727 <= NOT((fsm_output(4)) OR mux_tmp_2325);
  and_396_nl <= (fsm_output(3)) AND (fsm_output(2)) AND (fsm_output(1)) AND (fsm_output(6))
      AND (fsm_output(7));
  mux_2357_nl <= MUX_s_1_2_2(and_396_nl, nor_tmp_509, fsm_output(0));
  mux_2358_nl <= MUX_s_1_2_2((NOT mux_tmp_2325), mux_2357_nl, fsm_output(4));
  mux_2359_nl <= MUX_s_1_2_2(mux_2358_nl, nor_tmp_47, fsm_output(5));
  and_dcpl_270 <= NOT(mux_2359_nl OR (fsm_output(8)));
  nor_tmp_515 <= ((fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(7))) AND (fsm_output(8));
  mux_2362_nl <= MUX_s_1_2_2(mux_tmp_439, nor_tmp_115, or_2259_cse_1);
  mux_2361_nl <= MUX_s_1_2_2(mux_tmp_439, nor_tmp_115, or_36_cse);
  mux_tmp_2344 <= MUX_s_1_2_2(mux_2362_nl, mux_2361_nl, fsm_output(0));
  and_566_nl <= (and_674_cse OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")))
      AND (fsm_output(8));
  mux_tmp_2347 <= MUX_s_1_2_2(and_566_nl, (fsm_output(8)), fsm_output(3));
  mux_tmp_2348 <= MUX_s_1_2_2(nor_tmp_515, mux_tmp_2347, fsm_output(0));
  mux_tmp_2351 <= MUX_s_1_2_2(nor_tmp_115, and_728_cse, fsm_output(3));
  and_392_nl <= (fsm_output(4)) AND (fsm_output(3)) AND (fsm_output(2)) AND (fsm_output(6))
      AND (fsm_output(7));
  mux_2374_nl <= MUX_s_1_2_2(not_tmp_727, and_392_nl, fsm_output(5));
  and_dcpl_271 <= NOT(mux_2374_nl OR (fsm_output(8)));
  mux_tmp_2357 <= MUX_s_1_2_2(mux_tmp_2344, nor_tmp_115, fsm_output(4));
  and_388_nl <= or_2621_cse AND (fsm_output(8));
  mux_2381_nl <= MUX_s_1_2_2(and_388_nl, mux_tmp_2351, fsm_output(0));
  mux_2382_nl <= MUX_s_1_2_2(mux_tmp_2344, mux_2381_nl, fsm_output(4));
  mux_2383_itm <= MUX_s_1_2_2(mux_2382_nl, (fsm_output(8)), fsm_output(5));
  mux_tmp_2365 <= MUX_s_1_2_2(and_655_cse, nor_tmp_115, fsm_output(3));
  mux_2387_nl <= MUX_s_1_2_2(mux_464_cse, and_733_cse, or_2487_cse);
  mux_2386_nl <= MUX_s_1_2_2(mux_464_cse, and_733_cse, or_2486_cse);
  mux_tmp_2369 <= MUX_s_1_2_2(mux_2387_nl, mux_2386_nl, fsm_output(0));
  nor_tmp_528 <= ((or_2259_cse_1 AND (fsm_output(6))) OR (fsm_output(7))) AND (fsm_output(8));
  nor_tmp_530 <= (((fsm_output(3)) AND (fsm_output(6))) OR (fsm_output(7))) AND (fsm_output(8));
  mux_2397_nl <= MUX_s_1_2_2(nor_tmp_115, and_728_cse, and_407_cse);
  mux_2398_itm <= MUX_s_1_2_2(mux_tmp_2357, mux_2397_nl, fsm_output(5));
  mux_tmp_2384 <= MUX_s_1_2_2(mux_tmp_2369, and_733_cse, fsm_output(4));
  and_376_nl <= ((or_432_cse AND (fsm_output(6))) OR (fsm_output(7))) AND (fsm_output(8));
  mux_2407_nl <= MUX_s_1_2_2(and_733_cse, and_376_nl, fsm_output(3));
  mux_2408_nl <= MUX_s_1_2_2(mux_2407_nl, nor_tmp_530, fsm_output(0));
  mux_2409_nl <= MUX_s_1_2_2(mux_tmp_2369, mux_2408_nl, fsm_output(4));
  mux_2410_itm <= MUX_s_1_2_2(mux_2409_nl, nor_tmp_115, fsm_output(5));
  nor_tmp_537 <= or_2487_cse AND CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11"));
  mux_tmp_2392 <= MUX_s_1_2_2(nor_1630_cse, and_733_cse, fsm_output(6));
  mux_2413_nl <= MUX_s_1_2_2(mux_tmp_2392, and_dcpl_57, or_2259_cse_1);
  mux_2412_nl <= MUX_s_1_2_2(mux_tmp_2392, and_dcpl_57, or_36_cse);
  mux_tmp_2395 <= MUX_s_1_2_2(mux_2413_nl, mux_2412_nl, fsm_output(0));
  nor_tmp_538 <= or_2486_cse AND CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11"));
  and_372_nl <= or_tmp_29 AND CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11"));
  mux_tmp_2401 <= MUX_s_1_2_2(and_372_nl, and_733_cse, fsm_output(3));
  and_370_nl <= (((fsm_output(3)) AND (fsm_output(4)) AND (fsm_output(6))) OR (fsm_output(7)))
      AND (fsm_output(8));
  mux_2424_itm <= MUX_s_1_2_2(mux_tmp_2384, and_370_nl, fsm_output(5));
  nor_tmp_544 <= (fsm_output(4)) AND (fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(8));
  mux_tmp_2410 <= MUX_s_1_2_2(mux_tmp_2395, and_dcpl_57, fsm_output(4));
  or_2635_cse <= (fsm_output(3)) OR (fsm_output(6));
  and_366_nl <= or_2635_cse AND CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11"));
  mux_2433_nl <= MUX_s_1_2_2(and_366_nl, mux_tmp_2401, fsm_output(0));
  mux_2434_nl <= MUX_s_1_2_2(mux_tmp_2395, mux_2433_nl, fsm_output(4));
  mux_2435_itm <= MUX_s_1_2_2(mux_2434_nl, and_733_cse, fsm_output(5));
  nor_tmp_547 <= or_36_cse AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111"));
  nor_tmp_548 <= or_2612_cse AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111"));
  mux_2440_nl <= MUX_s_1_2_2(nor_tmp_339, nor_tmp_547, fsm_output(0));
  mux_2441_nl <= MUX_s_1_2_2((NOT mux_tmp_2282), mux_2440_nl, fsm_output(4));
  mux_2442_itm <= MUX_s_1_2_2(mux_2441_nl, and_dcpl_57, fsm_output(5));
  mux_2443_nl <= MUX_s_1_2_2(and_dcpl_57, mux_tmp_2401, fsm_output(4));
  mux_2444_itm <= MUX_s_1_2_2(mux_tmp_2410, mux_2443_nl, fsm_output(5));
  not_tmp_762 <= NOT((fsm_output(4)) OR mux_tmp_2282);
  mux_2448_nl <= MUX_s_1_2_2((NOT mux_tmp_2282), mux_tmp_1062, fsm_output(4));
  mux_2449_itm <= MUX_s_1_2_2(mux_2448_nl, and_dcpl_57, fsm_output(5));
  or_dcpl_207 <= (fsm_output(3)) OR (NOT (fsm_output(0))) OR or_2589_cse;
  and_dcpl_277 <= nor_1630_cse AND (NOT (fsm_output(6))) AND (fsm_output(1)) AND
      (fsm_output(2)) AND (NOT (fsm_output(0))) AND and_dcpl_45;
  or_tmp_2358 <= (NOT (fsm_output(8))) OR (fsm_output(4));
  or_427_nl <= (fsm_output(4)) OR (fsm_output(8));
  mux_tmp_2447 <= MUX_s_1_2_2(or_tmp_2358, or_427_nl, fsm_output(3));
  nand_tmp_100 <= NOT((fsm_output(7)) AND (NOT mux_tmp_2447));
  mux_2468_nl <= MUX_s_1_2_2(or_610_cse, or_tmp_2358, fsm_output(3));
  or_2571_nl <= (fsm_output(7)) OR mux_2468_nl;
  mux_tmp_2450 <= MUX_s_1_2_2(or_2571_nl, nand_tmp_100, fsm_output(2));
  or_tmp_2362 <= (fsm_output(6)) OR mux_tmp_2450;
  and_dcpl_286 <= and_dcpl_82 AND and_dcpl_66;
  or_tmp_2384 <= (fsm_output(3)) OR or_tmp_29;
  STAGE_LOOP_i_3_0_sva_mx0c1 <= and_dcpl_58 AND and_dcpl_54;
  VEC_LOOP_j_10_0_sva_9_0_mx0c0 <= and_dcpl_51 AND and_dcpl_64;
  and_361_nl <= (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(7)) AND (fsm_output(8));
  nor_577_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(8)));
  mux_2465_cse <= MUX_s_1_2_2(and_361_nl, nor_577_nl, fsm_output(4));
  COMP_LOOP_10_acc_8_itm_mx0c2 <= mux_2465_cse AND nor_1624_cse AND and_dcpl_171;
  nand_103_nl <= NOT((fsm_output(6)) AND (NOT mux_tmp_2450));
  mux_2471_nl <= MUX_s_1_2_2(nand_103_nl, or_tmp_2362, fsm_output(1));
  nor_576_nl <= NOT((fsm_output(5)) OR mux_2471_nl);
  or_2569_nl <= (fsm_output(7)) OR mux_tmp_2447;
  mux_2467_nl <= MUX_s_1_2_2(nand_tmp_100, or_2569_nl, fsm_output(2));
  nand_101_nl <= NOT((fsm_output(6)) AND (NOT mux_2467_nl));
  mux_2470_nl <= MUX_s_1_2_2(or_tmp_2362, nand_101_nl, fsm_output(1));
  and_360_nl <= (fsm_output(5)) AND (NOT mux_2470_nl);
  COMP_LOOP_10_acc_8_itm_mx0c3 <= MUX_s_1_2_2(nor_576_nl, and_360_nl, fsm_output(0));
  COMP_LOOP_10_acc_8_itm_mx0c6 <= and_dcpl_51 AND and_dcpl_54;
  COMP_LOOP_10_acc_8_itm_mx0c9 <= and_dcpl_79 AND and_dcpl_196;
  COMP_LOOP_10_acc_8_itm_mx0c12 <= and_dcpl_79 AND and_dcpl_286;
  COMP_LOOP_10_acc_8_itm_mx0c15 <= and_dcpl_89 AND and_dcpl_196;
  COMP_LOOP_10_acc_8_itm_mx0c18 <= and_dcpl_89 AND and_dcpl_286;
  COMP_LOOP_10_acc_8_itm_mx0c21 <= and_dcpl_97 AND and_dcpl_196;
  COMP_LOOP_10_acc_8_itm_mx0c24 <= and_dcpl_97 AND and_dcpl_286;
  COMP_LOOP_10_acc_8_itm_mx0c27 <= and_dcpl_105 AND and_dcpl_196;
  COMP_LOOP_10_acc_8_itm_mx0c30 <= and_dcpl_105 AND and_dcpl_286;
  COMP_LOOP_10_acc_8_itm_mx0c33 <= and_dcpl_113 AND and_dcpl_64;
  COMP_LOOP_10_acc_8_itm_mx0c36 <= and_dcpl_113 AND and_dcpl_69;
  COMP_LOOP_10_acc_8_itm_mx0c39 <= and_dcpl_121 AND and_dcpl_64;
  COMP_LOOP_10_acc_8_itm_mx0c42 <= and_dcpl_121 AND and_dcpl_69;
  COMP_LOOP_10_acc_8_itm_mx0c47 <= and_dcpl_128 AND and_dcpl_69;
  STAGE_LOOP_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT z_out_4)) +
      SIGNED'( "00001"), 5));
  STAGE_LOOP_acc_itm_4_1 <= STAGE_LOOP_acc_nl(4);
  or_44_nl <= (fsm_output(3)) OR and_674_cse;
  mux_27_nl <= MUX_s_1_2_2(or_44_nl, or_2259_cse_1, fsm_output(0));
  nor_575_nl <= NOT((fsm_output(4)) OR mux_27_nl);
  mux_2498_nl <= MUX_s_1_2_2(nor_575_nl, (fsm_output(4)), fsm_output(5));
  and_332_tmp <= (NOT mux_2498_nl) AND and_dcpl_5;
  nand_107_nl <= NOT((fsm_output(2)) AND (fsm_output(1)) AND (fsm_output(6)));
  mux_2507_nl <= MUX_s_1_2_2(or_tmp_29, nand_107_nl, fsm_output(3));
  mux_2508_nl <= MUX_s_1_2_2(or_tmp_2384, mux_2507_nl, fsm_output(0));
  mux_2509_nl <= MUX_s_1_2_2(mux_2508_nl, (NOT (fsm_output(6))), or_2589_cse);
  and_341_tmp <= mux_2509_nl AND nor_1630_cse;
  mux_2511_nl <= MUX_s_1_2_2(or_2635_cse, or_tmp_2384, fsm_output(0));
  nor_570_nl <= NOT((fsm_output(4)) OR mux_2511_nl);
  mux_2510_nl <= MUX_s_1_2_2(nor_tmp_10, (fsm_output(6)), fsm_output(4));
  mux_2512_nl <= MUX_s_1_2_2(nor_570_nl, mux_2510_nl, fsm_output(5));
  and_342_tmp <= (NOT mux_2512_nl) AND nor_1630_cse;
  and_354_nl <= or_tmp_29 AND (fsm_output(7));
  mux_2523_nl <= MUX_s_1_2_2(mux_228_cse, and_354_nl, fsm_output(3));
  and_356_nl <= or_2697_cse AND (fsm_output(7));
  mux_2522_nl <= MUX_s_1_2_2(mux_228_cse, and_356_nl, fsm_output(3));
  mux_2524_nl <= MUX_s_1_2_2(mux_2523_nl, mux_2522_nl, fsm_output(0));
  mux_2525_nl <= MUX_s_1_2_2(mux_2524_nl, (fsm_output(7)), or_2589_cse);
  nor_1798_tmp <= NOT(mux_2525_nl OR (fsm_output(8)));
  nor_1750_nl <= NOT((fsm_output(6)) OR (fsm_output(1)) OR (fsm_output(7)));
  mux_234_nl <= MUX_s_1_2_2(nor_1750_nl, nor_tmp_47, fsm_output(2));
  mux_2536_nl <= MUX_s_1_2_2(nor_572_cse, mux_234_nl, fsm_output(3));
  mux_232_nl <= MUX_s_1_2_2(nor_572_cse, nor_tmp_47, or_432_cse);
  mux_233_nl <= MUX_s_1_2_2(nor_572_cse, mux_232_nl, fsm_output(3));
  mux_2537_nl <= MUX_s_1_2_2(mux_2536_nl, mux_233_nl, fsm_output(0));
  mux_2538_nl <= MUX_s_1_2_2(mux_2537_nl, nor_tmp_47, or_2589_cse);
  nor_1796_tmp <= NOT(mux_2538_nl OR (fsm_output(8)));
  or_715_nl <= (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(5))) OR (fsm_output(4))
      OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(6));
  mux_1088_nl <= MUX_s_1_2_2(or_715_nl, mux_tmp_1067, fsm_output(8));
  or_711_nl <= (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(5)) OR (NOT (fsm_output(4)))
      OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(6));
  mux_1087_nl <= MUX_s_1_2_2(mux_tmp_1067, or_711_nl, fsm_output(8));
  mux_1089_nl <= MUX_s_1_2_2(mux_1088_nl, mux_1087_nl, fsm_output(3));
  vec_rsc_0_0_i_d_d_pff <= MUX_v_64_2_2(COMP_LOOP_10_acc_8_itm, COMP_LOOP_1_modulo_cmp_return_rsc_z,
      mux_1089_nl);
  and_94_nl <= and_dcpl_51 AND and_dcpl_67;
  and_99_nl <= and_dcpl_72 AND and_dcpl_47;
  and_106_nl <= and_dcpl_79 AND and_dcpl_77;
  and_110_nl <= and_dcpl_79 AND and_dcpl_83;
  and_116_nl <= and_dcpl_89 AND and_dcpl_77;
  and_120_nl <= and_dcpl_89 AND and_dcpl_83;
  and_124_nl <= and_dcpl_97 AND and_dcpl_77;
  and_127_nl <= and_dcpl_97 AND and_dcpl_83;
  and_132_nl <= and_dcpl_105 AND and_dcpl_77;
  and_135_nl <= and_dcpl_105 AND and_dcpl_83;
  and_140_nl <= and_dcpl_113 AND and_dcpl_111;
  and_143_nl <= and_dcpl_113 AND and_dcpl_54;
  and_148_nl <= and_dcpl_121 AND and_dcpl_111;
  and_152_nl <= and_dcpl_121 AND and_dcpl_54;
  and_155_nl <= and_dcpl_128 AND and_dcpl_111;
  vec_rsc_0_0_i_radr_d_pff <= MUX1HOT_v_6_32_2((COMP_LOOP_1_acc_10_itm_10_1_1(9 DOWNTO
      4)), COMP_LOOP_acc_psp_sva, (COMP_LOOP_acc_1_cse_2_sva(9 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_2_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_11_psp_sva(8 DOWNTO 3)), (COMP_LOOP_acc_10_cse_10_1_3_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_1_cse_4_sva(9 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_4_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_13_psp_sva(7 DOWNTO 2)), (COMP_LOOP_acc_10_cse_10_1_5_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_1_cse_6_sva(9 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_6_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_14_psp_sva(8 DOWNTO 3)), (COMP_LOOP_acc_10_cse_10_1_7_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_1_cse_8_sva(9 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_8_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_16_psp_sva(6 DOWNTO 1)), (COMP_LOOP_acc_10_cse_10_1_9_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_1_cse_10_sva(9 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_10_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_17_psp_sva(8 DOWNTO 3)), (COMP_LOOP_acc_10_cse_10_1_11_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_1_cse_12_sva(9 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_12_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_19_psp_sva(7 DOWNTO 2)), (COMP_LOOP_acc_10_cse_10_1_13_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_1_cse_14_sva(9 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_14_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_20_psp_sva(8 DOWNTO 3)), (COMP_LOOP_acc_10_cse_10_1_15_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_1_cse_sva(9 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_sva(9
      DOWNTO 4)), STD_LOGIC_VECTOR'( and_dcpl_62 & and_dcpl_65 & and_94_nl & and_dcpl_70
      & and_99_nl & and_dcpl_74 & and_106_nl & and_dcpl_81 & and_110_nl & and_dcpl_86
      & and_116_nl & and_dcpl_93 & and_120_nl & and_dcpl_95 & and_124_nl & and_dcpl_100
      & and_127_nl & and_dcpl_102 & and_132_nl & and_dcpl_108 & and_135_nl & and_dcpl_110
      & and_140_nl & and_dcpl_116 & and_143_nl & and_dcpl_119 & and_148_nl & and_dcpl_125
      & and_152_nl & and_dcpl_127 & and_155_nl & and_dcpl_130));
  and_158_nl <= and_dcpl_131 AND and_dcpl_77;
  and_159_nl <= and_dcpl_51 AND and_dcpl_69;
  and_160_nl <= and_dcpl_131 AND and_dcpl_83;
  and_161_nl <= and_dcpl_131 AND and_dcpl_85;
  and_163_nl <= and_dcpl_136 AND and_dcpl_77;
  and_164_nl <= and_dcpl_79 AND and_dcpl_91;
  and_165_nl <= and_dcpl_136 AND and_dcpl_83;
  and_166_nl <= and_dcpl_136 AND and_dcpl_85;
  and_168_nl <= and_dcpl_141 AND and_dcpl_77;
  and_169_nl <= and_dcpl_89 AND and_dcpl_91;
  and_170_nl <= and_dcpl_141 AND and_dcpl_83;
  and_171_nl <= and_dcpl_141 AND and_dcpl_85;
  and_173_nl <= and_dcpl_146 AND and_dcpl_77;
  and_174_nl <= and_dcpl_97 AND and_dcpl_91;
  and_175_nl <= and_dcpl_146 AND and_dcpl_83;
  and_176_nl <= and_dcpl_146 AND and_dcpl_85;
  and_178_nl <= and_dcpl_151 AND and_dcpl_111;
  and_179_nl <= and_dcpl_105 AND and_dcpl_91;
  and_180_nl <= and_dcpl_151 AND and_dcpl_54;
  and_181_nl <= and_dcpl_151 AND and_dcpl_118;
  and_183_nl <= and_dcpl_156 AND and_dcpl_111;
  and_184_nl <= and_dcpl_113 AND and_dcpl_123;
  and_185_nl <= and_dcpl_156 AND and_dcpl_54;
  and_186_nl <= and_dcpl_156 AND and_dcpl_118;
  and_188_nl <= and_dcpl_161 AND and_dcpl_111;
  and_189_nl <= and_dcpl_121 AND and_dcpl_123;
  and_190_nl <= and_dcpl_161 AND and_dcpl_54;
  and_191_nl <= and_dcpl_161 AND and_dcpl_118;
  and_193_nl <= and_dcpl_166 AND and_dcpl_111;
  and_194_nl <= and_dcpl_128 AND and_dcpl_123;
  and_195_nl <= and_dcpl_166 AND and_dcpl_54;
  and_196_nl <= and_dcpl_166 AND and_dcpl_118;
  vec_rsc_0_0_i_wadr_d_pff <= MUX1HOT_v_6_32_2((COMP_LOOP_acc_10_cse_10_1_1_sva(9
      DOWNTO 4)), COMP_LOOP_acc_psp_sva, (COMP_LOOP_acc_10_cse_10_1_2_sva(9 DOWNTO
      4)), (COMP_LOOP_acc_1_cse_2_sva(9 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_3_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_11_psp_sva(8 DOWNTO 3)), (COMP_LOOP_acc_10_cse_10_1_4_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_1_cse_4_sva(9 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_5_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_13_psp_sva(7 DOWNTO 2)), (COMP_LOOP_acc_10_cse_10_1_6_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_1_cse_6_sva(9 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_7_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_14_psp_sva(8 DOWNTO 3)), (COMP_LOOP_acc_10_cse_10_1_8_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_1_cse_8_sva(9 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_9_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_16_psp_sva(6 DOWNTO 1)), (COMP_LOOP_acc_10_cse_10_1_10_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_1_cse_10_sva(9 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_11_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_17_psp_sva(8 DOWNTO 3)), (COMP_LOOP_acc_10_cse_10_1_12_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_1_cse_12_sva(9 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_13_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_19_psp_sva(7 DOWNTO 2)), (COMP_LOOP_acc_10_cse_10_1_14_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_1_cse_14_sva(9 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_15_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_20_psp_sva(8 DOWNTO 3)), (COMP_LOOP_acc_10_cse_10_1_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_1_cse_sva(9 DOWNTO 4)), STD_LOGIC_VECTOR'( and_158_nl
      & and_159_nl & and_160_nl & and_161_nl & and_163_nl & and_164_nl & and_165_nl
      & and_166_nl & and_168_nl & and_169_nl & and_170_nl & and_171_nl & and_173_nl
      & and_174_nl & and_175_nl & and_176_nl & and_178_nl & and_179_nl & and_180_nl
      & and_181_nl & and_183_nl & and_184_nl & and_185_nl & and_186_nl & and_188_nl
      & and_189_nl & and_190_nl & and_191_nl & and_193_nl & and_194_nl & and_195_nl
      & and_196_nl));
  nor_1596_nl <= NOT((NOT (fsm_output(5))) OR (VEC_LOOP_j_10_0_sva_9_0(3)) OR (fsm_output(0))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(1)) OR (VEC_LOOP_j_10_0_sva_9_0(1))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")) OR (VEC_LOOP_j_10_0_sva_9_0(2))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  or_763_nl <= (VEC_LOOP_j_10_0_sva_9_0(1)) OR mux_1116_cse;
  or_757_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR nand_324_cse;
  or_755_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(7)) OR not_tmp_395;
  mux_1113_nl <= MUX_s_1_2_2(or_757_nl, or_755_nl, fsm_output(2));
  or_753_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011"));
  or_752_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001"));
  mux_1112_nl <= MUX_s_1_2_2(or_753_nl, or_752_nl, fsm_output(2));
  mux_1114_nl <= MUX_s_1_2_2(mux_1113_nl, mux_1112_nl, fsm_output(3));
  mux_1117_nl <= MUX_s_1_2_2(or_763_nl, mux_1114_nl, fsm_output(1));
  nor_1597_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1117_nl);
  nor_1598_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR nand_324_cse);
  nor_1599_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1109_nl <= MUX_s_1_2_2(nor_1598_nl, nor_1599_nl, fsm_output(2));
  nor_1600_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1601_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1108_nl <= MUX_s_1_2_2(nor_1600_nl, nor_1601_nl, fsm_output(2));
  mux_1110_nl <= MUX_s_1_2_2(mux_1109_nl, mux_1108_nl, fsm_output(3));
  nor_1602_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1603_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1106_nl <= MUX_s_1_2_2(nor_1602_nl, nor_1603_nl, fsm_output(2));
  nor_1604_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1605_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1105_nl <= MUX_s_1_2_2(nor_1604_nl, nor_1605_nl, fsm_output(2));
  mux_1107_nl <= MUX_s_1_2_2(mux_1106_nl, mux_1105_nl, fsm_output(3));
  mux_1111_nl <= MUX_s_1_2_2(mux_1110_nl, mux_1107_nl, fsm_output(1));
  mux_1118_nl <= MUX_s_1_2_2(nor_1597_nl, mux_1111_nl, fsm_output(0));
  nor_1606_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR nand_324_cse);
  nor_1607_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1101_nl <= MUX_s_1_2_2(nor_1606_nl, nor_1607_nl, fsm_output(2));
  nor_1608_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1609_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1100_nl <= MUX_s_1_2_2(nor_1608_nl, nor_1609_nl, fsm_output(2));
  mux_1102_nl <= MUX_s_1_2_2(mux_1101_nl, mux_1100_nl, fsm_output(3));
  nor_1610_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1611_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1098_nl <= MUX_s_1_2_2(nor_1610_nl, nor_1611_nl, fsm_output(2));
  nor_1612_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1613_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1097_nl <= MUX_s_1_2_2(nor_1612_nl, nor_1613_nl, fsm_output(2));
  mux_1099_nl <= MUX_s_1_2_2(mux_1098_nl, mux_1097_nl, fsm_output(3));
  mux_1103_nl <= MUX_s_1_2_2(mux_1102_nl, mux_1099_nl, fsm_output(1));
  nor_1614_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR nand_324_cse);
  nor_1615_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1094_nl <= MUX_s_1_2_2(nor_1614_nl, nor_1615_nl, fsm_output(2));
  nor_1616_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1617_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1093_nl <= MUX_s_1_2_2(nor_1616_nl, nor_1617_nl, fsm_output(2));
  mux_1095_nl <= MUX_s_1_2_2(mux_1094_nl, mux_1093_nl, fsm_output(3));
  nor_1618_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1619_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1091_nl <= MUX_s_1_2_2(nor_1618_nl, nor_1619_nl, fsm_output(2));
  nor_1620_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1621_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1090_nl <= MUX_s_1_2_2(nor_1620_nl, nor_1621_nl, fsm_output(2));
  mux_1092_nl <= MUX_s_1_2_2(mux_1091_nl, mux_1090_nl, fsm_output(3));
  mux_1096_nl <= MUX_s_1_2_2(mux_1095_nl, mux_1092_nl, fsm_output(1));
  mux_1104_nl <= MUX_s_1_2_2(mux_1103_nl, mux_1096_nl, fsm_output(0));
  mux_1119_nl <= MUX_s_1_2_2(mux_1118_nl, mux_1104_nl, fsm_output(5));
  vec_rsc_0_0_i_we_d_pff <= MUX_s_1_2_2(nor_1596_nl, mux_1119_nl, fsm_output(4));
  nor_1569_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(2))) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm) OR nand_301_cse);
  nor_1570_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1571_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR nand_301_cse);
  mux_1146_nl <= MUX_s_1_2_2(nor_1570_nl, nor_1571_nl, fsm_output(2));
  nor_1572_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1147_nl <= MUX_s_1_2_2(mux_1146_nl, nor_1572_nl, fsm_output(5));
  mux_1148_nl <= MUX_s_1_2_2(nor_1569_nl, mux_1147_nl, fsm_output(6));
  nor_1573_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1574_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR nand_301_cse);
  mux_1143_nl <= MUX_s_1_2_2(nor_1573_nl, nor_1574_nl, fsm_output(2));
  nor_1575_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1144_nl <= MUX_s_1_2_2(mux_1143_nl, nor_1575_nl, fsm_output(5));
  nor_1576_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) OR (NOT (fsm_output(5))) OR (NOT
      (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR not_tmp_399);
  mux_1145_nl <= MUX_s_1_2_2(mux_1144_nl, nor_1576_nl, fsm_output(6));
  mux_1149_nl <= MUX_s_1_2_2(mux_1148_nl, mux_1145_nl, fsm_output(1));
  nor_1577_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (NOT COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm)
      OR nand_301_cse);
  nor_1578_nl <= NOT((NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(7)) OR (fsm_output(4))
      OR (fsm_output(8)));
  nor_1579_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR nand_301_cse);
  mux_1139_nl <= MUX_s_1_2_2(nor_1578_nl, nor_1579_nl, fsm_output(2));
  mux_1140_nl <= MUX_s_1_2_2(nor_1577_nl, mux_1139_nl, fsm_output(5));
  nor_1580_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4))
      OR (fsm_output(8)));
  mux_1141_nl <= MUX_s_1_2_2(mux_1140_nl, nor_1580_nl, fsm_output(6));
  nor_1581_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) OR (VEC_LOOP_j_10_0_sva_9_0(3))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (VEC_LOOP_j_10_0_sva_9_0(2)) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1582_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR nand_301_cse);
  nor_1583_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm) OR (fsm_output(7)) OR not_tmp_399);
  mux_1136_nl <= MUX_s_1_2_2(nor_1582_nl, nor_1583_nl, fsm_output(2));
  nor_1584_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR not_tmp_399);
  mux_1137_nl <= MUX_s_1_2_2(mux_1136_nl, nor_1584_nl, fsm_output(5));
  mux_1138_nl <= MUX_s_1_2_2(nor_1581_nl, mux_1137_nl, fsm_output(6));
  mux_1142_nl <= MUX_s_1_2_2(mux_1141_nl, mux_1138_nl, fsm_output(1));
  mux_1150_nl <= MUX_s_1_2_2(mux_1149_nl, mux_1142_nl, fsm_output(0));
  nor_1585_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR not_tmp_399);
  nor_1586_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1132_nl <= MUX_s_1_2_2(nor_1585_nl, nor_1586_nl, fsm_output(2));
  and_561_nl <= (fsm_output(5)) AND mux_1132_nl;
  or_785_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_783_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1131_nl <= MUX_s_1_2_2(or_785_nl, or_783_nl, fsm_output(2));
  nor_1587_nl <= NOT((fsm_output(5)) OR mux_1131_nl);
  mux_1133_nl <= MUX_s_1_2_2(and_561_nl, nor_1587_nl, fsm_output(6));
  or_781_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_779_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1129_nl <= MUX_s_1_2_2(or_781_nl, or_779_nl, fsm_output(2));
  nor_1588_nl <= NOT((fsm_output(5)) OR mux_1129_nl);
  and_562_nl <= nor_346_cse AND mux_1128_cse;
  mux_1130_nl <= MUX_s_1_2_2(nor_1588_nl, and_562_nl, fsm_output(6));
  mux_1134_nl <= MUX_s_1_2_2(mux_1133_nl, mux_1130_nl, fsm_output(1));
  or_775_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm) OR (fsm_output(7)) OR not_tmp_399;
  or_773_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(4))) OR (fsm_output(8));
  mux_1125_nl <= MUX_s_1_2_2(or_775_nl, or_773_nl, fsm_output(2));
  or_772_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_770_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1124_nl <= MUX_s_1_2_2(or_772_nl, or_770_nl, fsm_output(2));
  mux_1126_nl <= MUX_s_1_2_2(mux_1125_nl, mux_1124_nl, fsm_output(5));
  nor_1591_nl <= NOT((fsm_output(6)) OR mux_1126_nl);
  nor_1592_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(4))) OR (fsm_output(8)));
  nor_1593_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR (fsm_output(7)) OR (NOT (fsm_output(4)))
      OR (fsm_output(8)));
  mux_1122_nl <= MUX_s_1_2_2(nor_1592_nl, nor_1593_nl, fsm_output(2));
  nor_1594_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  nor_1595_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(7)) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1121_nl <= MUX_s_1_2_2(nor_1594_nl, nor_1595_nl, fsm_output(2));
  mux_1123_nl <= MUX_s_1_2_2(mux_1122_nl, mux_1121_nl, fsm_output(5));
  and_563_nl <= (fsm_output(6)) AND mux_1123_nl;
  mux_1127_nl <= MUX_s_1_2_2(nor_1591_nl, and_563_nl, fsm_output(1));
  mux_1135_nl <= MUX_s_1_2_2(mux_1134_nl, mux_1127_nl, fsm_output(0));
  vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1150_nl, mux_1135_nl,
      fsm_output(3));
  nor_1539_nl <= NOT((NOT (fsm_output(5))) OR (VEC_LOOP_j_10_0_sva_9_0(3)) OR (fsm_output(0))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(1)) OR (VEC_LOOP_j_10_0_sva_9_0(1))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")) OR (VEC_LOOP_j_10_0_sva_9_0(2))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  nor_1540_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) OR mux_1116_cse);
  nor_1541_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR nand_324_cse);
  nor_1542_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1175_nl <= MUX_s_1_2_2(nor_1541_nl, nor_1542_nl, fsm_output(2));
  nor_1543_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1544_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1174_nl <= MUX_s_1_2_2(nor_1543_nl, nor_1544_nl, fsm_output(2));
  mux_1176_nl <= MUX_s_1_2_2(mux_1175_nl, mux_1174_nl, fsm_output(3));
  mux_1179_nl <= MUX_s_1_2_2(nor_1540_nl, mux_1176_nl, fsm_output(1));
  and_560_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1179_nl;
  nor_1545_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR nand_324_cse);
  nor_1546_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1171_nl <= MUX_s_1_2_2(nor_1545_nl, nor_1546_nl, fsm_output(2));
  nor_1547_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1548_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1170_nl <= MUX_s_1_2_2(nor_1547_nl, nor_1548_nl, fsm_output(2));
  mux_1172_nl <= MUX_s_1_2_2(mux_1171_nl, mux_1170_nl, fsm_output(3));
  nor_1549_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1550_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1168_nl <= MUX_s_1_2_2(nor_1549_nl, nor_1550_nl, fsm_output(2));
  nor_1551_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1552_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1167_nl <= MUX_s_1_2_2(nor_1551_nl, nor_1552_nl, fsm_output(2));
  mux_1169_nl <= MUX_s_1_2_2(mux_1168_nl, mux_1167_nl, fsm_output(3));
  mux_1173_nl <= MUX_s_1_2_2(mux_1172_nl, mux_1169_nl, fsm_output(1));
  mux_1180_nl <= MUX_s_1_2_2(and_560_nl, mux_1173_nl, fsm_output(0));
  nor_1553_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR nand_324_cse);
  mux_1163_nl <= MUX_s_1_2_2(nor_1553_nl, nor_1554_cse, fsm_output(2));
  nor_1556_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1162_nl <= MUX_s_1_2_2(nor_1523_cse, nor_1556_nl, fsm_output(2));
  mux_1164_nl <= MUX_s_1_2_2(mux_1163_nl, mux_1162_nl, fsm_output(3));
  nor_1557_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  mux_1160_nl <= MUX_s_1_2_2(nor_1557_nl, nor_1526_cse, fsm_output(2));
  nor_1560_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1159_nl <= MUX_s_1_2_2(nor_1527_cse, nor_1560_nl, fsm_output(2));
  mux_1161_nl <= MUX_s_1_2_2(mux_1160_nl, mux_1159_nl, fsm_output(3));
  mux_1165_nl <= MUX_s_1_2_2(mux_1164_nl, mux_1161_nl, fsm_output(1));
  nor_1561_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000"))
      OR nand_272_cse);
  nor_1562_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1156_nl <= MUX_s_1_2_2(nor_1561_nl, nor_1562_nl, fsm_output(2));
  nor_1563_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1564_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1155_nl <= MUX_s_1_2_2(nor_1563_nl, nor_1564_nl, fsm_output(2));
  mux_1157_nl <= MUX_s_1_2_2(mux_1156_nl, mux_1155_nl, fsm_output(3));
  nor_1565_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1566_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1153_nl <= MUX_s_1_2_2(nor_1565_nl, nor_1566_nl, fsm_output(2));
  nor_1567_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1568_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1152_nl <= MUX_s_1_2_2(nor_1567_nl, nor_1568_nl, fsm_output(2));
  mux_1154_nl <= MUX_s_1_2_2(mux_1153_nl, mux_1152_nl, fsm_output(3));
  mux_1158_nl <= MUX_s_1_2_2(mux_1157_nl, mux_1154_nl, fsm_output(1));
  mux_1166_nl <= MUX_s_1_2_2(mux_1165_nl, mux_1158_nl, fsm_output(0));
  mux_1181_nl <= MUX_s_1_2_2(mux_1180_nl, mux_1166_nl, fsm_output(5));
  vec_rsc_0_1_i_we_d_pff <= MUX_s_1_2_2(nor_1539_nl, mux_1181_nl, fsm_output(4));
  nor_1506_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_1507_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  mux_1210_nl <= MUX_s_1_2_2(nor_1506_nl, nor_1507_nl, fsm_output(5));
  nor_1508_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(8)));
  nor_1509_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1209_nl <= MUX_s_1_2_2(nor_1508_nl, nor_1509_nl, fsm_output(5));
  mux_1211_nl <= MUX_s_1_2_2(mux_1210_nl, mux_1209_nl, fsm_output(1));
  nor_1510_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_1511_nl <= NOT((NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1207_nl <= MUX_s_1_2_2(nor_1510_nl, nor_1511_nl, fsm_output(5));
  nor_1512_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(3)) OR (fsm_output(5)) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1208_nl <= MUX_s_1_2_2(mux_1207_nl, nor_1512_nl, fsm_output(1));
  mux_1212_nl <= MUX_s_1_2_2(mux_1211_nl, mux_1208_nl, fsm_output(0));
  nor_1513_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR nand_271_cse);
  nor_1514_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  mux_1204_nl <= MUX_s_1_2_2(nor_1513_nl, nor_1514_nl, fsm_output(5));
  nor_1515_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT
      (fsm_output(8))));
  nor_1516_nl <= NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm) OR (fsm_output(7)) OR not_tmp_395);
  mux_1203_nl <= MUX_s_1_2_2(nor_1515_nl, nor_1516_nl, fsm_output(5));
  mux_1205_nl <= MUX_s_1_2_2(mux_1204_nl, mux_1203_nl, fsm_output(1));
  nor_1517_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm) OR (NOT (fsm_output(2))) OR
      (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT (fsm_output(8))));
  nor_1518_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT
      (fsm_output(8))));
  mux_1201_nl <= MUX_s_1_2_2(nor_1517_nl, nor_1518_nl, fsm_output(5));
  nor_1519_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3
      DOWNTO 1)/=STD_LOGIC_VECTOR'("000")) OR nand_272_cse);
  nor_1520_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm) OR (fsm_output(7)) OR not_tmp_395);
  mux_1199_nl <= MUX_s_1_2_2(nor_1519_nl, nor_1520_nl, fsm_output(2));
  nor_1521_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR not_tmp_395);
  mux_1200_nl <= MUX_s_1_2_2(mux_1199_nl, nor_1521_nl, fsm_output(5));
  mux_1202_nl <= MUX_s_1_2_2(mux_1201_nl, mux_1200_nl, fsm_output(1));
  mux_1206_nl <= MUX_s_1_2_2(mux_1205_nl, mux_1202_nl, fsm_output(0));
  mux_1213_nl <= MUX_s_1_2_2(mux_1212_nl, mux_1206_nl, fsm_output(4));
  mux_1195_nl <= MUX_s_1_2_2(nor_1554_cse, nor_1523_cse, fsm_output(2));
  nor_1524_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1525_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("010")));
  mux_1194_nl <= MUX_s_1_2_2(nor_1524_nl, nor_1525_nl, fsm_output(2));
  and_558_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1194_nl;
  mux_1196_nl <= MUX_s_1_2_2(mux_1195_nl, and_558_nl, fsm_output(5));
  mux_1192_nl <= MUX_s_1_2_2(nor_1526_cse, nor_1527_cse, fsm_output(2));
  and_559_nl <= nor_351_cse AND mux_1191_cse;
  mux_1193_nl <= MUX_s_1_2_2(mux_1192_nl, and_559_nl, fsm_output(5));
  mux_1197_nl <= MUX_s_1_2_2(mux_1196_nl, mux_1193_nl, fsm_output(1));
  nor_1531_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1532_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("010")));
  mux_1187_nl <= MUX_s_1_2_2(nor_1531_nl, nor_1532_nl, fsm_output(2));
  nor_1533_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1534_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  mux_1186_nl <= MUX_s_1_2_2(nor_1533_nl, nor_1534_nl, fsm_output(2));
  mux_1188_nl <= MUX_s_1_2_2(mux_1187_nl, mux_1186_nl, fsm_output(5));
  nor_1535_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("011")));
  nor_1536_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("001")));
  mux_1184_nl <= MUX_s_1_2_2(nor_1535_nl, nor_1536_nl, fsm_output(2));
  nor_1537_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1538_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1183_nl <= MUX_s_1_2_2(nor_1537_nl, nor_1538_nl, fsm_output(2));
  mux_1185_nl <= MUX_s_1_2_2(mux_1184_nl, mux_1183_nl, fsm_output(5));
  mux_1189_nl <= MUX_s_1_2_2(mux_1188_nl, mux_1185_nl, fsm_output(1));
  mux_1198_nl <= MUX_s_1_2_2(mux_1197_nl, mux_1189_nl, fsm_output(0));
  and_557_nl <= (fsm_output(4)) AND mux_1198_nl;
  vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1213_nl, and_557_nl,
      fsm_output(3));
  nor_1477_nl <= NOT((NOT (fsm_output(5))) OR (VEC_LOOP_j_10_0_sva_9_0(3)) OR (fsm_output(0))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(1)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(1)))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")) OR (VEC_LOOP_j_10_0_sva_9_0(2))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  nand_31_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) AND mux_1241_cse);
  or_952_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR nand_324_cse;
  or_950_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(7)) OR not_tmp_395;
  mux_1238_nl <= MUX_s_1_2_2(or_952_nl, or_950_nl, fsm_output(2));
  or_948_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011"));
  or_947_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001"));
  mux_1237_nl <= MUX_s_1_2_2(or_948_nl, or_947_nl, fsm_output(2));
  mux_1239_nl <= MUX_s_1_2_2(mux_1238_nl, mux_1237_nl, fsm_output(3));
  mux_1242_nl <= MUX_s_1_2_2(nand_31_nl, mux_1239_nl, fsm_output(1));
  nor_1478_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1242_nl);
  nor_1482_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_15_sva(2)) OR (COMP_LOOP_acc_10_cse_10_1_15_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_15_sva(0)) OR nand_268_cse);
  nor_1483_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1234_nl <= MUX_s_1_2_2(nor_1482_nl, nor_1483_nl, fsm_output(2));
  nor_1484_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1485_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1233_nl <= MUX_s_1_2_2(nor_1484_nl, nor_1485_nl, fsm_output(2));
  mux_1235_nl <= MUX_s_1_2_2(mux_1234_nl, mux_1233_nl, fsm_output(3));
  nor_1486_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1487_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1231_nl <= MUX_s_1_2_2(nor_1486_nl, nor_1487_nl, fsm_output(2));
  nor_1488_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1489_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1230_nl <= MUX_s_1_2_2(nor_1488_nl, nor_1489_nl, fsm_output(2));
  mux_1232_nl <= MUX_s_1_2_2(mux_1231_nl, mux_1230_nl, fsm_output(3));
  mux_1236_nl <= MUX_s_1_2_2(mux_1235_nl, mux_1232_nl, fsm_output(1));
  mux_1243_nl <= MUX_s_1_2_2(nor_1478_nl, mux_1236_nl, fsm_output(0));
  nor_1490_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR nand_324_cse);
  nor_1491_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1226_nl <= MUX_s_1_2_2(nor_1490_nl, nor_1491_nl, fsm_output(2));
  nor_1492_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1493_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1225_nl <= MUX_s_1_2_2(nor_1492_nl, nor_1493_nl, fsm_output(2));
  mux_1227_nl <= MUX_s_1_2_2(mux_1226_nl, mux_1225_nl, fsm_output(3));
  nor_1494_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1495_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1223_nl <= MUX_s_1_2_2(nor_1494_nl, nor_1495_nl, fsm_output(2));
  nor_1496_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1497_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1222_nl <= MUX_s_1_2_2(nor_1496_nl, nor_1497_nl, fsm_output(2));
  mux_1224_nl <= MUX_s_1_2_2(mux_1223_nl, mux_1222_nl, fsm_output(3));
  mux_1228_nl <= MUX_s_1_2_2(mux_1227_nl, mux_1224_nl, fsm_output(1));
  nor_1498_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR nand_324_cse);
  nor_1499_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1219_nl <= MUX_s_1_2_2(nor_1498_nl, nor_1499_nl, fsm_output(2));
  nor_1500_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1501_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1218_nl <= MUX_s_1_2_2(nor_1500_nl, nor_1501_nl, fsm_output(2));
  mux_1220_nl <= MUX_s_1_2_2(mux_1219_nl, mux_1218_nl, fsm_output(3));
  nor_1502_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1503_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1216_nl <= MUX_s_1_2_2(nor_1502_nl, nor_1503_nl, fsm_output(2));
  nor_1504_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1505_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1215_nl <= MUX_s_1_2_2(nor_1504_nl, nor_1505_nl, fsm_output(2));
  mux_1217_nl <= MUX_s_1_2_2(mux_1216_nl, mux_1215_nl, fsm_output(3));
  mux_1221_nl <= MUX_s_1_2_2(mux_1220_nl, mux_1217_nl, fsm_output(1));
  mux_1229_nl <= MUX_s_1_2_2(mux_1228_nl, mux_1221_nl, fsm_output(0));
  mux_1244_nl <= MUX_s_1_2_2(mux_1243_nl, mux_1229_nl, fsm_output(5));
  vec_rsc_0_2_i_we_d_pff <= MUX_s_1_2_2(nor_1477_nl, mux_1244_nl, fsm_output(4));
  nor_1450_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(2))) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm) OR nand_301_cse);
  nor_1451_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1452_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR nand_301_cse);
  mux_1271_nl <= MUX_s_1_2_2(nor_1451_nl, nor_1452_nl, fsm_output(2));
  nor_1453_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1272_nl <= MUX_s_1_2_2(mux_1271_nl, nor_1453_nl, fsm_output(5));
  mux_1273_nl <= MUX_s_1_2_2(nor_1450_nl, mux_1272_nl, fsm_output(6));
  nor_1454_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1455_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR nand_301_cse);
  mux_1268_nl <= MUX_s_1_2_2(nor_1454_nl, nor_1455_nl, fsm_output(2));
  nor_1456_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1269_nl <= MUX_s_1_2_2(mux_1268_nl, nor_1456_nl, fsm_output(5));
  nor_1457_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(1))) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR not_tmp_399);
  mux_1270_nl <= MUX_s_1_2_2(mux_1269_nl, nor_1457_nl, fsm_output(6));
  mux_1274_nl <= MUX_s_1_2_2(mux_1273_nl, mux_1270_nl, fsm_output(1));
  nor_1458_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm)
      OR nand_301_cse);
  nor_1459_nl <= NOT((NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(7)) OR (fsm_output(4))
      OR (fsm_output(8)));
  nor_1460_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_15_sva(2)) OR (COMP_LOOP_acc_10_cse_10_1_15_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_15_sva(0)) OR nand_265_cse);
  mux_1264_nl <= MUX_s_1_2_2(nor_1459_nl, nor_1460_nl, fsm_output(2));
  mux_1265_nl <= MUX_s_1_2_2(nor_1458_nl, mux_1264_nl, fsm_output(5));
  nor_1461_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4))
      OR (fsm_output(8)));
  mux_1266_nl <= MUX_s_1_2_2(mux_1265_nl, nor_1461_nl, fsm_output(6));
  nor_1462_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(1))) OR (VEC_LOOP_j_10_0_sva_9_0(3))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (VEC_LOOP_j_10_0_sva_9_0(2)) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1463_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR nand_301_cse);
  nor_1464_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm) OR (fsm_output(7)) OR not_tmp_399);
  mux_1261_nl <= MUX_s_1_2_2(nor_1463_nl, nor_1464_nl, fsm_output(2));
  nor_1465_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR not_tmp_399);
  mux_1262_nl <= MUX_s_1_2_2(mux_1261_nl, nor_1465_nl, fsm_output(5));
  mux_1263_nl <= MUX_s_1_2_2(nor_1462_nl, mux_1262_nl, fsm_output(6));
  mux_1267_nl <= MUX_s_1_2_2(mux_1266_nl, mux_1263_nl, fsm_output(1));
  mux_1275_nl <= MUX_s_1_2_2(mux_1274_nl, mux_1267_nl, fsm_output(0));
  nor_1466_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR not_tmp_399);
  nor_1467_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1257_nl <= MUX_s_1_2_2(nor_1466_nl, nor_1467_nl, fsm_output(2));
  and_554_nl <= (fsm_output(5)) AND mux_1257_nl;
  or_979_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_977_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1256_nl <= MUX_s_1_2_2(or_979_nl, or_977_nl, fsm_output(2));
  nor_1468_nl <= NOT((fsm_output(5)) OR mux_1256_nl);
  mux_1258_nl <= MUX_s_1_2_2(and_554_nl, nor_1468_nl, fsm_output(6));
  or_975_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_973_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1254_nl <= MUX_s_1_2_2(or_975_nl, or_973_nl, fsm_output(2));
  nor_1469_nl <= NOT((fsm_output(5)) OR mux_1254_nl);
  and_555_nl <= (VEC_LOOP_j_10_0_sva_9_0(1)) AND (fsm_output(5)) AND mux_1128_cse;
  mux_1255_nl <= MUX_s_1_2_2(nor_1469_nl, and_555_nl, fsm_output(6));
  mux_1259_nl <= MUX_s_1_2_2(mux_1258_nl, mux_1255_nl, fsm_output(1));
  or_969_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm) OR (fsm_output(7)) OR not_tmp_399;
  or_967_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(4))) OR (fsm_output(8));
  mux_1250_nl <= MUX_s_1_2_2(or_969_nl, or_967_nl, fsm_output(2));
  or_966_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_964_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1249_nl <= MUX_s_1_2_2(or_966_nl, or_964_nl, fsm_output(2));
  mux_1251_nl <= MUX_s_1_2_2(mux_1250_nl, mux_1249_nl, fsm_output(5));
  nor_1472_nl <= NOT((fsm_output(6)) OR mux_1251_nl);
  nor_1473_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(4))) OR (fsm_output(8)));
  nor_1474_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR (fsm_output(7)) OR (NOT (fsm_output(4)))
      OR (fsm_output(8)));
  mux_1247_nl <= MUX_s_1_2_2(nor_1473_nl, nor_1474_nl, fsm_output(2));
  nor_1475_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  nor_1476_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(7)) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1246_nl <= MUX_s_1_2_2(nor_1475_nl, nor_1476_nl, fsm_output(2));
  mux_1248_nl <= MUX_s_1_2_2(mux_1247_nl, mux_1246_nl, fsm_output(5));
  and_556_nl <= (fsm_output(6)) AND mux_1248_nl;
  mux_1252_nl <= MUX_s_1_2_2(nor_1472_nl, and_556_nl, fsm_output(1));
  mux_1260_nl <= MUX_s_1_2_2(mux_1259_nl, mux_1252_nl, fsm_output(0));
  vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1275_nl, mux_1260_nl,
      fsm_output(3));
  nor_1418_nl <= NOT((NOT (fsm_output(5))) OR (VEC_LOOP_j_10_0_sva_9_0(3)) OR (fsm_output(0))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(1)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(1)))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")) OR (VEC_LOOP_j_10_0_sva_9_0(2))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  and_553_nl <= (VEC_LOOP_j_10_0_sva_9_0(1)) AND mux_1241_cse;
  nor_1422_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR nand_324_cse);
  nor_1423_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1300_nl <= MUX_s_1_2_2(nor_1422_nl, nor_1423_nl, fsm_output(2));
  nor_1424_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1425_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1299_nl <= MUX_s_1_2_2(nor_1424_nl, nor_1425_nl, fsm_output(2));
  mux_1301_nl <= MUX_s_1_2_2(mux_1300_nl, mux_1299_nl, fsm_output(3));
  mux_1304_nl <= MUX_s_1_2_2(and_553_nl, mux_1301_nl, fsm_output(1));
  and_552_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1304_nl;
  nor_1426_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR nand_261_cse);
  nor_1427_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1296_nl <= MUX_s_1_2_2(nor_1426_nl, nor_1427_nl, fsm_output(2));
  nor_1428_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1429_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1295_nl <= MUX_s_1_2_2(nor_1428_nl, nor_1429_nl, fsm_output(2));
  mux_1297_nl <= MUX_s_1_2_2(mux_1296_nl, mux_1295_nl, fsm_output(3));
  nor_1430_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1431_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1293_nl <= MUX_s_1_2_2(nor_1430_nl, nor_1431_nl, fsm_output(2));
  nor_1432_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1433_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1292_nl <= MUX_s_1_2_2(nor_1432_nl, nor_1433_nl, fsm_output(2));
  mux_1294_nl <= MUX_s_1_2_2(mux_1293_nl, mux_1292_nl, fsm_output(3));
  mux_1298_nl <= MUX_s_1_2_2(mux_1297_nl, mux_1294_nl, fsm_output(1));
  mux_1305_nl <= MUX_s_1_2_2(and_552_nl, mux_1298_nl, fsm_output(0));
  nor_1434_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR nand_324_cse);
  mux_1288_nl <= MUX_s_1_2_2(nor_1434_nl, nor_1435_cse, fsm_output(2));
  nor_1437_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1287_nl <= MUX_s_1_2_2(nor_1402_cse, nor_1437_nl, fsm_output(2));
  mux_1289_nl <= MUX_s_1_2_2(mux_1288_nl, mux_1287_nl, fsm_output(3));
  nor_1438_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  mux_1285_nl <= MUX_s_1_2_2(nor_1438_nl, nor_1405_cse, fsm_output(2));
  nor_1441_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1284_nl <= MUX_s_1_2_2(nor_1406_cse, nor_1441_nl, fsm_output(2));
  mux_1286_nl <= MUX_s_1_2_2(mux_1285_nl, mux_1284_nl, fsm_output(3));
  mux_1290_nl <= MUX_s_1_2_2(mux_1289_nl, mux_1286_nl, fsm_output(1));
  nor_1442_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("001"))
      OR nand_272_cse);
  nor_1443_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1281_nl <= MUX_s_1_2_2(nor_1442_nl, nor_1443_nl, fsm_output(2));
  nor_1444_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1445_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1280_nl <= MUX_s_1_2_2(nor_1444_nl, nor_1445_nl, fsm_output(2));
  mux_1282_nl <= MUX_s_1_2_2(mux_1281_nl, mux_1280_nl, fsm_output(3));
  nor_1446_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1447_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1278_nl <= MUX_s_1_2_2(nor_1446_nl, nor_1447_nl, fsm_output(2));
  nor_1448_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1449_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1277_nl <= MUX_s_1_2_2(nor_1448_nl, nor_1449_nl, fsm_output(2));
  mux_1279_nl <= MUX_s_1_2_2(mux_1278_nl, mux_1277_nl, fsm_output(3));
  mux_1283_nl <= MUX_s_1_2_2(mux_1282_nl, mux_1279_nl, fsm_output(1));
  mux_1291_nl <= MUX_s_1_2_2(mux_1290_nl, mux_1283_nl, fsm_output(0));
  mux_1306_nl <= MUX_s_1_2_2(mux_1305_nl, mux_1291_nl, fsm_output(5));
  vec_rsc_0_3_i_we_d_pff <= MUX_s_1_2_2(nor_1418_nl, mux_1306_nl, fsm_output(4));
  nor_1385_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_1386_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  mux_1335_nl <= MUX_s_1_2_2(nor_1385_nl, nor_1386_nl, fsm_output(5));
  nor_1387_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(8)));
  nor_1388_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1334_nl <= MUX_s_1_2_2(nor_1387_nl, nor_1388_nl, fsm_output(5));
  mux_1336_nl <= MUX_s_1_2_2(mux_1335_nl, mux_1334_nl, fsm_output(1));
  nor_1389_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_1390_nl <= NOT((NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1332_nl <= MUX_s_1_2_2(nor_1389_nl, nor_1390_nl, fsm_output(5));
  nor_1391_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(3)) OR (fsm_output(5)) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1333_nl <= MUX_s_1_2_2(mux_1332_nl, nor_1391_nl, fsm_output(1));
  mux_1337_nl <= MUX_s_1_2_2(mux_1336_nl, mux_1333_nl, fsm_output(0));
  nor_1392_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR nand_271_cse);
  nor_1393_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  mux_1329_nl <= MUX_s_1_2_2(nor_1392_nl, nor_1393_nl, fsm_output(5));
  nor_1394_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT
      (fsm_output(8))));
  nor_1395_nl <= NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm) OR (fsm_output(7)) OR not_tmp_395);
  mux_1328_nl <= MUX_s_1_2_2(nor_1394_nl, nor_1395_nl, fsm_output(5));
  mux_1330_nl <= MUX_s_1_2_2(mux_1329_nl, mux_1328_nl, fsm_output(1));
  nor_1396_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm) OR (NOT (fsm_output(2))) OR
      (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT (fsm_output(8))));
  nor_1397_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT
      (fsm_output(8))));
  mux_1326_nl <= MUX_s_1_2_2(nor_1396_nl, nor_1397_nl, fsm_output(5));
  nor_1398_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3
      DOWNTO 1)/=STD_LOGIC_VECTOR'("001")) OR nand_272_cse);
  nor_1399_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm) OR (fsm_output(7)) OR not_tmp_395);
  mux_1324_nl <= MUX_s_1_2_2(nor_1398_nl, nor_1399_nl, fsm_output(2));
  nor_1400_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR not_tmp_395);
  mux_1325_nl <= MUX_s_1_2_2(mux_1324_nl, nor_1400_nl, fsm_output(5));
  mux_1327_nl <= MUX_s_1_2_2(mux_1326_nl, mux_1325_nl, fsm_output(1));
  mux_1331_nl <= MUX_s_1_2_2(mux_1330_nl, mux_1327_nl, fsm_output(0));
  mux_1338_nl <= MUX_s_1_2_2(mux_1337_nl, mux_1331_nl, fsm_output(4));
  mux_1320_nl <= MUX_s_1_2_2(nor_1435_cse, nor_1402_cse, fsm_output(2));
  nor_1403_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1404_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("010")));
  mux_1319_nl <= MUX_s_1_2_2(nor_1403_nl, nor_1404_nl, fsm_output(2));
  and_550_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1319_nl;
  mux_1321_nl <= MUX_s_1_2_2(mux_1320_nl, and_550_nl, fsm_output(5));
  mux_1317_nl <= MUX_s_1_2_2(nor_1405_cse, nor_1406_cse, fsm_output(2));
  and_551_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND mux_1191_cse;
  mux_1318_nl <= MUX_s_1_2_2(mux_1317_nl, and_551_nl, fsm_output(5));
  mux_1322_nl <= MUX_s_1_2_2(mux_1321_nl, mux_1318_nl, fsm_output(1));
  nor_1410_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1411_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("010")));
  mux_1312_nl <= MUX_s_1_2_2(nor_1410_nl, nor_1411_nl, fsm_output(2));
  nor_1412_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1413_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  mux_1311_nl <= MUX_s_1_2_2(nor_1412_nl, nor_1413_nl, fsm_output(2));
  mux_1313_nl <= MUX_s_1_2_2(mux_1312_nl, mux_1311_nl, fsm_output(5));
  nor_1414_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("011")));
  nor_1415_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("001")));
  mux_1309_nl <= MUX_s_1_2_2(nor_1414_nl, nor_1415_nl, fsm_output(2));
  nor_1416_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1417_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1308_nl <= MUX_s_1_2_2(nor_1416_nl, nor_1417_nl, fsm_output(2));
  mux_1310_nl <= MUX_s_1_2_2(mux_1309_nl, mux_1308_nl, fsm_output(5));
  mux_1314_nl <= MUX_s_1_2_2(mux_1313_nl, mux_1310_nl, fsm_output(1));
  mux_1323_nl <= MUX_s_1_2_2(mux_1322_nl, mux_1314_nl, fsm_output(0));
  and_549_nl <= (fsm_output(4)) AND mux_1323_nl;
  vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1338_nl, and_549_nl,
      fsm_output(3));
  nor_1359_nl <= NOT((NOT (fsm_output(5))) OR (VEC_LOOP_j_10_0_sva_9_0(3)) OR (fsm_output(0))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(1)) OR (VEC_LOOP_j_10_0_sva_9_0(1))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  or_1151_nl <= (VEC_LOOP_j_10_0_sva_9_0(1)) OR mux_1366_cse;
  or_1145_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR nand_324_cse;
  or_1143_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(7)) OR not_tmp_395;
  mux_1363_nl <= MUX_s_1_2_2(or_1145_nl, or_1143_nl, fsm_output(2));
  or_1141_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011"));
  or_1140_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001"));
  mux_1362_nl <= MUX_s_1_2_2(or_1141_nl, or_1140_nl, fsm_output(2));
  mux_1364_nl <= MUX_s_1_2_2(mux_1363_nl, mux_1362_nl, fsm_output(3));
  mux_1367_nl <= MUX_s_1_2_2(or_1151_nl, mux_1364_nl, fsm_output(1));
  nor_1360_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1367_nl);
  nor_1361_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR nand_324_cse);
  nor_1362_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1359_nl <= MUX_s_1_2_2(nor_1361_nl, nor_1362_nl, fsm_output(2));
  nor_1363_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1364_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1358_nl <= MUX_s_1_2_2(nor_1363_nl, nor_1364_nl, fsm_output(2));
  mux_1360_nl <= MUX_s_1_2_2(mux_1359_nl, mux_1358_nl, fsm_output(3));
  nor_1365_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1366_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1356_nl <= MUX_s_1_2_2(nor_1365_nl, nor_1366_nl, fsm_output(2));
  nor_1367_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1368_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1355_nl <= MUX_s_1_2_2(nor_1367_nl, nor_1368_nl, fsm_output(2));
  mux_1357_nl <= MUX_s_1_2_2(mux_1356_nl, mux_1355_nl, fsm_output(3));
  mux_1361_nl <= MUX_s_1_2_2(mux_1360_nl, mux_1357_nl, fsm_output(1));
  mux_1368_nl <= MUX_s_1_2_2(nor_1360_nl, mux_1361_nl, fsm_output(0));
  nor_1369_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR nand_324_cse);
  nor_1370_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1351_nl <= MUX_s_1_2_2(nor_1369_nl, nor_1370_nl, fsm_output(2));
  nor_1371_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1372_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1350_nl <= MUX_s_1_2_2(nor_1371_nl, nor_1372_nl, fsm_output(2));
  mux_1352_nl <= MUX_s_1_2_2(mux_1351_nl, mux_1350_nl, fsm_output(3));
  nor_1373_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1374_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1348_nl <= MUX_s_1_2_2(nor_1373_nl, nor_1374_nl, fsm_output(2));
  nor_1375_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1376_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1347_nl <= MUX_s_1_2_2(nor_1375_nl, nor_1376_nl, fsm_output(2));
  mux_1349_nl <= MUX_s_1_2_2(mux_1348_nl, mux_1347_nl, fsm_output(3));
  mux_1353_nl <= MUX_s_1_2_2(mux_1352_nl, mux_1349_nl, fsm_output(1));
  nor_1377_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR nand_324_cse);
  nor_1378_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1344_nl <= MUX_s_1_2_2(nor_1377_nl, nor_1378_nl, fsm_output(2));
  nor_1379_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1380_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1343_nl <= MUX_s_1_2_2(nor_1379_nl, nor_1380_nl, fsm_output(2));
  mux_1345_nl <= MUX_s_1_2_2(mux_1344_nl, mux_1343_nl, fsm_output(3));
  nor_1381_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1382_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1341_nl <= MUX_s_1_2_2(nor_1381_nl, nor_1382_nl, fsm_output(2));
  nor_1383_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1384_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1340_nl <= MUX_s_1_2_2(nor_1383_nl, nor_1384_nl, fsm_output(2));
  mux_1342_nl <= MUX_s_1_2_2(mux_1341_nl, mux_1340_nl, fsm_output(3));
  mux_1346_nl <= MUX_s_1_2_2(mux_1345_nl, mux_1342_nl, fsm_output(1));
  mux_1354_nl <= MUX_s_1_2_2(mux_1353_nl, mux_1346_nl, fsm_output(0));
  mux_1369_nl <= MUX_s_1_2_2(mux_1368_nl, mux_1354_nl, fsm_output(5));
  vec_rsc_0_4_i_we_d_pff <= MUX_s_1_2_2(nor_1359_nl, mux_1369_nl, fsm_output(4));
  nor_1332_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(2))) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm) OR nand_301_cse);
  nor_1333_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1334_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR nand_301_cse);
  mux_1396_nl <= MUX_s_1_2_2(nor_1333_nl, nor_1334_nl, fsm_output(2));
  nor_1335_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1397_nl <= MUX_s_1_2_2(mux_1396_nl, nor_1335_nl, fsm_output(5));
  mux_1398_nl <= MUX_s_1_2_2(nor_1332_nl, mux_1397_nl, fsm_output(6));
  nor_1336_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1337_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR nand_301_cse);
  mux_1393_nl <= MUX_s_1_2_2(nor_1336_nl, nor_1337_nl, fsm_output(2));
  nor_1338_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1394_nl <= MUX_s_1_2_2(mux_1393_nl, nor_1338_nl, fsm_output(5));
  nor_1339_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) OR (NOT (fsm_output(5))) OR (NOT
      (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR not_tmp_399);
  mux_1395_nl <= MUX_s_1_2_2(mux_1394_nl, nor_1339_nl, fsm_output(6));
  mux_1399_nl <= MUX_s_1_2_2(mux_1398_nl, mux_1395_nl, fsm_output(1));
  nor_1340_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm)
      OR nand_301_cse);
  nor_1341_nl <= NOT((NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(7)) OR (fsm_output(4))
      OR (fsm_output(8)));
  nor_1342_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR nand_301_cse);
  mux_1389_nl <= MUX_s_1_2_2(nor_1341_nl, nor_1342_nl, fsm_output(2));
  mux_1390_nl <= MUX_s_1_2_2(nor_1340_nl, mux_1389_nl, fsm_output(5));
  nor_1343_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4))
      OR (fsm_output(8)));
  mux_1391_nl <= MUX_s_1_2_2(mux_1390_nl, nor_1343_nl, fsm_output(6));
  nor_1344_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) OR (VEC_LOOP_j_10_0_sva_9_0(3))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1345_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR nand_301_cse);
  nor_1346_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm) OR (fsm_output(7)) OR not_tmp_399);
  mux_1386_nl <= MUX_s_1_2_2(nor_1345_nl, nor_1346_nl, fsm_output(2));
  nor_1347_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR not_tmp_399);
  mux_1387_nl <= MUX_s_1_2_2(mux_1386_nl, nor_1347_nl, fsm_output(5));
  mux_1388_nl <= MUX_s_1_2_2(nor_1344_nl, mux_1387_nl, fsm_output(6));
  mux_1392_nl <= MUX_s_1_2_2(mux_1391_nl, mux_1388_nl, fsm_output(1));
  mux_1400_nl <= MUX_s_1_2_2(mux_1399_nl, mux_1392_nl, fsm_output(0));
  nor_1348_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR not_tmp_399);
  nor_1349_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1382_nl <= MUX_s_1_2_2(nor_1348_nl, nor_1349_nl, fsm_output(2));
  and_546_nl <= (fsm_output(5)) AND mux_1382_nl;
  or_1173_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_1171_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1381_nl <= MUX_s_1_2_2(or_1173_nl, or_1171_nl, fsm_output(2));
  nor_1350_nl <= NOT((fsm_output(5)) OR mux_1381_nl);
  mux_1383_nl <= MUX_s_1_2_2(and_546_nl, nor_1350_nl, fsm_output(6));
  or_1169_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_1167_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1379_nl <= MUX_s_1_2_2(or_1169_nl, or_1167_nl, fsm_output(2));
  nor_1351_nl <= NOT((fsm_output(5)) OR mux_1379_nl);
  and_547_nl <= nor_346_cse AND mux_1378_cse;
  mux_1380_nl <= MUX_s_1_2_2(nor_1351_nl, and_547_nl, fsm_output(6));
  mux_1384_nl <= MUX_s_1_2_2(mux_1383_nl, mux_1380_nl, fsm_output(1));
  or_1163_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm) OR (fsm_output(7)) OR not_tmp_399;
  or_1161_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(4))) OR (fsm_output(8));
  mux_1375_nl <= MUX_s_1_2_2(or_1163_nl, or_1161_nl, fsm_output(2));
  or_1160_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_1158_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1374_nl <= MUX_s_1_2_2(or_1160_nl, or_1158_nl, fsm_output(2));
  mux_1376_nl <= MUX_s_1_2_2(mux_1375_nl, mux_1374_nl, fsm_output(5));
  nor_1354_nl <= NOT((fsm_output(6)) OR mux_1376_nl);
  nor_1355_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(4))) OR (fsm_output(8)));
  nor_1356_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR (fsm_output(7)) OR (NOT (fsm_output(4)))
      OR (fsm_output(8)));
  mux_1372_nl <= MUX_s_1_2_2(nor_1355_nl, nor_1356_nl, fsm_output(2));
  nor_1357_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  nor_1358_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(7)) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1371_nl <= MUX_s_1_2_2(nor_1357_nl, nor_1358_nl, fsm_output(2));
  mux_1373_nl <= MUX_s_1_2_2(mux_1372_nl, mux_1371_nl, fsm_output(5));
  and_548_nl <= (fsm_output(6)) AND mux_1373_nl;
  mux_1377_nl <= MUX_s_1_2_2(nor_1354_nl, and_548_nl, fsm_output(1));
  mux_1385_nl <= MUX_s_1_2_2(mux_1384_nl, mux_1377_nl, fsm_output(0));
  vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1400_nl, mux_1385_nl,
      fsm_output(3));
  nor_1302_nl <= NOT((NOT (fsm_output(5))) OR (VEC_LOOP_j_10_0_sva_9_0(3)) OR (fsm_output(0))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(1)) OR (VEC_LOOP_j_10_0_sva_9_0(1))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  nor_1303_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) OR mux_1366_cse);
  nor_1304_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR nand_324_cse);
  nor_1305_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1425_nl <= MUX_s_1_2_2(nor_1304_nl, nor_1305_nl, fsm_output(2));
  nor_1306_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1307_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1424_nl <= MUX_s_1_2_2(nor_1306_nl, nor_1307_nl, fsm_output(2));
  mux_1426_nl <= MUX_s_1_2_2(mux_1425_nl, mux_1424_nl, fsm_output(3));
  mux_1429_nl <= MUX_s_1_2_2(nor_1303_nl, mux_1426_nl, fsm_output(1));
  and_545_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1429_nl;
  nor_1308_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR nand_324_cse);
  nor_1309_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1421_nl <= MUX_s_1_2_2(nor_1308_nl, nor_1309_nl, fsm_output(2));
  nor_1310_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1311_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1420_nl <= MUX_s_1_2_2(nor_1310_nl, nor_1311_nl, fsm_output(2));
  mux_1422_nl <= MUX_s_1_2_2(mux_1421_nl, mux_1420_nl, fsm_output(3));
  nor_1312_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1313_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1418_nl <= MUX_s_1_2_2(nor_1312_nl, nor_1313_nl, fsm_output(2));
  nor_1314_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1315_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1417_nl <= MUX_s_1_2_2(nor_1314_nl, nor_1315_nl, fsm_output(2));
  mux_1419_nl <= MUX_s_1_2_2(mux_1418_nl, mux_1417_nl, fsm_output(3));
  mux_1423_nl <= MUX_s_1_2_2(mux_1422_nl, mux_1419_nl, fsm_output(1));
  mux_1430_nl <= MUX_s_1_2_2(and_545_nl, mux_1423_nl, fsm_output(0));
  nor_1316_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR nand_324_cse);
  mux_1413_nl <= MUX_s_1_2_2(nor_1316_nl, nor_1317_cse, fsm_output(2));
  nor_1319_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1412_nl <= MUX_s_1_2_2(nor_1286_cse, nor_1319_nl, fsm_output(2));
  mux_1414_nl <= MUX_s_1_2_2(mux_1413_nl, mux_1412_nl, fsm_output(3));
  nor_1320_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  mux_1410_nl <= MUX_s_1_2_2(nor_1320_nl, nor_1289_cse, fsm_output(2));
  nor_1323_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1409_nl <= MUX_s_1_2_2(nor_1290_cse, nor_1323_nl, fsm_output(2));
  mux_1411_nl <= MUX_s_1_2_2(mux_1410_nl, mux_1409_nl, fsm_output(3));
  mux_1415_nl <= MUX_s_1_2_2(mux_1414_nl, mux_1411_nl, fsm_output(1));
  nor_1324_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010"))
      OR nand_272_cse);
  nor_1325_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1406_nl <= MUX_s_1_2_2(nor_1324_nl, nor_1325_nl, fsm_output(2));
  nor_1326_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1327_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1405_nl <= MUX_s_1_2_2(nor_1326_nl, nor_1327_nl, fsm_output(2));
  mux_1407_nl <= MUX_s_1_2_2(mux_1406_nl, mux_1405_nl, fsm_output(3));
  nor_1328_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1329_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1403_nl <= MUX_s_1_2_2(nor_1328_nl, nor_1329_nl, fsm_output(2));
  nor_1330_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1331_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1402_nl <= MUX_s_1_2_2(nor_1330_nl, nor_1331_nl, fsm_output(2));
  mux_1404_nl <= MUX_s_1_2_2(mux_1403_nl, mux_1402_nl, fsm_output(3));
  mux_1408_nl <= MUX_s_1_2_2(mux_1407_nl, mux_1404_nl, fsm_output(1));
  mux_1416_nl <= MUX_s_1_2_2(mux_1415_nl, mux_1408_nl, fsm_output(0));
  mux_1431_nl <= MUX_s_1_2_2(mux_1430_nl, mux_1416_nl, fsm_output(5));
  vec_rsc_0_5_i_we_d_pff <= MUX_s_1_2_2(nor_1302_nl, mux_1431_nl, fsm_output(4));
  nor_1269_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_1270_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  mux_1460_nl <= MUX_s_1_2_2(nor_1269_nl, nor_1270_nl, fsm_output(5));
  nor_1271_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(8)));
  nor_1272_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1459_nl <= MUX_s_1_2_2(nor_1271_nl, nor_1272_nl, fsm_output(5));
  mux_1461_nl <= MUX_s_1_2_2(mux_1460_nl, mux_1459_nl, fsm_output(1));
  nor_1273_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_1274_nl <= NOT((NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1457_nl <= MUX_s_1_2_2(nor_1273_nl, nor_1274_nl, fsm_output(5));
  nor_1275_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(3)) OR (fsm_output(5)) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1458_nl <= MUX_s_1_2_2(mux_1457_nl, nor_1275_nl, fsm_output(1));
  mux_1462_nl <= MUX_s_1_2_2(mux_1461_nl, mux_1458_nl, fsm_output(0));
  nor_1276_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR nand_271_cse);
  nor_1277_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  mux_1454_nl <= MUX_s_1_2_2(nor_1276_nl, nor_1277_nl, fsm_output(5));
  nor_1278_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT
      (fsm_output(8))));
  nor_1279_nl <= NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm) OR (fsm_output(7)) OR not_tmp_395);
  mux_1453_nl <= MUX_s_1_2_2(nor_1278_nl, nor_1279_nl, fsm_output(5));
  mux_1455_nl <= MUX_s_1_2_2(mux_1454_nl, mux_1453_nl, fsm_output(1));
  nor_1280_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm) OR (NOT (fsm_output(2))) OR
      (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT (fsm_output(8))));
  nor_1281_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT
      (fsm_output(8))));
  mux_1451_nl <= MUX_s_1_2_2(nor_1280_nl, nor_1281_nl, fsm_output(5));
  nor_1282_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3
      DOWNTO 1)/=STD_LOGIC_VECTOR'("010")) OR nand_272_cse);
  nor_1283_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm) OR (fsm_output(7)) OR not_tmp_395);
  mux_1449_nl <= MUX_s_1_2_2(nor_1282_nl, nor_1283_nl, fsm_output(2));
  nor_1284_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR not_tmp_395);
  mux_1450_nl <= MUX_s_1_2_2(mux_1449_nl, nor_1284_nl, fsm_output(5));
  mux_1452_nl <= MUX_s_1_2_2(mux_1451_nl, mux_1450_nl, fsm_output(1));
  mux_1456_nl <= MUX_s_1_2_2(mux_1455_nl, mux_1452_nl, fsm_output(0));
  mux_1463_nl <= MUX_s_1_2_2(mux_1462_nl, mux_1456_nl, fsm_output(4));
  mux_1445_nl <= MUX_s_1_2_2(nor_1317_cse, nor_1286_cse, fsm_output(2));
  nor_1287_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1288_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("010")));
  mux_1444_nl <= MUX_s_1_2_2(nor_1287_nl, nor_1288_nl, fsm_output(2));
  and_543_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1444_nl;
  mux_1446_nl <= MUX_s_1_2_2(mux_1445_nl, and_543_nl, fsm_output(5));
  mux_1442_nl <= MUX_s_1_2_2(nor_1289_cse, nor_1290_cse, fsm_output(2));
  and_544_nl <= nor_351_cse AND mux_1441_cse;
  mux_1443_nl <= MUX_s_1_2_2(mux_1442_nl, and_544_nl, fsm_output(5));
  mux_1447_nl <= MUX_s_1_2_2(mux_1446_nl, mux_1443_nl, fsm_output(1));
  nor_1294_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1295_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("010")));
  mux_1437_nl <= MUX_s_1_2_2(nor_1294_nl, nor_1295_nl, fsm_output(2));
  nor_1296_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1297_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  mux_1436_nl <= MUX_s_1_2_2(nor_1296_nl, nor_1297_nl, fsm_output(2));
  mux_1438_nl <= MUX_s_1_2_2(mux_1437_nl, mux_1436_nl, fsm_output(5));
  nor_1298_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("011")));
  nor_1299_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("001")));
  mux_1434_nl <= MUX_s_1_2_2(nor_1298_nl, nor_1299_nl, fsm_output(2));
  nor_1300_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1301_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1433_nl <= MUX_s_1_2_2(nor_1300_nl, nor_1301_nl, fsm_output(2));
  mux_1435_nl <= MUX_s_1_2_2(mux_1434_nl, mux_1433_nl, fsm_output(5));
  mux_1439_nl <= MUX_s_1_2_2(mux_1438_nl, mux_1435_nl, fsm_output(1));
  mux_1448_nl <= MUX_s_1_2_2(mux_1447_nl, mux_1439_nl, fsm_output(0));
  and_542_nl <= (fsm_output(4)) AND mux_1448_nl;
  vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1463_nl, and_542_nl,
      fsm_output(3));
  nor_1240_nl <= NOT((NOT (fsm_output(5))) OR (VEC_LOOP_j_10_0_sva_9_0(3)) OR (fsm_output(0))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(1)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(1)))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  nand_47_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) AND mux_1491_cse);
  or_1340_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR nand_324_cse;
  or_1338_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(7)) OR not_tmp_395;
  mux_1488_nl <= MUX_s_1_2_2(or_1340_nl, or_1338_nl, fsm_output(2));
  or_1336_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011"));
  or_1335_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001"));
  mux_1487_nl <= MUX_s_1_2_2(or_1336_nl, or_1335_nl, fsm_output(2));
  mux_1489_nl <= MUX_s_1_2_2(mux_1488_nl, mux_1487_nl, fsm_output(3));
  mux_1492_nl <= MUX_s_1_2_2(nand_47_nl, mux_1489_nl, fsm_output(1));
  nor_1241_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1492_nl);
  nor_1245_nl <= NOT((NOT (COMP_LOOP_acc_10_cse_10_1_15_sva(2))) OR (COMP_LOOP_acc_10_cse_10_1_15_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_15_sva(0)) OR nand_268_cse);
  nor_1246_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1484_nl <= MUX_s_1_2_2(nor_1245_nl, nor_1246_nl, fsm_output(2));
  nor_1247_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1248_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1483_nl <= MUX_s_1_2_2(nor_1247_nl, nor_1248_nl, fsm_output(2));
  mux_1485_nl <= MUX_s_1_2_2(mux_1484_nl, mux_1483_nl, fsm_output(3));
  nor_1249_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1250_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1481_nl <= MUX_s_1_2_2(nor_1249_nl, nor_1250_nl, fsm_output(2));
  nor_1251_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1252_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1480_nl <= MUX_s_1_2_2(nor_1251_nl, nor_1252_nl, fsm_output(2));
  mux_1482_nl <= MUX_s_1_2_2(mux_1481_nl, mux_1480_nl, fsm_output(3));
  mux_1486_nl <= MUX_s_1_2_2(mux_1485_nl, mux_1482_nl, fsm_output(1));
  mux_1493_nl <= MUX_s_1_2_2(nor_1241_nl, mux_1486_nl, fsm_output(0));
  nor_1253_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR nand_324_cse);
  nor_1254_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1476_nl <= MUX_s_1_2_2(nor_1253_nl, nor_1254_nl, fsm_output(2));
  nor_1255_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1256_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1475_nl <= MUX_s_1_2_2(nor_1255_nl, nor_1256_nl, fsm_output(2));
  mux_1477_nl <= MUX_s_1_2_2(mux_1476_nl, mux_1475_nl, fsm_output(3));
  nor_1257_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1258_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1473_nl <= MUX_s_1_2_2(nor_1257_nl, nor_1258_nl, fsm_output(2));
  nor_1259_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1260_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1472_nl <= MUX_s_1_2_2(nor_1259_nl, nor_1260_nl, fsm_output(2));
  mux_1474_nl <= MUX_s_1_2_2(mux_1473_nl, mux_1472_nl, fsm_output(3));
  mux_1478_nl <= MUX_s_1_2_2(mux_1477_nl, mux_1474_nl, fsm_output(1));
  nor_1261_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR nand_324_cse);
  nor_1262_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1469_nl <= MUX_s_1_2_2(nor_1261_nl, nor_1262_nl, fsm_output(2));
  nor_1263_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1264_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1468_nl <= MUX_s_1_2_2(nor_1263_nl, nor_1264_nl, fsm_output(2));
  mux_1470_nl <= MUX_s_1_2_2(mux_1469_nl, mux_1468_nl, fsm_output(3));
  nor_1265_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1266_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1466_nl <= MUX_s_1_2_2(nor_1265_nl, nor_1266_nl, fsm_output(2));
  nor_1267_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1268_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1465_nl <= MUX_s_1_2_2(nor_1267_nl, nor_1268_nl, fsm_output(2));
  mux_1467_nl <= MUX_s_1_2_2(mux_1466_nl, mux_1465_nl, fsm_output(3));
  mux_1471_nl <= MUX_s_1_2_2(mux_1470_nl, mux_1467_nl, fsm_output(1));
  mux_1479_nl <= MUX_s_1_2_2(mux_1478_nl, mux_1471_nl, fsm_output(0));
  mux_1494_nl <= MUX_s_1_2_2(mux_1493_nl, mux_1479_nl, fsm_output(5));
  vec_rsc_0_6_i_we_d_pff <= MUX_s_1_2_2(nor_1240_nl, mux_1494_nl, fsm_output(4));
  nor_1213_nl <= NOT((NOT((fsm_output(5)) AND (fsm_output(2)) AND (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      AND CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))
      AND COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm)) OR nand_301_cse);
  nor_1214_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1215_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR nand_301_cse);
  mux_1521_nl <= MUX_s_1_2_2(nor_1214_nl, nor_1215_nl, fsm_output(2));
  nor_1216_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1522_nl <= MUX_s_1_2_2(mux_1521_nl, nor_1216_nl, fsm_output(5));
  mux_1523_nl <= MUX_s_1_2_2(nor_1213_nl, mux_1522_nl, fsm_output(6));
  nor_1217_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1218_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR nand_301_cse);
  mux_1518_nl <= MUX_s_1_2_2(nor_1217_nl, nor_1218_nl, fsm_output(2));
  nor_1219_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1519_nl <= MUX_s_1_2_2(mux_1518_nl, nor_1219_nl, fsm_output(5));
  nor_1220_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(1))) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR not_tmp_399);
  mux_1520_nl <= MUX_s_1_2_2(mux_1519_nl, nor_1220_nl, fsm_output(6));
  mux_1524_nl <= MUX_s_1_2_2(mux_1523_nl, mux_1520_nl, fsm_output(1));
  nor_1221_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (NOT COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm)
      OR nand_301_cse);
  nor_1222_nl <= NOT((NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(7)) OR (fsm_output(4))
      OR (fsm_output(8)));
  nor_1223_nl <= NOT((NOT (COMP_LOOP_acc_10_cse_10_1_15_sva(2))) OR (COMP_LOOP_acc_10_cse_10_1_15_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_15_sva(0)) OR nand_265_cse);
  mux_1514_nl <= MUX_s_1_2_2(nor_1222_nl, nor_1223_nl, fsm_output(2));
  mux_1515_nl <= MUX_s_1_2_2(nor_1221_nl, mux_1514_nl, fsm_output(5));
  nor_1224_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4))
      OR (fsm_output(8)));
  mux_1516_nl <= MUX_s_1_2_2(mux_1515_nl, nor_1224_nl, fsm_output(6));
  nor_1225_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(1))) OR (VEC_LOOP_j_10_0_sva_9_0(3))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1226_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR nand_301_cse);
  nor_1227_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm) OR (fsm_output(7)) OR not_tmp_399);
  mux_1511_nl <= MUX_s_1_2_2(nor_1226_nl, nor_1227_nl, fsm_output(2));
  nor_1228_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR not_tmp_399);
  mux_1512_nl <= MUX_s_1_2_2(mux_1511_nl, nor_1228_nl, fsm_output(5));
  mux_1513_nl <= MUX_s_1_2_2(nor_1225_nl, mux_1512_nl, fsm_output(6));
  mux_1517_nl <= MUX_s_1_2_2(mux_1516_nl, mux_1513_nl, fsm_output(1));
  mux_1525_nl <= MUX_s_1_2_2(mux_1524_nl, mux_1517_nl, fsm_output(0));
  nor_1229_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR not_tmp_399);
  nor_1230_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1507_nl <= MUX_s_1_2_2(nor_1229_nl, nor_1230_nl, fsm_output(2));
  and_539_nl <= (fsm_output(5)) AND mux_1507_nl;
  or_1367_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_1365_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1506_nl <= MUX_s_1_2_2(or_1367_nl, or_1365_nl, fsm_output(2));
  nor_1231_nl <= NOT((fsm_output(5)) OR mux_1506_nl);
  mux_1508_nl <= MUX_s_1_2_2(and_539_nl, nor_1231_nl, fsm_output(6));
  or_1363_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_1361_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1504_nl <= MUX_s_1_2_2(or_1363_nl, or_1361_nl, fsm_output(2));
  nor_1232_nl <= NOT((fsm_output(5)) OR mux_1504_nl);
  and_540_nl <= (VEC_LOOP_j_10_0_sva_9_0(1)) AND (fsm_output(5)) AND mux_1378_cse;
  mux_1505_nl <= MUX_s_1_2_2(nor_1232_nl, and_540_nl, fsm_output(6));
  mux_1509_nl <= MUX_s_1_2_2(mux_1508_nl, mux_1505_nl, fsm_output(1));
  or_1357_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm) OR (fsm_output(7)) OR not_tmp_399;
  or_1355_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(4))) OR (fsm_output(8));
  mux_1500_nl <= MUX_s_1_2_2(or_1357_nl, or_1355_nl, fsm_output(2));
  or_1354_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_1352_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1499_nl <= MUX_s_1_2_2(or_1354_nl, or_1352_nl, fsm_output(2));
  mux_1501_nl <= MUX_s_1_2_2(mux_1500_nl, mux_1499_nl, fsm_output(5));
  nor_1235_nl <= NOT((fsm_output(6)) OR mux_1501_nl);
  nor_1236_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(4))) OR (fsm_output(8)));
  nor_1237_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR (fsm_output(7)) OR (NOT (fsm_output(4)))
      OR (fsm_output(8)));
  mux_1497_nl <= MUX_s_1_2_2(nor_1236_nl, nor_1237_nl, fsm_output(2));
  nor_1238_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  nor_1239_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(7)) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1496_nl <= MUX_s_1_2_2(nor_1238_nl, nor_1239_nl, fsm_output(2));
  mux_1498_nl <= MUX_s_1_2_2(mux_1497_nl, mux_1496_nl, fsm_output(5));
  and_541_nl <= (fsm_output(6)) AND mux_1498_nl;
  mux_1502_nl <= MUX_s_1_2_2(nor_1235_nl, and_541_nl, fsm_output(1));
  mux_1510_nl <= MUX_s_1_2_2(mux_1509_nl, mux_1502_nl, fsm_output(0));
  vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1525_nl, mux_1510_nl,
      fsm_output(3));
  nor_1184_nl <= NOT((NOT (fsm_output(5))) OR (VEC_LOOP_j_10_0_sva_9_0(3)) OR (fsm_output(0))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(1)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(1)))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  and_535_nl <= (VEC_LOOP_j_10_0_sva_9_0(1)) AND mux_1491_cse;
  nor_1188_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR nand_324_cse);
  nor_1189_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1550_nl <= MUX_s_1_2_2(nor_1188_nl, nor_1189_nl, fsm_output(2));
  nor_1190_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1191_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1549_nl <= MUX_s_1_2_2(nor_1190_nl, nor_1191_nl, fsm_output(2));
  mux_1551_nl <= MUX_s_1_2_2(mux_1550_nl, mux_1549_nl, fsm_output(3));
  mux_1554_nl <= MUX_s_1_2_2(and_535_nl, mux_1551_nl, fsm_output(1));
  and_534_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1554_nl;
  nor_1192_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"))
      OR nand_261_cse);
  nor_1193_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1546_nl <= MUX_s_1_2_2(nor_1192_nl, nor_1193_nl, fsm_output(2));
  and_536_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_1194_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1545_nl <= MUX_s_1_2_2(and_536_nl, nor_1194_nl, fsm_output(2));
  mux_1547_nl <= MUX_s_1_2_2(mux_1546_nl, mux_1545_nl, fsm_output(3));
  and_842_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  nor_1196_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1543_nl <= MUX_s_1_2_2(and_842_nl, nor_1196_nl, fsm_output(2));
  nor_1197_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1198_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1542_nl <= MUX_s_1_2_2(nor_1197_nl, nor_1198_nl, fsm_output(2));
  mux_1544_nl <= MUX_s_1_2_2(mux_1543_nl, mux_1542_nl, fsm_output(3));
  mux_1548_nl <= MUX_s_1_2_2(mux_1547_nl, mux_1544_nl, fsm_output(1));
  mux_1555_nl <= MUX_s_1_2_2(and_534_nl, mux_1548_nl, fsm_output(0));
  nor_1199_nl <= NOT(nand_226_cse OR nand_324_cse);
  mux_1538_nl <= MUX_s_1_2_2(nor_1199_nl, nor_1200_cse, fsm_output(2));
  nor_1201_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1537_nl <= MUX_s_1_2_2(and_529_cse, nor_1201_nl, fsm_output(2));
  mux_1539_nl <= MUX_s_1_2_2(mux_1538_nl, mux_1537_nl, fsm_output(3));
  and_853_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  mux_1535_nl <= MUX_s_1_2_2(and_853_nl, nor_1173_cse, fsm_output(2));
  nor_1205_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1534_nl <= MUX_s_1_2_2(nor_1174_cse, nor_1205_nl, fsm_output(2));
  mux_1536_nl <= MUX_s_1_2_2(mux_1535_nl, mux_1534_nl, fsm_output(3));
  mux_1540_nl <= MUX_s_1_2_2(mux_1539_nl, mux_1536_nl, fsm_output(1));
  nor_1206_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("011"))
      OR nand_272_cse);
  nor_1207_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1531_nl <= MUX_s_1_2_2(nor_1206_nl, nor_1207_nl, fsm_output(2));
  and_538_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_1208_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1530_nl <= MUX_s_1_2_2(and_538_nl, nor_1208_nl, fsm_output(2));
  mux_1532_nl <= MUX_s_1_2_2(mux_1531_nl, mux_1530_nl, fsm_output(3));
  and_872_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  nor_1210_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1528_nl <= MUX_s_1_2_2(and_872_nl, nor_1210_nl, fsm_output(2));
  nor_1211_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1212_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1527_nl <= MUX_s_1_2_2(nor_1211_nl, nor_1212_nl, fsm_output(2));
  mux_1529_nl <= MUX_s_1_2_2(mux_1528_nl, mux_1527_nl, fsm_output(3));
  mux_1533_nl <= MUX_s_1_2_2(mux_1532_nl, mux_1529_nl, fsm_output(1));
  mux_1541_nl <= MUX_s_1_2_2(mux_1540_nl, mux_1533_nl, fsm_output(0));
  mux_1556_nl <= MUX_s_1_2_2(mux_1555_nl, mux_1541_nl, fsm_output(5));
  vec_rsc_0_7_i_we_d_pff <= MUX_s_1_2_2(nor_1184_nl, mux_1556_nl, fsm_output(4));
  nor_1154_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_1155_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  mux_1585_nl <= MUX_s_1_2_2(nor_1154_nl, nor_1155_nl, fsm_output(5));
  nor_1156_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(8)));
  nor_1157_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1584_nl <= MUX_s_1_2_2(nor_1156_nl, nor_1157_nl, fsm_output(5));
  mux_1586_nl <= MUX_s_1_2_2(mux_1585_nl, mux_1584_nl, fsm_output(1));
  nor_1158_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_1159_nl <= NOT((NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1582_nl <= MUX_s_1_2_2(nor_1158_nl, nor_1159_nl, fsm_output(5));
  nor_1160_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(3)) OR (fsm_output(5)) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111")) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1583_nl <= MUX_s_1_2_2(mux_1582_nl, nor_1160_nl, fsm_output(1));
  mux_1587_nl <= MUX_s_1_2_2(mux_1586_nl, mux_1583_nl, fsm_output(0));
  nor_1161_nl <= NOT(nand_226_cse OR nand_271_cse);
  and_852_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (fsm_output(2)) AND CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("011")) AND COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  mux_1579_nl <= MUX_s_1_2_2(nor_1161_nl, and_852_nl, fsm_output(5));
  and_858_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (NOT (fsm_output(6))) AND (fsm_output(8));
  nor_1164_nl <= NOT((NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(2)) AND CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm AND (NOT (fsm_output(7))))) OR not_tmp_395);
  mux_1578_nl <= MUX_s_1_2_2(and_858_nl, nor_1164_nl, fsm_output(5));
  mux_1580_nl <= MUX_s_1_2_2(mux_1579_nl, mux_1578_nl, fsm_output(1));
  and_870_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm AND (fsm_output(2)) AND (fsm_output(7))
      AND (NOT (fsm_output(6))) AND (fsm_output(8));
  and_871_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (NOT (fsm_output(6))) AND (fsm_output(8));
  mux_1576_nl <= MUX_s_1_2_2(and_870_nl, and_871_nl, fsm_output(5));
  nor_1167_nl <= NOT((NOT(COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3
      DOWNTO 1)=STD_LOGIC_VECTOR'("011")))) OR nand_272_cse);
  nor_1168_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm) OR (fsm_output(7)) OR not_tmp_395);
  mux_1574_nl <= MUX_s_1_2_2(nor_1167_nl, nor_1168_nl, fsm_output(2));
  nor_1169_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR not_tmp_395);
  mux_1575_nl <= MUX_s_1_2_2(mux_1574_nl, nor_1169_nl, fsm_output(5));
  mux_1577_nl <= MUX_s_1_2_2(mux_1576_nl, mux_1575_nl, fsm_output(1));
  mux_1581_nl <= MUX_s_1_2_2(mux_1580_nl, mux_1577_nl, fsm_output(0));
  mux_1588_nl <= MUX_s_1_2_2(mux_1587_nl, mux_1581_nl, fsm_output(4));
  mux_1570_nl <= MUX_s_1_2_2(nor_1200_cse, and_529_cse, fsm_output(2));
  nor_1171_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1172_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("010")));
  mux_1569_nl <= MUX_s_1_2_2(nor_1171_nl, nor_1172_nl, fsm_output(2));
  and_530_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1569_nl;
  mux_1571_nl <= MUX_s_1_2_2(mux_1570_nl, and_530_nl, fsm_output(5));
  mux_1567_nl <= MUX_s_1_2_2(nor_1173_cse, nor_1174_cse, fsm_output(2));
  and_531_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND mux_1441_cse;
  mux_1568_nl <= MUX_s_1_2_2(mux_1567_nl, and_531_nl, fsm_output(5));
  mux_1572_nl <= MUX_s_1_2_2(mux_1571_nl, mux_1568_nl, fsm_output(1));
  nor_1178_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1179_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("010")));
  mux_1562_nl <= MUX_s_1_2_2(nor_1178_nl, nor_1179_nl, fsm_output(2));
  nor_1180_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1181_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  mux_1561_nl <= MUX_s_1_2_2(nor_1180_nl, nor_1181_nl, fsm_output(2));
  mux_1563_nl <= MUX_s_1_2_2(mux_1562_nl, mux_1561_nl, fsm_output(5));
  and_532_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm AND CONV_SL_1_1(fsm_output(8 DOWNTO
      6)=STD_LOGIC_VECTOR'("011"));
  nor_1182_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("001")));
  mux_1559_nl <= MUX_s_1_2_2(and_532_nl, nor_1182_nl, fsm_output(2));
  and_533_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_1183_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1558_nl <= MUX_s_1_2_2(and_533_nl, nor_1183_nl, fsm_output(2));
  mux_1560_nl <= MUX_s_1_2_2(mux_1559_nl, mux_1558_nl, fsm_output(5));
  mux_1564_nl <= MUX_s_1_2_2(mux_1563_nl, mux_1560_nl, fsm_output(1));
  mux_1573_nl <= MUX_s_1_2_2(mux_1572_nl, mux_1564_nl, fsm_output(0));
  and_528_nl <= (fsm_output(4)) AND mux_1573_nl;
  vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1588_nl, and_528_nl,
      fsm_output(3));
  nor_1128_nl <= NOT((NOT (fsm_output(5))) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(3)))
      OR (fsm_output(0)) OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(1)) OR (VEC_LOOP_j_10_0_sva_9_0(1))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")) OR (VEC_LOOP_j_10_0_sva_9_0(2))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  or_1539_nl <= (VEC_LOOP_j_10_0_sva_9_0(1)) OR mux_1616_cse;
  or_1533_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR nand_222_cse;
  or_1531_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(7)) OR not_tmp_395;
  mux_1613_nl <= MUX_s_1_2_2(or_1533_nl, or_1531_nl, fsm_output(2));
  or_1529_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011"));
  or_1528_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001"));
  mux_1612_nl <= MUX_s_1_2_2(or_1529_nl, or_1528_nl, fsm_output(2));
  mux_1614_nl <= MUX_s_1_2_2(mux_1613_nl, mux_1612_nl, fsm_output(3));
  mux_1617_nl <= MUX_s_1_2_2(or_1539_nl, mux_1614_nl, fsm_output(1));
  nor_1129_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1617_nl);
  nor_1130_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR nand_324_cse);
  nor_1131_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1609_nl <= MUX_s_1_2_2(nor_1130_nl, nor_1131_nl, fsm_output(2));
  nor_1132_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1133_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1608_nl <= MUX_s_1_2_2(nor_1132_nl, nor_1133_nl, fsm_output(2));
  mux_1610_nl <= MUX_s_1_2_2(mux_1609_nl, mux_1608_nl, fsm_output(3));
  nor_1134_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1135_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1606_nl <= MUX_s_1_2_2(nor_1134_nl, nor_1135_nl, fsm_output(2));
  nor_1136_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1137_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1605_nl <= MUX_s_1_2_2(nor_1136_nl, nor_1137_nl, fsm_output(2));
  mux_1607_nl <= MUX_s_1_2_2(mux_1606_nl, mux_1605_nl, fsm_output(3));
  mux_1611_nl <= MUX_s_1_2_2(mux_1610_nl, mux_1607_nl, fsm_output(1));
  mux_1618_nl <= MUX_s_1_2_2(nor_1129_nl, mux_1611_nl, fsm_output(0));
  nor_1138_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR nand_223_cse);
  nor_1139_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1601_nl <= MUX_s_1_2_2(nor_1138_nl, nor_1139_nl, fsm_output(2));
  nor_1140_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1141_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1600_nl <= MUX_s_1_2_2(nor_1140_nl, nor_1141_nl, fsm_output(2));
  mux_1602_nl <= MUX_s_1_2_2(mux_1601_nl, mux_1600_nl, fsm_output(3));
  nor_1142_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1143_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1598_nl <= MUX_s_1_2_2(nor_1142_nl, nor_1143_nl, fsm_output(2));
  nor_1144_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1145_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1597_nl <= MUX_s_1_2_2(nor_1144_nl, nor_1145_nl, fsm_output(2));
  mux_1599_nl <= MUX_s_1_2_2(mux_1598_nl, mux_1597_nl, fsm_output(3));
  mux_1603_nl <= MUX_s_1_2_2(mux_1602_nl, mux_1599_nl, fsm_output(1));
  nor_1146_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR nand_324_cse);
  nor_1147_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1594_nl <= MUX_s_1_2_2(nor_1146_nl, nor_1147_nl, fsm_output(2));
  nor_1148_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1149_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1593_nl <= MUX_s_1_2_2(nor_1148_nl, nor_1149_nl, fsm_output(2));
  mux_1595_nl <= MUX_s_1_2_2(mux_1594_nl, mux_1593_nl, fsm_output(3));
  nor_1150_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1151_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1591_nl <= MUX_s_1_2_2(nor_1150_nl, nor_1151_nl, fsm_output(2));
  nor_1152_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1153_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1590_nl <= MUX_s_1_2_2(nor_1152_nl, nor_1153_nl, fsm_output(2));
  mux_1592_nl <= MUX_s_1_2_2(mux_1591_nl, mux_1590_nl, fsm_output(3));
  mux_1596_nl <= MUX_s_1_2_2(mux_1595_nl, mux_1592_nl, fsm_output(1));
  mux_1604_nl <= MUX_s_1_2_2(mux_1603_nl, mux_1596_nl, fsm_output(0));
  mux_1619_nl <= MUX_s_1_2_2(mux_1618_nl, mux_1604_nl, fsm_output(5));
  vec_rsc_0_8_i_we_d_pff <= MUX_s_1_2_2(nor_1128_nl, mux_1619_nl, fsm_output(4));
  nor_1101_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(2))) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm) OR nand_301_cse);
  nor_1102_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1103_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR nand_219_cse);
  mux_1646_nl <= MUX_s_1_2_2(nor_1102_nl, nor_1103_nl, fsm_output(2));
  nor_1104_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1647_nl <= MUX_s_1_2_2(mux_1646_nl, nor_1104_nl, fsm_output(5));
  mux_1648_nl <= MUX_s_1_2_2(nor_1101_nl, mux_1647_nl, fsm_output(6));
  nor_1105_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1106_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR nand_301_cse);
  mux_1643_nl <= MUX_s_1_2_2(nor_1105_nl, nor_1106_nl, fsm_output(2));
  nor_1107_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1644_nl <= MUX_s_1_2_2(mux_1643_nl, nor_1107_nl, fsm_output(5));
  nor_1108_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) OR (NOT (fsm_output(5))) OR (NOT
      (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR not_tmp_399);
  mux_1645_nl <= MUX_s_1_2_2(mux_1644_nl, nor_1108_nl, fsm_output(6));
  mux_1649_nl <= MUX_s_1_2_2(mux_1648_nl, mux_1645_nl, fsm_output(1));
  nor_1109_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (NOT COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm)
      OR nand_301_cse);
  nor_1110_nl <= NOT((NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(7)) OR (fsm_output(4))
      OR (fsm_output(8)));
  nor_1111_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR nand_301_cse);
  mux_1639_nl <= MUX_s_1_2_2(nor_1110_nl, nor_1111_nl, fsm_output(2));
  mux_1640_nl <= MUX_s_1_2_2(nor_1109_nl, mux_1639_nl, fsm_output(5));
  nor_1112_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4))
      OR (fsm_output(8)));
  mux_1641_nl <= MUX_s_1_2_2(mux_1640_nl, nor_1112_nl, fsm_output(6));
  nor_1113_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(3)))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (VEC_LOOP_j_10_0_sva_9_0(2)) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_1114_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR nand_301_cse);
  nor_1115_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm) OR (fsm_output(7)) OR not_tmp_399);
  mux_1636_nl <= MUX_s_1_2_2(nor_1114_nl, nor_1115_nl, fsm_output(2));
  nor_1116_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR not_tmp_399);
  mux_1637_nl <= MUX_s_1_2_2(mux_1636_nl, nor_1116_nl, fsm_output(5));
  mux_1638_nl <= MUX_s_1_2_2(nor_1113_nl, mux_1637_nl, fsm_output(6));
  mux_1642_nl <= MUX_s_1_2_2(mux_1641_nl, mux_1638_nl, fsm_output(1));
  mux_1650_nl <= MUX_s_1_2_2(mux_1649_nl, mux_1642_nl, fsm_output(0));
  nor_1117_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR not_tmp_399);
  nor_1118_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1632_nl <= MUX_s_1_2_2(nor_1117_nl, nor_1118_nl, fsm_output(2));
  and_525_nl <= (fsm_output(5)) AND mux_1632_nl;
  or_1561_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_1559_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1631_nl <= MUX_s_1_2_2(or_1561_nl, or_1559_nl, fsm_output(2));
  nor_1119_nl <= NOT((fsm_output(5)) OR mux_1631_nl);
  mux_1633_nl <= MUX_s_1_2_2(and_525_nl, nor_1119_nl, fsm_output(6));
  or_1557_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_1555_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1629_nl <= MUX_s_1_2_2(or_1557_nl, or_1555_nl, fsm_output(2));
  nor_1120_nl <= NOT((fsm_output(5)) OR mux_1629_nl);
  and_526_nl <= nor_346_cse AND mux_1628_cse;
  mux_1630_nl <= MUX_s_1_2_2(nor_1120_nl, and_526_nl, fsm_output(6));
  mux_1634_nl <= MUX_s_1_2_2(mux_1633_nl, mux_1630_nl, fsm_output(1));
  or_1551_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm) OR (fsm_output(7)) OR not_tmp_399;
  or_1549_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(4))) OR (fsm_output(8));
  mux_1625_nl <= MUX_s_1_2_2(or_1551_nl, or_1549_nl, fsm_output(2));
  or_1548_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_1546_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1624_nl <= MUX_s_1_2_2(or_1548_nl, or_1546_nl, fsm_output(2));
  mux_1626_nl <= MUX_s_1_2_2(mux_1625_nl, mux_1624_nl, fsm_output(5));
  nor_1123_nl <= NOT((fsm_output(6)) OR mux_1626_nl);
  nor_1124_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(4))) OR (fsm_output(8)));
  nor_1125_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR (fsm_output(7)) OR (NOT (fsm_output(4)))
      OR (fsm_output(8)));
  mux_1622_nl <= MUX_s_1_2_2(nor_1124_nl, nor_1125_nl, fsm_output(2));
  nor_1126_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  nor_1127_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(7)) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1621_nl <= MUX_s_1_2_2(nor_1126_nl, nor_1127_nl, fsm_output(2));
  mux_1623_nl <= MUX_s_1_2_2(mux_1622_nl, mux_1621_nl, fsm_output(5));
  and_527_nl <= (fsm_output(6)) AND mux_1623_nl;
  mux_1627_nl <= MUX_s_1_2_2(nor_1123_nl, and_527_nl, fsm_output(1));
  mux_1635_nl <= MUX_s_1_2_2(mux_1634_nl, mux_1627_nl, fsm_output(0));
  vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1650_nl, mux_1635_nl,
      fsm_output(3));
  nor_1071_nl <= NOT((NOT (fsm_output(5))) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(3)))
      OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(1))
      OR (VEC_LOOP_j_10_0_sva_9_0(1)) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR (VEC_LOOP_j_10_0_sva_9_0(2)) OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  nor_1072_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) OR mux_1616_cse);
  nor_1073_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR nand_222_cse);
  nor_1074_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1675_nl <= MUX_s_1_2_2(nor_1073_nl, nor_1074_nl, fsm_output(2));
  nor_1075_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1076_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1674_nl <= MUX_s_1_2_2(nor_1075_nl, nor_1076_nl, fsm_output(2));
  mux_1676_nl <= MUX_s_1_2_2(mux_1675_nl, mux_1674_nl, fsm_output(3));
  mux_1679_nl <= MUX_s_1_2_2(nor_1072_nl, mux_1676_nl, fsm_output(1));
  and_524_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1679_nl;
  nor_1077_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR nand_324_cse);
  nor_1078_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1671_nl <= MUX_s_1_2_2(nor_1077_nl, nor_1078_nl, fsm_output(2));
  nor_1079_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1080_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1670_nl <= MUX_s_1_2_2(nor_1079_nl, nor_1080_nl, fsm_output(2));
  mux_1672_nl <= MUX_s_1_2_2(mux_1671_nl, mux_1670_nl, fsm_output(3));
  nor_1081_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1082_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1668_nl <= MUX_s_1_2_2(nor_1081_nl, nor_1082_nl, fsm_output(2));
  nor_1083_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1084_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1667_nl <= MUX_s_1_2_2(nor_1083_nl, nor_1084_nl, fsm_output(2));
  mux_1669_nl <= MUX_s_1_2_2(mux_1668_nl, mux_1667_nl, fsm_output(3));
  mux_1673_nl <= MUX_s_1_2_2(mux_1672_nl, mux_1669_nl, fsm_output(1));
  mux_1680_nl <= MUX_s_1_2_2(and_524_nl, mux_1673_nl, fsm_output(0));
  nor_1085_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR nand_223_cse);
  mux_1663_nl <= MUX_s_1_2_2(nor_1085_nl, nor_1086_cse, fsm_output(2));
  nor_1088_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1662_nl <= MUX_s_1_2_2(nor_1056_cse, nor_1088_nl, fsm_output(2));
  mux_1664_nl <= MUX_s_1_2_2(mux_1663_nl, mux_1662_nl, fsm_output(3));
  nor_1089_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  mux_1660_nl <= MUX_s_1_2_2(nor_1089_nl, nor_1059_cse, fsm_output(2));
  nor_1092_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1659_nl <= MUX_s_1_2_2(nor_1060_cse, nor_1092_nl, fsm_output(2));
  mux_1661_nl <= MUX_s_1_2_2(mux_1660_nl, mux_1659_nl, fsm_output(3));
  mux_1665_nl <= MUX_s_1_2_2(mux_1664_nl, mux_1661_nl, fsm_output(1));
  nor_1093_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))
      OR nand_212_cse);
  nor_1094_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1656_nl <= MUX_s_1_2_2(nor_1093_nl, nor_1094_nl, fsm_output(2));
  nor_1095_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1096_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1655_nl <= MUX_s_1_2_2(nor_1095_nl, nor_1096_nl, fsm_output(2));
  mux_1657_nl <= MUX_s_1_2_2(mux_1656_nl, mux_1655_nl, fsm_output(3));
  nor_1097_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1098_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1653_nl <= MUX_s_1_2_2(nor_1097_nl, nor_1098_nl, fsm_output(2));
  nor_1099_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1100_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1652_nl <= MUX_s_1_2_2(nor_1099_nl, nor_1100_nl, fsm_output(2));
  mux_1654_nl <= MUX_s_1_2_2(mux_1653_nl, mux_1652_nl, fsm_output(3));
  mux_1658_nl <= MUX_s_1_2_2(mux_1657_nl, mux_1654_nl, fsm_output(1));
  mux_1666_nl <= MUX_s_1_2_2(mux_1665_nl, mux_1658_nl, fsm_output(0));
  mux_1681_nl <= MUX_s_1_2_2(mux_1680_nl, mux_1666_nl, fsm_output(5));
  vec_rsc_0_9_i_we_d_pff <= MUX_s_1_2_2(nor_1071_nl, mux_1681_nl, fsm_output(4));
  nor_1039_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_1040_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  mux_1710_nl <= MUX_s_1_2_2(nor_1039_nl, nor_1040_nl, fsm_output(5));
  nor_1041_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(8)));
  nor_1042_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1709_nl <= MUX_s_1_2_2(nor_1041_nl, nor_1042_nl, fsm_output(5));
  mux_1711_nl <= MUX_s_1_2_2(mux_1710_nl, mux_1709_nl, fsm_output(1));
  nor_1043_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_1044_nl <= NOT((NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1707_nl <= MUX_s_1_2_2(nor_1043_nl, nor_1044_nl, fsm_output(5));
  nor_1045_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(3))) OR (fsm_output(5)) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1708_nl <= MUX_s_1_2_2(mux_1707_nl, nor_1045_nl, fsm_output(1));
  mux_1712_nl <= MUX_s_1_2_2(mux_1711_nl, mux_1708_nl, fsm_output(0));
  nor_1046_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR nand_211_cse);
  nor_1047_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  mux_1704_nl <= MUX_s_1_2_2(nor_1046_nl, nor_1047_nl, fsm_output(5));
  nor_1048_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT
      (fsm_output(8))));
  nor_1049_nl <= NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm) OR (fsm_output(7)) OR not_tmp_395);
  mux_1703_nl <= MUX_s_1_2_2(nor_1048_nl, nor_1049_nl, fsm_output(5));
  mux_1705_nl <= MUX_s_1_2_2(mux_1704_nl, mux_1703_nl, fsm_output(1));
  nor_1050_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm) OR (NOT (fsm_output(2))) OR
      (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT (fsm_output(8))));
  nor_1051_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT
      (fsm_output(8))));
  mux_1701_nl <= MUX_s_1_2_2(nor_1050_nl, nor_1051_nl, fsm_output(5));
  nor_1052_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2
      DOWNTO 1)/=STD_LOGIC_VECTOR'("00")) OR nand_212_cse);
  nor_1053_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm) OR (fsm_output(7)) OR not_tmp_395);
  mux_1699_nl <= MUX_s_1_2_2(nor_1052_nl, nor_1053_nl, fsm_output(2));
  nor_1054_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR not_tmp_395);
  mux_1700_nl <= MUX_s_1_2_2(mux_1699_nl, nor_1054_nl, fsm_output(5));
  mux_1702_nl <= MUX_s_1_2_2(mux_1701_nl, mux_1700_nl, fsm_output(1));
  mux_1706_nl <= MUX_s_1_2_2(mux_1705_nl, mux_1702_nl, fsm_output(0));
  mux_1713_nl <= MUX_s_1_2_2(mux_1712_nl, mux_1706_nl, fsm_output(4));
  mux_1695_nl <= MUX_s_1_2_2(nor_1086_cse, nor_1056_cse, fsm_output(2));
  nor_1057_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1058_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("010")));
  mux_1694_nl <= MUX_s_1_2_2(nor_1057_nl, nor_1058_nl, fsm_output(2));
  and_521_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1694_nl;
  mux_1696_nl <= MUX_s_1_2_2(mux_1695_nl, and_521_nl, fsm_output(5));
  mux_1692_nl <= MUX_s_1_2_2(nor_1059_cse, nor_1060_cse, fsm_output(2));
  and_522_nl <= nor_351_cse AND mux_1691_cse;
  mux_1693_nl <= MUX_s_1_2_2(mux_1692_nl, and_522_nl, fsm_output(5));
  mux_1697_nl <= MUX_s_1_2_2(mux_1696_nl, mux_1693_nl, fsm_output(1));
  nor_1063_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1064_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("010")));
  mux_1687_nl <= MUX_s_1_2_2(nor_1063_nl, nor_1064_nl, fsm_output(2));
  nor_1065_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_1066_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  mux_1686_nl <= MUX_s_1_2_2(nor_1065_nl, nor_1066_nl, fsm_output(2));
  mux_1688_nl <= MUX_s_1_2_2(mux_1687_nl, mux_1686_nl, fsm_output(5));
  nor_1067_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("011")));
  nor_1068_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("001")));
  mux_1684_nl <= MUX_s_1_2_2(nor_1067_nl, nor_1068_nl, fsm_output(2));
  nor_1069_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1070_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1683_nl <= MUX_s_1_2_2(nor_1069_nl, nor_1070_nl, fsm_output(2));
  mux_1685_nl <= MUX_s_1_2_2(mux_1684_nl, mux_1683_nl, fsm_output(5));
  mux_1689_nl <= MUX_s_1_2_2(mux_1688_nl, mux_1685_nl, fsm_output(1));
  mux_1698_nl <= MUX_s_1_2_2(mux_1697_nl, mux_1689_nl, fsm_output(0));
  and_520_nl <= (fsm_output(4)) AND mux_1698_nl;
  vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1713_nl, and_520_nl,
      fsm_output(3));
  nor_1010_nl <= NOT((NOT (fsm_output(5))) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(3)))
      OR (fsm_output(0)) OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(1)) OR (NOT
      (VEC_LOOP_j_10_0_sva_9_0(1))) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR (VEC_LOOP_j_10_0_sva_9_0(2)) OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  nand_63_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) AND mux_1741_cse);
  or_1728_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR nand_222_cse;
  or_1726_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(7)) OR not_tmp_395;
  mux_1738_nl <= MUX_s_1_2_2(or_1728_nl, or_1726_nl, fsm_output(2));
  or_1724_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011"));
  or_1723_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001"));
  mux_1737_nl <= MUX_s_1_2_2(or_1724_nl, or_1723_nl, fsm_output(2));
  mux_1739_nl <= MUX_s_1_2_2(mux_1738_nl, mux_1737_nl, fsm_output(3));
  mux_1742_nl <= MUX_s_1_2_2(nand_63_nl, mux_1739_nl, fsm_output(1));
  nor_1011_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1742_nl);
  nor_1015_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_15_sva(2)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_15_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_15_sva(0)) OR nand_268_cse);
  nor_1016_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1734_nl <= MUX_s_1_2_2(nor_1015_nl, nor_1016_nl, fsm_output(2));
  nor_1017_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1018_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1733_nl <= MUX_s_1_2_2(nor_1017_nl, nor_1018_nl, fsm_output(2));
  mux_1735_nl <= MUX_s_1_2_2(mux_1734_nl, mux_1733_nl, fsm_output(3));
  nor_1019_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1020_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1731_nl <= MUX_s_1_2_2(nor_1019_nl, nor_1020_nl, fsm_output(2));
  nor_1021_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1022_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1730_nl <= MUX_s_1_2_2(nor_1021_nl, nor_1022_nl, fsm_output(2));
  mux_1732_nl <= MUX_s_1_2_2(mux_1731_nl, mux_1730_nl, fsm_output(3));
  mux_1736_nl <= MUX_s_1_2_2(mux_1735_nl, mux_1732_nl, fsm_output(1));
  mux_1743_nl <= MUX_s_1_2_2(nor_1011_nl, mux_1736_nl, fsm_output(0));
  nor_1023_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR nand_223_cse);
  nor_1024_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1726_nl <= MUX_s_1_2_2(nor_1023_nl, nor_1024_nl, fsm_output(2));
  nor_1025_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1026_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1725_nl <= MUX_s_1_2_2(nor_1025_nl, nor_1026_nl, fsm_output(2));
  mux_1727_nl <= MUX_s_1_2_2(mux_1726_nl, mux_1725_nl, fsm_output(3));
  nor_1027_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1028_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1723_nl <= MUX_s_1_2_2(nor_1027_nl, nor_1028_nl, fsm_output(2));
  nor_1029_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1030_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1722_nl <= MUX_s_1_2_2(nor_1029_nl, nor_1030_nl, fsm_output(2));
  mux_1724_nl <= MUX_s_1_2_2(mux_1723_nl, mux_1722_nl, fsm_output(3));
  mux_1728_nl <= MUX_s_1_2_2(mux_1727_nl, mux_1724_nl, fsm_output(1));
  nor_1031_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR nand_324_cse);
  nor_1032_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1719_nl <= MUX_s_1_2_2(nor_1031_nl, nor_1032_nl, fsm_output(2));
  nor_1033_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_1034_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1718_nl <= MUX_s_1_2_2(nor_1033_nl, nor_1034_nl, fsm_output(2));
  mux_1720_nl <= MUX_s_1_2_2(mux_1719_nl, mux_1718_nl, fsm_output(3));
  nor_1035_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_1036_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1716_nl <= MUX_s_1_2_2(nor_1035_nl, nor_1036_nl, fsm_output(2));
  nor_1037_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_1038_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1715_nl <= MUX_s_1_2_2(nor_1037_nl, nor_1038_nl, fsm_output(2));
  mux_1717_nl <= MUX_s_1_2_2(mux_1716_nl, mux_1715_nl, fsm_output(3));
  mux_1721_nl <= MUX_s_1_2_2(mux_1720_nl, mux_1717_nl, fsm_output(1));
  mux_1729_nl <= MUX_s_1_2_2(mux_1728_nl, mux_1721_nl, fsm_output(0));
  mux_1744_nl <= MUX_s_1_2_2(mux_1743_nl, mux_1729_nl, fsm_output(5));
  vec_rsc_0_10_i_we_d_pff <= MUX_s_1_2_2(nor_1010_nl, mux_1744_nl, fsm_output(4));
  nor_983_nl <= NOT((NOT((fsm_output(5)) AND (fsm_output(2)) AND (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      AND CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("101"))
      AND COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm)) OR nand_301_cse);
  nor_984_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_985_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR nand_219_cse);
  mux_1771_nl <= MUX_s_1_2_2(nor_984_nl, nor_985_nl, fsm_output(2));
  nor_986_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1772_nl <= MUX_s_1_2_2(mux_1771_nl, nor_986_nl, fsm_output(5));
  mux_1773_nl <= MUX_s_1_2_2(nor_983_nl, mux_1772_nl, fsm_output(6));
  nor_987_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_988_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR nand_301_cse);
  mux_1768_nl <= MUX_s_1_2_2(nor_987_nl, nor_988_nl, fsm_output(2));
  nor_989_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1769_nl <= MUX_s_1_2_2(mux_1768_nl, nor_989_nl, fsm_output(5));
  nor_990_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(1))) OR (NOT (fsm_output(5))) OR
      (NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR not_tmp_399);
  mux_1770_nl <= MUX_s_1_2_2(mux_1769_nl, nor_990_nl, fsm_output(6));
  mux_1774_nl <= MUX_s_1_2_2(mux_1773_nl, mux_1770_nl, fsm_output(1));
  nor_991_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (NOT COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm)
      OR nand_301_cse);
  nor_992_nl <= NOT((NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(7)) OR (fsm_output(4))
      OR (fsm_output(8)));
  nor_993_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_15_sva(2)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_15_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_15_sva(0)) OR nand_265_cse);
  mux_1764_nl <= MUX_s_1_2_2(nor_992_nl, nor_993_nl, fsm_output(2));
  mux_1765_nl <= MUX_s_1_2_2(nor_991_nl, mux_1764_nl, fsm_output(5));
  nor_994_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4))
      OR (fsm_output(8)));
  mux_1766_nl <= MUX_s_1_2_2(mux_1765_nl, nor_994_nl, fsm_output(6));
  nor_995_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(1))) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(3)))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (VEC_LOOP_j_10_0_sva_9_0(2)) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_996_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR nand_301_cse);
  nor_997_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm) OR (fsm_output(7)) OR not_tmp_399);
  mux_1761_nl <= MUX_s_1_2_2(nor_996_nl, nor_997_nl, fsm_output(2));
  nor_998_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR not_tmp_399);
  mux_1762_nl <= MUX_s_1_2_2(mux_1761_nl, nor_998_nl, fsm_output(5));
  mux_1763_nl <= MUX_s_1_2_2(nor_995_nl, mux_1762_nl, fsm_output(6));
  mux_1767_nl <= MUX_s_1_2_2(mux_1766_nl, mux_1763_nl, fsm_output(1));
  mux_1775_nl <= MUX_s_1_2_2(mux_1774_nl, mux_1767_nl, fsm_output(0));
  nor_999_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR not_tmp_399);
  nor_1000_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1757_nl <= MUX_s_1_2_2(nor_999_nl, nor_1000_nl, fsm_output(2));
  and_517_nl <= (fsm_output(5)) AND mux_1757_nl;
  or_1755_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_1753_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1756_nl <= MUX_s_1_2_2(or_1755_nl, or_1753_nl, fsm_output(2));
  nor_1001_nl <= NOT((fsm_output(5)) OR mux_1756_nl);
  mux_1758_nl <= MUX_s_1_2_2(and_517_nl, nor_1001_nl, fsm_output(6));
  or_1751_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_1749_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1754_nl <= MUX_s_1_2_2(or_1751_nl, or_1749_nl, fsm_output(2));
  nor_1002_nl <= NOT((fsm_output(5)) OR mux_1754_nl);
  and_518_nl <= (VEC_LOOP_j_10_0_sva_9_0(1)) AND (fsm_output(5)) AND mux_1628_cse;
  mux_1755_nl <= MUX_s_1_2_2(nor_1002_nl, and_518_nl, fsm_output(6));
  mux_1759_nl <= MUX_s_1_2_2(mux_1758_nl, mux_1755_nl, fsm_output(1));
  or_1745_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm) OR (fsm_output(7)) OR not_tmp_399;
  or_1743_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(4))) OR (fsm_output(8));
  mux_1750_nl <= MUX_s_1_2_2(or_1745_nl, or_1743_nl, fsm_output(2));
  or_1742_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_1740_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1749_nl <= MUX_s_1_2_2(or_1742_nl, or_1740_nl, fsm_output(2));
  mux_1751_nl <= MUX_s_1_2_2(mux_1750_nl, mux_1749_nl, fsm_output(5));
  nor_1005_nl <= NOT((fsm_output(6)) OR mux_1751_nl);
  nor_1006_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(4))) OR (fsm_output(8)));
  nor_1007_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR (fsm_output(7)) OR (NOT (fsm_output(4)))
      OR (fsm_output(8)));
  mux_1747_nl <= MUX_s_1_2_2(nor_1006_nl, nor_1007_nl, fsm_output(2));
  nor_1008_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  nor_1009_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(7)) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1746_nl <= MUX_s_1_2_2(nor_1008_nl, nor_1009_nl, fsm_output(2));
  mux_1748_nl <= MUX_s_1_2_2(mux_1747_nl, mux_1746_nl, fsm_output(5));
  and_519_nl <= (fsm_output(6)) AND mux_1748_nl;
  mux_1752_nl <= MUX_s_1_2_2(nor_1005_nl, and_519_nl, fsm_output(1));
  mux_1760_nl <= MUX_s_1_2_2(mux_1759_nl, mux_1752_nl, fsm_output(0));
  vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1775_nl, mux_1760_nl,
      fsm_output(3));
  nor_954_nl <= NOT((NOT (fsm_output(5))) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(3))) OR
      (fsm_output(0)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(1)) OR
      (NOT (VEC_LOOP_j_10_0_sva_9_0(1))) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR (VEC_LOOP_j_10_0_sva_9_0(2)) OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  and_513_nl <= (VEC_LOOP_j_10_0_sva_9_0(1)) AND mux_1741_cse;
  nor_958_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR nand_222_cse);
  nor_959_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1800_nl <= MUX_s_1_2_2(nor_958_nl, nor_959_nl, fsm_output(2));
  nor_960_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_961_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1799_nl <= MUX_s_1_2_2(nor_960_nl, nor_961_nl, fsm_output(2));
  mux_1801_nl <= MUX_s_1_2_2(mux_1800_nl, mux_1799_nl, fsm_output(3));
  mux_1804_nl <= MUX_s_1_2_2(and_513_nl, mux_1801_nl, fsm_output(1));
  and_512_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1804_nl;
  nor_962_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_15_sva(2)) OR (NOT((COMP_LOOP_acc_10_cse_10_1_15_sva(3))
      AND (COMP_LOOP_acc_10_cse_10_1_15_sva(0)) AND (COMP_LOOP_acc_10_cse_10_1_15_sva(1))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111")))));
  nor_963_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1796_nl <= MUX_s_1_2_2(nor_962_nl, nor_963_nl, fsm_output(2));
  and_514_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_964_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1795_nl <= MUX_s_1_2_2(and_514_nl, nor_964_nl, fsm_output(2));
  mux_1797_nl <= MUX_s_1_2_2(mux_1796_nl, mux_1795_nl, fsm_output(3));
  and_841_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  nor_966_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1793_nl <= MUX_s_1_2_2(and_841_nl, nor_966_nl, fsm_output(2));
  nor_967_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_968_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1792_nl <= MUX_s_1_2_2(nor_967_nl, nor_968_nl, fsm_output(2));
  mux_1794_nl <= MUX_s_1_2_2(mux_1793_nl, mux_1792_nl, fsm_output(3));
  mux_1798_nl <= MUX_s_1_2_2(mux_1797_nl, mux_1794_nl, fsm_output(1));
  mux_1805_nl <= MUX_s_1_2_2(and_512_nl, mux_1798_nl, fsm_output(0));
  nor_969_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR nand_223_cse);
  mux_1788_nl <= MUX_s_1_2_2(nor_969_nl, nor_970_cse, fsm_output(2));
  nor_971_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1787_nl <= MUX_s_1_2_2(and_506_cse, nor_971_nl, fsm_output(2));
  mux_1789_nl <= MUX_s_1_2_2(mux_1788_nl, mux_1787_nl, fsm_output(3));
  and_851_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  mux_1785_nl <= MUX_s_1_2_2(and_851_nl, nor_944_cse, fsm_output(2));
  nor_975_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1784_nl <= MUX_s_1_2_2(nor_945_cse, nor_975_nl, fsm_output(2));
  mux_1786_nl <= MUX_s_1_2_2(mux_1785_nl, mux_1784_nl, fsm_output(3));
  mux_1790_nl <= MUX_s_1_2_2(mux_1789_nl, mux_1786_nl, fsm_output(1));
  nor_976_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01"))
      OR nand_212_cse);
  nor_977_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1781_nl <= MUX_s_1_2_2(nor_976_nl, nor_977_nl, fsm_output(2));
  and_516_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_978_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1780_nl <= MUX_s_1_2_2(and_516_nl, nor_978_nl, fsm_output(2));
  mux_1782_nl <= MUX_s_1_2_2(mux_1781_nl, mux_1780_nl, fsm_output(3));
  and_869_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  nor_980_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1778_nl <= MUX_s_1_2_2(and_869_nl, nor_980_nl, fsm_output(2));
  nor_981_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_982_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1777_nl <= MUX_s_1_2_2(nor_981_nl, nor_982_nl, fsm_output(2));
  mux_1779_nl <= MUX_s_1_2_2(mux_1778_nl, mux_1777_nl, fsm_output(3));
  mux_1783_nl <= MUX_s_1_2_2(mux_1782_nl, mux_1779_nl, fsm_output(1));
  mux_1791_nl <= MUX_s_1_2_2(mux_1790_nl, mux_1783_nl, fsm_output(0));
  mux_1806_nl <= MUX_s_1_2_2(mux_1805_nl, mux_1791_nl, fsm_output(5));
  vec_rsc_0_11_i_we_d_pff <= MUX_s_1_2_2(nor_954_nl, mux_1806_nl, fsm_output(4));
  nor_925_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_926_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  mux_1835_nl <= MUX_s_1_2_2(nor_925_nl, nor_926_nl, fsm_output(5));
  nor_927_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(8)));
  nor_928_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1834_nl <= MUX_s_1_2_2(nor_927_nl, nor_928_nl, fsm_output(5));
  mux_1836_nl <= MUX_s_1_2_2(mux_1835_nl, mux_1834_nl, fsm_output(1));
  nor_929_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_930_nl <= NOT((NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1832_nl <= MUX_s_1_2_2(nor_929_nl, nor_930_nl, fsm_output(5));
  nor_931_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(3))) OR (fsm_output(5)) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1833_nl <= MUX_s_1_2_2(mux_1832_nl, nor_931_nl, fsm_output(1));
  mux_1837_nl <= MUX_s_1_2_2(mux_1836_nl, mux_1833_nl, fsm_output(0));
  nor_932_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR nand_211_cse);
  and_850_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (fsm_output(2)) AND CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("101")) AND COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  mux_1829_nl <= MUX_s_1_2_2(nor_932_nl, and_850_nl, fsm_output(5));
  and_857_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (NOT (fsm_output(6))) AND (fsm_output(8));
  nor_935_nl <= NOT((NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(2)) AND CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm AND (NOT (fsm_output(7))))) OR not_tmp_395);
  mux_1828_nl <= MUX_s_1_2_2(and_857_nl, nor_935_nl, fsm_output(5));
  mux_1830_nl <= MUX_s_1_2_2(mux_1829_nl, mux_1828_nl, fsm_output(1));
  and_867_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm AND (fsm_output(2)) AND (fsm_output(7))
      AND (NOT (fsm_output(6))) AND (fsm_output(8));
  and_868_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (NOT (fsm_output(6))) AND (fsm_output(8));
  mux_1826_nl <= MUX_s_1_2_2(and_867_nl, and_868_nl, fsm_output(5));
  nor_938_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2
      DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR nand_212_cse);
  nor_939_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm) OR (fsm_output(7)) OR not_tmp_395);
  mux_1824_nl <= MUX_s_1_2_2(nor_938_nl, nor_939_nl, fsm_output(2));
  nor_940_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR not_tmp_395);
  mux_1825_nl <= MUX_s_1_2_2(mux_1824_nl, nor_940_nl, fsm_output(5));
  mux_1827_nl <= MUX_s_1_2_2(mux_1826_nl, mux_1825_nl, fsm_output(1));
  mux_1831_nl <= MUX_s_1_2_2(mux_1830_nl, mux_1827_nl, fsm_output(0));
  mux_1838_nl <= MUX_s_1_2_2(mux_1837_nl, mux_1831_nl, fsm_output(4));
  mux_1820_nl <= MUX_s_1_2_2(nor_970_cse, and_506_cse, fsm_output(2));
  nor_942_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_943_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("010")));
  mux_1819_nl <= MUX_s_1_2_2(nor_942_nl, nor_943_nl, fsm_output(2));
  and_507_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1819_nl;
  mux_1821_nl <= MUX_s_1_2_2(mux_1820_nl, and_507_nl, fsm_output(5));
  mux_1817_nl <= MUX_s_1_2_2(nor_944_cse, nor_945_cse, fsm_output(2));
  and_508_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND mux_1691_cse;
  mux_1818_nl <= MUX_s_1_2_2(mux_1817_nl, and_508_nl, fsm_output(5));
  mux_1822_nl <= MUX_s_1_2_2(mux_1821_nl, mux_1818_nl, fsm_output(1));
  nor_948_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_949_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("010")));
  mux_1812_nl <= MUX_s_1_2_2(nor_948_nl, nor_949_nl, fsm_output(2));
  nor_950_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_951_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  mux_1811_nl <= MUX_s_1_2_2(nor_950_nl, nor_951_nl, fsm_output(2));
  mux_1813_nl <= MUX_s_1_2_2(mux_1812_nl, mux_1811_nl, fsm_output(5));
  and_510_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm AND CONV_SL_1_1(fsm_output(8 DOWNTO
      6)=STD_LOGIC_VECTOR'("011"));
  nor_952_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("001")));
  mux_1809_nl <= MUX_s_1_2_2(and_510_nl, nor_952_nl, fsm_output(2));
  and_511_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_953_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1808_nl <= MUX_s_1_2_2(and_511_nl, nor_953_nl, fsm_output(2));
  mux_1810_nl <= MUX_s_1_2_2(mux_1809_nl, mux_1808_nl, fsm_output(5));
  mux_1814_nl <= MUX_s_1_2_2(mux_1813_nl, mux_1810_nl, fsm_output(1));
  mux_1823_nl <= MUX_s_1_2_2(mux_1822_nl, mux_1814_nl, fsm_output(0));
  and_505_nl <= (fsm_output(4)) AND mux_1823_nl;
  vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1838_nl, and_505_nl,
      fsm_output(3));
  nor_899_nl <= NOT((NOT (fsm_output(5))) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(3))) OR
      (fsm_output(0)) OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(1)) OR (VEC_LOOP_j_10_0_sva_9_0(1))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  or_1925_nl <= (VEC_LOOP_j_10_0_sva_9_0(1)) OR mux_1866_cse;
  or_1919_nl <= (COMP_LOOP_acc_20_psp_sva(0)) OR nand_184_cse;
  or_1918_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(7)) OR not_tmp_395;
  mux_1863_nl <= MUX_s_1_2_2(or_1919_nl, or_1918_nl, fsm_output(2));
  or_1916_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011"));
  or_1915_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001"));
  mux_1862_nl <= MUX_s_1_2_2(or_1916_nl, or_1915_nl, fsm_output(2));
  mux_1864_nl <= MUX_s_1_2_2(mux_1863_nl, mux_1862_nl, fsm_output(3));
  mux_1867_nl <= MUX_s_1_2_2(or_1925_nl, mux_1864_nl, fsm_output(1));
  nor_900_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1867_nl);
  nor_901_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR nand_324_cse);
  nor_902_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1859_nl <= MUX_s_1_2_2(nor_901_nl, nor_902_nl, fsm_output(2));
  nor_903_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_904_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1858_nl <= MUX_s_1_2_2(nor_903_nl, nor_904_nl, fsm_output(2));
  mux_1860_nl <= MUX_s_1_2_2(mux_1859_nl, mux_1858_nl, fsm_output(3));
  nor_905_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_906_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1856_nl <= MUX_s_1_2_2(nor_905_nl, nor_906_nl, fsm_output(2));
  nor_907_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_908_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1855_nl <= MUX_s_1_2_2(nor_907_nl, nor_908_nl, fsm_output(2));
  mux_1857_nl <= MUX_s_1_2_2(mux_1856_nl, mux_1855_nl, fsm_output(3));
  mux_1861_nl <= MUX_s_1_2_2(mux_1860_nl, mux_1857_nl, fsm_output(1));
  mux_1868_nl <= MUX_s_1_2_2(nor_900_nl, mux_1861_nl, fsm_output(0));
  nor_909_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR nand_185_cse);
  nor_910_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1851_nl <= MUX_s_1_2_2(nor_909_nl, nor_910_nl, fsm_output(2));
  nor_911_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_912_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1850_nl <= MUX_s_1_2_2(nor_911_nl, nor_912_nl, fsm_output(2));
  mux_1852_nl <= MUX_s_1_2_2(mux_1851_nl, mux_1850_nl, fsm_output(3));
  nor_913_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_914_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1848_nl <= MUX_s_1_2_2(nor_913_nl, nor_914_nl, fsm_output(2));
  nor_915_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_916_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1847_nl <= MUX_s_1_2_2(nor_915_nl, nor_916_nl, fsm_output(2));
  mux_1849_nl <= MUX_s_1_2_2(mux_1848_nl, mux_1847_nl, fsm_output(3));
  mux_1853_nl <= MUX_s_1_2_2(mux_1852_nl, mux_1849_nl, fsm_output(1));
  nor_917_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR nand_324_cse);
  nor_918_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1844_nl <= MUX_s_1_2_2(nor_917_nl, nor_918_nl, fsm_output(2));
  nor_919_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_920_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1843_nl <= MUX_s_1_2_2(nor_919_nl, nor_920_nl, fsm_output(2));
  mux_1845_nl <= MUX_s_1_2_2(mux_1844_nl, mux_1843_nl, fsm_output(3));
  nor_921_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("110")));
  nor_922_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1841_nl <= MUX_s_1_2_2(nor_921_nl, nor_922_nl, fsm_output(2));
  nor_923_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_924_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1840_nl <= MUX_s_1_2_2(nor_923_nl, nor_924_nl, fsm_output(2));
  mux_1842_nl <= MUX_s_1_2_2(mux_1841_nl, mux_1840_nl, fsm_output(3));
  mux_1846_nl <= MUX_s_1_2_2(mux_1845_nl, mux_1842_nl, fsm_output(1));
  mux_1854_nl <= MUX_s_1_2_2(mux_1853_nl, mux_1846_nl, fsm_output(0));
  mux_1869_nl <= MUX_s_1_2_2(mux_1868_nl, mux_1854_nl, fsm_output(5));
  vec_rsc_0_12_i_we_d_pff <= MUX_s_1_2_2(nor_899_nl, mux_1869_nl, fsm_output(4));
  nor_873_nl <= NOT((NOT((fsm_output(5)) AND (fsm_output(2)) AND (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      AND CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("110"))
      AND COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm)) OR nand_301_cse);
  nor_874_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_875_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(7)) AND (fsm_output(4)) AND (fsm_output(8)))));
  mux_1896_nl <= MUX_s_1_2_2(nor_874_nl, nor_875_nl, fsm_output(2));
  nor_876_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1897_nl <= MUX_s_1_2_2(mux_1896_nl, nor_876_nl, fsm_output(5));
  mux_1898_nl <= MUX_s_1_2_2(nor_873_nl, mux_1897_nl, fsm_output(6));
  nor_877_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_878_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR nand_301_cse);
  mux_1893_nl <= MUX_s_1_2_2(nor_877_nl, nor_878_nl, fsm_output(2));
  nor_879_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_1894_nl <= MUX_s_1_2_2(mux_1893_nl, nor_879_nl, fsm_output(5));
  nor_880_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) OR (NOT (fsm_output(5))) OR (NOT
      (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR not_tmp_399);
  mux_1895_nl <= MUX_s_1_2_2(mux_1894_nl, nor_880_nl, fsm_output(6));
  mux_1899_nl <= MUX_s_1_2_2(mux_1898_nl, mux_1895_nl, fsm_output(1));
  nor_881_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (NOT COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm)
      OR nand_301_cse);
  nor_882_nl <= NOT((NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(7)) OR (fsm_output(4))
      OR (fsm_output(8)));
  nor_883_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR nand_301_cse);
  mux_1889_nl <= MUX_s_1_2_2(nor_882_nl, nor_883_nl, fsm_output(2));
  mux_1890_nl <= MUX_s_1_2_2(nor_881_nl, mux_1889_nl, fsm_output(5));
  nor_884_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4))
      OR (fsm_output(8)));
  mux_1891_nl <= MUX_s_1_2_2(mux_1890_nl, nor_884_nl, fsm_output(6));
  nor_885_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(3)))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_886_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR nand_301_cse);
  nor_887_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm) OR (fsm_output(7)) OR not_tmp_399);
  mux_1886_nl <= MUX_s_1_2_2(nor_886_nl, nor_887_nl, fsm_output(2));
  nor_888_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR not_tmp_399);
  mux_1887_nl <= MUX_s_1_2_2(mux_1886_nl, nor_888_nl, fsm_output(5));
  mux_1888_nl <= MUX_s_1_2_2(nor_885_nl, mux_1887_nl, fsm_output(6));
  mux_1892_nl <= MUX_s_1_2_2(mux_1891_nl, mux_1888_nl, fsm_output(1));
  mux_1900_nl <= MUX_s_1_2_2(mux_1899_nl, mux_1892_nl, fsm_output(0));
  nor_889_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR not_tmp_399);
  nor_890_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1882_nl <= MUX_s_1_2_2(nor_889_nl, nor_890_nl, fsm_output(2));
  and_501_nl <= (fsm_output(5)) AND mux_1882_nl;
  or_1947_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_1945_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1881_nl <= MUX_s_1_2_2(or_1947_nl, or_1945_nl, fsm_output(2));
  nor_891_nl <= NOT((fsm_output(5)) OR mux_1881_nl);
  mux_1883_nl <= MUX_s_1_2_2(and_501_nl, nor_891_nl, fsm_output(6));
  or_1943_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_1941_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1879_nl <= MUX_s_1_2_2(or_1943_nl, or_1941_nl, fsm_output(2));
  nor_892_nl <= NOT((fsm_output(5)) OR mux_1879_nl);
  and_502_nl <= nor_346_cse AND mux_1878_cse;
  mux_1880_nl <= MUX_s_1_2_2(nor_892_nl, and_502_nl, fsm_output(6));
  mux_1884_nl <= MUX_s_1_2_2(mux_1883_nl, mux_1880_nl, fsm_output(1));
  or_1937_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm) OR (fsm_output(7)) OR not_tmp_399;
  or_1935_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(4))) OR (fsm_output(8));
  mux_1875_nl <= MUX_s_1_2_2(or_1937_nl, or_1935_nl, fsm_output(2));
  or_1934_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(7)) OR not_tmp_399;
  or_1932_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8));
  mux_1874_nl <= MUX_s_1_2_2(or_1934_nl, or_1932_nl, fsm_output(2));
  mux_1876_nl <= MUX_s_1_2_2(mux_1875_nl, mux_1874_nl, fsm_output(5));
  nor_894_nl <= NOT((fsm_output(6)) OR mux_1876_nl);
  nor_895_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(4))) OR (fsm_output(8)));
  nor_896_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR (fsm_output(7)) OR (NOT (fsm_output(4)))
      OR (fsm_output(8)));
  mux_1872_nl <= MUX_s_1_2_2(nor_895_nl, nor_896_nl, fsm_output(2));
  nor_897_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  nor_898_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(7)) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1871_nl <= MUX_s_1_2_2(nor_897_nl, nor_898_nl, fsm_output(2));
  mux_1873_nl <= MUX_s_1_2_2(mux_1872_nl, mux_1871_nl, fsm_output(5));
  and_504_nl <= (fsm_output(6)) AND mux_1873_nl;
  mux_1877_nl <= MUX_s_1_2_2(nor_894_nl, and_504_nl, fsm_output(1));
  mux_1885_nl <= MUX_s_1_2_2(mux_1884_nl, mux_1877_nl, fsm_output(0));
  vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1900_nl, mux_1885_nl,
      fsm_output(3));
  nor_846_nl <= NOT((NOT (fsm_output(5))) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(3))) OR
      (fsm_output(0)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(1)) OR
      (VEC_LOOP_j_10_0_sva_9_0(1)) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2))) OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  nor_847_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) OR mux_1866_cse);
  nor_848_nl <= NOT((COMP_LOOP_acc_20_psp_sva(0)) OR nand_184_cse);
  nor_849_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1925_nl <= MUX_s_1_2_2(nor_848_nl, nor_849_nl, fsm_output(2));
  nor_850_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("011")));
  nor_851_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1924_nl <= MUX_s_1_2_2(nor_850_nl, nor_851_nl, fsm_output(2));
  mux_1926_nl <= MUX_s_1_2_2(mux_1925_nl, mux_1924_nl, fsm_output(3));
  mux_1929_nl <= MUX_s_1_2_2(nor_847_nl, mux_1926_nl, fsm_output(1));
  and_497_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1929_nl;
  nor_852_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))))
      OR nand_324_cse);
  nor_853_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1921_nl <= MUX_s_1_2_2(nor_852_nl, nor_853_nl, fsm_output(2));
  and_498_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_854_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1920_nl <= MUX_s_1_2_2(and_498_nl, nor_854_nl, fsm_output(2));
  mux_1922_nl <= MUX_s_1_2_2(mux_1921_nl, mux_1920_nl, fsm_output(3));
  and_840_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  nor_856_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1918_nl <= MUX_s_1_2_2(and_840_nl, nor_856_nl, fsm_output(2));
  nor_857_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_858_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1917_nl <= MUX_s_1_2_2(nor_857_nl, nor_858_nl, fsm_output(2));
  mux_1919_nl <= MUX_s_1_2_2(mux_1918_nl, mux_1917_nl, fsm_output(3));
  mux_1923_nl <= MUX_s_1_2_2(mux_1922_nl, mux_1919_nl, fsm_output(1));
  mux_1930_nl <= MUX_s_1_2_2(and_497_nl, mux_1923_nl, fsm_output(0));
  nor_859_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR nand_185_cse);
  mux_1913_nl <= MUX_s_1_2_2(nor_859_nl, nor_860_cse, fsm_output(2));
  nor_861_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1912_nl <= MUX_s_1_2_2(and_490_cse, nor_861_nl, fsm_output(2));
  mux_1914_nl <= MUX_s_1_2_2(mux_1913_nl, mux_1912_nl, fsm_output(3));
  and_849_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  mux_1910_nl <= MUX_s_1_2_2(and_849_nl, nor_837_cse, fsm_output(2));
  nor_865_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1909_nl <= MUX_s_1_2_2(nor_838_cse, nor_865_nl, fsm_output(2));
  mux_1911_nl <= MUX_s_1_2_2(mux_1910_nl, mux_1909_nl, fsm_output(3));
  mux_1915_nl <= MUX_s_1_2_2(mux_1914_nl, mux_1911_nl, fsm_output(1));
  nor_866_nl <= NOT((COMP_LOOP_acc_1_cse_sva(1)) OR nand_170_cse);
  nor_867_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1906_nl <= MUX_s_1_2_2(nor_866_nl, nor_867_nl, fsm_output(2));
  and_500_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_868_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1905_nl <= MUX_s_1_2_2(and_500_nl, nor_868_nl, fsm_output(2));
  mux_1907_nl <= MUX_s_1_2_2(mux_1906_nl, mux_1905_nl, fsm_output(3));
  and_866_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  nor_870_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1903_nl <= MUX_s_1_2_2(and_866_nl, nor_870_nl, fsm_output(2));
  nor_871_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_872_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1902_nl <= MUX_s_1_2_2(nor_871_nl, nor_872_nl, fsm_output(2));
  mux_1904_nl <= MUX_s_1_2_2(mux_1903_nl, mux_1902_nl, fsm_output(3));
  mux_1908_nl <= MUX_s_1_2_2(mux_1907_nl, mux_1904_nl, fsm_output(1));
  mux_1916_nl <= MUX_s_1_2_2(mux_1915_nl, mux_1908_nl, fsm_output(0));
  mux_1931_nl <= MUX_s_1_2_2(mux_1930_nl, mux_1916_nl, fsm_output(5));
  vec_rsc_0_13_i_we_d_pff <= MUX_s_1_2_2(nor_846_nl, mux_1931_nl, fsm_output(4));
  nor_818_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_819_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  mux_1960_nl <= MUX_s_1_2_2(nor_818_nl, nor_819_nl, fsm_output(5));
  nor_820_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(8)));
  nor_821_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1959_nl <= MUX_s_1_2_2(nor_820_nl, nor_821_nl, fsm_output(5));
  mux_1961_nl <= MUX_s_1_2_2(mux_1960_nl, mux_1959_nl, fsm_output(1));
  nor_822_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_823_nl <= NOT((NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1957_nl <= MUX_s_1_2_2(nor_822_nl, nor_823_nl, fsm_output(5));
  nor_824_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(3))) OR (fsm_output(5)) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(8)));
  mux_1958_nl <= MUX_s_1_2_2(mux_1957_nl, nor_824_nl, fsm_output(1));
  mux_1962_nl <= MUX_s_1_2_2(mux_1961_nl, mux_1958_nl, fsm_output(0));
  nor_825_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (fsm_output(6)) AND (fsm_output(8)))));
  and_848_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (fsm_output(2)) AND CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("110")) AND COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  mux_1954_nl <= MUX_s_1_2_2(nor_825_nl, and_848_nl, fsm_output(5));
  and_856_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (NOT (fsm_output(6))) AND (fsm_output(8));
  nor_828_nl <= NOT((NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND (fsm_output(2)) AND CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm AND (NOT (fsm_output(7))))) OR not_tmp_395);
  mux_1953_nl <= MUX_s_1_2_2(and_856_nl, nor_828_nl, fsm_output(5));
  mux_1955_nl <= MUX_s_1_2_2(mux_1954_nl, mux_1953_nl, fsm_output(1));
  and_864_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm AND (fsm_output(2)) AND (fsm_output(7))
      AND (NOT (fsm_output(6))) AND (fsm_output(8));
  and_865_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (NOT (fsm_output(6))) AND (fsm_output(8));
  mux_1951_nl <= MUX_s_1_2_2(and_864_nl, and_865_nl, fsm_output(5));
  nor_831_nl <= NOT((NOT COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm) OR (COMP_LOOP_acc_1_cse_sva(1))
      OR nand_170_cse);
  nor_832_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm) OR (fsm_output(7)) OR not_tmp_395);
  mux_1949_nl <= MUX_s_1_2_2(nor_831_nl, nor_832_nl, fsm_output(2));
  nor_833_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR not_tmp_395);
  mux_1950_nl <= MUX_s_1_2_2(mux_1949_nl, nor_833_nl, fsm_output(5));
  mux_1952_nl <= MUX_s_1_2_2(mux_1951_nl, mux_1950_nl, fsm_output(1));
  mux_1956_nl <= MUX_s_1_2_2(mux_1955_nl, mux_1952_nl, fsm_output(0));
  mux_1963_nl <= MUX_s_1_2_2(mux_1962_nl, mux_1956_nl, fsm_output(4));
  mux_1945_nl <= MUX_s_1_2_2(nor_860_cse, and_490_cse, fsm_output(2));
  nor_835_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_836_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("010")));
  mux_1944_nl <= MUX_s_1_2_2(nor_835_nl, nor_836_nl, fsm_output(2));
  and_491_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1944_nl;
  mux_1946_nl <= MUX_s_1_2_2(mux_1945_nl, and_491_nl, fsm_output(5));
  mux_1942_nl <= MUX_s_1_2_2(nor_837_cse, nor_838_cse, fsm_output(2));
  and_492_nl <= nor_351_cse AND mux_1941_cse;
  mux_1943_nl <= MUX_s_1_2_2(mux_1942_nl, and_492_nl, fsm_output(5));
  mux_1947_nl <= MUX_s_1_2_2(mux_1946_nl, mux_1943_nl, fsm_output(1));
  nor_840_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8
      DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_841_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("010")));
  mux_1937_nl <= MUX_s_1_2_2(nor_840_nl, nor_841_nl, fsm_output(2));
  nor_842_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  nor_843_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  mux_1936_nl <= MUX_s_1_2_2(nor_842_nl, nor_843_nl, fsm_output(2));
  mux_1938_nl <= MUX_s_1_2_2(mux_1937_nl, mux_1936_nl, fsm_output(5));
  and_495_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm AND CONV_SL_1_1(fsm_output(8 DOWNTO
      6)=STD_LOGIC_VECTOR'("011"));
  nor_844_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("001")));
  mux_1934_nl <= MUX_s_1_2_2(and_495_nl, nor_844_nl, fsm_output(2));
  and_496_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_845_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1933_nl <= MUX_s_1_2_2(and_496_nl, nor_845_nl, fsm_output(2));
  mux_1935_nl <= MUX_s_1_2_2(mux_1934_nl, mux_1933_nl, fsm_output(5));
  mux_1939_nl <= MUX_s_1_2_2(mux_1938_nl, mux_1935_nl, fsm_output(1));
  mux_1948_nl <= MUX_s_1_2_2(mux_1947_nl, mux_1939_nl, fsm_output(0));
  and_489_nl <= (fsm_output(4)) AND mux_1948_nl;
  vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1963_nl, and_489_nl,
      fsm_output(3));
  nor_792_nl <= NOT((NOT (fsm_output(5))) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(3))) OR
      (fsm_output(0)) OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(1)) OR (NOT
      (VEC_LOOP_j_10_0_sva_9_0(1))) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2))) OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  nand_79_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(1)) AND mux_1991_cse);
  nand_156_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111")));
  or_2109_nl <= nand_157_cse OR not_tmp_395;
  mux_1988_nl <= MUX_s_1_2_2(nand_156_nl, or_2109_nl, fsm_output(2));
  nand_158_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011")));
  or_2106_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001"));
  mux_1987_nl <= MUX_s_1_2_2(nand_158_nl, or_2106_nl, fsm_output(2));
  mux_1989_nl <= MUX_s_1_2_2(mux_1988_nl, mux_1987_nl, fsm_output(3));
  mux_1992_nl <= MUX_s_1_2_2(nand_79_nl, mux_1989_nl, fsm_output(1));
  nor_793_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1992_nl);
  nor_797_nl <= NOT((NOT (COMP_LOOP_acc_10_cse_10_1_15_sva(2))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_15_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_15_sva(0)) OR nand_268_cse);
  nor_798_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1984_nl <= MUX_s_1_2_2(nor_797_nl, nor_798_nl, fsm_output(2));
  and_486_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_799_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1983_nl <= MUX_s_1_2_2(and_486_nl, nor_799_nl, fsm_output(2));
  mux_1985_nl <= MUX_s_1_2_2(mux_1984_nl, mux_1983_nl, fsm_output(3));
  and_839_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  nor_801_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1981_nl <= MUX_s_1_2_2(and_839_nl, nor_801_nl, fsm_output(2));
  nor_802_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_803_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1980_nl <= MUX_s_1_2_2(nor_802_nl, nor_803_nl, fsm_output(2));
  mux_1982_nl <= MUX_s_1_2_2(mux_1981_nl, mux_1980_nl, fsm_output(3));
  mux_1986_nl <= MUX_s_1_2_2(mux_1985_nl, mux_1982_nl, fsm_output(1));
  mux_1993_nl <= MUX_s_1_2_2(nor_793_nl, mux_1986_nl, fsm_output(0));
  nor_804_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_sva(0)) OR (NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3
      DOWNTO 1)=STD_LOGIC_VECTOR'("111")) AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111")))));
  nor_805_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1976_nl <= MUX_s_1_2_2(nor_804_nl, nor_805_nl, fsm_output(2));
  and_487_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_806_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1975_nl <= MUX_s_1_2_2(and_487_nl, nor_806_nl, fsm_output(2));
  mux_1977_nl <= MUX_s_1_2_2(mux_1976_nl, mux_1975_nl, fsm_output(3));
  and_847_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  nor_808_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1973_nl <= MUX_s_1_2_2(and_847_nl, nor_808_nl, fsm_output(2));
  nor_809_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_810_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1972_nl <= MUX_s_1_2_2(nor_809_nl, nor_810_nl, fsm_output(2));
  mux_1974_nl <= MUX_s_1_2_2(mux_1973_nl, mux_1972_nl, fsm_output(3));
  mux_1978_nl <= MUX_s_1_2_2(mux_1977_nl, mux_1974_nl, fsm_output(1));
  nor_811_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))))
      OR nand_324_cse);
  nor_812_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(7)) OR not_tmp_395);
  mux_1969_nl <= MUX_s_1_2_2(nor_811_nl, nor_812_nl, fsm_output(2));
  and_488_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_813_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_1968_nl <= MUX_s_1_2_2(and_488_nl, nor_813_nl, fsm_output(2));
  mux_1970_nl <= MUX_s_1_2_2(mux_1969_nl, mux_1968_nl, fsm_output(3));
  and_863_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  nor_815_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("100")));
  mux_1966_nl <= MUX_s_1_2_2(and_863_nl, nor_815_nl, fsm_output(2));
  nor_816_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("010")));
  nor_817_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_1965_nl <= MUX_s_1_2_2(nor_816_nl, nor_817_nl, fsm_output(2));
  mux_1967_nl <= MUX_s_1_2_2(mux_1966_nl, mux_1965_nl, fsm_output(3));
  mux_1971_nl <= MUX_s_1_2_2(mux_1970_nl, mux_1967_nl, fsm_output(1));
  mux_1979_nl <= MUX_s_1_2_2(mux_1978_nl, mux_1971_nl, fsm_output(0));
  mux_1994_nl <= MUX_s_1_2_2(mux_1993_nl, mux_1979_nl, fsm_output(5));
  vec_rsc_0_14_i_we_d_pff <= MUX_s_1_2_2(nor_792_nl, mux_1994_nl, fsm_output(4));
  nor_769_nl <= NOT((NOT((fsm_output(5)) AND (fsm_output(2)) AND (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      AND CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm)) OR nand_301_cse);
  nor_770_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_771_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_sva(0)) OR (NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3
      DOWNTO 1)=STD_LOGIC_VECTOR'("111")) AND (fsm_output(7)) AND (fsm_output(4))
      AND (fsm_output(8)))));
  mux_2021_nl <= MUX_s_1_2_2(nor_770_nl, nor_771_nl, fsm_output(2));
  nor_772_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_2022_nl <= MUX_s_1_2_2(mux_2021_nl, nor_772_nl, fsm_output(5));
  mux_2023_nl <= MUX_s_1_2_2(nor_769_nl, mux_2022_nl, fsm_output(6));
  nor_773_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_774_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))))
      OR nand_301_cse);
  mux_2018_nl <= MUX_s_1_2_2(nor_773_nl, nor_774_nl, fsm_output(2));
  nor_775_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  mux_2019_nl <= MUX_s_1_2_2(mux_2018_nl, nor_775_nl, fsm_output(5));
  nor_776_nl <= NOT((NOT((VEC_LOOP_j_10_0_sva_9_0(1)) AND (fsm_output(5)) AND (fsm_output(2))
      AND CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm AND (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      AND (NOT (fsm_output(7))))) OR not_tmp_399);
  mux_2020_nl <= MUX_s_1_2_2(mux_2019_nl, nor_776_nl, fsm_output(6));
  mux_2024_nl <= MUX_s_1_2_2(mux_2023_nl, mux_2020_nl, fsm_output(1));
  nor_777_nl <= NOT((NOT((fsm_output(2)) AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1110")) AND COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm))
      OR nand_301_cse);
  nor_778_nl <= NOT((NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(7)) OR (fsm_output(4))
      OR (fsm_output(8)));
  nor_779_nl <= NOT((NOT (COMP_LOOP_acc_10_cse_10_1_15_sva(2))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_15_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_15_sva(0)) OR nand_265_cse);
  mux_2014_nl <= MUX_s_1_2_2(nor_778_nl, nor_779_nl, fsm_output(2));
  mux_2015_nl <= MUX_s_1_2_2(nor_777_nl, mux_2014_nl, fsm_output(5));
  nor_780_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(4))
      OR (fsm_output(8)));
  mux_2016_nl <= MUX_s_1_2_2(mux_2015_nl, nor_780_nl, fsm_output(6));
  nor_781_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(1))) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(3)))
      OR (fsm_output(5)) OR (fsm_output(2)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  nor_782_nl <= NOT((NOT(COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1110")))) OR nand_301_cse);
  nor_783_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm) OR (fsm_output(7)) OR not_tmp_399);
  mux_2011_nl <= MUX_s_1_2_2(nor_782_nl, nor_783_nl, fsm_output(2));
  nor_784_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR not_tmp_399);
  mux_2012_nl <= MUX_s_1_2_2(mux_2011_nl, nor_784_nl, fsm_output(5));
  mux_2013_nl <= MUX_s_1_2_2(nor_781_nl, mux_2012_nl, fsm_output(6));
  mux_2017_nl <= MUX_s_1_2_2(mux_2016_nl, mux_2013_nl, fsm_output(1));
  mux_2025_nl <= MUX_s_1_2_2(mux_2024_nl, mux_2017_nl, fsm_output(0));
  nor_785_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (NOT COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (fsm_output(7)) OR not_tmp_399);
  and_480_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm AND (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      AND (fsm_output(7)) AND (fsm_output(4)) AND (NOT (fsm_output(8)));
  mux_2007_nl <= MUX_s_1_2_2(nor_785_nl, and_480_nl, fsm_output(2));
  and_479_nl <= (fsm_output(5)) AND mux_2007_nl;
  or_2136_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(7)) OR not_tmp_399;
  nand_149_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(7)) AND (fsm_output(4)) AND (NOT (fsm_output(8))));
  mux_2006_nl <= MUX_s_1_2_2(or_2136_nl, nand_149_nl, fsm_output(2));
  nor_786_nl <= NOT((fsm_output(5)) OR mux_2006_nl);
  mux_2008_nl <= MUX_s_1_2_2(and_479_nl, nor_786_nl, fsm_output(6));
  or_2132_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(7)) OR not_tmp_399;
  nand_150_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(7)) AND (fsm_output(4)) AND (NOT (fsm_output(8))));
  mux_2004_nl <= MUX_s_1_2_2(or_2132_nl, nand_150_nl, fsm_output(2));
  nor_787_nl <= NOT((fsm_output(5)) OR mux_2004_nl);
  and_481_nl <= (VEC_LOOP_j_10_0_sva_9_0(1)) AND (fsm_output(5)) AND mux_1878_cse;
  mux_2005_nl <= MUX_s_1_2_2(nor_787_nl, and_481_nl, fsm_output(6));
  mux_2009_nl <= MUX_s_1_2_2(mux_2008_nl, mux_2005_nl, fsm_output(1));
  or_2126_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm) OR (fsm_output(7)) OR not_tmp_399;
  nand_151_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND (fsm_output(7)) AND (fsm_output(4))
      AND (NOT (fsm_output(8))));
  mux_2000_nl <= MUX_s_1_2_2(or_2126_nl, nand_151_nl, fsm_output(2));
  or_2123_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(7)) OR not_tmp_399;
  nand_152_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(7)) AND (fsm_output(4)) AND (NOT (fsm_output(8))));
  mux_1999_nl <= MUX_s_1_2_2(or_2123_nl, nand_152_nl, fsm_output(2));
  mux_2001_nl <= MUX_s_1_2_2(mux_2000_nl, mux_1999_nl, fsm_output(5));
  nor_789_nl <= NOT((fsm_output(6)) OR mux_2001_nl);
  and_484_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm AND (fsm_output(7)) AND (fsm_output(4))
      AND (NOT (fsm_output(8)));
  nor_790_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR (fsm_output(7)) OR (NOT (fsm_output(4)))
      OR (fsm_output(8)));
  mux_1997_nl <= MUX_s_1_2_2(and_484_nl, nor_790_nl, fsm_output(2));
  and_485_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(7)) AND (fsm_output(4)) AND (NOT (fsm_output(8)));
  nor_791_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(7)) OR (NOT (fsm_output(4))) OR (fsm_output(8)));
  mux_1996_nl <= MUX_s_1_2_2(and_485_nl, nor_791_nl, fsm_output(2));
  mux_1998_nl <= MUX_s_1_2_2(mux_1997_nl, mux_1996_nl, fsm_output(5));
  and_483_nl <= (fsm_output(6)) AND mux_1998_nl;
  mux_2002_nl <= MUX_s_1_2_2(nor_789_nl, and_483_nl, fsm_output(1));
  mux_2010_nl <= MUX_s_1_2_2(mux_2009_nl, mux_2002_nl, fsm_output(0));
  vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_2025_nl, mux_2010_nl,
      fsm_output(3));
  nor_751_nl <= NOT((NOT (fsm_output(5))) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(3))) OR
      (fsm_output(0)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(1)) OR
      (NOT (VEC_LOOP_j_10_0_sva_9_0(1))) OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2))) OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  and_464_nl <= (VEC_LOOP_j_10_0_sva_9_0(1)) AND mux_1991_cse;
  and_465_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111"));
  nor_755_nl <= NOT(nand_157_cse OR not_tmp_395);
  mux_2050_nl <= MUX_s_1_2_2(and_465_nl, nor_755_nl, fsm_output(2));
  and_466_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  nor_756_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("001")));
  mux_2049_nl <= MUX_s_1_2_2(and_466_nl, nor_756_nl, fsm_output(2));
  mux_2051_nl <= MUX_s_1_2_2(mux_2050_nl, mux_2049_nl, fsm_output(3));
  mux_2054_nl <= MUX_s_1_2_2(and_464_nl, mux_2051_nl, fsm_output(1));
  and_463_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_2054_nl;
  and_467_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111"));
  nor_757_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(7))))) OR not_tmp_395);
  mux_2046_nl <= MUX_s_1_2_2(and_467_nl, nor_757_nl, fsm_output(2));
  and_468_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  and_469_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("001"));
  mux_2045_nl <= MUX_s_1_2_2(and_468_nl, and_469_nl, fsm_output(2));
  mux_2047_nl <= MUX_s_1_2_2(mux_2046_nl, mux_2045_nl, fsm_output(3));
  and_838_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  and_844_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("100"));
  mux_2043_nl <= MUX_s_1_2_2(and_838_nl, and_844_nl, fsm_output(2));
  and_470_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("010"));
  nor_760_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_2042_nl <= MUX_s_1_2_2(and_470_nl, nor_760_nl, fsm_output(2));
  mux_2044_nl <= MUX_s_1_2_2(mux_2043_nl, mux_2042_nl, fsm_output(3));
  mux_2048_nl <= MUX_s_1_2_2(mux_2047_nl, mux_2044_nl, fsm_output(1));
  mux_2055_nl <= MUX_s_1_2_2(and_463_nl, mux_2048_nl, fsm_output(0));
  and_471_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111"));
  mux_2038_nl <= MUX_s_1_2_2(and_471_nl, nor_761_cse, fsm_output(2));
  and_473_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("001"));
  mux_2037_nl <= MUX_s_1_2_2(and_450_cse, and_473_nl, fsm_output(2));
  mux_2039_nl <= MUX_s_1_2_2(mux_2038_nl, mux_2037_nl, fsm_output(3));
  and_846_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  mux_2035_nl <= MUX_s_1_2_2(and_846_nl, and_836_cse, fsm_output(2));
  nor_764_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_2034_nl <= MUX_s_1_2_2(and_453_cse, nor_764_nl, fsm_output(2));
  mux_2036_nl <= MUX_s_1_2_2(mux_2035_nl, mux_2034_nl, fsm_output(3));
  mux_2040_nl <= MUX_s_1_2_2(mux_2039_nl, mux_2036_nl, fsm_output(1));
  and_475_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111"));
  nor_765_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(7))))) OR not_tmp_395);
  mux_2031_nl <= MUX_s_1_2_2(and_475_nl, nor_765_nl, fsm_output(2));
  and_476_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  and_477_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("001"));
  mux_2030_nl <= MUX_s_1_2_2(and_476_nl, and_477_nl, fsm_output(2));
  mux_2032_nl <= MUX_s_1_2_2(mux_2031_nl, mux_2030_nl, fsm_output(3));
  and_861_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  and_862_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("100"));
  mux_2028_nl <= MUX_s_1_2_2(and_861_nl, and_862_nl, fsm_output(2));
  and_478_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("010"));
  nor_768_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  mux_2027_nl <= MUX_s_1_2_2(and_478_nl, nor_768_nl, fsm_output(2));
  mux_2029_nl <= MUX_s_1_2_2(mux_2028_nl, mux_2027_nl, fsm_output(3));
  mux_2033_nl <= MUX_s_1_2_2(mux_2032_nl, mux_2029_nl, fsm_output(1));
  mux_2041_nl <= MUX_s_1_2_2(mux_2040_nl, mux_2033_nl, fsm_output(0));
  mux_2056_nl <= MUX_s_1_2_2(mux_2055_nl, mux_2041_nl, fsm_output(5));
  vec_rsc_0_15_i_we_d_pff <= MUX_s_1_2_2(nor_751_nl, mux_2056_nl, fsm_output(4));
  nor_731_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111")) OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_732_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  mux_2085_nl <= MUX_s_1_2_2(nor_731_nl, nor_732_nl, fsm_output(5));
  nor_733_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(8)));
  nor_734_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(8)));
  mux_2084_nl <= MUX_s_1_2_2(nor_733_nl, nor_734_nl, fsm_output(5));
  mux_2086_nl <= MUX_s_1_2_2(mux_2085_nl, mux_2084_nl, fsm_output(1));
  nor_735_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(8)));
  nor_736_nl <= NOT((NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1111")) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(8)));
  mux_2082_nl <= MUX_s_1_2_2(nor_735_nl, nor_736_nl, fsm_output(5));
  nor_737_nl <= NOT((NOT (VEC_LOOP_j_10_0_sva_9_0(3))) OR (fsm_output(5)) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111")) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(8)));
  mux_2083_nl <= MUX_s_1_2_2(mux_2082_nl, nor_737_nl, fsm_output(1));
  mux_2087_nl <= MUX_s_1_2_2(mux_2086_nl, mux_2083_nl, fsm_output(0));
  and_447_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (fsm_output(6)) AND (fsm_output(8));
  and_845_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (fsm_output(2)) AND CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("110"));
  mux_2079_nl <= MUX_s_1_2_2(and_447_nl, and_845_nl, fsm_output(5));
  and_854_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (NOT (fsm_output(6))) AND (fsm_output(8));
  nor_740_nl <= NOT((NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(2)) AND CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm AND (NOT (fsm_output(7))))) OR not_tmp_395);
  mux_2078_nl <= MUX_s_1_2_2(and_854_nl, nor_740_nl, fsm_output(5));
  mux_2080_nl <= MUX_s_1_2_2(mux_2079_nl, mux_2078_nl, fsm_output(1));
  and_859_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm AND (fsm_output(2)) AND (fsm_output(7))
      AND (NOT (fsm_output(6))) AND (fsm_output(8));
  and_860_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_15_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(2)) AND (fsm_output(7)) AND (NOT (fsm_output(6))) AND (fsm_output(8));
  mux_2076_nl <= MUX_s_1_2_2(and_859_nl, and_860_nl, fsm_output(5));
  and_448_nl <= COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111"));
  nor_743_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm AND (NOT (fsm_output(7))))) OR not_tmp_395);
  mux_2074_nl <= MUX_s_1_2_2(and_448_nl, nor_743_nl, fsm_output(2));
  nor_744_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_13_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(2)) AND (NOT (fsm_output(7))))) OR not_tmp_395);
  mux_2075_nl <= MUX_s_1_2_2(mux_2074_nl, nor_744_nl, fsm_output(5));
  mux_2077_nl <= MUX_s_1_2_2(mux_2076_nl, mux_2075_nl, fsm_output(1));
  mux_2081_nl <= MUX_s_1_2_2(mux_2080_nl, mux_2077_nl, fsm_output(0));
  mux_2088_nl <= MUX_s_1_2_2(mux_2087_nl, mux_2081_nl, fsm_output(4));
  mux_2070_nl <= MUX_s_1_2_2(nor_761_cse, and_450_cse, fsm_output(2));
  and_833_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(8 DOWNTO
      6)=STD_LOGIC_VECTOR'("100"));
  and_452_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(8 DOWNTO
      6)=STD_LOGIC_VECTOR'("010"));
  mux_2069_nl <= MUX_s_1_2_2(and_833_nl, and_452_nl, fsm_output(2));
  and_451_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_2069_nl;
  mux_2071_nl <= MUX_s_1_2_2(mux_2070_nl, and_451_nl, fsm_output(5));
  mux_2067_nl <= MUX_s_1_2_2(and_836_cse, and_453_cse, fsm_output(2));
  and_454_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND mux_1941_cse;
  mux_2068_nl <= MUX_s_1_2_2(mux_2067_nl, and_454_nl, fsm_output(5));
  mux_2072_nl <= MUX_s_1_2_2(mux_2071_nl, mux_2068_nl, fsm_output(1));
  and_837_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(8 DOWNTO
      6)=STD_LOGIC_VECTOR'("100"));
  and_457_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(8 DOWNTO
      6)=STD_LOGIC_VECTOR'("010"));
  mux_2062_nl <= MUX_s_1_2_2(and_837_nl, and_457_nl, fsm_output(2));
  and_843_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_11_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("100"));
  and_458_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("010"));
  mux_2061_nl <= MUX_s_1_2_2(and_843_nl, and_458_nl, fsm_output(2));
  mux_2063_nl <= MUX_s_1_2_2(mux_2062_nl, mux_2061_nl, fsm_output(5));
  and_459_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm AND CONV_SL_1_1(fsm_output(8 DOWNTO
      6)=STD_LOGIC_VECTOR'("011"));
  and_460_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm AND CONV_SL_1_1(fsm_output(8 DOWNTO
      6)=STD_LOGIC_VECTOR'("001"));
  mux_2059_nl <= MUX_s_1_2_2(and_459_nl, and_460_nl, fsm_output(2));
  and_461_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_9_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("011"));
  and_462_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("001"));
  mux_2058_nl <= MUX_s_1_2_2(and_461_nl, and_462_nl, fsm_output(2));
  mux_2060_nl <= MUX_s_1_2_2(mux_2059_nl, mux_2058_nl, fsm_output(5));
  mux_2064_nl <= MUX_s_1_2_2(mux_2063_nl, mux_2060_nl, fsm_output(1));
  mux_2073_nl <= MUX_s_1_2_2(mux_2072_nl, mux_2064_nl, fsm_output(0));
  and_449_nl <= (fsm_output(4)) AND mux_2073_nl;
  vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_2088_nl, and_449_nl,
      fsm_output(3));
  COMP_LOOP_1_tmp_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( UNSIGNED(COMP_LOOP_1_tmp_lshift_itm)
      * UNSIGNED(COMP_LOOP_k_10_4_sva_5_0)), 6));
  twiddle_rsc_0_0_i_radr_d <= MUX1HOT_v_6_6_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_1_tmp_mul_nl),
      6)), (COMP_LOOP_10_tmp_mul_idiv_sva(9 DOWNTO 4)), (COMP_LOOP_11_tmp_mul_idiv_sva(8
      DOWNTO 3)), (COMP_LOOP_5_tmp_mul_idiv_sva(7 DOWNTO 2)), (COMP_LOOP_9_tmp_lshift_itm(6
      DOWNTO 1)), (COMP_LOOP_13_tmp_mul_idiv_sva(7 DOWNTO 2)), STD_LOGIC_VECTOR'(
      and_dcpl_62 & and_dcpl_175 & and_dcpl_180 & and_dcpl_181 & and_dcpl_183 & and_dcpl_184));
  mux_2095_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), (fsm_output(4)), or_2259_cse_1);
  or_2260_nl <= CONV_SL_1_1(COMP_LOOP_11_tmp_mul_idiv_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR mux_2095_nl;
  or_2257_nl <= (NOT (fsm_output(4))) OR CONV_SL_1_1(COMP_LOOP_10_tmp_mul_idiv_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"));
  mux_2094_nl <= MUX_s_1_2_2(or_2257_nl, or_tmp_2077, or_2259_cse_1);
  mux_2096_nl <= MUX_s_1_2_2(or_2260_nl, mux_2094_nl, fsm_output(0));
  or_2255_nl <= CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(4));
  mux_2091_nl <= MUX_s_1_2_2((fsm_output(4)), or_2255_nl, fsm_output(2));
  or_2254_nl <= (COMP_LOOP_9_tmp_lshift_itm(0)) OR (fsm_output(4));
  or_2253_nl <= CONV_SL_1_1(COMP_LOOP_13_tmp_mul_idiv_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(4));
  mux_2090_nl <= MUX_s_1_2_2(or_2254_nl, or_2253_nl, fsm_output(2));
  mux_2092_nl <= MUX_s_1_2_2(mux_2091_nl, mux_2090_nl, fsm_output(3));
  mux_2093_nl <= MUX_s_1_2_2(mux_2092_nl, or_tmp_2077, fsm_output(0));
  mux_2097_nl <= MUX_s_1_2_2(mux_2096_nl, mux_2093_nl, fsm_output(1));
  twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2097_nl) AND and_dcpl_186;
  twiddle_rsc_0_1_i_radr_d_pff <= z_out_3(9 DOWNTO 4);
  nor_724_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(4)));
  nor_723_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")) OR
      nand_122_cse);
  mux_2102_nl <= MUX_s_1_2_2(nor_723_nl, nor_724_cse, fsm_output(1));
  mux_2103_nl <= MUX_s_1_2_2(mux_2102_nl, nor_724_cse, fsm_output(2));
  mux_2104_nl <= MUX_s_1_2_2(mux_2103_nl, nor_724_cse, fsm_output(3));
  twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2104_nl AND and_dcpl_193;
  twiddle_rsc_0_2_i_radr_d_pff <= MUX_v_6_2_2((z_out_3(9 DOWNTO 4)), (z_out_3(8 DOWNTO
      3)), COMP_LOOP_tmp_or_19_cse);
  nor_712_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(4)));
  nor_711_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR
      (NOT (fsm_output(4))));
  mux_2112_nl <= MUX_s_1_2_2(nor_711_nl, nor_712_cse, fsm_output(2));
  mux_2113_nl <= MUX_s_1_2_2(mux_2112_nl, nor_712_cse, fsm_output(1));
  mux_2114_nl <= MUX_s_1_2_2(mux_2113_nl, nor_712_cse, fsm_output(3));
  and_445_nl <= (fsm_output(1)) AND (NOT(CONV_SL_1_1(z_out_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(4))));
  mux_2115_nl <= MUX_s_1_2_2(mux_2114_nl, and_445_nl, fsm_output(0));
  twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2115_nl AND and_dcpl_186;
  nor_704_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(4)));
  nor_703_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")) OR
      nand_121_cse);
  mux_2120_nl <= MUX_s_1_2_2(nor_703_nl, nor_704_cse, fsm_output(1));
  mux_2121_nl <= MUX_s_1_2_2(mux_2120_nl, nor_704_cse, fsm_output(2));
  mux_2122_nl <= MUX_s_1_2_2(mux_2121_nl, nor_704_cse, fsm_output(3));
  twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2122_nl AND and_dcpl_193;
  COMP_LOOP_tmp_or_46_cse <= (and_dcpl_188 AND and_dcpl_64) OR and_dcpl_202;
  twiddle_rsc_0_4_i_radr_d_pff <= MUX1HOT_v_6_3_2((z_out_3(9 DOWNTO 4)), (z_out_3(8
      DOWNTO 3)), (z_out_3(7 DOWNTO 2)), STD_LOGIC_VECTOR'( COMP_LOOP_tmp_or_1_cse
      & COMP_LOOP_tmp_or_19_cse & COMP_LOOP_tmp_or_46_cse));
  nor_691_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(4)));
  nor_692_nl <= NOT(CONV_SL_1_1(z_out_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR
      (fsm_output(4)));
  mux_2131_cse <= MUX_s_1_2_2(nor_691_cse, nor_692_nl, fsm_output(0));
  nor_689_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR
      (fsm_output(0)) OR (NOT (fsm_output(4))));
  nor_690_nl <= NOT((fsm_output(0)) OR CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(4)));
  mux_2133_nl <= MUX_s_1_2_2(nor_689_nl, nor_690_nl, fsm_output(3));
  mux_2134_nl <= MUX_s_1_2_2(mux_2133_nl, mux_2131_cse, fsm_output(1));
  nor_696_nl <= NOT(CONV_SL_1_1(z_out_3(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (fsm_output(4)));
  mux_2127_nl <= MUX_s_1_2_2(nor_691_cse, nor_696_nl, fsm_output(0));
  mux_2129_nl <= MUX_s_1_2_2(mux_2127_nl, mux_2131_cse, fsm_output(1));
  mux_2135_nl <= MUX_s_1_2_2(mux_2134_nl, mux_2129_nl, fsm_output(2));
  twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2135_nl AND and_dcpl_186;
  nor_682_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(4)));
  nor_681_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010")) OR
      nand_122_cse);
  mux_2140_nl <= MUX_s_1_2_2(nor_681_nl, nor_682_cse, fsm_output(1));
  mux_2141_nl <= MUX_s_1_2_2(mux_2140_nl, nor_682_cse, fsm_output(2));
  mux_2142_nl <= MUX_s_1_2_2(mux_2141_nl, nor_682_cse, fsm_output(3));
  twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2142_nl AND and_dcpl_193;
  nor_670_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(4)));
  nor_669_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR
      (NOT (fsm_output(4))));
  mux_2150_nl <= MUX_s_1_2_2(nor_669_nl, nor_670_cse, fsm_output(2));
  mux_2151_nl <= MUX_s_1_2_2(mux_2150_nl, nor_670_cse, fsm_output(1));
  mux_2152_nl <= MUX_s_1_2_2(mux_2151_nl, nor_670_cse, fsm_output(3));
  and_443_nl <= (fsm_output(1)) AND (NOT(CONV_SL_1_1(z_out_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(4))));
  mux_2153_nl <= MUX_s_1_2_2(mux_2152_nl, and_443_nl, fsm_output(0));
  twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2153_nl AND and_dcpl_186;
  nor_662_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(4)));
  nor_661_nl <= NOT((z_out_3(3)) OR (NOT(CONV_SL_1_1(z_out_3(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(4)))));
  mux_2158_nl <= MUX_s_1_2_2(nor_661_nl, nor_662_cse, fsm_output(1));
  mux_2159_nl <= MUX_s_1_2_2(mux_2158_nl, nor_662_cse, fsm_output(2));
  mux_2160_nl <= MUX_s_1_2_2(mux_2159_nl, nor_662_cse, fsm_output(3));
  twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2160_nl AND and_dcpl_193;
  twiddle_rsc_0_8_i_radr_d <= MUX1HOT_v_6_4_2((z_out_3(9 DOWNTO 4)), (z_out_3(8 DOWNTO
      3)), (z_out_3(7 DOWNTO 2)), (z_out_3(6 DOWNTO 1)), STD_LOGIC_VECTOR'( COMP_LOOP_tmp_or_1_cse
      & COMP_LOOP_tmp_or_19_cse & COMP_LOOP_tmp_or_46_cse & and_dcpl_207));
  nor_647_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(4)));
  nor_650_nl <= NOT(CONV_SL_1_1(z_out_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR
      (fsm_output(4)));
  mux_2169_cse <= MUX_s_1_2_2(nor_647_cse, nor_650_nl, fsm_output(0));
  nor_646_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR
      (fsm_output(0)) OR (NOT (fsm_output(4))));
  nor_648_nl <= NOT((NOT (z_out_3(0))) OR (fsm_output(4)));
  mux_2171_nl <= MUX_s_1_2_2(nor_647_cse, nor_648_nl, fsm_output(0));
  mux_2172_nl <= MUX_s_1_2_2(nor_646_nl, mux_2171_nl, fsm_output(3));
  mux_2173_nl <= MUX_s_1_2_2(mux_2172_nl, mux_2169_cse, fsm_output(1));
  nor_654_nl <= NOT(CONV_SL_1_1(z_out_3(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (fsm_output(4)));
  mux_2165_nl <= MUX_s_1_2_2(nor_647_cse, nor_654_nl, fsm_output(0));
  mux_2167_nl <= MUX_s_1_2_2(mux_2165_nl, mux_2169_cse, fsm_output(1));
  mux_2174_nl <= MUX_s_1_2_2(mux_2173_nl, mux_2167_nl, fsm_output(2));
  twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2174_nl AND and_dcpl_186;
  nor_639_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(4)));
  nor_638_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("100")) OR
      nand_122_cse);
  mux_2179_nl <= MUX_s_1_2_2(nor_638_nl, nor_639_cse, fsm_output(1));
  mux_2180_nl <= MUX_s_1_2_2(mux_2179_nl, nor_639_cse, fsm_output(2));
  mux_2181_nl <= MUX_s_1_2_2(mux_2180_nl, nor_639_cse, fsm_output(3));
  twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2181_nl AND and_dcpl_193;
  nor_627_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(4)));
  nor_626_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR
      (NOT (fsm_output(4))));
  mux_2189_nl <= MUX_s_1_2_2(nor_626_nl, nor_627_cse, fsm_output(2));
  mux_2190_nl <= MUX_s_1_2_2(mux_2189_nl, nor_627_cse, fsm_output(1));
  mux_2191_nl <= MUX_s_1_2_2(mux_2190_nl, nor_627_cse, fsm_output(3));
  and_441_nl <= (fsm_output(1)) AND (NOT(CONV_SL_1_1(z_out_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(4))));
  mux_2192_nl <= MUX_s_1_2_2(mux_2191_nl, and_441_nl, fsm_output(0));
  twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2192_nl AND and_dcpl_186;
  nor_619_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(4)));
  nor_618_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10")) OR
      nand_121_cse);
  mux_2197_nl <= MUX_s_1_2_2(nor_618_nl, nor_619_cse, fsm_output(1));
  mux_2198_nl <= MUX_s_1_2_2(mux_2197_nl, nor_619_cse, fsm_output(2));
  mux_2199_nl <= MUX_s_1_2_2(mux_2198_nl, nor_619_cse, fsm_output(3));
  twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2199_nl AND and_dcpl_193;
  nor_606_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(4)));
  nor_607_nl <= NOT(CONV_SL_1_1(z_out_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR
      (fsm_output(4)));
  mux_2208_cse <= MUX_s_1_2_2(nor_606_cse, nor_607_nl, fsm_output(0));
  nor_604_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR
      (fsm_output(0)) OR (NOT (fsm_output(4))));
  nor_605_nl <= NOT((fsm_output(0)) OR CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(4)));
  mux_2210_nl <= MUX_s_1_2_2(nor_604_nl, nor_605_nl, fsm_output(3));
  mux_2211_nl <= MUX_s_1_2_2(mux_2210_nl, mux_2208_cse, fsm_output(1));
  nor_611_nl <= NOT(CONV_SL_1_1(z_out_3(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (fsm_output(4)));
  mux_2204_nl <= MUX_s_1_2_2(nor_606_cse, nor_611_nl, fsm_output(0));
  mux_2206_nl <= MUX_s_1_2_2(mux_2204_nl, mux_2208_cse, fsm_output(1));
  mux_2212_nl <= MUX_s_1_2_2(mux_2211_nl, mux_2206_nl, fsm_output(2));
  twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2212_nl AND and_dcpl_186;
  nor_597_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(4)));
  nor_596_nl <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("110")) OR
      nand_122_cse);
  mux_2217_nl <= MUX_s_1_2_2(nor_596_nl, nor_597_cse, fsm_output(1));
  mux_2218_nl <= MUX_s_1_2_2(mux_2217_nl, nor_597_cse, fsm_output(2));
  mux_2219_nl <= MUX_s_1_2_2(mux_2218_nl, nor_597_cse, fsm_output(3));
  twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2219_nl AND and_dcpl_193;
  nor_589_cse <= NOT(CONV_SL_1_1(z_out_3(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(4)));
  and_434_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110")) AND (fsm_output(4));
  mux_2227_nl <= MUX_s_1_2_2(and_434_nl, nor_589_cse, fsm_output(2));
  mux_2228_nl <= MUX_s_1_2_2(mux_2227_nl, nor_589_cse, fsm_output(1));
  mux_2229_nl <= MUX_s_1_2_2(mux_2228_nl, nor_589_cse, fsm_output(3));
  and_435_nl <= (fsm_output(1)) AND CONV_SL_1_1(z_out_3(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (NOT (fsm_output(4)));
  mux_2230_nl <= MUX_s_1_2_2(mux_2229_nl, and_435_nl, fsm_output(0));
  twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2230_nl AND and_dcpl_186;
  and_427_cse <= CONV_SL_1_1(z_out_3(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND (NOT
      (fsm_output(4)));
  and_426_nl <= CONV_SL_1_1(z_out_3(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(4));
  mux_2235_nl <= MUX_s_1_2_2(and_426_nl, and_427_cse, fsm_output(1));
  mux_2236_nl <= MUX_s_1_2_2(mux_2235_nl, and_427_cse, fsm_output(2));
  mux_2237_nl <= MUX_s_1_2_2(mux_2236_nl, and_427_cse, fsm_output(3));
  twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2237_nl AND and_dcpl_193;
  and_dcpl_356 <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111")) AND
      nor_1624_cse AND (fsm_output(1)) AND (fsm_output(0)) AND (fsm_output(4)) AND
      (fsm_output(5));
  and_dcpl_360 <= mux_2465_cse AND nor_1624_cse AND (fsm_output(0)) AND (NOT (fsm_output(5)));
  and_dcpl_362 <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_366 <= and_dcpl_5 AND nor_1624_cse;
  and_dcpl_367 <= and_dcpl_366 AND and_dcpl_362 AND CONV_SL_1_1(fsm_output(5 DOWNTO
      4)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_370 <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      and_dcpl_45;
  and_dcpl_373 <= nor_1630_cse AND (fsm_output(6)) AND and_570_cse;
  and_dcpl_374 <= and_dcpl_373 AND and_dcpl_370;
  and_dcpl_376 <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_377 <= and_dcpl_376 AND and_dcpl_66;
  and_dcpl_378 <= and_dcpl_373 AND and_dcpl_377;
  and_dcpl_380 <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01")) AND
      and_dcpl_45;
  and_dcpl_383 <= and_dcpl_87 AND (NOT (fsm_output(6))) AND and_570_cse;
  and_dcpl_384 <= and_dcpl_383 AND and_dcpl_380;
  and_dcpl_385 <= and_dcpl_362 AND and_dcpl_66;
  and_dcpl_386 <= and_dcpl_383 AND and_dcpl_385;
  and_dcpl_387 <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_389 <= and_dcpl_87 AND (fsm_output(6)) AND and_dcpl_387;
  and_dcpl_390 <= and_dcpl_389 AND and_dcpl_370;
  and_dcpl_391 <= and_dcpl_389 AND and_dcpl_377;
  and_dcpl_394 <= and_dcpl_103 AND (NOT (fsm_output(6))) AND and_dcpl_387;
  and_dcpl_395 <= and_dcpl_394 AND and_dcpl_380;
  and_dcpl_396 <= and_dcpl_394 AND and_dcpl_385;
  and_dcpl_397 <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_399 <= and_dcpl_103 AND (fsm_output(6)) AND and_dcpl_397;
  and_dcpl_400 <= and_dcpl_399 AND and_dcpl_370;
  and_dcpl_401 <= and_dcpl_399 AND and_dcpl_377;
  and_dcpl_404 <= and_733_cse AND (NOT (fsm_output(6))) AND and_dcpl_397;
  and_dcpl_405 <= and_dcpl_404 AND and_dcpl_380;
  and_dcpl_406 <= and_dcpl_404 AND and_dcpl_385;
  and_dcpl_409 <= and_733_cse AND (fsm_output(6)) AND nor_1624_cse AND and_dcpl_377;
  and_dcpl_410 <= and_dcpl_376 AND and_dcpl_45;
  and_dcpl_411 <= and_dcpl_366 AND and_dcpl_410;
  and_dcpl_412 <= and_dcpl_5 AND and_dcpl_387;
  and_dcpl_413 <= and_dcpl_412 AND and_dcpl_380;
  and_dcpl_414 <= and_dcpl_362 AND and_dcpl_45;
  and_dcpl_415 <= and_dcpl_5 AND and_dcpl_397;
  and_dcpl_416 <= and_dcpl_415 AND and_dcpl_414;
  and_dcpl_417 <= and_dcpl_415 AND and_dcpl_410;
  and_dcpl_418 <= and_dcpl_412 AND and_dcpl_414;
  and_dcpl_419 <= and_dcpl_412 AND and_dcpl_410;
  and_dcpl_420 <= and_dcpl_5 AND and_570_cse;
  and_dcpl_421 <= and_dcpl_420 AND and_dcpl_414;
  and_dcpl_422 <= and_dcpl_420 AND and_dcpl_410;
  and_dcpl_425 <= and_dcpl_366 AND and_dcpl_362 AND CONV_SL_1_1(fsm_output(5 DOWNTO
      4)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_426 <= and_dcpl_366 AND and_dcpl_370;
  and_dcpl_427 <= and_dcpl_415 AND and_dcpl_370;
  and_dcpl_428 <= and_dcpl_412 AND and_dcpl_370;
  and_dcpl_429 <= and_dcpl_420 AND and_dcpl_370;
  and_dcpl_430 <= and_dcpl_420 AND and_dcpl_380;
  and_dcpl_431 <= and_dcpl_415 AND and_dcpl_380;
  and_dcpl_447 <= NOT(CONV_SL_1_1(fsm_output/=STD_LOGIC_VECTOR'("000000010")));
  and_dcpl_465 <= nor_1630_cse AND (fsm_output(6)) AND nor_1624_cse;
  and_1025_cse <= and_dcpl_465 AND and_dcpl_376 AND and_dcpl_45;
  and_dcpl_467 <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  and_1028_cse <= and_dcpl_465 AND and_dcpl_467 AND and_dcpl_66;
  and_dcpl_475 <= and_1189_cse AND and_dcpl_75;
  and_dcpl_477 <= and_dcpl_88 AND and_570_cse;
  and_1037_cse <= and_dcpl_477 AND and_dcpl_475;
  and_dcpl_480 <= and_dcpl_376 AND and_dcpl_53;
  and_1040_cse <= and_dcpl_477 AND and_dcpl_480;
  and_dcpl_482 <= and_dcpl_467 AND and_dcpl_75;
  and_dcpl_484 <= and_dcpl_87 AND (fsm_output(6)) AND and_570_cse;
  and_1044_cse <= and_dcpl_484 AND and_dcpl_482;
  and_dcpl_486 <= and_dcpl_362 AND and_dcpl_53;
  and_1046_cse <= and_dcpl_484 AND and_dcpl_486;
  and_1051_cse <= and_dcpl_394 AND and_dcpl_475;
  and_1052_cse <= and_dcpl_394 AND and_dcpl_480;
  and_dcpl_495 <= and_dcpl_103 AND (fsm_output(6)) AND and_dcpl_387;
  and_1055_cse <= and_dcpl_495 AND and_dcpl_482;
  and_1056_cse <= and_dcpl_495 AND and_dcpl_486;
  and_1060_cse <= and_dcpl_404 AND and_dcpl_475;
  and_1061_cse <= and_dcpl_404 AND and_dcpl_480;
  and_1064_cse <= and_733_cse AND (fsm_output(6)) AND and_dcpl_397 AND and_dcpl_482;
  and_dcpl_571 <= and_dcpl_5 AND and_dcpl_397 AND and_dcpl_414;
  and_dcpl_577 <= and_dcpl_5 AND nor_1624_cse AND and_1189_cse AND and_dcpl_66;
  and_dcpl_589 <= and_dcpl_88 AND nor_1624_cse AND and_dcpl_414;
  COMP_LOOP_or_17_ssc <= and_dcpl_360 OR and_dcpl_367 OR and_dcpl_374 OR and_dcpl_378
      OR and_dcpl_384 OR and_dcpl_386 OR and_dcpl_390 OR and_dcpl_391 OR and_dcpl_395
      OR and_dcpl_396 OR and_dcpl_400 OR and_dcpl_401 OR and_dcpl_405 OR and_dcpl_406
      OR and_dcpl_409;
  or_tmp_2410 <= (fsm_output(3)) OR (fsm_output(0)) OR (fsm_output(2));
  COMP_LOOP_nor_itm <= NOT(and_dcpl_411 OR and_dcpl_413 OR and_dcpl_416 OR and_dcpl_417
      OR and_dcpl_418 OR and_dcpl_419 OR and_dcpl_421 OR and_dcpl_422 OR and_dcpl_425
      OR and_dcpl_426 OR and_dcpl_427 OR and_dcpl_428 OR and_dcpl_429 OR and_dcpl_430
      OR and_dcpl_431);
  COMP_LOOP_or_40_itm <= and_dcpl_416 OR and_dcpl_417 OR and_dcpl_418 OR and_dcpl_419
      OR and_dcpl_421 OR and_dcpl_422 OR and_dcpl_425;
  COMP_LOOP_nor_621_itm <= NOT(and_dcpl_413 OR and_dcpl_426 OR and_dcpl_427 OR and_dcpl_428
      OR and_dcpl_429 OR and_dcpl_430 OR and_dcpl_431);
  COMP_LOOP_or_41_itm <= and_dcpl_411 OR and_dcpl_426;
  COMP_LOOP_or_43_itm <= and_dcpl_427 OR and_dcpl_428 OR and_dcpl_429;
  COMP_LOOP_nor_622_itm <= NOT(and_dcpl_413 OR and_dcpl_430 OR and_dcpl_431);
  COMP_LOOP_or_47_itm <= and_dcpl_430 OR and_dcpl_431;
  COMP_LOOP_or_52_itm <= and_dcpl_411 OR and_dcpl_416 OR and_dcpl_417 OR and_dcpl_418
      OR and_dcpl_419 OR and_dcpl_421 OR and_dcpl_422 OR and_dcpl_425;
  COMP_LOOP_or_54_itm <= and_dcpl_426 OR and_dcpl_427 OR and_dcpl_428 OR and_dcpl_429;
  COMP_LOOP_or_18_itm <= (nor_1630_cse AND (NOT (fsm_output(6))) AND nor_1624_cse
      AND and_1189_cse AND and_dcpl_66) OR and_1025_cse OR and_1028_cse OR (and_dcpl_88
      AND nor_1624_cse AND and_dcpl_362 AND and_dcpl_45) OR and_1037_cse OR and_1040_cse
      OR and_1044_cse OR and_1046_cse OR and_1051_cse OR and_1052_cse OR and_1055_cse
      OR and_1056_cse OR and_1060_cse OR and_1061_cse OR and_1064_cse;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( ((and_dcpl_51 AND and_dcpl_47) OR STAGE_LOOP_i_3_0_sva_mx0c1) = '1' )
          THEN
        STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'( "1010"), z_out_4,
            STAGE_LOOP_i_3_0_sva_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(nor_1871_nl, and_1183_nl, fsm_output(5))) = '1' ) THEN
        p_sva <= p_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_vec_rsc_triosy_0_15_obj_ld_cse <= '0';
        reg_ensig_cgo_cse <= '0';
      ELSE
        reg_vec_rsc_triosy_0_15_obj_ld_cse <= and_dcpl_58 AND and_dcpl_46 AND CONV_SL_1_1(fsm_output(5
            DOWNTO 4)=STD_LOGIC_VECTOR'("11")) AND (NOT STAGE_LOOP_acc_itm_4_1);
        reg_ensig_cgo_cse <= mux_2255_rmff;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      tmp_33_sva_6 <= twiddle_rsc_0_6_i_q_d;
      tmp_33_sva_8 <= twiddle_rsc_0_8_i_q_d;
      tmp_33_sva_11 <= MUX_v_64_2_2(twiddle_rsc_0_11_i_q_d, twiddle_rsc_0_12_i_q_d,
          and_dcpl_180);
      tmp_33_sva_12 <= MUX_v_64_2_2(twiddle_rsc_0_12_i_q_d, twiddle_rsc_0_14_i_q_d,
          and_dcpl_180);
      tmp_33_sva_13 <= MUX_v_64_2_2(twiddle_rsc_0_13_i_q_d, tmp_33_sva_13_mx0w1,
          and_dcpl_192);
      tmp_33_sva_14 <= twiddle_rsc_0_14_i_q_d;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        VEC_LOOP_j_10_0_sva_9_0 <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (VEC_LOOP_j_10_0_sva_9_0_mx0c0 OR (and_dcpl_128 AND and_dcpl_118))
          = '1' ) THEN
        VEC_LOOP_j_10_0_sva_9_0 <= MUX_v_10_2_2(STD_LOGIC_VECTOR'("0000000000"),
            (z_out_2(9 DOWNTO 0)), VEC_LOOP_j_not_1_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(nor_1870_nl, and_nl, fsm_output(5))) = '1' ) THEN
        STAGE_LOOP_lshift_psp_sva <= z_out;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_2558_nl, mux_nl, fsm_output(4))) = '1' ) THEN
        COMP_LOOP_k_10_4_sva_5_0 <= MUX_v_6_2_2(STD_LOGIC_VECTOR'("000000"), reg_COMP_LOOP_k_10_4_ftd,
            nand_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_1_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_acc_10_cse_10_1_1_sva <= COMP_LOOP_1_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_acc_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0(9
            DOWNTO 4)) + UNSIGNED(COMP_LOOP_k_10_4_sva_5_0), 6));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm <= z_out_2(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_2_tmp_lshift_ncse_sva <= z_out_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_9_tmp_lshift_itm <= STD_LOGIC_VECTOR'( "0000000");
      ELSIF ( (and_dcpl_62 OR and_dcpl_207) = '1' ) THEN
        COMP_LOOP_9_tmp_lshift_itm <= MUX_v_7_2_2((z_out(6 DOWNTO 0)), (z_out_3(6
            DOWNTO 0)), and_dcpl_207);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_1_tmp_acc_cse_sva <= z_out_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_244_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_62_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_185_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_64_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_65_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_66_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_6_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_68_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_69_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_70_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_10_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_72_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_12_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_13_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_14_itm <= '0';
      ELSIF ( mux_2303_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_itm <= NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_COMP_LOOP_and_244_itm <= (COMP_LOOP_acc_13_psp_sva_1(0)) AND (VEC_LOOP_j_10_0_sva_9_0(0))
            AND (NOT((COMP_LOOP_acc_13_psp_sva_1(1)) OR (VEC_LOOP_j_10_0_sva_9_0(1))));
        COMP_LOOP_COMP_LOOP_and_62_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_COMP_LOOP_and_185_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_64_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_65_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_66_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_COMP_LOOP_and_6_itm <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_COMP_LOOP_and_68_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_69_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_70_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_10_itm <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_72_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_12_itm <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_13_itm <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_14_itm <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_13_psp_sva <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( (mux_2309_nl OR (fsm_output(8))) = '1' ) THEN
        COMP_LOOP_acc_13_psp_sva <= COMP_LOOP_acc_13_psp_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_4_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (NOT((NOT mux_2312_nl) AND nor_1630_cse)) = '1' ) THEN
        COMP_LOOP_acc_1_cse_4_sva <= COMP_LOOP_acc_1_cse_4_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_2_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (NOT(mux_2314_nl AND and_dcpl_5)) = '1' ) THEN
        COMP_LOOP_acc_1_cse_2_sva <= COMP_LOOP_acc_1_cse_2_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_2_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (NOT(mux_2315_nl AND and_dcpl_5)) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_2_sva <= COMP_LOOP_2_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (NOT((and_1189_cse OR (fsm_output(2)) OR or_dcpl_190) AND and_dcpl_5))
          = '1' ) THEN
        COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_3_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_5_itm <= '0';
      ELSIF ( and_dcpl_248 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_5_itm <= NOT(CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_51_itm <= '0';
      ELSIF ( and_dcpl_248 = '0' ) THEN
        COMP_LOOP_nor_51_itm <= NOT(CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(3 DOWNTO
            1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_52_itm <= '0';
      ELSIF ( and_dcpl_248 = '0' ) THEN
        COMP_LOOP_nor_52_itm <= NOT((COMP_LOOP_2_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_77_itm <= '0';
      ELSIF ( and_dcpl_248 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_77_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_54_itm <= '0';
      ELSIF ( and_dcpl_248 = '0' ) THEN
        COMP_LOOP_nor_54_itm <= NOT((COMP_LOOP_2_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_79_itm <= '0';
      ELSIF ( and_dcpl_248 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_79_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_80_itm <= '0';
      ELSIF ( and_dcpl_248 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_80_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_81_itm <= '0';
      ELSIF ( and_dcpl_248 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_81_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_57_itm <= '0';
      ELSIF ( and_dcpl_248 = '0' ) THEN
        COMP_LOOP_nor_57_itm <= NOT(CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(2 DOWNTO
            0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_83_itm <= '0';
      ELSIF ( and_dcpl_248 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_83_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_84_itm <= '0';
      ELSIF ( and_dcpl_248 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_84_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_85_itm <= '0';
      ELSIF ( and_dcpl_248 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_85_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_86_itm <= '0';
      ELSIF ( and_dcpl_248 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_86_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_87_itm <= '0';
      ELSIF ( and_dcpl_248 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_87_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_88_itm <= '0';
      ELSIF ( and_dcpl_248 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_88_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_89_itm <= '0';
      ELSIF ( and_dcpl_248 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_89_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_itm <= '0';
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_nor_itm <= '0';
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_tmp_nor_itm <= COMP_LOOP_tmp_nor_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_nor_1_itm <= '0';
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_tmp_nor_1_itm <= COMP_LOOP_tmp_nor_1_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_itm <= '0';
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_nor_3_itm <= '0';
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_tmp_nor_3_itm <= COMP_LOOP_tmp_nor_3_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_itm <= '0';
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_itm <= '0';
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_itm <= '0';
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_nor_6_itm <= '0';
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_tmp_nor_6_itm <= COMP_LOOP_tmp_nor_6_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_itm <= '0';
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_itm <= '0';
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_itm <= '0';
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_itm <= '0';
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_itm <= '0';
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_itm <= '0';
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_itm <= '0';
      ELSIF ( or_dcpl_184 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_11_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( (NOT((NOT mux_2317_nl) AND nor_1630_cse)) = '1' ) THEN
        COMP_LOOP_acc_11_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0(9
            DOWNTO 1)) + UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 & STD_LOGIC_VECTOR'( "001")),
            9));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_3_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (NOT((NOT mux_2319_nl) AND nor_1630_cse)) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_3_sva <= COMP_LOOP_3_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (NOT(mux_2321_nl AND nor_1630_cse)) = '1' ) THEN
        COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm <= COMP_LOOP_acc_12_nl(8);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_9_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_9_itm <= NOT(CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_91_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_nor_91_itm <= NOT(CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(3 DOWNTO
            1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_92_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_nor_92_itm <= NOT((COMP_LOOP_3_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_3_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_137_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_137_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_94_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_nor_94_itm <= NOT((COMP_LOOP_3_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_3_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_139_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_139_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_140_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_140_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_141_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_141_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_97_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_nor_97_itm <= NOT(CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(2 DOWNTO
            0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_143_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_143_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_144_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_144_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_145_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_145_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_146_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_146_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_147_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_147_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_148_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_148_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_149_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_149_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_4_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (NOT((NOT mux_2326_nl) AND nor_1630_cse)) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_4_sva <= COMP_LOOP_4_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (NOT((NOT mux_2327_nl) AND nor_1630_cse)) = '1' ) THEN
        COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_5_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_13_itm <= '0';
      ELSIF ( and_dcpl_255 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_13_itm <= NOT(CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_131_itm <= '0';
      ELSIF ( and_dcpl_255 = '0' ) THEN
        COMP_LOOP_nor_131_itm <= NOT(CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_132_itm <= '0';
      ELSIF ( and_dcpl_255 = '0' ) THEN
        COMP_LOOP_nor_132_itm <= NOT((COMP_LOOP_4_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_4_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_197_itm <= '0';
      ELSIF ( and_dcpl_255 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_197_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_134_itm <= '0';
      ELSIF ( and_dcpl_255 = '0' ) THEN
        COMP_LOOP_nor_134_itm <= NOT((COMP_LOOP_4_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_4_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_199_itm <= '0';
      ELSIF ( and_dcpl_255 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_199_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_200_itm <= '0';
      ELSIF ( and_dcpl_255 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_200_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_201_itm <= '0';
      ELSIF ( and_dcpl_255 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_201_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_137_itm <= '0';
      ELSIF ( and_dcpl_255 = '0' ) THEN
        COMP_LOOP_nor_137_itm <= NOT(CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_203_itm <= '0';
      ELSIF ( and_dcpl_255 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_203_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_204_itm <= '0';
      ELSIF ( and_dcpl_255 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_204_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_205_itm <= '0';
      ELSIF ( and_dcpl_255 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_205_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_206_itm <= '0';
      ELSIF ( and_dcpl_255 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_206_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_207_itm <= '0';
      ELSIF ( and_dcpl_255 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_207_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_208_itm <= '0';
      ELSIF ( and_dcpl_255 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_208_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_209_itm <= '0';
      ELSIF ( and_dcpl_255 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_209_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_5_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_2332_nl OR (fsm_output(8))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_5_sva <= COMP_LOOP_5_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_2335_nl OR (fsm_output(8))) = '1' ) THEN
        COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_6_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_17_itm <= '0';
      ELSIF ( and_dcpl_258 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_17_itm <= NOT(CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_171_itm <= '0';
      ELSIF ( and_dcpl_258 = '0' ) THEN
        COMP_LOOP_nor_171_itm <= NOT(CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_172_itm <= '0';
      ELSIF ( and_dcpl_258 = '0' ) THEN
        COMP_LOOP_nor_172_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_257_itm <= '0';
      ELSIF ( and_dcpl_258 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_257_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_174_itm <= '0';
      ELSIF ( and_dcpl_258 = '0' ) THEN
        COMP_LOOP_nor_174_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_259_itm <= '0';
      ELSIF ( and_dcpl_258 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_259_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_260_itm <= '0';
      ELSIF ( and_dcpl_258 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_260_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_261_itm <= '0';
      ELSIF ( and_dcpl_258 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_261_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_177_itm <= '0';
      ELSIF ( and_dcpl_258 = '0' ) THEN
        COMP_LOOP_nor_177_itm <= NOT(CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_263_itm <= '0';
      ELSIF ( and_dcpl_258 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_263_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_264_itm <= '0';
      ELSIF ( and_dcpl_258 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_264_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_265_itm <= '0';
      ELSIF ( and_dcpl_258 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_265_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_266_itm <= '0';
      ELSIF ( and_dcpl_258 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_266_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_267_itm <= '0';
      ELSIF ( and_dcpl_258 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_267_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_268_itm <= '0';
      ELSIF ( and_dcpl_258 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_268_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_269_itm <= '0';
      ELSIF ( and_dcpl_258 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_269_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_6_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_2338_nl OR (fsm_output(8))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_6_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0)
            + UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 & STD_LOGIC_VECTOR'( "0101")), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_6_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_2340_nl OR (fsm_output(8))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_6_sva <= COMP_LOOP_6_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_2341_nl OR (fsm_output(8))) = '1' ) THEN
        COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_7_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_21_itm <= '0';
      ELSIF ( and_dcpl_262 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_21_itm <= NOT(CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_211_itm <= '0';
      ELSIF ( and_dcpl_262 = '0' ) THEN
        COMP_LOOP_nor_211_itm <= NOT(CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_212_itm <= '0';
      ELSIF ( and_dcpl_262 = '0' ) THEN
        COMP_LOOP_nor_212_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_317_itm <= '0';
      ELSIF ( and_dcpl_262 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_317_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_214_itm <= '0';
      ELSIF ( and_dcpl_262 = '0' ) THEN
        COMP_LOOP_nor_214_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_319_itm <= '0';
      ELSIF ( and_dcpl_262 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_319_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_320_itm <= '0';
      ELSIF ( and_dcpl_262 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_320_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_321_itm <= '0';
      ELSIF ( and_dcpl_262 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_321_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_217_itm <= '0';
      ELSIF ( and_dcpl_262 = '0' ) THEN
        COMP_LOOP_nor_217_itm <= NOT(CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_323_itm <= '0';
      ELSIF ( and_dcpl_262 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_323_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_324_itm <= '0';
      ELSIF ( and_dcpl_262 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_324_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_325_itm <= '0';
      ELSIF ( and_dcpl_262 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_325_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_326_itm <= '0';
      ELSIF ( and_dcpl_262 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_326_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_327_itm <= '0';
      ELSIF ( and_dcpl_262 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_327_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_328_itm <= '0';
      ELSIF ( and_dcpl_262 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_328_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_329_itm <= '0';
      ELSIF ( and_dcpl_262 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_329_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_14_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( (mux_2346_nl OR (fsm_output(8))) = '1' ) THEN
        COMP_LOOP_acc_14_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0(9
            DOWNTO 1)) + UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 & STD_LOGIC_VECTOR'( "011")),
            9));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_7_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_2349_nl OR (fsm_output(8))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_7_sva <= COMP_LOOP_7_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_2352_nl OR (fsm_output(8))) = '1' ) THEN
        COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm <= COMP_LOOP_acc_15_nl(7);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_25_itm <= '0';
      ELSIF ( and_dcpl_266 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_25_itm <= NOT(CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_251_itm <= '0';
      ELSIF ( and_dcpl_266 = '0' ) THEN
        COMP_LOOP_nor_251_itm <= NOT(CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_252_itm <= '0';
      ELSIF ( and_dcpl_266 = '0' ) THEN
        COMP_LOOP_nor_252_itm <= NOT((COMP_LOOP_7_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_377_itm <= '0';
      ELSIF ( and_dcpl_266 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_377_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_254_itm <= '0';
      ELSIF ( and_dcpl_266 = '0' ) THEN
        COMP_LOOP_nor_254_itm <= NOT((COMP_LOOP_7_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_379_itm <= '0';
      ELSIF ( and_dcpl_266 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_379_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_380_itm <= '0';
      ELSIF ( and_dcpl_266 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_380_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_381_itm <= '0';
      ELSIF ( and_dcpl_266 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_381_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_257_itm <= '0';
      ELSIF ( and_dcpl_266 = '0' ) THEN
        COMP_LOOP_nor_257_itm <= NOT(CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_383_itm <= '0';
      ELSIF ( and_dcpl_266 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_383_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_384_itm <= '0';
      ELSIF ( and_dcpl_266 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_384_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_385_itm <= '0';
      ELSIF ( and_dcpl_266 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_385_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_386_itm <= '0';
      ELSIF ( and_dcpl_266 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_386_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_387_itm <= '0';
      ELSIF ( and_dcpl_266 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_387_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_388_itm <= '0';
      ELSIF ( and_dcpl_266 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_388_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_389_itm <= '0';
      ELSIF ( and_dcpl_266 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_389_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_8_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_2354_nl OR (fsm_output(8))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_8_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0)
            + UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 & STD_LOGIC_VECTOR'( "0111")), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_8_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_2355_nl OR (fsm_output(8))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_8_sva <= COMP_LOOP_8_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_2356_nl OR (fsm_output(8))) = '1' ) THEN
        COMP_LOOP_9_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_9_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_29_itm <= '0';
      ELSIF ( and_dcpl_270 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_29_itm <= NOT(CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_291_itm <= '0';
      ELSIF ( and_dcpl_270 = '0' ) THEN
        COMP_LOOP_nor_291_itm <= NOT(CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_292_itm <= '0';
      ELSIF ( and_dcpl_270 = '0' ) THEN
        COMP_LOOP_nor_292_itm <= NOT((COMP_LOOP_8_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_437_itm <= '0';
      ELSIF ( and_dcpl_270 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_437_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_294_itm <= '0';
      ELSIF ( and_dcpl_270 = '0' ) THEN
        COMP_LOOP_nor_294_itm <= NOT((COMP_LOOP_8_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_439_itm <= '0';
      ELSIF ( and_dcpl_270 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_439_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_440_itm <= '0';
      ELSIF ( and_dcpl_270 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_440_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_441_itm <= '0';
      ELSIF ( and_dcpl_270 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_441_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_297_itm <= '0';
      ELSIF ( and_dcpl_270 = '0' ) THEN
        COMP_LOOP_nor_297_itm <= NOT(CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_443_itm <= '0';
      ELSIF ( and_dcpl_270 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_443_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_444_itm <= '0';
      ELSIF ( and_dcpl_270 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_444_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_445_itm <= '0';
      ELSIF ( and_dcpl_270 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_445_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_446_itm <= '0';
      ELSIF ( and_dcpl_270 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_446_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_447_itm <= '0';
      ELSIF ( and_dcpl_270 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_447_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_448_itm <= '0';
      ELSIF ( and_dcpl_270 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_448_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_449_itm <= '0';
      ELSIF ( and_dcpl_270 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_449_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_16_psp_sva <= STD_LOGIC_VECTOR'( "0000000");
      ELSIF ( (MUX_s_1_2_2(mux_2364_nl, (fsm_output(8)), fsm_output(5))) = '1' )
          THEN
        COMP_LOOP_acc_16_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0(9
            DOWNTO 3)) + UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 & '1'), 7));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_9_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_2368_nl, (fsm_output(8)), fsm_output(5))) = '1' )
          THEN
        COMP_LOOP_acc_10_cse_10_1_9_sva <= COMP_LOOP_9_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_2372_nl, (fsm_output(8)), fsm_output(5))) = '1' ) THEN
        COMP_LOOP_10_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_10_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_33_itm <= '0';
      ELSIF ( and_dcpl_271 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_33_itm <= NOT(CONV_SL_1_1(COMP_LOOP_9_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_331_itm <= '0';
      ELSIF ( and_dcpl_271 = '0' ) THEN
        COMP_LOOP_nor_331_itm <= NOT(CONV_SL_1_1(COMP_LOOP_9_acc_10_itm_10_1_1(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_332_itm <= '0';
      ELSIF ( and_dcpl_271 = '0' ) THEN
        COMP_LOOP_nor_332_itm <= NOT((COMP_LOOP_9_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_9_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_9_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_497_itm <= '0';
      ELSIF ( and_dcpl_271 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_497_itm <= CONV_SL_1_1(COMP_LOOP_9_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_334_itm <= '0';
      ELSIF ( and_dcpl_271 = '0' ) THEN
        COMP_LOOP_nor_334_itm <= NOT((COMP_LOOP_9_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_9_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_9_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_499_itm <= '0';
      ELSIF ( and_dcpl_271 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_499_itm <= CONV_SL_1_1(COMP_LOOP_9_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_500_itm <= '0';
      ELSIF ( and_dcpl_271 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_500_itm <= CONV_SL_1_1(COMP_LOOP_9_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_501_itm <= '0';
      ELSIF ( and_dcpl_271 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_501_itm <= CONV_SL_1_1(COMP_LOOP_9_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_337_itm <= '0';
      ELSIF ( and_dcpl_271 = '0' ) THEN
        COMP_LOOP_nor_337_itm <= NOT(CONV_SL_1_1(COMP_LOOP_9_acc_10_itm_10_1_1(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_503_itm <= '0';
      ELSIF ( and_dcpl_271 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_503_itm <= CONV_SL_1_1(COMP_LOOP_9_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_504_itm <= '0';
      ELSIF ( and_dcpl_271 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_504_itm <= CONV_SL_1_1(COMP_LOOP_9_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_505_itm <= '0';
      ELSIF ( and_dcpl_271 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_505_itm <= CONV_SL_1_1(COMP_LOOP_9_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_506_itm <= '0';
      ELSIF ( and_dcpl_271 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_506_itm <= CONV_SL_1_1(COMP_LOOP_9_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_507_itm <= '0';
      ELSIF ( and_dcpl_271 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_507_itm <= CONV_SL_1_1(COMP_LOOP_9_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_508_itm <= '0';
      ELSIF ( and_dcpl_271 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_508_itm <= CONV_SL_1_1(COMP_LOOP_9_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_509_itm <= '0';
      ELSIF ( and_dcpl_271 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_509_itm <= CONV_SL_1_1(COMP_LOOP_9_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_10_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_tmp_2357, mux_2375_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_10_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0)
            + UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 & STD_LOGIC_VECTOR'( "1001")), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_10_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_tmp_2357, mux_2378_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_10_sva <= COMP_LOOP_10_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_tmp_2357, and_390_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_11_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_11_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_37_itm <= '0';
        COMP_LOOP_nor_371_itm <= '0';
        COMP_LOOP_nor_372_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_557_itm <= '0';
        COMP_LOOP_nor_374_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_559_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_560_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_561_itm <= '0';
        COMP_LOOP_nor_377_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_563_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_564_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_565_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_566_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_567_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_568_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_569_itm <= '0';
      ELSIF ( mux_2383_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_37_itm <= NOT(CONV_SL_1_1(COMP_LOOP_10_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_371_itm <= NOT(CONV_SL_1_1(COMP_LOOP_10_acc_10_itm_10_1_1(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_nor_372_itm <= NOT((COMP_LOOP_10_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_10_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_10_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_557_itm <= CONV_SL_1_1(COMP_LOOP_10_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_nor_374_itm <= NOT((COMP_LOOP_10_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_10_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_10_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_559_itm <= CONV_SL_1_1(COMP_LOOP_10_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_560_itm <= CONV_SL_1_1(COMP_LOOP_10_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_561_itm <= CONV_SL_1_1(COMP_LOOP_10_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_nor_377_itm <= NOT(CONV_SL_1_1(COMP_LOOP_10_acc_10_itm_10_1_1(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_563_itm <= CONV_SL_1_1(COMP_LOOP_10_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_564_itm <= CONV_SL_1_1(COMP_LOOP_10_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_565_itm <= CONV_SL_1_1(COMP_LOOP_10_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_566_itm <= CONV_SL_1_1(COMP_LOOP_10_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_567_itm <= CONV_SL_1_1(COMP_LOOP_10_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_568_itm <= CONV_SL_1_1(COMP_LOOP_10_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_569_itm <= CONV_SL_1_1(COMP_LOOP_10_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_17_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( (MUX_s_1_2_2(mux_2389_nl, nor_tmp_115, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_17_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0(9
            DOWNTO 1)) + UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 & STD_LOGIC_VECTOR'( "101")),
            9));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_11_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_2392_nl, nor_tmp_115, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_11_sva <= COMP_LOOP_11_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_2395_nl, nor_tmp_115, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_slc_COMP_LOOP_acc_18_8_itm <= COMP_LOOP_acc_18_nl(8);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_41_itm <= '0';
        COMP_LOOP_nor_411_itm <= '0';
        COMP_LOOP_nor_412_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_617_itm <= '0';
        COMP_LOOP_nor_414_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_619_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_620_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_621_itm <= '0';
        COMP_LOOP_nor_417_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_623_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_624_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_625_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_626_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_627_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_628_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_629_itm <= '0';
      ELSIF ( mux_2398_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_41_itm <= NOT(CONV_SL_1_1(COMP_LOOP_11_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_411_itm <= NOT(CONV_SL_1_1(COMP_LOOP_11_acc_10_itm_10_1_1(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_nor_412_itm <= NOT((COMP_LOOP_11_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_11_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_11_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_617_itm <= CONV_SL_1_1(COMP_LOOP_11_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_nor_414_itm <= NOT((COMP_LOOP_11_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_11_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_11_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_619_itm <= CONV_SL_1_1(COMP_LOOP_11_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_620_itm <= CONV_SL_1_1(COMP_LOOP_11_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_621_itm <= CONV_SL_1_1(COMP_LOOP_11_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_nor_417_itm <= NOT(CONV_SL_1_1(COMP_LOOP_11_acc_10_itm_10_1_1(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_623_itm <= CONV_SL_1_1(COMP_LOOP_11_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_624_itm <= CONV_SL_1_1(COMP_LOOP_11_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_625_itm <= CONV_SL_1_1(COMP_LOOP_11_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_626_itm <= CONV_SL_1_1(COMP_LOOP_11_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_627_itm <= CONV_SL_1_1(COMP_LOOP_11_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_628_itm <= CONV_SL_1_1(COMP_LOOP_11_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_629_itm <= CONV_SL_1_1(COMP_LOOP_11_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_12_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_2400_nl, (fsm_output(8)), fsm_output(7))) = '1' )
          THEN
        COMP_LOOP_acc_1_cse_12_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0)
            + UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 & STD_LOGIC_VECTOR'( "1011")), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_12_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_tmp_2384, mux_2402_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_12_sva <= COMP_LOOP_12_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_tmp_2384, mux_2405_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_13_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_13_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_45_itm <= '0';
        COMP_LOOP_nor_451_itm <= '0';
        COMP_LOOP_nor_452_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_677_itm <= '0';
        COMP_LOOP_nor_454_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_679_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_680_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_681_itm <= '0';
        COMP_LOOP_nor_457_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_683_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_684_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_685_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_686_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_687_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_688_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_689_itm <= '0';
      ELSIF ( mux_2410_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_45_itm <= NOT(CONV_SL_1_1(COMP_LOOP_12_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_451_itm <= NOT(CONV_SL_1_1(COMP_LOOP_12_acc_10_itm_10_1_1(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_nor_452_itm <= NOT((COMP_LOOP_12_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_12_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_12_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_677_itm <= CONV_SL_1_1(COMP_LOOP_12_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_nor_454_itm <= NOT((COMP_LOOP_12_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_12_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_12_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_679_itm <= CONV_SL_1_1(COMP_LOOP_12_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_680_itm <= CONV_SL_1_1(COMP_LOOP_12_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_681_itm <= CONV_SL_1_1(COMP_LOOP_12_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_nor_457_itm <= NOT(CONV_SL_1_1(COMP_LOOP_12_acc_10_itm_10_1_1(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_683_itm <= CONV_SL_1_1(COMP_LOOP_12_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_684_itm <= CONV_SL_1_1(COMP_LOOP_12_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_685_itm <= CONV_SL_1_1(COMP_LOOP_12_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_686_itm <= CONV_SL_1_1(COMP_LOOP_12_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_687_itm <= CONV_SL_1_1(COMP_LOOP_12_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_688_itm <= CONV_SL_1_1(COMP_LOOP_12_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_689_itm <= CONV_SL_1_1(COMP_LOOP_12_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_19_psp_sva <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( (MUX_s_1_2_2(mux_2415_nl, and_733_cse, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_19_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0(9
            DOWNTO 2)) + UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 & STD_LOGIC_VECTOR'( "11")),
            8));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_13_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_2418_nl, and_733_cse, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_13_sva <= COMP_LOOP_13_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_2422_nl, and_733_cse, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_14_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_14_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_49_itm <= '0';
        COMP_LOOP_nor_491_itm <= '0';
        COMP_LOOP_nor_492_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_737_itm <= '0';
        COMP_LOOP_nor_494_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_739_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_740_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_741_itm <= '0';
        COMP_LOOP_nor_497_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_743_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_744_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_745_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_746_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_747_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_748_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_749_itm <= '0';
      ELSIF ( mux_2424_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_49_itm <= NOT(CONV_SL_1_1(COMP_LOOP_13_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_491_itm <= NOT(CONV_SL_1_1(COMP_LOOP_13_acc_10_itm_10_1_1(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_nor_492_itm <= NOT((COMP_LOOP_13_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_13_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_13_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_737_itm <= CONV_SL_1_1(COMP_LOOP_13_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_nor_494_itm <= NOT((COMP_LOOP_13_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_13_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_13_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_739_itm <= CONV_SL_1_1(COMP_LOOP_13_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_740_itm <= CONV_SL_1_1(COMP_LOOP_13_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_741_itm <= CONV_SL_1_1(COMP_LOOP_13_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_nor_497_itm <= NOT(CONV_SL_1_1(COMP_LOOP_13_acc_10_itm_10_1_1(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_743_itm <= CONV_SL_1_1(COMP_LOOP_13_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_744_itm <= CONV_SL_1_1(COMP_LOOP_13_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_745_itm <= CONV_SL_1_1(COMP_LOOP_13_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_746_itm <= CONV_SL_1_1(COMP_LOOP_13_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_747_itm <= CONV_SL_1_1(COMP_LOOP_13_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_748_itm <= CONV_SL_1_1(COMP_LOOP_13_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_749_itm <= CONV_SL_1_1(COMP_LOOP_13_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_14_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_2426_nl, and_733_cse, fsm_output(6))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_14_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0)
            + UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 & STD_LOGIC_VECTOR'( "1101")), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_14_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_tmp_2410, mux_2428_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_14_sva <= COMP_LOOP_14_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_tmp_2410, mux_2431_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_15_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_15_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_53_itm <= '0';
        COMP_LOOP_nor_531_itm <= '0';
        COMP_LOOP_nor_532_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_797_itm <= '0';
        COMP_LOOP_nor_534_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_799_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_800_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_801_itm <= '0';
        COMP_LOOP_nor_537_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_803_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_804_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_805_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_806_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_807_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_808_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_809_itm <= '0';
      ELSIF ( mux_2435_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_53_itm <= NOT(CONV_SL_1_1(COMP_LOOP_14_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_531_itm <= NOT(CONV_SL_1_1(COMP_LOOP_14_acc_10_itm_10_1_1(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_nor_532_itm <= NOT((COMP_LOOP_14_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_14_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_14_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_797_itm <= CONV_SL_1_1(COMP_LOOP_14_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_nor_534_itm <= NOT((COMP_LOOP_14_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_14_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_14_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_799_itm <= CONV_SL_1_1(COMP_LOOP_14_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_800_itm <= CONV_SL_1_1(COMP_LOOP_14_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_801_itm <= CONV_SL_1_1(COMP_LOOP_14_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_nor_537_itm <= NOT(CONV_SL_1_1(COMP_LOOP_14_acc_10_itm_10_1_1(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_803_itm <= CONV_SL_1_1(COMP_LOOP_14_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_804_itm <= CONV_SL_1_1(COMP_LOOP_14_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_805_itm <= CONV_SL_1_1(COMP_LOOP_14_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_806_itm <= CONV_SL_1_1(COMP_LOOP_14_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_807_itm <= CONV_SL_1_1(COMP_LOOP_14_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_808_itm <= CONV_SL_1_1(COMP_LOOP_14_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_809_itm <= CONV_SL_1_1(COMP_LOOP_14_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_20_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( (MUX_s_1_2_2(mux_2436_nl, and_dcpl_57, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_20_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0(9
            DOWNTO 1)) + UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 & STD_LOGIC_VECTOR'( "111")),
            9));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_15_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_2438_nl, and_dcpl_57, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_15_sva <= COMP_LOOP_15_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mux_2442_itm = '1' ) THEN
        COMP_LOOP_slc_COMP_LOOP_acc_21_6_itm <= COMP_LOOP_acc_21_nl(6);
        reg_COMP_LOOP_k_10_4_ftd <= COMP_LOOP_k_10_4_sva_2(5 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_57_itm <= '0';
        COMP_LOOP_nor_571_itm <= '0';
        COMP_LOOP_nor_572_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_857_itm <= '0';
        COMP_LOOP_nor_574_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_859_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_860_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_861_itm <= '0';
        COMP_LOOP_nor_577_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_863_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_864_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_865_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_866_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_867_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_868_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_869_itm <= '0';
      ELSIF ( mux_2444_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_57_itm <= NOT(CONV_SL_1_1(COMP_LOOP_15_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_571_itm <= NOT(CONV_SL_1_1(COMP_LOOP_15_acc_10_itm_10_1_1(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_nor_572_itm <= NOT((COMP_LOOP_15_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_15_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_15_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_857_itm <= CONV_SL_1_1(COMP_LOOP_15_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_nor_574_itm <= NOT((COMP_LOOP_15_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_15_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_15_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_859_itm <= CONV_SL_1_1(COMP_LOOP_15_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_860_itm <= CONV_SL_1_1(COMP_LOOP_15_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_861_itm <= CONV_SL_1_1(COMP_LOOP_15_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_nor_577_itm <= NOT(CONV_SL_1_1(COMP_LOOP_15_acc_10_itm_10_1_1(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_863_itm <= CONV_SL_1_1(COMP_LOOP_15_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_864_itm <= CONV_SL_1_1(COMP_LOOP_15_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_865_itm <= CONV_SL_1_1(COMP_LOOP_15_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_866_itm <= CONV_SL_1_1(COMP_LOOP_15_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_867_itm <= CONV_SL_1_1(COMP_LOOP_15_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_868_itm <= CONV_SL_1_1(COMP_LOOP_15_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_869_itm <= CONV_SL_1_1(COMP_LOOP_15_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(not_tmp_762, and_303_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0)
            + UNSIGNED(COMP_LOOP_k_10_4_sva_5_0 & STD_LOGIC_VECTOR'( "1111")), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(not_tmp_762, and_363_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_sva <= COMP_LOOP_16_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(not_tmp_762, and_304_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_1_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_61_itm <= '0';
        COMP_LOOP_nor_611_itm <= '0';
        COMP_LOOP_nor_612_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_917_itm <= '0';
        COMP_LOOP_nor_614_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_919_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_920_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_921_itm <= '0';
        COMP_LOOP_nor_617_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_923_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_924_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_925_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_926_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_927_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_928_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_929_itm <= '0';
      ELSIF ( mux_2449_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_61_itm <= NOT(CONV_SL_1_1(COMP_LOOP_16_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_611_itm <= NOT(CONV_SL_1_1(COMP_LOOP_16_acc_10_itm_10_1_1(3
            DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_nor_612_itm <= NOT((COMP_LOOP_16_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_16_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_16_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_917_itm <= CONV_SL_1_1(COMP_LOOP_16_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_nor_614_itm <= NOT((COMP_LOOP_16_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_16_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_16_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_919_itm <= CONV_SL_1_1(COMP_LOOP_16_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_920_itm <= CONV_SL_1_1(COMP_LOOP_16_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_921_itm <= CONV_SL_1_1(COMP_LOOP_16_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_nor_617_itm <= NOT(CONV_SL_1_1(COMP_LOOP_16_acc_10_itm_10_1_1(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_923_itm <= CONV_SL_1_1(COMP_LOOP_16_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_924_itm <= CONV_SL_1_1(COMP_LOOP_16_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_925_itm <= CONV_SL_1_1(COMP_LOOP_16_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_926_itm <= CONV_SL_1_1(COMP_LOOP_16_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_927_itm <= CONV_SL_1_1(COMP_LOOP_16_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_928_itm <= CONV_SL_1_1(COMP_LOOP_16_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_929_itm <= CONV_SL_1_1(COMP_LOOP_16_acc_10_itm_10_1_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_10_tmp_mul_idiv_sva <= STD_LOGIC_VECTOR'( "0000000000");
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm <= '0';
        COMP_LOOP_tmp_nor_13_itm <= '0';
        COMP_LOOP_tmp_nor_14_itm <= '0';
        COMP_LOOP_tmp_nor_16_itm <= '0';
        COMP_LOOP_tmp_nor_19_itm <= '0';
      ELSIF ( COMP_LOOP_tmp_or_1_cse = '1' ) THEN
        COMP_LOOP_10_tmp_mul_idiv_sva <= z_out_3(9 DOWNTO 0);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_23_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_cse,
            STD_LOGIC_VECTOR'( and_dcpl_62 & and_dcpl_189 & COMP_LOOP_or_27_cse));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_24_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_cse,
            STD_LOGIC_VECTOR'( and_dcpl_62 & and_dcpl_189 & COMP_LOOP_or_27_cse));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_25_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_cse,
            STD_LOGIC_VECTOR'( and_dcpl_62 & and_dcpl_189 & COMP_LOOP_or_27_cse));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_26_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse,
            STD_LOGIC_VECTOR'( and_dcpl_62 & and_dcpl_189 & COMP_LOOP_or_27_cse));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_27_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse,
            STD_LOGIC_VECTOR'( and_dcpl_62 & and_dcpl_189 & COMP_LOOP_or_27_cse));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_28_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse,
            STD_LOGIC_VECTOR'( and_dcpl_62 & and_dcpl_189 & COMP_LOOP_or_27_cse));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_29_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse,
            STD_LOGIC_VECTOR'( and_dcpl_62 & and_dcpl_189 & COMP_LOOP_or_27_cse));
        COMP_LOOP_tmp_nor_13_itm <= MUX_s_1_2_2(COMP_LOOP_nor_11_nl, COMP_LOOP_tmp_nor_cse,
            COMP_LOOP_or_23_cse);
        COMP_LOOP_tmp_nor_14_itm <= MUX_s_1_2_2(COMP_LOOP_nor_12_nl, COMP_LOOP_tmp_nor_1_cse,
            COMP_LOOP_or_23_cse);
        COMP_LOOP_tmp_nor_16_itm <= MUX_s_1_2_2(COMP_LOOP_nor_14_nl, COMP_LOOP_tmp_nor_3_cse,
            COMP_LOOP_or_23_cse);
        COMP_LOOP_tmp_nor_19_itm <= MUX_s_1_2_2(COMP_LOOP_nor_17_nl, COMP_LOOP_tmp_nor_6_cse,
            COMP_LOOP_or_23_cse);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm <= '0';
      ELSIF ( COMP_LOOP_tmp_or_2_cse = '1' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_17_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_17_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_cse,
            STD_LOGIC_VECTOR'( and_dcpl_62 & and_dcpl_65 & COMP_LOOP_or_27_cse));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_19_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_19_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_cse,
            STD_LOGIC_VECTOR'( and_dcpl_62 & and_dcpl_65 & COMP_LOOP_or_27_cse));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_20_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_20_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_cse,
            STD_LOGIC_VECTOR'( and_dcpl_62 & and_dcpl_65 & COMP_LOOP_or_27_cse));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_21_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_21_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_cse,
            STD_LOGIC_VECTOR'( and_dcpl_62 & and_dcpl_65 & COMP_LOOP_or_27_cse));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm <= '0';
      ELSIF ( (and_dcpl_62 OR and_dcpl_189 OR and_dcpl_195 OR and_dcpl_197 OR and_dcpl_198)
          = '1' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_nor_1_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_17_cse,
            STD_LOGIC_VECTOR'( and_dcpl_62 & and_dcpl_189 & COMP_LOOP_or_31_cse));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (NOT(or_dcpl_183 OR or_dcpl_207)) = '1' ) THEN
        COMP_LOOP_3_tmp_lshift_ncse_sva <= z_out_1(8 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_2565_nl AND CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("00"))
          AND nor_1630_cse) = '1' ) THEN
        tmp_33_sva_1 <= MUX1HOT_v_64_4_2(twiddle_rsc_0_1_i_q_d, twiddle_rsc_0_6_i_q_d,
            twiddle_rsc_0_12_i_q_d, COMP_LOOP_tmp_mux1h_4_itm_mx0w3, STD_LOGIC_VECTOR'(
            and_dcpl_175 & and_dcpl_180 & and_dcpl_277 & and_311_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( ((COMP_LOOP_tmp_nor_1_itm OR COMP_LOOP_tmp_nor_14_itm) AND (COMP_LOOP_10_tmp_mul_idiv_sva(1)))
          = '1' ) THEN
        tmp_33_sva_2 <= twiddle_rsc_0_2_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm) = '1' ) THEN
        tmp_33_sva_3 <= twiddle_rsc_0_3_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( ((COMP_LOOP_tmp_nor_3_itm OR COMP_LOOP_tmp_nor_16_itm) AND (COMP_LOOP_10_tmp_mul_idiv_sva(2)))
          = '1' ) THEN
        tmp_33_sva_4 <= twiddle_rsc_0_4_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_5 OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_itm) = '1' ) THEN
        tmp_33_sva_5 <= twiddle_rsc_0_5_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm) = '1' ) THEN
        tmp_33_sva_7 <= twiddle_rsc_0_7_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm) = '1' ) THEN
        tmp_33_sva_9 <= twiddle_rsc_0_9_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_5 OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm) = '1' ) THEN
        tmp_33_sva_10 <= twiddle_rsc_0_10_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm) = '1' ) THEN
        tmp_33_sva_15 <= twiddle_rsc_0_15_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_itm <= '0';
      ELSIF ( (and_dcpl_65 OR and_dcpl_181 OR and_dcpl_190 OR and_dcpl_183 OR and_dcpl_191
          OR and_dcpl_184 OR and_dcpl_192) = '1' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_nor_6_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_nor_cse, COMP_LOOP_or_27_cse);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_2463_nl, and_dcpl_57, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_tmp_mux1h_12_itm <= MUX1HOT_v_64_6_2(twiddle_rsc_0_0_i_q_d, tmp_33_sva_13,
            tmp_33_sva_1, tmp_33_sva_10, tmp_33_sva_11, tmp_33_sva_12, STD_LOGIC_VECTOR'(
            COMP_LOOP_tmp_or_33_nl & COMP_LOOP_tmp_and_55_nl & COMP_LOOP_tmp_and_56_nl
            & COMP_LOOP_tmp_and_57_nl & COMP_LOOP_tmp_and_58_nl & COMP_LOOP_tmp_and_59_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (and_dcpl_65 OR and_dcpl_189 OR COMP_LOOP_10_acc_8_itm_mx0c2 OR COMP_LOOP_10_acc_8_itm_mx0c3
          OR and_dcpl_70 OR and_dcpl_220 OR COMP_LOOP_10_acc_8_itm_mx0c6 OR and_dcpl_74
          OR and_dcpl_222 OR COMP_LOOP_10_acc_8_itm_mx0c9 OR and_dcpl_81 OR and_dcpl_223
          OR COMP_LOOP_10_acc_8_itm_mx0c12 OR and_dcpl_86 OR and_dcpl_225 OR COMP_LOOP_10_acc_8_itm_mx0c15
          OR and_dcpl_93 OR and_dcpl_226 OR COMP_LOOP_10_acc_8_itm_mx0c18 OR and_dcpl_95
          OR and_dcpl_227 OR COMP_LOOP_10_acc_8_itm_mx0c21 OR and_dcpl_100 OR and_dcpl_228
          OR COMP_LOOP_10_acc_8_itm_mx0c24 OR and_dcpl_102 OR and_dcpl_229 OR COMP_LOOP_10_acc_8_itm_mx0c27
          OR and_dcpl_108 OR and_dcpl_230 OR COMP_LOOP_10_acc_8_itm_mx0c30 OR and_dcpl_110
          OR and_dcpl_231 OR COMP_LOOP_10_acc_8_itm_mx0c33 OR and_dcpl_116 OR and_dcpl_232
          OR COMP_LOOP_10_acc_8_itm_mx0c36 OR and_dcpl_119 OR and_dcpl_233 OR COMP_LOOP_10_acc_8_itm_mx0c39
          OR and_dcpl_125 OR and_dcpl_234 OR COMP_LOOP_10_acc_8_itm_mx0c42 OR and_dcpl_127
          OR and_dcpl_235 OR and_dcpl_130 OR and_dcpl_236 OR COMP_LOOP_10_acc_8_itm_mx0c47)
          = '1' ) THEN
        COMP_LOOP_10_acc_8_itm <= MUX1HOT_v_64_19_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d,
            vec_rsc_0_2_i_q_d, vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d,
            vec_rsc_0_6_i_q_d, vec_rsc_0_7_i_q_d, vec_rsc_0_8_i_q_d, vec_rsc_0_9_i_q_d,
            vec_rsc_0_10_i_q_d, vec_rsc_0_11_i_q_d, vec_rsc_0_12_i_q_d, vec_rsc_0_13_i_q_d,
            vec_rsc_0_14_i_q_d, vec_rsc_0_15_i_q_d, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_acc_23_nl),
            64)), z_out_3, COMP_LOOP_1_modulo_cmp_return_rsc_z, STD_LOGIC_VECTOR'(
            COMP_LOOP_or_nl & COMP_LOOP_or_1_nl & COMP_LOOP_or_2_nl & COMP_LOOP_or_3_nl
            & COMP_LOOP_or_4_nl & COMP_LOOP_or_5_nl & COMP_LOOP_or_6_nl & COMP_LOOP_or_7_nl
            & COMP_LOOP_or_8_nl & COMP_LOOP_or_9_nl & COMP_LOOP_or_10_nl & COMP_LOOP_or_11_nl
            & COMP_LOOP_or_12_nl & COMP_LOOP_or_13_nl & COMP_LOOP_or_14_nl & COMP_LOOP_or_15_nl
            & COMP_LOOP_or_21_nl & COMP_LOOP_or_22_nl & COMP_LOOP_10_acc_8_itm_mx0c3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_11_tmp_mul_idiv_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( COMP_LOOP_tmp_or_19_cse = '1' ) THEN
        COMP_LOOP_11_tmp_mul_idiv_sva <= z_out_3(8 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( and_332_tmp = '0' ) THEN
        COMP_LOOP_tmp_mux1h_itm <= MUX1HOT_v_64_16_2(twiddle_rsc_0_0_i_q_d, tmp_33_sva_1,
            tmp_33_sva_2, tmp_33_sva_3, tmp_33_sva_4, tmp_33_sva_5, tmp_33_sva_6,
            tmp_33_sva_7, tmp_33_sva_8, tmp_33_sva_9, tmp_33_sva_10, tmp_33_sva_11,
            tmp_33_sva_12, tmp_33_sva_13, tmp_33_sva_14, tmp_33_sva_15, STD_LOGIC_VECTOR'(
            COMP_LOOP_tmp_and_42_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_1_nl
            & COMP_LOOP_tmp_and_43_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl & COMP_LOOP_tmp_and_44_nl
            & COMP_LOOP_tmp_and_45_nl & COMP_LOOP_tmp_and_46_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_7_nl
            & COMP_LOOP_tmp_and_47_nl & COMP_LOOP_tmp_and_48_nl & COMP_LOOP_tmp_and_49_nl
            & COMP_LOOP_tmp_and_50_nl & COMP_LOOP_tmp_and_51_nl & COMP_LOOP_tmp_and_52_nl
            & COMP_LOOP_tmp_and_53_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_2504_nl, (fsm_output(8)), or_2589_cse)) = '1' ) THEN
        COMP_LOOP_tmp_mux_itm <= MUX1HOT_v_64_3_2(tmp_33_sva_13_mx0w1, twiddle_rsc_0_8_i_q_d,
            twiddle_rsc_0_0_i_q_d, STD_LOGIC_VECTOR'( and_336_nl & and_dcpl_183 &
            and_340_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_13_tmp_mul_idiv_sva <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( (and_dcpl_189 OR and_dcpl_202) = '1' ) THEN
        COMP_LOOP_13_tmp_mul_idiv_sva <= MUX_v_8_2_2((z_out_1(7 DOWNTO 0)), (z_out_3(7
            DOWNTO 0)), and_dcpl_202);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_12_itm <= '0';
      ELSIF ( COMP_LOOP_tmp_or_21_cse = '1' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_19_cse, COMP_LOOP_or_31_cse);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_20_cse, COMP_LOOP_or_31_cse);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_21_cse, COMP_LOOP_or_31_cse);
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_12_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_nor_cse,
            COMP_LOOP_tmp_nor_6_cse, COMP_LOOP_or_31_cse);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_5_tmp_mul_idiv_sva <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( (NOT(or_dcpl_182 OR CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("10"))
          OR or_dcpl_207)) = '1' ) THEN
        COMP_LOOP_5_tmp_mul_idiv_sva <= z_out_3(7 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( and_341_tmp = '0' ) THEN
        COMP_LOOP_tmp_mux1h_1_itm <= MUX1HOT_v_64_6_2(twiddle_rsc_0_0_i_q_d, COMP_LOOP_tmp_mux_itm,
            tmp_33_sva_1, tmp_33_sva_10, tmp_33_sva_11, tmp_33_sva_12, STD_LOGIC_VECTOR'(
            COMP_LOOP_tmp_and_36_nl & COMP_LOOP_tmp_and_37_nl & COMP_LOOP_tmp_and_38_nl
            & COMP_LOOP_tmp_and_39_nl & COMP_LOOP_tmp_and_40_nl & COMP_LOOP_tmp_and_41_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( and_342_tmp = '0' ) THEN
        COMP_LOOP_tmp_mux1h_2_itm <= MUX1HOT_v_64_16_2(twiddle_rsc_0_0_i_q_d, tmp_33_sva_1,
            tmp_33_sva_2, tmp_33_sva_3, tmp_33_sva_4, tmp_33_sva_5, tmp_33_sva_6,
            tmp_33_sva_7, tmp_33_sva_8, tmp_33_sva_9, tmp_33_sva_10, tmp_33_sva_11,
            tmp_33_sva_12, tmp_33_sva_13, tmp_33_sva_14, tmp_33_sva_15, STD_LOGIC_VECTOR'(
            COMP_LOOP_tmp_and_20_nl & COMP_LOOP_tmp_and_21_nl & COMP_LOOP_tmp_and_22_nl
            & COMP_LOOP_tmp_and_23_nl & COMP_LOOP_tmp_and_24_nl & COMP_LOOP_tmp_and_25_nl
            & COMP_LOOP_tmp_and_26_nl & COMP_LOOP_tmp_and_27_nl & COMP_LOOP_tmp_and_28_nl
            & COMP_LOOP_tmp_and_29_nl & COMP_LOOP_tmp_and_30_nl & COMP_LOOP_tmp_and_31_nl
            & COMP_LOOP_tmp_and_32_nl & COMP_LOOP_tmp_and_33_nl & COMP_LOOP_tmp_and_34_nl
            & COMP_LOOP_tmp_and_35_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( ((COMP_LOOP_tmp_COMP_LOOP_tmp_nor_14_cse OR (CONV_SL_1_1(COMP_LOOP_13_tmp_mul_idiv_sva(1
          DOWNTO 0)=STD_LOGIC_VECTOR'("10"))) OR (CONV_SL_1_1(COMP_LOOP_13_tmp_mul_idiv_sva(1
          DOWNTO 0)=STD_LOGIC_VECTOR'("11"))) OR and_dcpl_277) AND mux_2518_nl) =
          '1' ) THEN
        tmp_36_sva_1 <= MUX1HOT_v_64_4_2(twiddle_rsc_0_4_i_q_d, twiddle_rsc_0_0_i_q_d,
            tmp_36_sva_2, tmp_33_sva_1, STD_LOGIC_VECTOR'( and_dcpl_277 & COMP_LOOP_tmp_and_nl
            & COMP_LOOP_tmp_and_17_nl & COMP_LOOP_tmp_and_18_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_2520_nl, and_357_nl, fsm_output(5))) = '1' ) THEN
        tmp_36_sva_2 <= MUX_v_64_2_2(twiddle_rsc_0_8_i_q_d, COMP_LOOP_tmp_mux1h_4_itm_mx0w3,
            and_dcpl_192);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_COMP_LOOP_tmp_nor_16_rgt OR COMP_LOOP_tmp_and_14_rgt OR
          COMP_LOOP_tmp_and_15_rgt OR COMP_LOOP_tmp_and_16_rgt) = '1' ) THEN
        COMP_LOOP_tmp_mux1h_3_itm <= MUX1HOT_v_64_4_2(twiddle_rsc_0_0_i_q_d, tmp_36_sva_1,
            tmp_36_sva_2, tmp_33_sva_1, STD_LOGIC_VECTOR'( COMP_LOOP_tmp_COMP_LOOP_tmp_nor_16_rgt
            & COMP_LOOP_tmp_and_14_rgt & COMP_LOOP_tmp_and_15_rgt & COMP_LOOP_tmp_and_16_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_2532_nl OR (fsm_output(8))) = '1' ) THEN
        COMP_LOOP_tmp_mux1h_4_itm <= COMP_LOOP_tmp_mux1h_4_itm_mx0w3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( nor_1796_tmp = '0' ) THEN
        COMP_LOOP_tmp_mux1h_5_itm <= MUX1HOT_v_64_6_2(twiddle_rsc_0_0_i_q_d, COMP_LOOP_tmp_mux_itm,
            tmp_33_sva_1, tmp_33_sva_10, tmp_33_sva_11, tmp_33_sva_12, STD_LOGIC_VECTOR'(
            COMP_LOOP_tmp_and_7_nl & COMP_LOOP_tmp_and_8_nl & COMP_LOOP_tmp_and_9_nl
            & COMP_LOOP_tmp_and_10_nl & COMP_LOOP_tmp_and_11_nl & COMP_LOOP_tmp_and_12_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_2542_nl OR (fsm_output(8))) = '1' ) THEN
        COMP_LOOP_tmp_mux1h_6_itm <= COMP_LOOP_tmp_mux1h_4_itm_mx0w3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_2546_nl, and_352_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_tmp_mux1h_7_itm <= COMP_LOOP_tmp_mux1h_4_itm_mx0w3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (((NOT(COMP_LOOP_tmp_COMP_LOOP_tmp_and_155 OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_157
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_159)) OR COMP_LOOP_tmp_COMP_LOOP_tmp_nor_12_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm
          OR and_dcpl_191) AND mux_2553_nl) = '1' ) THEN
        COMP_LOOP_tmp_mux1h_8_itm <= MUX1HOT_v_64_6_2(tmp_33_sva_13_mx0w1, twiddle_rsc_0_0_i_q_d,
            tmp_33_sva_1, tmp_33_sva_10, tmp_33_sva_11, tmp_33_sva_12, STD_LOGIC_VECTOR'(
            and_dcpl_191 & COMP_LOOP_tmp_and_2_nl & COMP_LOOP_tmp_and_3_nl & COMP_LOOP_tmp_and_4_nl
            & COMP_LOOP_tmp_and_5_nl & COMP_LOOP_tmp_and_6_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_2556_nl, mux_2554_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_tmp_mux1h_9_itm <= COMP_LOOP_tmp_mux1h_4_itm_mx0w3;
      END IF;
    END IF;
  END PROCESS;
  nor_1871_nl <= NOT((fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(2))
      OR (fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(8)));
  and_1183_nl <= (fsm_output(4)) AND mux_tmp_1062;
  VEC_LOOP_j_not_1_nl <= NOT VEC_LOOP_j_10_0_sva_9_0_mx0c0;
  nor_1870_nl <= NOT((fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(1))
      OR (fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(8)));
  and_nl <= (fsm_output(4)) AND nor_tmp_339;
  nor_1622_nl <= NOT((fsm_output(4)) OR (fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(7))
      OR (fsm_output(8)));
  and_568_nl <= (fsm_output(4)) AND (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(7))
      AND (fsm_output(8));
  mux_1074_nl <= MUX_s_1_2_2(nor_1622_nl, and_568_nl, fsm_output(5));
  nand_nl <= NOT(mux_1074_nl AND nor_1624_cse AND (fsm_output(0)));
  or_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")) OR (NOT(CONV_SL_1_1(fsm_output(3
      DOWNTO 1)/=STD_LOGIC_VECTOR'("000"))));
  mux_2558_nl <= MUX_s_1_2_2(or_nl, nand_324_cse, fsm_output(5));
  nand_325_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111"))
      AND or_2259_cse_1);
  nand_323_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 6)=STD_LOGIC_VECTOR'("111"))
      AND (NOT(and_1189_cse OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")))));
  mux_nl <= MUX_s_1_2_2(nand_325_nl, nand_323_nl, fsm_output(5));
  mux_2308_nl <= MUX_s_1_2_2(mux_tmp_2288, nor_tmp_489, fsm_output(4));
  mux_2309_nl <= MUX_s_1_2_2(mux_2308_nl, (fsm_output(7)), fsm_output(5));
  and_270_nl <= (fsm_output(4)) AND mux_tmp_2291;
  mux_2312_nl <= MUX_s_1_2_2(not_tmp_703, and_270_nl, fsm_output(5));
  nand_320_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111")));
  mux_2314_nl <= MUX_s_1_2_2(or_tmp_2300, nand_320_nl, fsm_output(5));
  nand_111_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1111")));
  mux_2315_nl <= MUX_s_1_2_2(or_tmp_2300, nand_111_nl, fsm_output(5));
  COMP_LOOP_3_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0
      & STD_LOGIC_VECTOR'( "0010")), 10), 11) + SIGNED'( "00000000001"), 11));
  mux_2316_nl <= MUX_s_1_2_2((NOT mux_tmp_2292), nor_tmp_10, fsm_output(4));
  mux_2317_nl <= MUX_s_1_2_2(mux_2316_nl, (fsm_output(6)), fsm_output(5));
  mux_2318_nl <= MUX_s_1_2_2((NOT mux_tmp_2292), mux_tmp_2291, fsm_output(4));
  mux_2319_nl <= MUX_s_1_2_2(mux_2318_nl, (fsm_output(6)), fsm_output(5));
  COMP_LOOP_acc_12_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 3)))) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0
      & STD_LOGIC_VECTOR'( "00")), 8), 9) + UNSIGNED'( "000000001"), 9));
  nand_110_nl <= NOT((fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(2)) AND
      (fsm_output(1)) AND (fsm_output(6)));
  mux_2320_nl <= MUX_s_1_2_2(mux_tmp_2292, nand_110_nl, fsm_output(4));
  mux_2321_nl <= MUX_s_1_2_2(mux_2320_nl, (NOT (fsm_output(6))), fsm_output(5));
  and_823_nl <= (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(4)) AND (fsm_output(6));
  mux_2326_nl <= MUX_s_1_2_2(not_tmp_703, and_823_nl, fsm_output(5));
  COMP_LOOP_5_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0
      & STD_LOGIC_VECTOR'( "0100")), 10), 11) + SIGNED'( "00000000001"), 11));
  and_412_nl <= (fsm_output(4)) AND (fsm_output(3)) AND (fsm_output(2)) AND (fsm_output(1))
      AND (fsm_output(6));
  mux_2327_nl <= MUX_s_1_2_2(not_tmp_703, and_412_nl, fsm_output(5));
  mux_2331_nl <= MUX_s_1_2_2(mux_tmp_2288, mux_tmp_2311, fsm_output(4));
  mux_2332_nl <= MUX_s_1_2_2(mux_2331_nl, (fsm_output(7)), fsm_output(5));
  COMP_LOOP_6_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0
      & STD_LOGIC_VECTOR'( "0101")), 10), 11) + SIGNED'( "00000000001"), 11));
  and_408_nl <= (and_831_cse OR (fsm_output(6))) AND (fsm_output(7));
  mux_2333_nl <= MUX_s_1_2_2(and_408_nl, nor_tmp_489, fsm_output(0));
  mux_2334_nl <= MUX_s_1_2_2(mux_tmp_2288, mux_2333_nl, fsm_output(4));
  mux_2335_nl <= MUX_s_1_2_2(mux_2334_nl, (fsm_output(7)), fsm_output(5));
  mux_2336_nl <= MUX_s_1_2_2(nor_tmp_47, mux_tmp_2311, fsm_output(4));
  mux_2338_nl <= MUX_s_1_2_2(mux_tmp_2318, mux_2336_nl, fsm_output(5));
  mux_2339_nl <= MUX_s_1_2_2(nor_tmp_47, nor_tmp_499, and_407_cse);
  mux_2340_nl <= MUX_s_1_2_2(mux_tmp_2318, mux_2339_nl, fsm_output(5));
  COMP_LOOP_7_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0
      & STD_LOGIC_VECTOR'( "0110")), 10), 11) + SIGNED'( "00000000001"), 11));
  and_405_nl <= ((CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111"))) OR
      (fsm_output(6))) AND (fsm_output(7));
  mux_2341_nl <= MUX_s_1_2_2(mux_tmp_2318, and_405_nl, fsm_output(5));
  mux_2345_nl <= MUX_s_1_2_2((NOT mux_tmp_2325), and_tmp_28, fsm_output(4));
  mux_2346_nl <= MUX_s_1_2_2(mux_2345_nl, nor_tmp_47, fsm_output(5));
  mux_2348_nl <= MUX_s_1_2_2((NOT mux_tmp_2325), mux_tmp_2328, fsm_output(4));
  mux_2349_nl <= MUX_s_1_2_2(mux_2348_nl, nor_tmp_47, fsm_output(5));
  COMP_LOOP_acc_15_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 4)))) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0
      & '0'), 7), 8) + UNSIGNED'( "00000001"), 8));
  mux_2350_nl <= MUX_s_1_2_2(nor_tmp_509, and_tmp_28, fsm_output(0));
  mux_2351_nl <= MUX_s_1_2_2((NOT mux_tmp_2325), mux_2350_nl, fsm_output(4));
  mux_2352_nl <= MUX_s_1_2_2(mux_2351_nl, nor_tmp_47, fsm_output(5));
  and_296_nl <= (fsm_output(4)) AND mux_tmp_2328;
  mux_2354_nl <= MUX_s_1_2_2(not_tmp_727, and_296_nl, fsm_output(5));
  and_397_nl <= (fsm_output(4)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(7));
  mux_2355_nl <= MUX_s_1_2_2(not_tmp_727, and_397_nl, fsm_output(5));
  COMP_LOOP_9_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0
      & STD_LOGIC_VECTOR'( "1000")), 10), 11) + SIGNED'( "00000000001"), 11));
  and_299_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11")) AND nor_tmp_507;
  mux_2356_nl <= MUX_s_1_2_2(not_tmp_727, and_299_nl, fsm_output(5));
  mux_2364_nl <= MUX_s_1_2_2(mux_tmp_2344, nor_tmp_515, fsm_output(4));
  mux_2368_nl <= MUX_s_1_2_2(mux_tmp_2344, mux_tmp_2348, fsm_output(4));
  COMP_LOOP_10_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0
      & STD_LOGIC_VECTOR'( "1001")), 10), 11) + SIGNED'( "00000000001"), 11));
  mux_2371_nl <= MUX_s_1_2_2(mux_tmp_2351, nor_tmp_515, fsm_output(0));
  mux_2372_nl <= MUX_s_1_2_2(mux_tmp_2344, mux_2371_nl, fsm_output(4));
  mux_2375_nl <= MUX_s_1_2_2(nor_tmp_115, mux_tmp_2348, fsm_output(4));
  mux_2378_nl <= MUX_s_1_2_2(nor_tmp_115, mux_tmp_2347, fsm_output(4));
  COMP_LOOP_11_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0
      & STD_LOGIC_VECTOR'( "1010")), 10), 11) + SIGNED'( "00000000001"), 11));
  and_390_nl <= (and_407_cse OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")))
      AND (fsm_output(8));
  mux_2389_nl <= MUX_s_1_2_2(mux_tmp_2369, mux_tmp_2365, fsm_output(4));
  mux_2391_nl <= MUX_s_1_2_2(mux_tmp_2365, nor_tmp_528, fsm_output(0));
  mux_2392_nl <= MUX_s_1_2_2(mux_tmp_2369, mux_2391_nl, fsm_output(4));
  COMP_LOOP_acc_18_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 3)))) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0
      & STD_LOGIC_VECTOR'( "10")), 8), 9) + UNSIGNED'( "000000001"), 9));
  mux_2394_nl <= MUX_s_1_2_2(nor_tmp_530, mux_tmp_2365, fsm_output(0));
  mux_2395_nl <= MUX_s_1_2_2(mux_tmp_2369, mux_2394_nl, fsm_output(4));
  nor_581_nl <= NOT(and_1189_cse OR (fsm_output(4)) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(8)));
  and_379_nl <= (CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))) AND
      (fsm_output(4)) AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(8));
  mux_2399_nl <= MUX_s_1_2_2(nor_581_nl, and_379_nl, fsm_output(2));
  and_380_nl <= (fsm_output(4)) AND (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(8));
  mux_2400_nl <= MUX_s_1_2_2(mux_2399_nl, and_380_nl, fsm_output(3));
  mux_2402_nl <= MUX_s_1_2_2(and_733_cse, nor_tmp_528, fsm_output(4));
  COMP_LOOP_13_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0
      & STD_LOGIC_VECTOR'( "1100")), 10), 11) + SIGNED'( "00000000001"), 11));
  mux_2405_nl <= MUX_s_1_2_2(and_733_cse, mux_tmp_2365, fsm_output(4));
  mux_2415_nl <= MUX_s_1_2_2(mux_tmp_2395, nor_tmp_537, fsm_output(4));
  mux_2417_nl <= MUX_s_1_2_2(nor_tmp_537, nor_tmp_538, fsm_output(0));
  mux_2418_nl <= MUX_s_1_2_2(mux_tmp_2395, mux_2417_nl, fsm_output(4));
  COMP_LOOP_14_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0
      & STD_LOGIC_VECTOR'( "1101")), 10), 11) + SIGNED'( "00000000001"), 11));
  mux_2421_nl <= MUX_s_1_2_2(mux_tmp_2401, nor_tmp_537, fsm_output(0));
  mux_2422_nl <= MUX_s_1_2_2(mux_tmp_2395, mux_2421_nl, fsm_output(4));
  nor_580_nl <= NOT((fsm_output(4)) OR (fsm_output(5)) OR (fsm_output(7)) OR (fsm_output(8)));
  mux_2425_nl <= MUX_s_1_2_2(nor_580_nl, nor_tmp_544, and_1189_cse);
  mux_2426_nl <= MUX_s_1_2_2(mux_2425_nl, nor_tmp_544, or_2259_cse_1);
  mux_2428_nl <= MUX_s_1_2_2(and_dcpl_57, nor_tmp_538, fsm_output(4));
  COMP_LOOP_15_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0
      & STD_LOGIC_VECTOR'( "1110")), 10), 11) + SIGNED'( "00000000001"), 11));
  mux_2431_nl <= MUX_s_1_2_2(and_dcpl_57, nor_tmp_537, fsm_output(4));
  mux_2436_nl <= MUX_s_1_2_2((NOT mux_tmp_2282), nor_tmp_547, fsm_output(4));
  mux_2438_nl <= MUX_s_1_2_2((NOT mux_tmp_2282), nor_tmp_548, fsm_output(4));
  COMP_LOOP_acc_21_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 5)))) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_4_sva_5_0),
      6), 7) + UNSIGNED'( "0000001"), 7));
  and_303_nl <= (fsm_output(4)) AND nor_tmp_548;
  and_363_nl <= (fsm_output(4)) AND (fsm_output(6)) AND (fsm_output(7)) AND (fsm_output(8));
  COMP_LOOP_1_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(COMP_LOOP_k_10_4_sva_2
      & STD_LOGIC_VECTOR'( "0000")) + SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + SIGNED'( "00000000001"), 11));
  and_304_nl <= (fsm_output(4)) AND nor_tmp_547;
  COMP_LOOP_COMP_LOOP_and_23_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO
      0)=STD_LOGIC_VECTOR'("1001"));
  COMP_LOOP_COMP_LOOP_and_24_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO
      0)=STD_LOGIC_VECTOR'("1010"));
  COMP_LOOP_COMP_LOOP_and_25_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO
      0)=STD_LOGIC_VECTOR'("1011"));
  COMP_LOOP_COMP_LOOP_and_26_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO
      0)=STD_LOGIC_VECTOR'("1100"));
  COMP_LOOP_COMP_LOOP_and_27_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO
      0)=STD_LOGIC_VECTOR'("1101"));
  COMP_LOOP_COMP_LOOP_and_28_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO
      0)=STD_LOGIC_VECTOR'("1110"));
  COMP_LOOP_COMP_LOOP_and_29_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO
      0)=STD_LOGIC_VECTOR'("1111"));
  COMP_LOOP_nor_11_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
  COMP_LOOP_nor_12_nl <= NOT((COMP_LOOP_1_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_1_acc_10_itm_10_1_1(2))
      OR (COMP_LOOP_1_acc_10_itm_10_1_1(0)));
  COMP_LOOP_nor_14_nl <= NOT((COMP_LOOP_1_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_1_acc_10_itm_10_1_1(1))
      OR (COMP_LOOP_1_acc_10_itm_10_1_1(0)));
  COMP_LOOP_nor_17_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
  COMP_LOOP_COMP_LOOP_and_17_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO
      0)=STD_LOGIC_VECTOR'("0011"));
  COMP_LOOP_COMP_LOOP_and_19_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO
      0)=STD_LOGIC_VECTOR'("0101"));
  COMP_LOOP_COMP_LOOP_and_20_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO
      0)=STD_LOGIC_VECTOR'("0110"));
  COMP_LOOP_COMP_LOOP_and_21_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO
      0)=STD_LOGIC_VECTOR'("0111"));
  COMP_LOOP_COMP_LOOP_nor_1_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
  and_311_nl <= and_dcpl_61 AND and_dcpl_123;
  or_2758_nl <= (fsm_output(0)) OR (fsm_output(2));
  mux_2564_nl <= MUX_s_1_2_2(or_2259_cse_1, or_2758_nl, fsm_output(1));
  or_2756_nl <= (NOT (COMP_LOOP_10_tmp_mul_idiv_sva(3))) OR (NOT COMP_LOOP_tmp_nor_19_itm)
      OR (fsm_output(3)) OR (fsm_output(0)) OR (fsm_output(2));
  mux_2560_nl <= MUX_s_1_2_2(or_2756_nl, or_tmp_2410, and_1190_cse);
  mux_2561_nl <= MUX_s_1_2_2(mux_2560_nl, or_tmp_2410, and_1191_cse);
  or_2754_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm
      OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm
      OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm
      OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm
      OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm
      OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm;
  mux_2562_nl <= MUX_s_1_2_2(mux_2561_nl, or_tmp_2410, or_2754_nl);
  mux_2563_nl <= MUX_s_1_2_2(or_2259_cse_1, mux_2562_nl, fsm_output(1));
  mux_2565_nl <= MUX_s_1_2_2(mux_2564_nl, (NOT mux_2563_nl), fsm_output(4));
  COMP_LOOP_tmp_or_33_nl <= and_dcpl_65 OR (COMP_LOOP_tmp_COMP_LOOP_tmp_nor_12_itm
      AND and_314_m1c);
  COMP_LOOP_tmp_and_55_nl <= COMP_LOOP_tmp_or_29_cse AND and_314_m1c;
  COMP_LOOP_tmp_and_56_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm AND and_314_m1c;
  COMP_LOOP_tmp_and_57_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm AND and_314_m1c;
  COMP_LOOP_tmp_and_58_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm AND and_314_m1c;
  COMP_LOOP_tmp_and_59_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm AND and_314_m1c;
  mux_2461_nl <= MUX_s_1_2_2(and_dcpl_5, and_dcpl_57, or_2259_cse_1);
  mux_2459_nl <= MUX_s_1_2_2(and_dcpl_5, mux_tmp_2392, fsm_output(1));
  mux_2460_nl <= MUX_s_1_2_2(mux_2459_nl, and_dcpl_57, or_2259_cse_1);
  mux_2462_nl <= MUX_s_1_2_2(mux_2461_nl, mux_2460_nl, fsm_output(0));
  or_2563_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"));
  mux_2458_nl <= MUX_s_1_2_2(mux_tmp_2392, and_dcpl_57, or_2563_nl);
  mux_2463_nl <= MUX_s_1_2_2(mux_2462_nl, mux_2458_nl, fsm_output(4));
  COMP_LOOP_COMP_LOOP_mux_9_nl <= MUX_v_64_2_2(COMP_LOOP_10_acc_8_itm, z_out_7, COMP_LOOP_or_18_itm);
  COMP_LOOP_acc_23_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_361_cse)
      + UNSIGNED(COMP_LOOP_COMP_LOOP_mux_9_nl), 64));
  COMP_LOOP_or_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm AND and_dcpl_65) OR
      (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_70) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_dcpl_74) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_81) OR (COMP_LOOP_COMP_LOOP_and_72_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_93) OR (COMP_LOOP_COMP_LOOP_and_70_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_69_itm AND and_dcpl_100) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_dcpl_102) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_108) OR (COMP_LOOP_COMP_LOOP_and_66_itm
      AND and_dcpl_110) OR (COMP_LOOP_COMP_LOOP_and_65_itm AND and_dcpl_116) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_dcpl_119) OR (COMP_LOOP_COMP_LOOP_and_185_itm AND and_dcpl_125) OR
      (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_127) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_130);
  COMP_LOOP_or_1_nl <= ((COMP_LOOP_acc_10_cse_10_1_1_sva(0)) AND COMP_LOOP_tmp_nor_13_itm
      AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_70) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_74) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_81) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_72_itm AND and_dcpl_93) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_70_itm AND and_dcpl_100) OR (COMP_LOOP_COMP_LOOP_and_69_itm
      AND and_dcpl_102) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_108) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_110) OR (COMP_LOOP_COMP_LOOP_and_66_itm AND and_dcpl_116) OR (COMP_LOOP_COMP_LOOP_and_65_itm
      AND and_dcpl_119) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_125) OR (COMP_LOOP_COMP_LOOP_and_185_itm
      AND and_dcpl_127) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_130);
  COMP_LOOP_or_2_nl <= ((COMP_LOOP_acc_10_cse_10_1_1_sva(1)) AND COMP_LOOP_tmp_nor_14_itm
      AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_dcpl_70) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_dcpl_74) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_81) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_93) OR (COMP_LOOP_COMP_LOOP_and_72_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_100) OR (COMP_LOOP_COMP_LOOP_and_70_itm
      AND and_dcpl_102) OR (COMP_LOOP_COMP_LOOP_and_69_itm AND and_dcpl_108) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_dcpl_110) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_116) OR (COMP_LOOP_COMP_LOOP_and_66_itm
      AND and_dcpl_119) OR (COMP_LOOP_COMP_LOOP_and_65_itm AND and_dcpl_125) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_dcpl_127) OR (COMP_LOOP_COMP_LOOP_and_185_itm AND and_dcpl_130);
  COMP_LOOP_or_3_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm AND and_dcpl_65)
      OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_70) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_74) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_81) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_93) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_72_itm AND and_dcpl_100) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_102) OR (COMP_LOOP_COMP_LOOP_and_70_itm AND and_dcpl_108) OR (COMP_LOOP_COMP_LOOP_and_69_itm
      AND and_dcpl_110) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_116) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_119) OR (COMP_LOOP_COMP_LOOP_and_66_itm AND and_dcpl_125) OR (COMP_LOOP_COMP_LOOP_and_65_itm
      AND and_dcpl_127) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_130);
  COMP_LOOP_or_4_nl <= ((COMP_LOOP_acc_10_cse_10_1_1_sva(2)) AND COMP_LOOP_tmp_nor_16_itm
      AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_185_itm AND and_dcpl_70) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_dcpl_74) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_dcpl_81) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_93) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_100) OR (COMP_LOOP_COMP_LOOP_and_72_itm
      AND and_dcpl_102) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_108) OR (COMP_LOOP_COMP_LOOP_and_70_itm
      AND and_dcpl_110) OR (COMP_LOOP_COMP_LOOP_and_69_itm AND and_dcpl_116) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_dcpl_119) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_125) OR (COMP_LOOP_COMP_LOOP_and_66_itm
      AND and_dcpl_127) OR (COMP_LOOP_COMP_LOOP_and_65_itm AND and_dcpl_130);
  COMP_LOOP_or_5_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm AND and_dcpl_65)
      OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_70) OR (COMP_LOOP_COMP_LOOP_and_185_itm
      AND and_dcpl_74) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_81) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_93) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_100) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_102) OR (COMP_LOOP_COMP_LOOP_and_72_itm AND and_dcpl_108) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_110) OR (COMP_LOOP_COMP_LOOP_and_70_itm AND and_dcpl_116) OR (COMP_LOOP_COMP_LOOP_and_69_itm
      AND and_dcpl_119) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_125) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_127) OR (COMP_LOOP_COMP_LOOP_and_66_itm AND and_dcpl_130);
  COMP_LOOP_or_6_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm AND and_dcpl_65)
      OR (COMP_LOOP_COMP_LOOP_and_65_itm AND and_dcpl_70) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_dcpl_74) OR (COMP_LOOP_COMP_LOOP_and_185_itm AND and_dcpl_81) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_dcpl_93) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_100) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_dcpl_102) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_108) OR (COMP_LOOP_COMP_LOOP_and_72_itm
      AND and_dcpl_110) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_116) OR (COMP_LOOP_COMP_LOOP_and_70_itm
      AND and_dcpl_119) OR (COMP_LOOP_COMP_LOOP_and_69_itm AND and_dcpl_125) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_dcpl_127) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_130);
  COMP_LOOP_or_7_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm AND and_dcpl_65)
      OR (COMP_LOOP_COMP_LOOP_and_66_itm AND and_dcpl_70) OR (COMP_LOOP_COMP_LOOP_and_65_itm
      AND and_dcpl_74) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_81) OR (COMP_LOOP_COMP_LOOP_and_185_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_93) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_100) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_102) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_108) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_110) OR (COMP_LOOP_COMP_LOOP_and_72_itm AND and_dcpl_116) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_119) OR (COMP_LOOP_COMP_LOOP_and_70_itm AND and_dcpl_125) OR (COMP_LOOP_COMP_LOOP_and_69_itm
      AND and_dcpl_127) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_130);
  COMP_LOOP_or_8_nl <= ((COMP_LOOP_acc_10_cse_10_1_1_sva(3)) AND COMP_LOOP_tmp_nor_19_itm
      AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_70) OR (COMP_LOOP_COMP_LOOP_and_66_itm
      AND and_dcpl_74) OR (COMP_LOOP_COMP_LOOP_and_65_itm AND and_dcpl_81) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_185_itm AND and_dcpl_93) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_dcpl_100) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_dcpl_102) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_108) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_dcpl_110) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_116) OR (COMP_LOOP_COMP_LOOP_and_72_itm
      AND and_dcpl_119) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_125) OR (COMP_LOOP_COMP_LOOP_and_70_itm
      AND and_dcpl_127) OR (COMP_LOOP_COMP_LOOP_and_69_itm AND and_dcpl_130);
  COMP_LOOP_or_9_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm AND and_dcpl_65)
      OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_70) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_74) OR (COMP_LOOP_COMP_LOOP_and_66_itm AND and_dcpl_81) OR (COMP_LOOP_COMP_LOOP_and_65_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_93) OR (COMP_LOOP_COMP_LOOP_and_185_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_100) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_102) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_108) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_110) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_116) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_119) OR (COMP_LOOP_COMP_LOOP_and_72_itm AND and_dcpl_125) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_127) OR (COMP_LOOP_COMP_LOOP_and_70_itm AND and_dcpl_130);
  COMP_LOOP_or_10_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm AND and_dcpl_65)
      OR (COMP_LOOP_COMP_LOOP_and_69_itm AND and_dcpl_70) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_dcpl_74) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_81) OR (COMP_LOOP_COMP_LOOP_and_66_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_65_itm AND and_dcpl_93) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_185_itm AND and_dcpl_100) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_dcpl_102) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_dcpl_108) OR
      (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_110) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_116) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_119) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_125) OR (COMP_LOOP_COMP_LOOP_and_72_itm AND and_dcpl_127) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_130);
  COMP_LOOP_or_11_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm AND and_dcpl_65)
      OR (COMP_LOOP_COMP_LOOP_and_70_itm AND and_dcpl_70) OR (COMP_LOOP_COMP_LOOP_and_69_itm
      AND and_dcpl_74) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_81) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_66_itm AND and_dcpl_93) OR (COMP_LOOP_COMP_LOOP_and_65_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_100) OR (COMP_LOOP_COMP_LOOP_and_185_itm
      AND and_dcpl_102) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_108) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_110) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_116) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_119) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_125) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_127) OR (COMP_LOOP_COMP_LOOP_and_72_itm AND and_dcpl_130);
  COMP_LOOP_or_12_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm AND and_dcpl_65)
      OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_70) OR (COMP_LOOP_COMP_LOOP_and_70_itm
      AND and_dcpl_74) OR (COMP_LOOP_COMP_LOOP_and_69_itm AND and_dcpl_81) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_93) OR (COMP_LOOP_COMP_LOOP_and_66_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_65_itm AND and_dcpl_100) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_dcpl_102) OR (COMP_LOOP_COMP_LOOP_and_185_itm AND and_dcpl_108) OR
      (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_110) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_116) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_119) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_125) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_127) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_130);
  COMP_LOOP_or_13_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm AND and_dcpl_65)
      OR (COMP_LOOP_COMP_LOOP_and_72_itm AND and_dcpl_70) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_74) OR (COMP_LOOP_COMP_LOOP_and_70_itm AND and_dcpl_81) OR (COMP_LOOP_COMP_LOOP_and_69_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_93) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_66_itm AND and_dcpl_100) OR (COMP_LOOP_COMP_LOOP_and_65_itm
      AND and_dcpl_102) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_108) OR (COMP_LOOP_COMP_LOOP_and_185_itm
      AND and_dcpl_110) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_116) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_119) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_125) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_127) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_130);
  COMP_LOOP_or_14_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm AND and_dcpl_65)
      OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_70) OR (COMP_LOOP_COMP_LOOP_and_72_itm
      AND and_dcpl_74) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_81) OR (COMP_LOOP_COMP_LOOP_and_70_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_69_itm AND and_dcpl_93) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_100) OR (COMP_LOOP_COMP_LOOP_and_66_itm
      AND and_dcpl_102) OR (COMP_LOOP_COMP_LOOP_and_65_itm AND and_dcpl_108) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_dcpl_110) OR (COMP_LOOP_COMP_LOOP_and_185_itm AND and_dcpl_116) OR
      (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_119) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_125) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_127) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_130);
  COMP_LOOP_or_15_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm AND and_dcpl_65)
      OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_70) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_74) OR (COMP_LOOP_COMP_LOOP_and_72_itm AND and_dcpl_81) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_70_itm AND and_dcpl_93) OR (COMP_LOOP_COMP_LOOP_and_69_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_100) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_102) OR (COMP_LOOP_COMP_LOOP_and_66_itm AND and_dcpl_108) OR (COMP_LOOP_COMP_LOOP_and_65_itm
      AND and_dcpl_110) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_116) OR (COMP_LOOP_COMP_LOOP_and_185_itm
      AND and_dcpl_119) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_125) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_127) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_130);
  COMP_LOOP_or_21_nl <= and_dcpl_189 OR and_dcpl_220 OR and_dcpl_222 OR and_dcpl_223
      OR and_dcpl_225 OR and_dcpl_226 OR and_dcpl_227 OR and_dcpl_228 OR and_dcpl_229
      OR and_dcpl_230 OR and_dcpl_231 OR and_dcpl_232 OR and_dcpl_233 OR and_dcpl_234
      OR and_dcpl_235 OR and_dcpl_236;
  COMP_LOOP_or_22_nl <= COMP_LOOP_10_acc_8_itm_mx0c2 OR COMP_LOOP_10_acc_8_itm_mx0c6
      OR COMP_LOOP_10_acc_8_itm_mx0c9 OR COMP_LOOP_10_acc_8_itm_mx0c12 OR COMP_LOOP_10_acc_8_itm_mx0c15
      OR COMP_LOOP_10_acc_8_itm_mx0c18 OR COMP_LOOP_10_acc_8_itm_mx0c21 OR COMP_LOOP_10_acc_8_itm_mx0c24
      OR COMP_LOOP_10_acc_8_itm_mx0c27 OR COMP_LOOP_10_acc_8_itm_mx0c30 OR COMP_LOOP_10_acc_8_itm_mx0c33
      OR COMP_LOOP_10_acc_8_itm_mx0c36 OR COMP_LOOP_10_acc_8_itm_mx0c39 OR COMP_LOOP_10_acc_8_itm_mx0c42
      OR COMP_LOOP_10_acc_8_itm_mx0c47;
  COMP_LOOP_tmp_and_42_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_itm AND (NOT and_332_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_nl <= (COMP_LOOP_10_tmp_mul_idiv_sva(0)) AND COMP_LOOP_tmp_nor_itm
      AND (NOT and_332_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_1_nl <= (COMP_LOOP_10_tmp_mul_idiv_sva(1)) AND
      COMP_LOOP_tmp_nor_1_itm AND (NOT and_332_tmp);
  COMP_LOOP_tmp_and_43_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_itm AND (NOT and_332_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl <= (COMP_LOOP_10_tmp_mul_idiv_sva(2)) AND
      COMP_LOOP_tmp_nor_3_itm AND (NOT and_332_tmp);
  COMP_LOOP_tmp_and_44_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_itm AND (NOT and_332_tmp);
  COMP_LOOP_tmp_and_45_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_itm AND (NOT and_332_tmp);
  COMP_LOOP_tmp_and_46_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_itm AND (NOT and_332_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_7_nl <= (COMP_LOOP_10_tmp_mul_idiv_sva(3)) AND
      COMP_LOOP_tmp_nor_6_itm AND (NOT and_332_tmp);
  COMP_LOOP_tmp_and_47_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_itm AND (NOT and_332_tmp);
  COMP_LOOP_tmp_and_48_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_9_itm AND (NOT and_332_tmp);
  COMP_LOOP_tmp_and_49_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_itm AND (NOT and_332_tmp);
  COMP_LOOP_tmp_and_50_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_itm AND (NOT and_332_tmp);
  COMP_LOOP_tmp_and_51_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_itm AND (NOT and_332_tmp);
  COMP_LOOP_tmp_and_52_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_itm AND (NOT and_332_tmp);
  COMP_LOOP_tmp_and_53_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_itm AND (NOT and_332_tmp);
  and_336_nl <= and_dcpl_5 AND ((fsm_output(2)) XOR (fsm_output(3))) AND CONV_SL_1_1(fsm_output(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("00")) AND and_dcpl_45;
  and_340_nl <= and_dcpl_61 AND (NOT (COMP_LOOP_9_tmp_lshift_itm(0))) AND (fsm_output(3))
      AND (fsm_output(0)) AND and_dcpl_45;
  or_2595_nl <= nor_572_cse OR (fsm_output(8));
  mux_2501_nl <= MUX_s_1_2_2(mux_tmp_439, or_2595_nl, fsm_output(1));
  mux_2502_nl <= MUX_s_1_2_2(mux_2501_nl, (fsm_output(8)), fsm_output(2));
  mux_2503_nl <= MUX_s_1_2_2(mux_tmp_439, mux_2502_nl, fsm_output(3));
  or_2593_nl <= (NOT((fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(7)))) OR (fsm_output(8));
  or_2591_nl <= (NOT((fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(7))))
      OR (fsm_output(8));
  mux_2499_nl <= MUX_s_1_2_2(or_2593_nl, or_2591_nl, COMP_LOOP_9_tmp_lshift_itm(0));
  mux_2500_nl <= MUX_s_1_2_2(mux_tmp_439, mux_2499_nl, fsm_output(3));
  mux_2504_nl <= MUX_s_1_2_2(mux_2503_nl, mux_2500_nl, fsm_output(0));
  COMP_LOOP_tmp_and_36_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_itm AND (NOT and_341_tmp);
  COMP_LOOP_tmp_and_37_nl <= COMP_LOOP_tmp_or_29_cse AND (NOT and_341_tmp);
  COMP_LOOP_tmp_and_38_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm AND (NOT and_341_tmp);
  COMP_LOOP_tmp_and_39_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm AND (NOT and_341_tmp);
  COMP_LOOP_tmp_and_40_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm AND (NOT and_341_tmp);
  COMP_LOOP_tmp_and_41_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm AND (NOT and_341_tmp);
  COMP_LOOP_tmp_and_20_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_12_itm AND (NOT and_342_tmp);
  COMP_LOOP_tmp_and_21_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_167 AND (NOT and_342_tmp);
  COMP_LOOP_tmp_and_22_nl <= and_1191_cse AND (NOT and_342_tmp);
  COMP_LOOP_tmp_and_23_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm AND (NOT and_342_tmp);
  COMP_LOOP_tmp_and_24_nl <= and_1190_cse AND (NOT and_342_tmp);
  COMP_LOOP_tmp_and_25_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm AND (NOT and_342_tmp);
  COMP_LOOP_tmp_and_26_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm AND (NOT and_342_tmp);
  COMP_LOOP_tmp_and_27_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm AND (NOT and_342_tmp);
  COMP_LOOP_tmp_and_28_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_161 AND (NOT and_342_tmp);
  COMP_LOOP_tmp_and_29_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm AND (NOT and_342_tmp);
  COMP_LOOP_tmp_and_30_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm AND (NOT and_342_tmp);
  COMP_LOOP_tmp_and_31_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm AND (NOT and_342_tmp);
  COMP_LOOP_tmp_and_32_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm AND (NOT and_342_tmp);
  COMP_LOOP_tmp_and_33_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm AND (NOT and_342_tmp);
  COMP_LOOP_tmp_and_34_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm AND (NOT and_342_tmp);
  COMP_LOOP_tmp_and_35_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm AND (NOT and_342_tmp);
  COMP_LOOP_tmp_and_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_14_cse AND and_dcpl_198;
  COMP_LOOP_tmp_and_17_nl <= CONV_SL_1_1(COMP_LOOP_13_tmp_mul_idiv_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND and_dcpl_198;
  COMP_LOOP_tmp_and_18_nl <= CONV_SL_1_1(COMP_LOOP_13_tmp_mul_idiv_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND and_dcpl_198;
  mux_2515_nl <= MUX_s_1_2_2(mux_tmp_2392, mux_559_cse, and_674_cse);
  mux_2516_nl <= MUX_s_1_2_2(mux_2515_nl, mux_559_cse, fsm_output(3));
  mux_2514_nl <= MUX_s_1_2_2(mux_tmp_2392, mux_559_cse, or_2259_cse_1);
  mux_2517_nl <= MUX_s_1_2_2(mux_2516_nl, mux_2514_nl, fsm_output(0));
  mux_2518_nl <= MUX_s_1_2_2(mux_2517_nl, and_733_cse, or_2589_cse);
  mux_2519_nl <= MUX_s_1_2_2(mux_tmp_2392, and_dcpl_57, or_2612_cse);
  mux_2520_nl <= MUX_s_1_2_2(mux_tmp_2392, mux_2519_nl, fsm_output(4));
  and_357_nl <= ((fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(6)))
      AND CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11"));
  mux_2528_nl <= MUX_s_1_2_2(mux_228_cse, nor_tmp_47, or_432_cse);
  mux_2529_nl <= MUX_s_1_2_2(mux_228_cse, mux_2528_nl, fsm_output(3));
  mux_2527_nl <= MUX_s_1_2_2(mux_228_cse, nor_tmp_47, fsm_output(3));
  mux_2530_nl <= MUX_s_1_2_2(mux_2529_nl, mux_2527_nl, fsm_output(0));
  mux_2531_nl <= MUX_s_1_2_2(mux_2530_nl, nor_tmp_47, fsm_output(4));
  mux_2526_nl <= MUX_s_1_2_2(nor_tmp_489, (fsm_output(7)), fsm_output(4));
  mux_2532_nl <= MUX_s_1_2_2(mux_2531_nl, mux_2526_nl, fsm_output(5));
  COMP_LOOP_tmp_and_7_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_12_itm AND (NOT nor_1796_tmp);
  COMP_LOOP_tmp_and_8_nl <= COMP_LOOP_tmp_or_29_cse AND (NOT nor_1796_tmp);
  COMP_LOOP_tmp_and_9_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm AND (NOT nor_1796_tmp);
  COMP_LOOP_tmp_and_10_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm AND (NOT nor_1796_tmp);
  COMP_LOOP_tmp_and_11_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm AND (NOT nor_1796_tmp);
  COMP_LOOP_tmp_and_12_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm AND (NOT nor_1796_tmp);
  mux_2540_nl <= MUX_s_1_2_2(or_2732_cse, or_2729_cse, fsm_output(3));
  mux_2541_nl <= MUX_s_1_2_2(or_2621_cse, mux_2540_nl, fsm_output(0));
  nor_568_nl <= NOT((fsm_output(4)) OR mux_2541_nl);
  mux_2539_nl <= MUX_s_1_2_2(and_tmp_28, nor_tmp_47, fsm_output(4));
  mux_2542_nl <= MUX_s_1_2_2(nor_568_nl, mux_2539_nl, fsm_output(5));
  mux_2544_nl <= MUX_s_1_2_2(mux_tmp_439, nor_tmp_115, and_831_cse);
  mux_2543_nl <= MUX_s_1_2_2(mux_tmp_439, nor_tmp_115, and_570_cse);
  mux_2545_nl <= MUX_s_1_2_2(mux_2544_nl, mux_2543_nl, fsm_output(0));
  mux_2546_nl <= MUX_s_1_2_2(mux_2545_nl, nor_tmp_115, fsm_output(4));
  and_352_nl <= ((fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(7)))
      AND (fsm_output(8));
  COMP_LOOP_tmp_and_2_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_12_itm AND and_dcpl_202;
  COMP_LOOP_tmp_and_3_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm AND and_dcpl_202;
  COMP_LOOP_tmp_and_4_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm AND and_dcpl_202;
  COMP_LOOP_tmp_and_5_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm AND and_dcpl_202;
  COMP_LOOP_tmp_and_6_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm AND and_dcpl_202;
  mux_2551_nl <= MUX_s_1_2_2(mux_559_cse, mux_tmp_538, fsm_output(3));
  mux_560_nl <= MUX_s_1_2_2(mux_559_cse, mux_tmp_439, and_674_cse);
  mux_561_nl <= MUX_s_1_2_2(mux_560_nl, mux_tmp_538, fsm_output(3));
  mux_2552_nl <= MUX_s_1_2_2(mux_2551_nl, mux_561_nl, fsm_output(0));
  mux_2553_nl <= MUX_s_1_2_2(mux_2552_nl, nor_tmp_115, or_2589_cse);
  mux_2555_nl <= MUX_s_1_2_2(mux_464_cse, and_733_cse, or_2626_cse);
  mux_2556_nl <= MUX_s_1_2_2(mux_2555_nl, and_733_cse, fsm_output(4));
  or_2625_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"));
  mux_2554_nl <= MUX_s_1_2_2(and_655_cse, nor_tmp_115, or_2625_nl);
  COMP_LOOP_mux_358_nl <= MUX_v_11_2_2(('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))), STAGE_LOOP_lshift_psp_sva, and_dcpl_356);
  COMP_LOOP_COMP_LOOP_nand_1_nl <= NOT(and_dcpl_356 AND (NOT(CONV_SL_1_1(fsm_output(8
      DOWNTO 6)=STD_LOGIC_VECTOR'("000")) AND nor_1624_cse AND CONV_SL_1_1(fsm_output(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("10")) AND and_dcpl_45)));
  COMP_LOOP_mux_359_nl <= MUX_v_10_2_2((COMP_LOOP_k_10_4_sva_5_0 & STD_LOGIC_VECTOR'(
      "0001")), VEC_LOOP_j_10_0_sva_9_0, and_dcpl_356);
  acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_358_nl & COMP_LOOP_COMP_LOOP_nand_1_nl)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_359_nl & '1'), 11), 12),
      12));
  z_out_2 <= acc_nl(11 DOWNTO 1);
  COMP_LOOP_mux1h_710_nl <= MUX1HOT_v_54_15_2((COMP_LOOP_tmp_mux1h_12_itm(63 DOWNTO
      10)), (COMP_LOOP_tmp_mux1h_itm(63 DOWNTO 10)), (COMP_LOOP_tmp_mux1h_1_itm(63
      DOWNTO 10)), (COMP_LOOP_tmp_mux1h_2_itm(63 DOWNTO 10)), (COMP_LOOP_tmp_mux1h_3_itm(63
      DOWNTO 10)), (COMP_LOOP_tmp_mux1h_4_itm(63 DOWNTO 10)), (COMP_LOOP_tmp_mux1h_5_itm(63
      DOWNTO 10)), (COMP_LOOP_tmp_mux1h_6_itm(63 DOWNTO 10)), (COMP_LOOP_tmp_mux_itm(63
      DOWNTO 10)), (COMP_LOOP_tmp_mux1h_7_itm(63 DOWNTO 10)), (COMP_LOOP_tmp_mux1h_8_itm(63
      DOWNTO 10)), (COMP_LOOP_tmp_mux1h_9_itm(63 DOWNTO 10)), (tmp_36_sva_1(63 DOWNTO
      10)), (tmp_36_sva_2(63 DOWNTO 10)), (tmp_33_sva_1(63 DOWNTO 10)), STD_LOGIC_VECTOR'(
      and_dcpl_360 & and_dcpl_367 & and_dcpl_374 & and_dcpl_378 & and_dcpl_384 &
      and_dcpl_386 & and_dcpl_390 & and_dcpl_391 & and_dcpl_395 & and_dcpl_396 &
      and_dcpl_400 & and_dcpl_401 & and_dcpl_405 & and_dcpl_406 & and_dcpl_409));
  COMP_LOOP_and_260_nl <= MUX_v_54_2_2(STD_LOGIC_VECTOR'("000000000000000000000000000000000000000000000000000000"),
      COMP_LOOP_mux1h_710_nl, COMP_LOOP_nor_itm);
  COMP_LOOP_mux1h_711_nl <= MUX1HOT_s_1_17_2((COMP_LOOP_tmp_mux1h_12_itm(9)), (COMP_LOOP_tmp_mux1h_itm(9)),
      (COMP_LOOP_tmp_mux1h_1_itm(9)), (COMP_LOOP_tmp_mux1h_2_itm(9)), (COMP_LOOP_tmp_mux1h_3_itm(9)),
      (COMP_LOOP_tmp_mux1h_4_itm(9)), (COMP_LOOP_tmp_mux1h_5_itm(9)), (COMP_LOOP_tmp_mux1h_6_itm(9)),
      (COMP_LOOP_tmp_mux_itm(9)), (COMP_LOOP_tmp_mux1h_7_itm(9)), (COMP_LOOP_tmp_mux1h_8_itm(9)),
      (COMP_LOOP_tmp_mux1h_9_itm(9)), (tmp_36_sva_1(9)), (tmp_36_sva_2(9)), (tmp_33_sva_1(9)),
      (z_out_1(9)), (COMP_LOOP_2_tmp_lshift_ncse_sva(9)), STD_LOGIC_VECTOR'( and_dcpl_360
      & and_dcpl_367 & and_dcpl_374 & and_dcpl_378 & and_dcpl_384 & and_dcpl_386
      & and_dcpl_390 & and_dcpl_391 & and_dcpl_395 & and_dcpl_396 & and_dcpl_400
      & and_dcpl_401 & and_dcpl_405 & and_dcpl_406 & and_dcpl_409 & and_dcpl_411
      & COMP_LOOP_or_40_itm));
  COMP_LOOP_and_261_nl <= COMP_LOOP_mux1h_711_nl AND COMP_LOOP_nor_621_itm;
  COMP_LOOP_mux1h_712_nl <= MUX1HOT_s_1_18_2((COMP_LOOP_tmp_mux1h_12_itm(8)), (COMP_LOOP_tmp_mux1h_itm(8)),
      (COMP_LOOP_tmp_mux1h_1_itm(8)), (COMP_LOOP_tmp_mux1h_2_itm(8)), (COMP_LOOP_tmp_mux1h_3_itm(8)),
      (COMP_LOOP_tmp_mux1h_4_itm(8)), (COMP_LOOP_tmp_mux1h_5_itm(8)), (COMP_LOOP_tmp_mux1h_6_itm(8)),
      (COMP_LOOP_tmp_mux_itm(8)), (COMP_LOOP_tmp_mux1h_7_itm(8)), (COMP_LOOP_tmp_mux1h_8_itm(8)),
      (COMP_LOOP_tmp_mux1h_9_itm(8)), (tmp_36_sva_1(8)), (tmp_36_sva_2(8)), (tmp_33_sva_1(8)),
      (z_out_1(8)), (COMP_LOOP_2_tmp_lshift_ncse_sva(8)), (COMP_LOOP_3_tmp_lshift_ncse_sva(8)),
      STD_LOGIC_VECTOR'( and_dcpl_360 & and_dcpl_367 & and_dcpl_374 & and_dcpl_378
      & and_dcpl_384 & and_dcpl_386 & and_dcpl_390 & and_dcpl_391 & and_dcpl_395
      & and_dcpl_396 & and_dcpl_400 & and_dcpl_401 & and_dcpl_405 & and_dcpl_406
      & and_dcpl_409 & COMP_LOOP_or_41_itm & COMP_LOOP_or_40_itm & COMP_LOOP_or_43_itm));
  COMP_LOOP_and_262_nl <= COMP_LOOP_mux1h_712_nl AND COMP_LOOP_nor_622_itm;
  COMP_LOOP_mux1h_713_nl <= MUX1HOT_v_8_20_2((COMP_LOOP_tmp_mux1h_12_itm(7 DOWNTO
      0)), (COMP_LOOP_tmp_mux1h_itm(7 DOWNTO 0)), (COMP_LOOP_tmp_mux1h_1_itm(7 DOWNTO
      0)), (COMP_LOOP_tmp_mux1h_2_itm(7 DOWNTO 0)), (COMP_LOOP_tmp_mux1h_3_itm(7
      DOWNTO 0)), (COMP_LOOP_tmp_mux1h_4_itm(7 DOWNTO 0)), (COMP_LOOP_tmp_mux1h_5_itm(7
      DOWNTO 0)), (COMP_LOOP_tmp_mux1h_6_itm(7 DOWNTO 0)), (COMP_LOOP_tmp_mux_itm(7
      DOWNTO 0)), (COMP_LOOP_tmp_mux1h_7_itm(7 DOWNTO 0)), (COMP_LOOP_tmp_mux1h_8_itm(7
      DOWNTO 0)), (COMP_LOOP_tmp_mux1h_9_itm(7 DOWNTO 0)), (tmp_36_sva_1(7 DOWNTO
      0)), (tmp_36_sva_2(7 DOWNTO 0)), (tmp_33_sva_1(7 DOWNTO 0)), (z_out_1(7 DOWNTO
      0)), ('0' & COMP_LOOP_9_tmp_lshift_itm), (COMP_LOOP_2_tmp_lshift_ncse_sva(7
      DOWNTO 0)), (COMP_LOOP_3_tmp_lshift_ncse_sva(7 DOWNTO 0)), COMP_LOOP_13_tmp_mul_idiv_sva,
      STD_LOGIC_VECTOR'( and_dcpl_360 & and_dcpl_367 & and_dcpl_374 & and_dcpl_378
      & and_dcpl_384 & and_dcpl_386 & and_dcpl_390 & and_dcpl_391 & and_dcpl_395
      & and_dcpl_396 & and_dcpl_400 & and_dcpl_401 & and_dcpl_405 & and_dcpl_406
      & and_dcpl_409 & COMP_LOOP_or_41_itm & and_dcpl_413 & COMP_LOOP_or_40_itm &
      COMP_LOOP_or_43_itm & COMP_LOOP_or_47_itm));
  COMP_LOOP_COMP_LOOP_and_983_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(63)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_984_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(62)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_985_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(61)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_986_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(60)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_987_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(59)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_988_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(58)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_989_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(57)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_990_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(56)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_991_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(55)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_992_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(54)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_993_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(53)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_994_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(52)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_995_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(51)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_996_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(50)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_997_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(49)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_998_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(48)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_999_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(47)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1000_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(46)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1001_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(45)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1002_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(44)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1003_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(43)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1004_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(42)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1005_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(41)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1006_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(40)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1007_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(39)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1008_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(38)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1009_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(37)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1010_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(36)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1011_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(35)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1012_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(34)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1013_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(33)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1014_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(32)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1015_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(31)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1016_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(30)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1017_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(29)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1018_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(28)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1019_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(27)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1020_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(26)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1021_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(25)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1022_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(24)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1023_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(23)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1024_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(22)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1025_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(21)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1026_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(20)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1027_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(19)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1028_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(18)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1029_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(17)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1030_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(16)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1031_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(15)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1032_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(14)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1033_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(13)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1034_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(12)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1035_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(11)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_and_1036_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(10)) AND
      COMP_LOOP_nor_itm;
  COMP_LOOP_COMP_LOOP_mux_8_nl <= MUX_s_1_2_2((COMP_LOOP_1_modulo_cmp_return_rsc_z(9)),
      (COMP_LOOP_k_10_4_sva_5_0(5)), COMP_LOOP_or_52_itm);
  COMP_LOOP_and_263_nl <= COMP_LOOP_COMP_LOOP_mux_8_nl AND COMP_LOOP_nor_621_itm;
  COMP_LOOP_mux1h_714_nl <= MUX1HOT_s_1_3_2((COMP_LOOP_1_modulo_cmp_return_rsc_z(8)),
      (COMP_LOOP_k_10_4_sva_5_0(4)), (COMP_LOOP_k_10_4_sva_5_0(5)), STD_LOGIC_VECTOR'(
      COMP_LOOP_or_17_ssc & COMP_LOOP_or_52_itm & COMP_LOOP_or_54_itm));
  COMP_LOOP_and_264_nl <= COMP_LOOP_mux1h_714_nl AND COMP_LOOP_nor_622_itm;
  COMP_LOOP_mux1h_715_nl <= MUX1HOT_v_4_5_2((COMP_LOOP_1_modulo_cmp_return_rsc_z(7
      DOWNTO 4)), (COMP_LOOP_k_10_4_sva_5_0(3 DOWNTO 0)), ('0' & (COMP_LOOP_k_10_4_sva_5_0(5
      DOWNTO 3))), (COMP_LOOP_k_10_4_sva_5_0(4 DOWNTO 1)), (COMP_LOOP_k_10_4_sva_5_0(5
      DOWNTO 2)), STD_LOGIC_VECTOR'( COMP_LOOP_or_17_ssc & COMP_LOOP_or_52_itm &
      and_dcpl_413 & COMP_LOOP_or_54_itm & COMP_LOOP_or_47_itm));
  COMP_LOOP_mux1h_716_nl <= MUX1HOT_s_1_4_2((COMP_LOOP_1_modulo_cmp_return_rsc_z(3)),
      (COMP_LOOP_k_10_4_sva_5_0(2)), (COMP_LOOP_k_10_4_sva_5_0(0)), (COMP_LOOP_k_10_4_sva_5_0(1)),
      STD_LOGIC_VECTOR'( COMP_LOOP_or_17_ssc & and_dcpl_413 & COMP_LOOP_or_54_itm
      & COMP_LOOP_or_47_itm));
  COMP_LOOP_or_61_nl <= (COMP_LOOP_mux1h_716_nl AND (NOT(and_dcpl_411 OR and_dcpl_416
      OR and_dcpl_417 OR and_dcpl_418))) OR and_dcpl_419 OR and_dcpl_421 OR and_dcpl_422
      OR and_dcpl_425;
  COMP_LOOP_mux1h_717_nl <= MUX1HOT_s_1_3_2((COMP_LOOP_1_modulo_cmp_return_rsc_z(2)),
      (COMP_LOOP_k_10_4_sva_5_0(1)), (COMP_LOOP_k_10_4_sva_5_0(0)), STD_LOGIC_VECTOR'(
      COMP_LOOP_or_17_ssc & and_dcpl_413 & COMP_LOOP_or_47_itm));
  COMP_LOOP_or_62_nl <= (COMP_LOOP_mux1h_717_nl AND (NOT(and_dcpl_411 OR and_dcpl_416
      OR and_dcpl_419 OR and_dcpl_421 OR and_dcpl_426 OR and_dcpl_427))) OR and_dcpl_417
      OR and_dcpl_418 OR and_dcpl_422 OR and_dcpl_425 OR and_dcpl_428 OR and_dcpl_429;
  COMP_LOOP_mux_360_nl <= MUX_s_1_2_2((COMP_LOOP_1_modulo_cmp_return_rsc_z(1)), (COMP_LOOP_k_10_4_sva_5_0(0)),
      and_dcpl_413);
  COMP_LOOP_COMP_LOOP_or_2_nl <= (COMP_LOOP_mux_360_nl AND (NOT(and_dcpl_411 OR and_dcpl_417
      OR and_dcpl_419 OR and_dcpl_422 OR and_dcpl_426 OR and_dcpl_428 OR and_dcpl_431)))
      OR and_dcpl_416 OR and_dcpl_418 OR and_dcpl_421 OR and_dcpl_425 OR and_dcpl_427
      OR and_dcpl_429 OR and_dcpl_430;
  COMP_LOOP_COMP_LOOP_or_3_nl <= (COMP_LOOP_1_modulo_cmp_return_rsc_z(0)) OR and_dcpl_411
      OR and_dcpl_416 OR and_dcpl_417 OR and_dcpl_418 OR and_dcpl_419 OR and_dcpl_421
      OR and_dcpl_422 OR and_dcpl_425 OR and_dcpl_426 OR and_dcpl_427 OR and_dcpl_428
      OR and_dcpl_429 OR and_dcpl_430 OR and_dcpl_431 OR and_dcpl_413;
  z_out_3 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( UNSIGNED(COMP_LOOP_and_260_nl
      & COMP_LOOP_and_261_nl & COMP_LOOP_and_262_nl & COMP_LOOP_mux1h_713_nl) * UNSIGNED(COMP_LOOP_COMP_LOOP_and_983_nl
      & COMP_LOOP_COMP_LOOP_and_984_nl & COMP_LOOP_COMP_LOOP_and_985_nl & COMP_LOOP_COMP_LOOP_and_986_nl
      & COMP_LOOP_COMP_LOOP_and_987_nl & COMP_LOOP_COMP_LOOP_and_988_nl & COMP_LOOP_COMP_LOOP_and_989_nl
      & COMP_LOOP_COMP_LOOP_and_990_nl & COMP_LOOP_COMP_LOOP_and_991_nl & COMP_LOOP_COMP_LOOP_and_992_nl
      & COMP_LOOP_COMP_LOOP_and_993_nl & COMP_LOOP_COMP_LOOP_and_994_nl & COMP_LOOP_COMP_LOOP_and_995_nl
      & COMP_LOOP_COMP_LOOP_and_996_nl & COMP_LOOP_COMP_LOOP_and_997_nl & COMP_LOOP_COMP_LOOP_and_998_nl
      & COMP_LOOP_COMP_LOOP_and_999_nl & COMP_LOOP_COMP_LOOP_and_1000_nl & COMP_LOOP_COMP_LOOP_and_1001_nl
      & COMP_LOOP_COMP_LOOP_and_1002_nl & COMP_LOOP_COMP_LOOP_and_1003_nl & COMP_LOOP_COMP_LOOP_and_1004_nl
      & COMP_LOOP_COMP_LOOP_and_1005_nl & COMP_LOOP_COMP_LOOP_and_1006_nl & COMP_LOOP_COMP_LOOP_and_1007_nl
      & COMP_LOOP_COMP_LOOP_and_1008_nl & COMP_LOOP_COMP_LOOP_and_1009_nl & COMP_LOOP_COMP_LOOP_and_1010_nl
      & COMP_LOOP_COMP_LOOP_and_1011_nl & COMP_LOOP_COMP_LOOP_and_1012_nl & COMP_LOOP_COMP_LOOP_and_1013_nl
      & COMP_LOOP_COMP_LOOP_and_1014_nl & COMP_LOOP_COMP_LOOP_and_1015_nl & COMP_LOOP_COMP_LOOP_and_1016_nl
      & COMP_LOOP_COMP_LOOP_and_1017_nl & COMP_LOOP_COMP_LOOP_and_1018_nl & COMP_LOOP_COMP_LOOP_and_1019_nl
      & COMP_LOOP_COMP_LOOP_and_1020_nl & COMP_LOOP_COMP_LOOP_and_1021_nl & COMP_LOOP_COMP_LOOP_and_1022_nl
      & COMP_LOOP_COMP_LOOP_and_1023_nl & COMP_LOOP_COMP_LOOP_and_1024_nl & COMP_LOOP_COMP_LOOP_and_1025_nl
      & COMP_LOOP_COMP_LOOP_and_1026_nl & COMP_LOOP_COMP_LOOP_and_1027_nl & COMP_LOOP_COMP_LOOP_and_1028_nl
      & COMP_LOOP_COMP_LOOP_and_1029_nl & COMP_LOOP_COMP_LOOP_and_1030_nl & COMP_LOOP_COMP_LOOP_and_1031_nl
      & COMP_LOOP_COMP_LOOP_and_1032_nl & COMP_LOOP_COMP_LOOP_and_1033_nl & COMP_LOOP_COMP_LOOP_and_1034_nl
      & COMP_LOOP_COMP_LOOP_and_1035_nl & COMP_LOOP_COMP_LOOP_and_1036_nl & COMP_LOOP_and_263_nl
      & COMP_LOOP_and_264_nl & COMP_LOOP_mux1h_715_nl & COMP_LOOP_or_61_nl & COMP_LOOP_or_62_nl
      & COMP_LOOP_COMP_LOOP_or_2_nl & COMP_LOOP_COMP_LOOP_or_3_nl)), 64));
  STAGE_LOOP_mux_4_nl <= MUX_v_4_2_2(STAGE_LOOP_i_3_0_sva, (NOT STAGE_LOOP_i_3_0_sva),
      and_dcpl_447);
  z_out_4 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_LOOP_mux_4_nl) + UNSIGNED('1'
      & (NOT and_dcpl_447) & STD_LOGIC_VECTOR'( "11")), 4));
  COMP_LOOP_mux_361_cse <= MUX_v_64_2_2(z_out_7, COMP_LOOP_10_acc_8_itm, COMP_LOOP_or_18_itm);
  COMP_LOOP_mux1h_718_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_nor_itm, COMP_LOOP_COMP_LOOP_nor_5_itm,
      COMP_LOOP_COMP_LOOP_nor_9_itm, COMP_LOOP_COMP_LOOP_nor_13_itm, COMP_LOOP_COMP_LOOP_nor_17_itm,
      COMP_LOOP_COMP_LOOP_nor_21_itm, COMP_LOOP_COMP_LOOP_nor_25_itm, COMP_LOOP_COMP_LOOP_nor_29_itm,
      COMP_LOOP_COMP_LOOP_nor_33_itm, COMP_LOOP_COMP_LOOP_nor_37_itm, COMP_LOOP_COMP_LOOP_nor_41_itm,
      COMP_LOOP_COMP_LOOP_nor_45_itm, COMP_LOOP_COMP_LOOP_nor_49_itm, COMP_LOOP_COMP_LOOP_nor_53_itm,
      COMP_LOOP_COMP_LOOP_nor_57_itm, COMP_LOOP_COMP_LOOP_nor_61_itm, STD_LOGIC_VECTOR'(
      and_dcpl_571 & and_dcpl_577 & and_1025_cse & and_1028_cse & and_dcpl_589 &
      and_1037_cse & and_1040_cse & and_1044_cse & and_1046_cse & and_1051_cse &
      and_1052_cse & and_1055_cse & and_1056_cse & and_1060_cse & and_1061_cse &
      and_1064_cse));
  COMP_LOOP_COMP_LOOP_and_1037_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(0)) AND COMP_LOOP_nor_51_itm;
  COMP_LOOP_COMP_LOOP_and_1038_nl <= (COMP_LOOP_acc_10_cse_10_1_3_sva(0)) AND COMP_LOOP_nor_91_itm;
  COMP_LOOP_COMP_LOOP_and_1039_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(0)) AND COMP_LOOP_nor_131_itm;
  COMP_LOOP_COMP_LOOP_and_1040_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(0)) AND COMP_LOOP_nor_171_itm;
  COMP_LOOP_COMP_LOOP_and_1041_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(0)) AND COMP_LOOP_nor_211_itm;
  COMP_LOOP_COMP_LOOP_and_1042_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) AND COMP_LOOP_nor_251_itm;
  COMP_LOOP_COMP_LOOP_and_1043_nl <= (COMP_LOOP_acc_10_cse_10_1_8_sva(0)) AND COMP_LOOP_nor_291_itm;
  COMP_LOOP_COMP_LOOP_and_1044_nl <= (COMP_LOOP_acc_10_cse_10_1_9_sva(0)) AND COMP_LOOP_nor_331_itm;
  COMP_LOOP_COMP_LOOP_and_1045_nl <= (COMP_LOOP_acc_10_cse_10_1_10_sva(0)) AND COMP_LOOP_nor_371_itm;
  COMP_LOOP_COMP_LOOP_and_1046_nl <= (COMP_LOOP_acc_10_cse_10_1_11_sva(0)) AND COMP_LOOP_nor_411_itm;
  COMP_LOOP_COMP_LOOP_and_1047_nl <= (COMP_LOOP_acc_10_cse_10_1_12_sva(0)) AND COMP_LOOP_nor_451_itm;
  COMP_LOOP_COMP_LOOP_and_1048_nl <= (COMP_LOOP_acc_10_cse_10_1_13_sva(0)) AND COMP_LOOP_nor_491_itm;
  COMP_LOOP_COMP_LOOP_and_1049_nl <= (COMP_LOOP_acc_10_cse_10_1_14_sva(0)) AND COMP_LOOP_nor_531_itm;
  COMP_LOOP_COMP_LOOP_and_1050_nl <= (COMP_LOOP_acc_10_cse_10_1_15_sva(0)) AND COMP_LOOP_nor_571_itm;
  COMP_LOOP_COMP_LOOP_and_1051_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(0)) AND COMP_LOOP_nor_611_itm;
  COMP_LOOP_mux1h_719_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_244_itm, COMP_LOOP_COMP_LOOP_and_1037_nl,
      COMP_LOOP_COMP_LOOP_and_1038_nl, COMP_LOOP_COMP_LOOP_and_1039_nl, COMP_LOOP_COMP_LOOP_and_1040_nl,
      COMP_LOOP_COMP_LOOP_and_1041_nl, COMP_LOOP_COMP_LOOP_and_1042_nl, COMP_LOOP_COMP_LOOP_and_1043_nl,
      COMP_LOOP_COMP_LOOP_and_1044_nl, COMP_LOOP_COMP_LOOP_and_1045_nl, COMP_LOOP_COMP_LOOP_and_1046_nl,
      COMP_LOOP_COMP_LOOP_and_1047_nl, COMP_LOOP_COMP_LOOP_and_1048_nl, COMP_LOOP_COMP_LOOP_and_1049_nl,
      COMP_LOOP_COMP_LOOP_and_1050_nl, COMP_LOOP_COMP_LOOP_and_1051_nl, STD_LOGIC_VECTOR'(
      and_dcpl_571 & and_dcpl_577 & and_1025_cse & and_1028_cse & and_dcpl_589 &
      and_1037_cse & and_1040_cse & and_1044_cse & and_1046_cse & and_1051_cse &
      and_1052_cse & and_1055_cse & and_1056_cse & and_1060_cse & and_1061_cse &
      and_1064_cse));
  COMP_LOOP_COMP_LOOP_and_1052_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(1)) AND COMP_LOOP_nor_52_itm;
  COMP_LOOP_COMP_LOOP_and_1053_nl <= (COMP_LOOP_acc_10_cse_10_1_3_sva(1)) AND COMP_LOOP_nor_92_itm;
  COMP_LOOP_COMP_LOOP_and_1054_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(1)) AND COMP_LOOP_nor_132_itm;
  COMP_LOOP_COMP_LOOP_and_1055_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(1)) AND COMP_LOOP_nor_172_itm;
  COMP_LOOP_COMP_LOOP_and_1056_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(1)) AND COMP_LOOP_nor_212_itm;
  COMP_LOOP_COMP_LOOP_and_1057_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(1)) AND COMP_LOOP_nor_252_itm;
  COMP_LOOP_COMP_LOOP_and_1058_nl <= (COMP_LOOP_acc_10_cse_10_1_8_sva(1)) AND COMP_LOOP_nor_292_itm;
  COMP_LOOP_COMP_LOOP_and_1059_nl <= (COMP_LOOP_acc_10_cse_10_1_9_sva(1)) AND COMP_LOOP_nor_332_itm;
  COMP_LOOP_COMP_LOOP_and_1060_nl <= (COMP_LOOP_acc_10_cse_10_1_10_sva(1)) AND COMP_LOOP_nor_372_itm;
  COMP_LOOP_COMP_LOOP_and_1061_nl <= (COMP_LOOP_acc_10_cse_10_1_11_sva(1)) AND COMP_LOOP_nor_412_itm;
  COMP_LOOP_COMP_LOOP_and_1062_nl <= (COMP_LOOP_acc_10_cse_10_1_12_sva(1)) AND COMP_LOOP_nor_452_itm;
  COMP_LOOP_COMP_LOOP_and_1063_nl <= (COMP_LOOP_acc_10_cse_10_1_13_sva(1)) AND COMP_LOOP_nor_492_itm;
  COMP_LOOP_COMP_LOOP_and_1064_nl <= (COMP_LOOP_acc_10_cse_10_1_14_sva(1)) AND COMP_LOOP_nor_532_itm;
  COMP_LOOP_COMP_LOOP_and_1065_nl <= (COMP_LOOP_acc_10_cse_10_1_15_sva(1)) AND COMP_LOOP_nor_572_itm;
  COMP_LOOP_COMP_LOOP_and_1066_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(1)) AND COMP_LOOP_nor_612_itm;
  COMP_LOOP_mux1h_720_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_62_itm, COMP_LOOP_COMP_LOOP_and_1052_nl,
      COMP_LOOP_COMP_LOOP_and_1053_nl, COMP_LOOP_COMP_LOOP_and_1054_nl, COMP_LOOP_COMP_LOOP_and_1055_nl,
      COMP_LOOP_COMP_LOOP_and_1056_nl, COMP_LOOP_COMP_LOOP_and_1057_nl, COMP_LOOP_COMP_LOOP_and_1058_nl,
      COMP_LOOP_COMP_LOOP_and_1059_nl, COMP_LOOP_COMP_LOOP_and_1060_nl, COMP_LOOP_COMP_LOOP_and_1061_nl,
      COMP_LOOP_COMP_LOOP_and_1062_nl, COMP_LOOP_COMP_LOOP_and_1063_nl, COMP_LOOP_COMP_LOOP_and_1064_nl,
      COMP_LOOP_COMP_LOOP_and_1065_nl, COMP_LOOP_COMP_LOOP_and_1066_nl, STD_LOGIC_VECTOR'(
      and_dcpl_571 & and_dcpl_577 & and_1025_cse & and_1028_cse & and_dcpl_589 &
      and_1037_cse & and_1040_cse & and_1044_cse & and_1046_cse & and_1051_cse &
      and_1052_cse & and_1055_cse & and_1056_cse & and_1060_cse & and_1061_cse &
      and_1064_cse));
  COMP_LOOP_mux1h_721_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_185_itm, COMP_LOOP_COMP_LOOP_and_77_itm,
      COMP_LOOP_COMP_LOOP_and_137_itm, COMP_LOOP_COMP_LOOP_and_197_itm, COMP_LOOP_COMP_LOOP_and_257_itm,
      COMP_LOOP_COMP_LOOP_and_317_itm, COMP_LOOP_COMP_LOOP_and_377_itm, COMP_LOOP_COMP_LOOP_and_437_itm,
      COMP_LOOP_COMP_LOOP_and_497_itm, COMP_LOOP_COMP_LOOP_and_557_itm, COMP_LOOP_COMP_LOOP_and_617_itm,
      COMP_LOOP_COMP_LOOP_and_677_itm, COMP_LOOP_COMP_LOOP_and_737_itm, COMP_LOOP_COMP_LOOP_and_797_itm,
      COMP_LOOP_COMP_LOOP_and_857_itm, COMP_LOOP_COMP_LOOP_and_917_itm, STD_LOGIC_VECTOR'(
      and_dcpl_571 & and_dcpl_577 & and_1025_cse & and_1028_cse & and_dcpl_589 &
      and_1037_cse & and_1040_cse & and_1044_cse & and_1046_cse & and_1051_cse &
      and_1052_cse & and_1055_cse & and_1056_cse & and_1060_cse & and_1061_cse &
      and_1064_cse));
  COMP_LOOP_COMP_LOOP_and_1067_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(2)) AND COMP_LOOP_nor_54_itm;
  COMP_LOOP_COMP_LOOP_and_1068_nl <= (COMP_LOOP_acc_10_cse_10_1_3_sva(2)) AND COMP_LOOP_nor_94_itm;
  COMP_LOOP_COMP_LOOP_and_1069_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(2)) AND COMP_LOOP_nor_134_itm;
  COMP_LOOP_COMP_LOOP_and_1070_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(2)) AND COMP_LOOP_nor_174_itm;
  COMP_LOOP_COMP_LOOP_and_1071_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(2)) AND COMP_LOOP_nor_214_itm;
  COMP_LOOP_COMP_LOOP_and_1072_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(2)) AND COMP_LOOP_nor_254_itm;
  COMP_LOOP_COMP_LOOP_and_1073_nl <= (COMP_LOOP_acc_10_cse_10_1_8_sva(2)) AND COMP_LOOP_nor_294_itm;
  COMP_LOOP_COMP_LOOP_and_1074_nl <= (COMP_LOOP_acc_10_cse_10_1_9_sva(2)) AND COMP_LOOP_nor_334_itm;
  COMP_LOOP_COMP_LOOP_and_1075_nl <= (COMP_LOOP_acc_10_cse_10_1_10_sva(2)) AND COMP_LOOP_nor_374_itm;
  COMP_LOOP_COMP_LOOP_and_1076_nl <= (COMP_LOOP_acc_10_cse_10_1_11_sva(2)) AND COMP_LOOP_nor_414_itm;
  COMP_LOOP_COMP_LOOP_and_1077_nl <= (COMP_LOOP_acc_10_cse_10_1_12_sva(2)) AND COMP_LOOP_nor_454_itm;
  COMP_LOOP_COMP_LOOP_and_1078_nl <= (COMP_LOOP_acc_10_cse_10_1_13_sva(2)) AND COMP_LOOP_nor_494_itm;
  COMP_LOOP_COMP_LOOP_and_1079_nl <= (COMP_LOOP_acc_10_cse_10_1_14_sva(2)) AND COMP_LOOP_nor_534_itm;
  COMP_LOOP_COMP_LOOP_and_1080_nl <= (COMP_LOOP_acc_10_cse_10_1_15_sva(2)) AND COMP_LOOP_nor_574_itm;
  COMP_LOOP_COMP_LOOP_and_1081_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(2)) AND COMP_LOOP_nor_614_itm;
  COMP_LOOP_mux1h_722_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_64_itm, COMP_LOOP_COMP_LOOP_and_1067_nl,
      COMP_LOOP_COMP_LOOP_and_1068_nl, COMP_LOOP_COMP_LOOP_and_1069_nl, COMP_LOOP_COMP_LOOP_and_1070_nl,
      COMP_LOOP_COMP_LOOP_and_1071_nl, COMP_LOOP_COMP_LOOP_and_1072_nl, COMP_LOOP_COMP_LOOP_and_1073_nl,
      COMP_LOOP_COMP_LOOP_and_1074_nl, COMP_LOOP_COMP_LOOP_and_1075_nl, COMP_LOOP_COMP_LOOP_and_1076_nl,
      COMP_LOOP_COMP_LOOP_and_1077_nl, COMP_LOOP_COMP_LOOP_and_1078_nl, COMP_LOOP_COMP_LOOP_and_1079_nl,
      COMP_LOOP_COMP_LOOP_and_1080_nl, COMP_LOOP_COMP_LOOP_and_1081_nl, STD_LOGIC_VECTOR'(
      and_dcpl_571 & and_dcpl_577 & and_1025_cse & and_1028_cse & and_dcpl_589 &
      and_1037_cse & and_1040_cse & and_1044_cse & and_1046_cse & and_1051_cse &
      and_1052_cse & and_1055_cse & and_1056_cse & and_1060_cse & and_1061_cse &
      and_1064_cse));
  COMP_LOOP_mux1h_723_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_65_itm, COMP_LOOP_COMP_LOOP_and_79_itm,
      COMP_LOOP_COMP_LOOP_and_139_itm, COMP_LOOP_COMP_LOOP_and_199_itm, COMP_LOOP_COMP_LOOP_and_259_itm,
      COMP_LOOP_COMP_LOOP_and_319_itm, COMP_LOOP_COMP_LOOP_and_379_itm, COMP_LOOP_COMP_LOOP_and_439_itm,
      COMP_LOOP_COMP_LOOP_and_499_itm, COMP_LOOP_COMP_LOOP_and_559_itm, COMP_LOOP_COMP_LOOP_and_619_itm,
      COMP_LOOP_COMP_LOOP_and_679_itm, COMP_LOOP_COMP_LOOP_and_739_itm, COMP_LOOP_COMP_LOOP_and_799_itm,
      COMP_LOOP_COMP_LOOP_and_859_itm, COMP_LOOP_COMP_LOOP_and_919_itm, STD_LOGIC_VECTOR'(
      and_dcpl_571 & and_dcpl_577 & and_1025_cse & and_1028_cse & and_dcpl_589 &
      and_1037_cse & and_1040_cse & and_1044_cse & and_1046_cse & and_1051_cse &
      and_1052_cse & and_1055_cse & and_1056_cse & and_1060_cse & and_1061_cse &
      and_1064_cse));
  COMP_LOOP_mux1h_724_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_66_itm, COMP_LOOP_COMP_LOOP_and_80_itm,
      COMP_LOOP_COMP_LOOP_and_140_itm, COMP_LOOP_COMP_LOOP_and_200_itm, COMP_LOOP_COMP_LOOP_and_260_itm,
      COMP_LOOP_COMP_LOOP_and_320_itm, COMP_LOOP_COMP_LOOP_and_380_itm, COMP_LOOP_COMP_LOOP_and_440_itm,
      COMP_LOOP_COMP_LOOP_and_500_itm, COMP_LOOP_COMP_LOOP_and_560_itm, COMP_LOOP_COMP_LOOP_and_620_itm,
      COMP_LOOP_COMP_LOOP_and_680_itm, COMP_LOOP_COMP_LOOP_and_740_itm, COMP_LOOP_COMP_LOOP_and_800_itm,
      COMP_LOOP_COMP_LOOP_and_860_itm, COMP_LOOP_COMP_LOOP_and_920_itm, STD_LOGIC_VECTOR'(
      and_dcpl_571 & and_dcpl_577 & and_1025_cse & and_1028_cse & and_dcpl_589 &
      and_1037_cse & and_1040_cse & and_1044_cse & and_1046_cse & and_1051_cse &
      and_1052_cse & and_1055_cse & and_1056_cse & and_1060_cse & and_1061_cse &
      and_1064_cse));
  COMP_LOOP_mux1h_725_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_6_itm, COMP_LOOP_COMP_LOOP_and_81_itm,
      COMP_LOOP_COMP_LOOP_and_141_itm, COMP_LOOP_COMP_LOOP_and_201_itm, COMP_LOOP_COMP_LOOP_and_261_itm,
      COMP_LOOP_COMP_LOOP_and_321_itm, COMP_LOOP_COMP_LOOP_and_381_itm, COMP_LOOP_COMP_LOOP_and_441_itm,
      COMP_LOOP_COMP_LOOP_and_501_itm, COMP_LOOP_COMP_LOOP_and_561_itm, COMP_LOOP_COMP_LOOP_and_621_itm,
      COMP_LOOP_COMP_LOOP_and_681_itm, COMP_LOOP_COMP_LOOP_and_741_itm, COMP_LOOP_COMP_LOOP_and_801_itm,
      COMP_LOOP_COMP_LOOP_and_861_itm, COMP_LOOP_COMP_LOOP_and_921_itm, STD_LOGIC_VECTOR'(
      and_dcpl_571 & and_dcpl_577 & and_1025_cse & and_1028_cse & and_dcpl_589 &
      and_1037_cse & and_1040_cse & and_1044_cse & and_1046_cse & and_1051_cse &
      and_1052_cse & and_1055_cse & and_1056_cse & and_1060_cse & and_1061_cse &
      and_1064_cse));
  COMP_LOOP_COMP_LOOP_and_1082_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(3)) AND COMP_LOOP_nor_57_itm;
  COMP_LOOP_COMP_LOOP_and_1083_nl <= (COMP_LOOP_acc_10_cse_10_1_3_sva(3)) AND COMP_LOOP_nor_97_itm;
  COMP_LOOP_COMP_LOOP_and_1084_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(3)) AND COMP_LOOP_nor_137_itm;
  COMP_LOOP_COMP_LOOP_and_1085_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(3)) AND COMP_LOOP_nor_177_itm;
  COMP_LOOP_COMP_LOOP_and_1086_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(3)) AND COMP_LOOP_nor_217_itm;
  COMP_LOOP_COMP_LOOP_and_1087_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(3)) AND COMP_LOOP_nor_257_itm;
  COMP_LOOP_COMP_LOOP_and_1088_nl <= (COMP_LOOP_acc_10_cse_10_1_8_sva(3)) AND COMP_LOOP_nor_297_itm;
  COMP_LOOP_COMP_LOOP_and_1089_nl <= (COMP_LOOP_acc_10_cse_10_1_9_sva(3)) AND COMP_LOOP_nor_337_itm;
  COMP_LOOP_COMP_LOOP_and_1090_nl <= (COMP_LOOP_acc_10_cse_10_1_10_sva(3)) AND COMP_LOOP_nor_377_itm;
  COMP_LOOP_COMP_LOOP_and_1091_nl <= (COMP_LOOP_acc_10_cse_10_1_11_sva(3)) AND COMP_LOOP_nor_417_itm;
  COMP_LOOP_COMP_LOOP_and_1092_nl <= (COMP_LOOP_acc_10_cse_10_1_12_sva(3)) AND COMP_LOOP_nor_457_itm;
  COMP_LOOP_COMP_LOOP_and_1093_nl <= (COMP_LOOP_acc_10_cse_10_1_13_sva(3)) AND COMP_LOOP_nor_497_itm;
  COMP_LOOP_COMP_LOOP_and_1094_nl <= (COMP_LOOP_acc_10_cse_10_1_14_sva(3)) AND COMP_LOOP_nor_537_itm;
  COMP_LOOP_COMP_LOOP_and_1095_nl <= (COMP_LOOP_acc_10_cse_10_1_15_sva(3)) AND COMP_LOOP_nor_577_itm;
  COMP_LOOP_COMP_LOOP_and_1096_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(3)) AND COMP_LOOP_nor_617_itm;
  COMP_LOOP_mux1h_726_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_68_itm, COMP_LOOP_COMP_LOOP_and_1082_nl,
      COMP_LOOP_COMP_LOOP_and_1083_nl, COMP_LOOP_COMP_LOOP_and_1084_nl, COMP_LOOP_COMP_LOOP_and_1085_nl,
      COMP_LOOP_COMP_LOOP_and_1086_nl, COMP_LOOP_COMP_LOOP_and_1087_nl, COMP_LOOP_COMP_LOOP_and_1088_nl,
      COMP_LOOP_COMP_LOOP_and_1089_nl, COMP_LOOP_COMP_LOOP_and_1090_nl, COMP_LOOP_COMP_LOOP_and_1091_nl,
      COMP_LOOP_COMP_LOOP_and_1092_nl, COMP_LOOP_COMP_LOOP_and_1093_nl, COMP_LOOP_COMP_LOOP_and_1094_nl,
      COMP_LOOP_COMP_LOOP_and_1095_nl, COMP_LOOP_COMP_LOOP_and_1096_nl, STD_LOGIC_VECTOR'(
      and_dcpl_571 & and_dcpl_577 & and_1025_cse & and_1028_cse & and_dcpl_589 &
      and_1037_cse & and_1040_cse & and_1044_cse & and_1046_cse & and_1051_cse &
      and_1052_cse & and_1055_cse & and_1056_cse & and_1060_cse & and_1061_cse &
      and_1064_cse));
  COMP_LOOP_mux1h_727_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_69_itm, COMP_LOOP_COMP_LOOP_and_83_itm,
      COMP_LOOP_COMP_LOOP_and_143_itm, COMP_LOOP_COMP_LOOP_and_203_itm, COMP_LOOP_COMP_LOOP_and_263_itm,
      COMP_LOOP_COMP_LOOP_and_323_itm, COMP_LOOP_COMP_LOOP_and_383_itm, COMP_LOOP_COMP_LOOP_and_443_itm,
      COMP_LOOP_COMP_LOOP_and_503_itm, COMP_LOOP_COMP_LOOP_and_563_itm, COMP_LOOP_COMP_LOOP_and_623_itm,
      COMP_LOOP_COMP_LOOP_and_683_itm, COMP_LOOP_COMP_LOOP_and_743_itm, COMP_LOOP_COMP_LOOP_and_803_itm,
      COMP_LOOP_COMP_LOOP_and_863_itm, COMP_LOOP_COMP_LOOP_and_923_itm, STD_LOGIC_VECTOR'(
      and_dcpl_571 & and_dcpl_577 & and_1025_cse & and_1028_cse & and_dcpl_589 &
      and_1037_cse & and_1040_cse & and_1044_cse & and_1046_cse & and_1051_cse &
      and_1052_cse & and_1055_cse & and_1056_cse & and_1060_cse & and_1061_cse &
      and_1064_cse));
  COMP_LOOP_mux1h_728_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_70_itm, COMP_LOOP_COMP_LOOP_and_84_itm,
      COMP_LOOP_COMP_LOOP_and_144_itm, COMP_LOOP_COMP_LOOP_and_204_itm, COMP_LOOP_COMP_LOOP_and_264_itm,
      COMP_LOOP_COMP_LOOP_and_324_itm, COMP_LOOP_COMP_LOOP_and_384_itm, COMP_LOOP_COMP_LOOP_and_444_itm,
      COMP_LOOP_COMP_LOOP_and_504_itm, COMP_LOOP_COMP_LOOP_and_564_itm, COMP_LOOP_COMP_LOOP_and_624_itm,
      COMP_LOOP_COMP_LOOP_and_684_itm, COMP_LOOP_COMP_LOOP_and_744_itm, COMP_LOOP_COMP_LOOP_and_804_itm,
      COMP_LOOP_COMP_LOOP_and_864_itm, COMP_LOOP_COMP_LOOP_and_924_itm, STD_LOGIC_VECTOR'(
      and_dcpl_571 & and_dcpl_577 & and_1025_cse & and_1028_cse & and_dcpl_589 &
      and_1037_cse & and_1040_cse & and_1044_cse & and_1046_cse & and_1051_cse &
      and_1052_cse & and_1055_cse & and_1056_cse & and_1060_cse & and_1061_cse &
      and_1064_cse));
  COMP_LOOP_mux1h_729_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_10_itm, COMP_LOOP_COMP_LOOP_and_85_itm,
      COMP_LOOP_COMP_LOOP_and_145_itm, COMP_LOOP_COMP_LOOP_and_205_itm, COMP_LOOP_COMP_LOOP_and_265_itm,
      COMP_LOOP_COMP_LOOP_and_325_itm, COMP_LOOP_COMP_LOOP_and_385_itm, COMP_LOOP_COMP_LOOP_and_445_itm,
      COMP_LOOP_COMP_LOOP_and_505_itm, COMP_LOOP_COMP_LOOP_and_565_itm, COMP_LOOP_COMP_LOOP_and_625_itm,
      COMP_LOOP_COMP_LOOP_and_685_itm, COMP_LOOP_COMP_LOOP_and_745_itm, COMP_LOOP_COMP_LOOP_and_805_itm,
      COMP_LOOP_COMP_LOOP_and_865_itm, COMP_LOOP_COMP_LOOP_and_925_itm, STD_LOGIC_VECTOR'(
      and_dcpl_571 & and_dcpl_577 & and_1025_cse & and_1028_cse & and_dcpl_589 &
      and_1037_cse & and_1040_cse & and_1044_cse & and_1046_cse & and_1051_cse &
      and_1052_cse & and_1055_cse & and_1056_cse & and_1060_cse & and_1061_cse &
      and_1064_cse));
  COMP_LOOP_mux1h_730_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_72_itm, COMP_LOOP_COMP_LOOP_and_86_itm,
      COMP_LOOP_COMP_LOOP_and_146_itm, COMP_LOOP_COMP_LOOP_and_206_itm, COMP_LOOP_COMP_LOOP_and_266_itm,
      COMP_LOOP_COMP_LOOP_and_326_itm, COMP_LOOP_COMP_LOOP_and_386_itm, COMP_LOOP_COMP_LOOP_and_446_itm,
      COMP_LOOP_COMP_LOOP_and_506_itm, COMP_LOOP_COMP_LOOP_and_566_itm, COMP_LOOP_COMP_LOOP_and_626_itm,
      COMP_LOOP_COMP_LOOP_and_686_itm, COMP_LOOP_COMP_LOOP_and_746_itm, COMP_LOOP_COMP_LOOP_and_806_itm,
      COMP_LOOP_COMP_LOOP_and_866_itm, COMP_LOOP_COMP_LOOP_and_926_itm, STD_LOGIC_VECTOR'(
      and_dcpl_571 & and_dcpl_577 & and_1025_cse & and_1028_cse & and_dcpl_589 &
      and_1037_cse & and_1040_cse & and_1044_cse & and_1046_cse & and_1051_cse &
      and_1052_cse & and_1055_cse & and_1056_cse & and_1060_cse & and_1061_cse &
      and_1064_cse));
  COMP_LOOP_mux1h_731_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_12_itm, COMP_LOOP_COMP_LOOP_and_87_itm,
      COMP_LOOP_COMP_LOOP_and_147_itm, COMP_LOOP_COMP_LOOP_and_207_itm, COMP_LOOP_COMP_LOOP_and_267_itm,
      COMP_LOOP_COMP_LOOP_and_327_itm, COMP_LOOP_COMP_LOOP_and_387_itm, COMP_LOOP_COMP_LOOP_and_447_itm,
      COMP_LOOP_COMP_LOOP_and_507_itm, COMP_LOOP_COMP_LOOP_and_567_itm, COMP_LOOP_COMP_LOOP_and_627_itm,
      COMP_LOOP_COMP_LOOP_and_687_itm, COMP_LOOP_COMP_LOOP_and_747_itm, COMP_LOOP_COMP_LOOP_and_807_itm,
      COMP_LOOP_COMP_LOOP_and_867_itm, COMP_LOOP_COMP_LOOP_and_927_itm, STD_LOGIC_VECTOR'(
      and_dcpl_571 & and_dcpl_577 & and_1025_cse & and_1028_cse & and_dcpl_589 &
      and_1037_cse & and_1040_cse & and_1044_cse & and_1046_cse & and_1051_cse &
      and_1052_cse & and_1055_cse & and_1056_cse & and_1060_cse & and_1061_cse &
      and_1064_cse));
  COMP_LOOP_mux1h_732_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_13_itm, COMP_LOOP_COMP_LOOP_and_88_itm,
      COMP_LOOP_COMP_LOOP_and_148_itm, COMP_LOOP_COMP_LOOP_and_208_itm, COMP_LOOP_COMP_LOOP_and_268_itm,
      COMP_LOOP_COMP_LOOP_and_328_itm, COMP_LOOP_COMP_LOOP_and_388_itm, COMP_LOOP_COMP_LOOP_and_448_itm,
      COMP_LOOP_COMP_LOOP_and_508_itm, COMP_LOOP_COMP_LOOP_and_568_itm, COMP_LOOP_COMP_LOOP_and_628_itm,
      COMP_LOOP_COMP_LOOP_and_688_itm, COMP_LOOP_COMP_LOOP_and_748_itm, COMP_LOOP_COMP_LOOP_and_808_itm,
      COMP_LOOP_COMP_LOOP_and_868_itm, COMP_LOOP_COMP_LOOP_and_928_itm, STD_LOGIC_VECTOR'(
      and_dcpl_571 & and_dcpl_577 & and_1025_cse & and_1028_cse & and_dcpl_589 &
      and_1037_cse & and_1040_cse & and_1044_cse & and_1046_cse & and_1051_cse &
      and_1052_cse & and_1055_cse & and_1056_cse & and_1060_cse & and_1061_cse &
      and_1064_cse));
  COMP_LOOP_mux1h_733_nl <= MUX1HOT_s_1_16_2(COMP_LOOP_COMP_LOOP_and_14_itm, COMP_LOOP_COMP_LOOP_and_89_itm,
      COMP_LOOP_COMP_LOOP_and_149_itm, COMP_LOOP_COMP_LOOP_and_209_itm, COMP_LOOP_COMP_LOOP_and_269_itm,
      COMP_LOOP_COMP_LOOP_and_329_itm, COMP_LOOP_COMP_LOOP_and_389_itm, COMP_LOOP_COMP_LOOP_and_449_itm,
      COMP_LOOP_COMP_LOOP_and_509_itm, COMP_LOOP_COMP_LOOP_and_569_itm, COMP_LOOP_COMP_LOOP_and_629_itm,
      COMP_LOOP_COMP_LOOP_and_689_itm, COMP_LOOP_COMP_LOOP_and_749_itm, COMP_LOOP_COMP_LOOP_and_809_itm,
      COMP_LOOP_COMP_LOOP_and_869_itm, COMP_LOOP_COMP_LOOP_and_929_itm, STD_LOGIC_VECTOR'(
      and_dcpl_571 & and_dcpl_577 & and_1025_cse & and_1028_cse & and_dcpl_589 &
      and_1037_cse & and_1040_cse & and_1044_cse & and_1046_cse & and_1051_cse &
      and_1052_cse & and_1055_cse & and_1056_cse & and_1060_cse & and_1061_cse &
      and_1064_cse));
  z_out_7 <= MUX1HOT_v_64_16_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d, vec_rsc_0_2_i_q_d,
      vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d, vec_rsc_0_6_i_q_d,
      vec_rsc_0_7_i_q_d, vec_rsc_0_8_i_q_d, vec_rsc_0_9_i_q_d, vec_rsc_0_10_i_q_d,
      vec_rsc_0_11_i_q_d, vec_rsc_0_12_i_q_d, vec_rsc_0_13_i_q_d, vec_rsc_0_14_i_q_d,
      vec_rsc_0_15_i_q_d, STD_LOGIC_VECTOR'( COMP_LOOP_mux1h_718_nl & COMP_LOOP_mux1h_719_nl
      & COMP_LOOP_mux1h_720_nl & COMP_LOOP_mux1h_721_nl & COMP_LOOP_mux1h_722_nl
      & COMP_LOOP_mux1h_723_nl & COMP_LOOP_mux1h_724_nl & COMP_LOOP_mux1h_725_nl
      & COMP_LOOP_mux1h_726_nl & COMP_LOOP_mux1h_727_nl & COMP_LOOP_mux1h_728_nl
      & COMP_LOOP_mux1h_729_nl & COMP_LOOP_mux1h_730_nl & COMP_LOOP_mux1h_731_nl
      & COMP_LOOP_mux1h_732_nl & COMP_LOOP_mux1h_733_nl));
END v7;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_0_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_0_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_we : OUT STD_LOGIC;
    vec_rsc_0_0_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_0_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_0_1_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_1_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_we : OUT STD_LOGIC;
    vec_rsc_0_1_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_1_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_0_2_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_2_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_we : OUT STD_LOGIC;
    vec_rsc_0_2_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_2_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_0_3_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_3_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_we : OUT STD_LOGIC;
    vec_rsc_0_3_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_3_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_0_4_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_4_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_we : OUT STD_LOGIC;
    vec_rsc_0_4_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_4_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_0_5_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_5_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_we : OUT STD_LOGIC;
    vec_rsc_0_5_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_5_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_0_6_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_6_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_we : OUT STD_LOGIC;
    vec_rsc_0_6_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_6_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_0_7_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_7_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_we : OUT STD_LOGIC;
    vec_rsc_0_7_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_7_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    vec_rsc_0_8_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_8_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_8_we : OUT STD_LOGIC;
    vec_rsc_0_8_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_8_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    vec_rsc_0_9_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_9_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_9_we : OUT STD_LOGIC;
    vec_rsc_0_9_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_9_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    vec_rsc_0_10_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_10_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_10_we : OUT STD_LOGIC;
    vec_rsc_0_10_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_10_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    vec_rsc_0_11_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_11_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_11_we : OUT STD_LOGIC;
    vec_rsc_0_11_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_11_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    vec_rsc_0_12_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_12_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_12_we : OUT STD_LOGIC;
    vec_rsc_0_12_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_12_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    vec_rsc_0_13_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_13_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_13_we : OUT STD_LOGIC;
    vec_rsc_0_13_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_13_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    vec_rsc_0_14_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_14_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_14_we : OUT STD_LOGIC;
    vec_rsc_0_14_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_14_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    vec_rsc_0_15_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_15_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_15_we : OUT STD_LOGIC;
    vec_rsc_0_15_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_15_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsc_0_0_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_0_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_rsc_0_1_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_1_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_rsc_0_2_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_2_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_rsc_0_3_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_3_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_rsc_0_4_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_4_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_rsc_0_5_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_5_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_rsc_0_6_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_6_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_rsc_0_7_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_7_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_rsc_0_8_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_8_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_rsc_0_9_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_9_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_rsc_0_10_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_10_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_rsc_0_11_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_11_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_rsc_0_12_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_12_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_rsc_0_13_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_13_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_rsc_0_14_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_14_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_rsc_0_15_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_15_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC
  );
END inPlaceNTT_DIF;

ARCHITECTURE v7 OF inPlaceNTT_DIF IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_0_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_8_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_9_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_10_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_11_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_12_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_13_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_14_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_15_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_0_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_1_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_2_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_3_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_4_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_5_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_6_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_7_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_8_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_9_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_10_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_11_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_12_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_13_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_14_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_15_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_d_d_iff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_radr_d_iff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wadr_d_iff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_8_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_9_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_10_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_11_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_12_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_13_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_14_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_15_i_we_d_iff : STD_LOGIC;
  SIGNAL twiddle_rsc_0_1_i_radr_d_iff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_radr_d_iff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_radr_d_iff : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_0_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_1_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_2_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_3_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_4_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_5_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_6_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_7_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_8_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_9_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_10_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_11_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_12_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_13_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_14_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_15_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_25_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_0_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_radr_d_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_26_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_1_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_27_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_2_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_28_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_3_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_29_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_4_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_30_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_5_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_31_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_6_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_32_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_7_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_33_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_8_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_radr_d_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_34_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_9_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_35_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_10_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_36_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_11_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_37_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_12_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_38_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_13_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_39_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_14_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_40_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_15_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      p_rsc_triosy_lz : OUT STD_LOGIC;
      r_rsc_triosy_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      vec_rsc_0_0_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_1_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_2_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_3_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_4_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_5_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_6_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_7_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_8_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_9_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_10_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_11_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_12_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_13_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_14_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_15_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_0_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_0_i_radr_d : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_1_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_2_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_3_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_4_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_5_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_6_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_7_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_8_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_8_i_radr_d : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_9_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_10_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_11_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_12_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_13_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_14_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_15_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_0_i_d_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_radr_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      vec_rsc_0_0_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      vec_rsc_0_0_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_1_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_2_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_3_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_4_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_5_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_6_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_7_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_8_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_9_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_10_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_11_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_12_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_13_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_14_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_15_i_we_d_pff : OUT STD_LOGIC;
      twiddle_rsc_0_1_i_radr_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_2_i_radr_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_4_i_radr_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_core_inst_p_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_1_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_2_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_3_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_4_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_5_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_6_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_7_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_8_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_9_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_10_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_11_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_12_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_13_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_14_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_15_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_radr_d : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_3_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_5_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_6_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_7_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_8_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_8_i_radr_d : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_9_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_10_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_11_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_12_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_13_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_14_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_15_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_d_d_pff : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_radr_d_pff : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_wadr_d_pff : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_radr_d_pff : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_radr_d_pff : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_radr_d_pff : STD_LOGIC_VECTOR
      (5 DOWNTO 0);

BEGIN
  vec_rsc_0_0_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_0_i_q,
      radr => vec_rsc_0_0_i_radr,
      we => vec_rsc_0_0_we,
      d => vec_rsc_0_0_i_d,
      wadr => vec_rsc_0_0_i_wadr,
      d_d => vec_rsc_0_0_i_d_d,
      q_d => vec_rsc_0_0_i_q_d_1,
      radr_d => vec_rsc_0_0_i_radr_d,
      wadr_d => vec_rsc_0_0_i_wadr_d,
      we_d => vec_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_0_i_q <= vec_rsc_0_0_q;
  vec_rsc_0_0_radr <= vec_rsc_0_0_i_radr;
  vec_rsc_0_0_d <= vec_rsc_0_0_i_d;
  vec_rsc_0_0_wadr <= vec_rsc_0_0_i_wadr;
  vec_rsc_0_0_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_0_i_q_d <= vec_rsc_0_0_i_q_d_1;
  vec_rsc_0_0_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_0_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_1_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_1_i_q,
      radr => vec_rsc_0_1_i_radr,
      we => vec_rsc_0_1_we,
      d => vec_rsc_0_1_i_d,
      wadr => vec_rsc_0_1_i_wadr,
      d_d => vec_rsc_0_1_i_d_d,
      q_d => vec_rsc_0_1_i_q_d_1,
      radr_d => vec_rsc_0_1_i_radr_d,
      wadr_d => vec_rsc_0_1_i_wadr_d,
      we_d => vec_rsc_0_1_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_1_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_1_i_q <= vec_rsc_0_1_q;
  vec_rsc_0_1_radr <= vec_rsc_0_1_i_radr;
  vec_rsc_0_1_d <= vec_rsc_0_1_i_d;
  vec_rsc_0_1_wadr <= vec_rsc_0_1_i_wadr;
  vec_rsc_0_1_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_1_i_q_d <= vec_rsc_0_1_i_q_d_1;
  vec_rsc_0_1_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_1_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_2_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_2_i_q,
      radr => vec_rsc_0_2_i_radr,
      we => vec_rsc_0_2_we,
      d => vec_rsc_0_2_i_d,
      wadr => vec_rsc_0_2_i_wadr,
      d_d => vec_rsc_0_2_i_d_d,
      q_d => vec_rsc_0_2_i_q_d_1,
      radr_d => vec_rsc_0_2_i_radr_d,
      wadr_d => vec_rsc_0_2_i_wadr_d,
      we_d => vec_rsc_0_2_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_2_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_2_i_q <= vec_rsc_0_2_q;
  vec_rsc_0_2_radr <= vec_rsc_0_2_i_radr;
  vec_rsc_0_2_d <= vec_rsc_0_2_i_d;
  vec_rsc_0_2_wadr <= vec_rsc_0_2_i_wadr;
  vec_rsc_0_2_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_2_i_q_d <= vec_rsc_0_2_i_q_d_1;
  vec_rsc_0_2_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_2_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_3_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_3_i_q,
      radr => vec_rsc_0_3_i_radr,
      we => vec_rsc_0_3_we,
      d => vec_rsc_0_3_i_d,
      wadr => vec_rsc_0_3_i_wadr,
      d_d => vec_rsc_0_3_i_d_d,
      q_d => vec_rsc_0_3_i_q_d_1,
      radr_d => vec_rsc_0_3_i_radr_d,
      wadr_d => vec_rsc_0_3_i_wadr_d,
      we_d => vec_rsc_0_3_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_3_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_3_i_q <= vec_rsc_0_3_q;
  vec_rsc_0_3_radr <= vec_rsc_0_3_i_radr;
  vec_rsc_0_3_d <= vec_rsc_0_3_i_d;
  vec_rsc_0_3_wadr <= vec_rsc_0_3_i_wadr;
  vec_rsc_0_3_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_3_i_q_d <= vec_rsc_0_3_i_q_d_1;
  vec_rsc_0_3_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_3_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_4_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_4_i_q,
      radr => vec_rsc_0_4_i_radr,
      we => vec_rsc_0_4_we,
      d => vec_rsc_0_4_i_d,
      wadr => vec_rsc_0_4_i_wadr,
      d_d => vec_rsc_0_4_i_d_d,
      q_d => vec_rsc_0_4_i_q_d_1,
      radr_d => vec_rsc_0_4_i_radr_d,
      wadr_d => vec_rsc_0_4_i_wadr_d,
      we_d => vec_rsc_0_4_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_4_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_4_i_q <= vec_rsc_0_4_q;
  vec_rsc_0_4_radr <= vec_rsc_0_4_i_radr;
  vec_rsc_0_4_d <= vec_rsc_0_4_i_d;
  vec_rsc_0_4_wadr <= vec_rsc_0_4_i_wadr;
  vec_rsc_0_4_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_4_i_q_d <= vec_rsc_0_4_i_q_d_1;
  vec_rsc_0_4_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_4_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_5_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_5_i_q,
      radr => vec_rsc_0_5_i_radr,
      we => vec_rsc_0_5_we,
      d => vec_rsc_0_5_i_d,
      wadr => vec_rsc_0_5_i_wadr,
      d_d => vec_rsc_0_5_i_d_d,
      q_d => vec_rsc_0_5_i_q_d_1,
      radr_d => vec_rsc_0_5_i_radr_d,
      wadr_d => vec_rsc_0_5_i_wadr_d,
      we_d => vec_rsc_0_5_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_5_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_5_i_q <= vec_rsc_0_5_q;
  vec_rsc_0_5_radr <= vec_rsc_0_5_i_radr;
  vec_rsc_0_5_d <= vec_rsc_0_5_i_d;
  vec_rsc_0_5_wadr <= vec_rsc_0_5_i_wadr;
  vec_rsc_0_5_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_5_i_q_d <= vec_rsc_0_5_i_q_d_1;
  vec_rsc_0_5_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_5_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_6_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_6_i_q,
      radr => vec_rsc_0_6_i_radr,
      we => vec_rsc_0_6_we,
      d => vec_rsc_0_6_i_d,
      wadr => vec_rsc_0_6_i_wadr,
      d_d => vec_rsc_0_6_i_d_d,
      q_d => vec_rsc_0_6_i_q_d_1,
      radr_d => vec_rsc_0_6_i_radr_d,
      wadr_d => vec_rsc_0_6_i_wadr_d,
      we_d => vec_rsc_0_6_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_6_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_6_i_q <= vec_rsc_0_6_q;
  vec_rsc_0_6_radr <= vec_rsc_0_6_i_radr;
  vec_rsc_0_6_d <= vec_rsc_0_6_i_d;
  vec_rsc_0_6_wadr <= vec_rsc_0_6_i_wadr;
  vec_rsc_0_6_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_6_i_q_d <= vec_rsc_0_6_i_q_d_1;
  vec_rsc_0_6_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_6_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_7_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_7_i_q,
      radr => vec_rsc_0_7_i_radr,
      we => vec_rsc_0_7_we,
      d => vec_rsc_0_7_i_d,
      wadr => vec_rsc_0_7_i_wadr,
      d_d => vec_rsc_0_7_i_d_d,
      q_d => vec_rsc_0_7_i_q_d_1,
      radr_d => vec_rsc_0_7_i_radr_d,
      wadr_d => vec_rsc_0_7_i_wadr_d,
      we_d => vec_rsc_0_7_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_7_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_7_i_q <= vec_rsc_0_7_q;
  vec_rsc_0_7_radr <= vec_rsc_0_7_i_radr;
  vec_rsc_0_7_d <= vec_rsc_0_7_i_d;
  vec_rsc_0_7_wadr <= vec_rsc_0_7_i_wadr;
  vec_rsc_0_7_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_7_i_q_d <= vec_rsc_0_7_i_q_d_1;
  vec_rsc_0_7_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_7_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_8_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_8_i_q,
      radr => vec_rsc_0_8_i_radr,
      we => vec_rsc_0_8_we,
      d => vec_rsc_0_8_i_d,
      wadr => vec_rsc_0_8_i_wadr,
      d_d => vec_rsc_0_8_i_d_d,
      q_d => vec_rsc_0_8_i_q_d_1,
      radr_d => vec_rsc_0_8_i_radr_d,
      wadr_d => vec_rsc_0_8_i_wadr_d,
      we_d => vec_rsc_0_8_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_8_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_8_i_q <= vec_rsc_0_8_q;
  vec_rsc_0_8_radr <= vec_rsc_0_8_i_radr;
  vec_rsc_0_8_d <= vec_rsc_0_8_i_d;
  vec_rsc_0_8_wadr <= vec_rsc_0_8_i_wadr;
  vec_rsc_0_8_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_8_i_q_d <= vec_rsc_0_8_i_q_d_1;
  vec_rsc_0_8_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_8_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_9_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_9_i_q,
      radr => vec_rsc_0_9_i_radr,
      we => vec_rsc_0_9_we,
      d => vec_rsc_0_9_i_d,
      wadr => vec_rsc_0_9_i_wadr,
      d_d => vec_rsc_0_9_i_d_d,
      q_d => vec_rsc_0_9_i_q_d_1,
      radr_d => vec_rsc_0_9_i_radr_d,
      wadr_d => vec_rsc_0_9_i_wadr_d,
      we_d => vec_rsc_0_9_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_9_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_9_i_q <= vec_rsc_0_9_q;
  vec_rsc_0_9_radr <= vec_rsc_0_9_i_radr;
  vec_rsc_0_9_d <= vec_rsc_0_9_i_d;
  vec_rsc_0_9_wadr <= vec_rsc_0_9_i_wadr;
  vec_rsc_0_9_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_9_i_q_d <= vec_rsc_0_9_i_q_d_1;
  vec_rsc_0_9_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_9_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_10_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_10_i_q,
      radr => vec_rsc_0_10_i_radr,
      we => vec_rsc_0_10_we,
      d => vec_rsc_0_10_i_d,
      wadr => vec_rsc_0_10_i_wadr,
      d_d => vec_rsc_0_10_i_d_d,
      q_d => vec_rsc_0_10_i_q_d_1,
      radr_d => vec_rsc_0_10_i_radr_d,
      wadr_d => vec_rsc_0_10_i_wadr_d,
      we_d => vec_rsc_0_10_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_10_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_10_i_q <= vec_rsc_0_10_q;
  vec_rsc_0_10_radr <= vec_rsc_0_10_i_radr;
  vec_rsc_0_10_d <= vec_rsc_0_10_i_d;
  vec_rsc_0_10_wadr <= vec_rsc_0_10_i_wadr;
  vec_rsc_0_10_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_10_i_q_d <= vec_rsc_0_10_i_q_d_1;
  vec_rsc_0_10_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_10_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_11_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_11_i_q,
      radr => vec_rsc_0_11_i_radr,
      we => vec_rsc_0_11_we,
      d => vec_rsc_0_11_i_d,
      wadr => vec_rsc_0_11_i_wadr,
      d_d => vec_rsc_0_11_i_d_d,
      q_d => vec_rsc_0_11_i_q_d_1,
      radr_d => vec_rsc_0_11_i_radr_d,
      wadr_d => vec_rsc_0_11_i_wadr_d,
      we_d => vec_rsc_0_11_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_11_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_11_i_q <= vec_rsc_0_11_q;
  vec_rsc_0_11_radr <= vec_rsc_0_11_i_radr;
  vec_rsc_0_11_d <= vec_rsc_0_11_i_d;
  vec_rsc_0_11_wadr <= vec_rsc_0_11_i_wadr;
  vec_rsc_0_11_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_11_i_q_d <= vec_rsc_0_11_i_q_d_1;
  vec_rsc_0_11_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_11_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_12_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_12_i_q,
      radr => vec_rsc_0_12_i_radr,
      we => vec_rsc_0_12_we,
      d => vec_rsc_0_12_i_d,
      wadr => vec_rsc_0_12_i_wadr,
      d_d => vec_rsc_0_12_i_d_d,
      q_d => vec_rsc_0_12_i_q_d_1,
      radr_d => vec_rsc_0_12_i_radr_d,
      wadr_d => vec_rsc_0_12_i_wadr_d,
      we_d => vec_rsc_0_12_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_12_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_12_i_q <= vec_rsc_0_12_q;
  vec_rsc_0_12_radr <= vec_rsc_0_12_i_radr;
  vec_rsc_0_12_d <= vec_rsc_0_12_i_d;
  vec_rsc_0_12_wadr <= vec_rsc_0_12_i_wadr;
  vec_rsc_0_12_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_12_i_q_d <= vec_rsc_0_12_i_q_d_1;
  vec_rsc_0_12_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_12_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_13_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_13_i_q,
      radr => vec_rsc_0_13_i_radr,
      we => vec_rsc_0_13_we,
      d => vec_rsc_0_13_i_d,
      wadr => vec_rsc_0_13_i_wadr,
      d_d => vec_rsc_0_13_i_d_d,
      q_d => vec_rsc_0_13_i_q_d_1,
      radr_d => vec_rsc_0_13_i_radr_d,
      wadr_d => vec_rsc_0_13_i_wadr_d,
      we_d => vec_rsc_0_13_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_13_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_13_i_q <= vec_rsc_0_13_q;
  vec_rsc_0_13_radr <= vec_rsc_0_13_i_radr;
  vec_rsc_0_13_d <= vec_rsc_0_13_i_d;
  vec_rsc_0_13_wadr <= vec_rsc_0_13_i_wadr;
  vec_rsc_0_13_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_13_i_q_d <= vec_rsc_0_13_i_q_d_1;
  vec_rsc_0_13_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_13_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_14_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_14_i_q,
      radr => vec_rsc_0_14_i_radr,
      we => vec_rsc_0_14_we,
      d => vec_rsc_0_14_i_d,
      wadr => vec_rsc_0_14_i_wadr,
      d_d => vec_rsc_0_14_i_d_d,
      q_d => vec_rsc_0_14_i_q_d_1,
      radr_d => vec_rsc_0_14_i_radr_d,
      wadr_d => vec_rsc_0_14_i_wadr_d,
      we_d => vec_rsc_0_14_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_14_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_14_i_q <= vec_rsc_0_14_q;
  vec_rsc_0_14_radr <= vec_rsc_0_14_i_radr;
  vec_rsc_0_14_d <= vec_rsc_0_14_i_d;
  vec_rsc_0_14_wadr <= vec_rsc_0_14_i_wadr;
  vec_rsc_0_14_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_14_i_q_d <= vec_rsc_0_14_i_q_d_1;
  vec_rsc_0_14_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_14_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_15_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_15_i_q,
      radr => vec_rsc_0_15_i_radr,
      we => vec_rsc_0_15_we,
      d => vec_rsc_0_15_i_d,
      wadr => vec_rsc_0_15_i_wadr,
      d_d => vec_rsc_0_15_i_d_d,
      q_d => vec_rsc_0_15_i_q_d_1,
      radr_d => vec_rsc_0_15_i_radr_d,
      wadr_d => vec_rsc_0_15_i_wadr_d,
      we_d => vec_rsc_0_15_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_15_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_15_i_q <= vec_rsc_0_15_q;
  vec_rsc_0_15_radr <= vec_rsc_0_15_i_radr;
  vec_rsc_0_15_d <= vec_rsc_0_15_i_d;
  vec_rsc_0_15_wadr <= vec_rsc_0_15_i_wadr;
  vec_rsc_0_15_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_15_i_q_d <= vec_rsc_0_15_i_q_d_1;
  vec_rsc_0_15_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_15_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  twiddle_rsc_0_0_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_25_6_64_64_64_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_0_i_q,
      radr => twiddle_rsc_0_0_i_radr,
      q_d => twiddle_rsc_0_0_i_q_d_1,
      radr_d => twiddle_rsc_0_0_i_radr_d_1,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_0_i_q <= twiddle_rsc_0_0_q;
  twiddle_rsc_0_0_radr <= twiddle_rsc_0_0_i_radr;
  twiddle_rsc_0_0_i_q_d <= twiddle_rsc_0_0_i_q_d_1;
  twiddle_rsc_0_0_i_radr_d_1 <= twiddle_rsc_0_0_i_radr_d;

  twiddle_rsc_0_1_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_26_6_64_64_64_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_1_i_q,
      radr => twiddle_rsc_0_1_i_radr,
      q_d => twiddle_rsc_0_1_i_q_d_1,
      radr_d => twiddle_rsc_0_1_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_1_i_q <= twiddle_rsc_0_1_q;
  twiddle_rsc_0_1_radr <= twiddle_rsc_0_1_i_radr;
  twiddle_rsc_0_1_i_q_d <= twiddle_rsc_0_1_i_q_d_1;
  twiddle_rsc_0_1_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_2_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_27_6_64_64_64_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_2_i_q,
      radr => twiddle_rsc_0_2_i_radr,
      q_d => twiddle_rsc_0_2_i_q_d_1,
      radr_d => twiddle_rsc_0_2_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_2_i_q <= twiddle_rsc_0_2_q;
  twiddle_rsc_0_2_radr <= twiddle_rsc_0_2_i_radr;
  twiddle_rsc_0_2_i_q_d <= twiddle_rsc_0_2_i_q_d_1;
  twiddle_rsc_0_2_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_3_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_28_6_64_64_64_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_3_i_q,
      radr => twiddle_rsc_0_3_i_radr,
      q_d => twiddle_rsc_0_3_i_q_d_1,
      radr_d => twiddle_rsc_0_3_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_3_i_q <= twiddle_rsc_0_3_q;
  twiddle_rsc_0_3_radr <= twiddle_rsc_0_3_i_radr;
  twiddle_rsc_0_3_i_q_d <= twiddle_rsc_0_3_i_q_d_1;
  twiddle_rsc_0_3_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_4_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_29_6_64_64_64_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_4_i_q,
      radr => twiddle_rsc_0_4_i_radr,
      q_d => twiddle_rsc_0_4_i_q_d_1,
      radr_d => twiddle_rsc_0_4_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_4_i_q <= twiddle_rsc_0_4_q;
  twiddle_rsc_0_4_radr <= twiddle_rsc_0_4_i_radr;
  twiddle_rsc_0_4_i_q_d <= twiddle_rsc_0_4_i_q_d_1;
  twiddle_rsc_0_4_i_radr_d <= twiddle_rsc_0_4_i_radr_d_iff;

  twiddle_rsc_0_5_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_30_6_64_64_64_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_5_i_q,
      radr => twiddle_rsc_0_5_i_radr,
      q_d => twiddle_rsc_0_5_i_q_d_1,
      radr_d => twiddle_rsc_0_5_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_5_i_q <= twiddle_rsc_0_5_q;
  twiddle_rsc_0_5_radr <= twiddle_rsc_0_5_i_radr;
  twiddle_rsc_0_5_i_q_d <= twiddle_rsc_0_5_i_q_d_1;
  twiddle_rsc_0_5_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_6_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_31_6_64_64_64_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_6_i_q,
      radr => twiddle_rsc_0_6_i_radr,
      q_d => twiddle_rsc_0_6_i_q_d_1,
      radr_d => twiddle_rsc_0_6_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_6_i_q <= twiddle_rsc_0_6_q;
  twiddle_rsc_0_6_radr <= twiddle_rsc_0_6_i_radr;
  twiddle_rsc_0_6_i_q_d <= twiddle_rsc_0_6_i_q_d_1;
  twiddle_rsc_0_6_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_7_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_32_6_64_64_64_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_7_i_q,
      radr => twiddle_rsc_0_7_i_radr,
      q_d => twiddle_rsc_0_7_i_q_d_1,
      radr_d => twiddle_rsc_0_7_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_7_i_q <= twiddle_rsc_0_7_q;
  twiddle_rsc_0_7_radr <= twiddle_rsc_0_7_i_radr;
  twiddle_rsc_0_7_i_q_d <= twiddle_rsc_0_7_i_q_d_1;
  twiddle_rsc_0_7_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_8_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_33_6_64_64_64_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_8_i_q,
      radr => twiddle_rsc_0_8_i_radr,
      q_d => twiddle_rsc_0_8_i_q_d_1,
      radr_d => twiddle_rsc_0_8_i_radr_d_1,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_8_i_q <= twiddle_rsc_0_8_q;
  twiddle_rsc_0_8_radr <= twiddle_rsc_0_8_i_radr;
  twiddle_rsc_0_8_i_q_d <= twiddle_rsc_0_8_i_q_d_1;
  twiddle_rsc_0_8_i_radr_d_1 <= twiddle_rsc_0_8_i_radr_d;

  twiddle_rsc_0_9_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_34_6_64_64_64_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_9_i_q,
      radr => twiddle_rsc_0_9_i_radr,
      q_d => twiddle_rsc_0_9_i_q_d_1,
      radr_d => twiddle_rsc_0_9_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_9_i_q <= twiddle_rsc_0_9_q;
  twiddle_rsc_0_9_radr <= twiddle_rsc_0_9_i_radr;
  twiddle_rsc_0_9_i_q_d <= twiddle_rsc_0_9_i_q_d_1;
  twiddle_rsc_0_9_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_10_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_35_6_64_64_64_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_10_i_q,
      radr => twiddle_rsc_0_10_i_radr,
      q_d => twiddle_rsc_0_10_i_q_d_1,
      radr_d => twiddle_rsc_0_10_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_10_i_q <= twiddle_rsc_0_10_q;
  twiddle_rsc_0_10_radr <= twiddle_rsc_0_10_i_radr;
  twiddle_rsc_0_10_i_q_d <= twiddle_rsc_0_10_i_q_d_1;
  twiddle_rsc_0_10_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_11_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_36_6_64_64_64_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_11_i_q,
      radr => twiddle_rsc_0_11_i_radr,
      q_d => twiddle_rsc_0_11_i_q_d_1,
      radr_d => twiddle_rsc_0_11_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_11_i_q <= twiddle_rsc_0_11_q;
  twiddle_rsc_0_11_radr <= twiddle_rsc_0_11_i_radr;
  twiddle_rsc_0_11_i_q_d <= twiddle_rsc_0_11_i_q_d_1;
  twiddle_rsc_0_11_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_12_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_37_6_64_64_64_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_12_i_q,
      radr => twiddle_rsc_0_12_i_radr,
      q_d => twiddle_rsc_0_12_i_q_d_1,
      radr_d => twiddle_rsc_0_12_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_12_i_q <= twiddle_rsc_0_12_q;
  twiddle_rsc_0_12_radr <= twiddle_rsc_0_12_i_radr;
  twiddle_rsc_0_12_i_q_d <= twiddle_rsc_0_12_i_q_d_1;
  twiddle_rsc_0_12_i_radr_d <= twiddle_rsc_0_4_i_radr_d_iff;

  twiddle_rsc_0_13_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_38_6_64_64_64_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_13_i_q,
      radr => twiddle_rsc_0_13_i_radr,
      q_d => twiddle_rsc_0_13_i_q_d_1,
      radr_d => twiddle_rsc_0_13_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_13_i_q <= twiddle_rsc_0_13_q;
  twiddle_rsc_0_13_radr <= twiddle_rsc_0_13_i_radr;
  twiddle_rsc_0_13_i_q_d <= twiddle_rsc_0_13_i_q_d_1;
  twiddle_rsc_0_13_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_14_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_39_6_64_64_64_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_14_i_q,
      radr => twiddle_rsc_0_14_i_radr,
      q_d => twiddle_rsc_0_14_i_q_d_1,
      radr_d => twiddle_rsc_0_14_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_14_i_q <= twiddle_rsc_0_14_q;
  twiddle_rsc_0_14_radr <= twiddle_rsc_0_14_i_radr;
  twiddle_rsc_0_14_i_q_d <= twiddle_rsc_0_14_i_q_d_1;
  twiddle_rsc_0_14_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_15_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_40_6_64_64_64_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_15_i_q,
      radr => twiddle_rsc_0_15_i_radr,
      q_d => twiddle_rsc_0_15_i_q_d_1,
      radr_d => twiddle_rsc_0_15_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_15_i_q <= twiddle_rsc_0_15_q;
  twiddle_rsc_0_15_radr <= twiddle_rsc_0_15_i_radr;
  twiddle_rsc_0_15_i_q_d <= twiddle_rsc_0_15_i_q_d_1;
  twiddle_rsc_0_15_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  inPlaceNTT_DIF_core_inst : inPlaceNTT_DIF_core
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_triosy_0_0_lz => vec_rsc_triosy_0_0_lz,
      vec_rsc_triosy_0_1_lz => vec_rsc_triosy_0_1_lz,
      vec_rsc_triosy_0_2_lz => vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz => vec_rsc_triosy_0_3_lz,
      vec_rsc_triosy_0_4_lz => vec_rsc_triosy_0_4_lz,
      vec_rsc_triosy_0_5_lz => vec_rsc_triosy_0_5_lz,
      vec_rsc_triosy_0_6_lz => vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz => vec_rsc_triosy_0_7_lz,
      vec_rsc_triosy_0_8_lz => vec_rsc_triosy_0_8_lz,
      vec_rsc_triosy_0_9_lz => vec_rsc_triosy_0_9_lz,
      vec_rsc_triosy_0_10_lz => vec_rsc_triosy_0_10_lz,
      vec_rsc_triosy_0_11_lz => vec_rsc_triosy_0_11_lz,
      vec_rsc_triosy_0_12_lz => vec_rsc_triosy_0_12_lz,
      vec_rsc_triosy_0_13_lz => vec_rsc_triosy_0_13_lz,
      vec_rsc_triosy_0_14_lz => vec_rsc_triosy_0_14_lz,
      vec_rsc_triosy_0_15_lz => vec_rsc_triosy_0_15_lz,
      p_rsc_dat => inPlaceNTT_DIF_core_inst_p_rsc_dat,
      p_rsc_triosy_lz => p_rsc_triosy_lz,
      r_rsc_triosy_lz => r_rsc_triosy_lz,
      twiddle_rsc_triosy_0_0_lz => twiddle_rsc_triosy_0_0_lz,
      twiddle_rsc_triosy_0_1_lz => twiddle_rsc_triosy_0_1_lz,
      twiddle_rsc_triosy_0_2_lz => twiddle_rsc_triosy_0_2_lz,
      twiddle_rsc_triosy_0_3_lz => twiddle_rsc_triosy_0_3_lz,
      twiddle_rsc_triosy_0_4_lz => twiddle_rsc_triosy_0_4_lz,
      twiddle_rsc_triosy_0_5_lz => twiddle_rsc_triosy_0_5_lz,
      twiddle_rsc_triosy_0_6_lz => twiddle_rsc_triosy_0_6_lz,
      twiddle_rsc_triosy_0_7_lz => twiddle_rsc_triosy_0_7_lz,
      twiddle_rsc_triosy_0_8_lz => twiddle_rsc_triosy_0_8_lz,
      twiddle_rsc_triosy_0_9_lz => twiddle_rsc_triosy_0_9_lz,
      twiddle_rsc_triosy_0_10_lz => twiddle_rsc_triosy_0_10_lz,
      twiddle_rsc_triosy_0_11_lz => twiddle_rsc_triosy_0_11_lz,
      twiddle_rsc_triosy_0_12_lz => twiddle_rsc_triosy_0_12_lz,
      twiddle_rsc_triosy_0_13_lz => twiddle_rsc_triosy_0_13_lz,
      twiddle_rsc_triosy_0_14_lz => twiddle_rsc_triosy_0_14_lz,
      twiddle_rsc_triosy_0_15_lz => twiddle_rsc_triosy_0_15_lz,
      vec_rsc_0_0_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_q_d,
      vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_1_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_1_i_q_d,
      vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_2_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_2_i_q_d,
      vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_3_i_q_d,
      vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_4_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_4_i_q_d,
      vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_5_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_5_i_q_d,
      vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_6_i_q_d,
      vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_7_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_7_i_q_d,
      vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_8_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_8_i_q_d,
      vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_9_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_9_i_q_d,
      vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_10_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_10_i_q_d,
      vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_11_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_11_i_q_d,
      vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_12_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_12_i_q_d,
      vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_13_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_13_i_q_d,
      vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_14_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_14_i_q_d,
      vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_15_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_15_i_q_d,
      vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_0_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_q_d,
      twiddle_rsc_0_0_i_radr_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_radr_d,
      twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_1_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_q_d,
      twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_2_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_q_d,
      twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_3_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_3_i_q_d,
      twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_4_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_q_d,
      twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_5_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_5_i_q_d,
      twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_6_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_6_i_q_d,
      twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_7_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_7_i_q_d,
      twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_8_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_8_i_q_d,
      twiddle_rsc_0_8_i_radr_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_8_i_radr_d,
      twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_9_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_9_i_q_d,
      twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_10_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_10_i_q_d,
      twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_11_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_11_i_q_d,
      twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_12_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_12_i_q_d,
      twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_13_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_13_i_q_d,
      twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_14_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_14_i_q_d,
      twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_15_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_15_i_q_d,
      twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_0_i_d_d_pff => inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_d_d_pff,
      vec_rsc_0_0_i_radr_d_pff => inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_radr_d_pff,
      vec_rsc_0_0_i_wadr_d_pff => inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_wadr_d_pff,
      vec_rsc_0_0_i_we_d_pff => vec_rsc_0_0_i_we_d_iff,
      vec_rsc_0_1_i_we_d_pff => vec_rsc_0_1_i_we_d_iff,
      vec_rsc_0_2_i_we_d_pff => vec_rsc_0_2_i_we_d_iff,
      vec_rsc_0_3_i_we_d_pff => vec_rsc_0_3_i_we_d_iff,
      vec_rsc_0_4_i_we_d_pff => vec_rsc_0_4_i_we_d_iff,
      vec_rsc_0_5_i_we_d_pff => vec_rsc_0_5_i_we_d_iff,
      vec_rsc_0_6_i_we_d_pff => vec_rsc_0_6_i_we_d_iff,
      vec_rsc_0_7_i_we_d_pff => vec_rsc_0_7_i_we_d_iff,
      vec_rsc_0_8_i_we_d_pff => vec_rsc_0_8_i_we_d_iff,
      vec_rsc_0_9_i_we_d_pff => vec_rsc_0_9_i_we_d_iff,
      vec_rsc_0_10_i_we_d_pff => vec_rsc_0_10_i_we_d_iff,
      vec_rsc_0_11_i_we_d_pff => vec_rsc_0_11_i_we_d_iff,
      vec_rsc_0_12_i_we_d_pff => vec_rsc_0_12_i_we_d_iff,
      vec_rsc_0_13_i_we_d_pff => vec_rsc_0_13_i_we_d_iff,
      vec_rsc_0_14_i_we_d_pff => vec_rsc_0_14_i_we_d_iff,
      vec_rsc_0_15_i_we_d_pff => vec_rsc_0_15_i_we_d_iff,
      twiddle_rsc_0_1_i_radr_d_pff => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_radr_d_pff,
      twiddle_rsc_0_2_i_radr_d_pff => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_radr_d_pff,
      twiddle_rsc_0_4_i_radr_d_pff => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_radr_d_pff
    );
  inPlaceNTT_DIF_core_inst_p_rsc_dat <= p_rsc_dat;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_q_d <= vec_rsc_0_0_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_1_i_q_d <= vec_rsc_0_1_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_2_i_q_d <= vec_rsc_0_2_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_3_i_q_d <= vec_rsc_0_3_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_4_i_q_d <= vec_rsc_0_4_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_5_i_q_d <= vec_rsc_0_5_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_6_i_q_d <= vec_rsc_0_6_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_7_i_q_d <= vec_rsc_0_7_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_8_i_q_d <= vec_rsc_0_8_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_9_i_q_d <= vec_rsc_0_9_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_10_i_q_d <= vec_rsc_0_10_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_11_i_q_d <= vec_rsc_0_11_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_12_i_q_d <= vec_rsc_0_12_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_13_i_q_d <= vec_rsc_0_13_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_14_i_q_d <= vec_rsc_0_14_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_15_i_q_d <= vec_rsc_0_15_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_q_d <= twiddle_rsc_0_0_i_q_d;
  twiddle_rsc_0_0_i_radr_d <= inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_radr_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_q_d <= twiddle_rsc_0_1_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_q_d <= twiddle_rsc_0_2_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_3_i_q_d <= twiddle_rsc_0_3_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_q_d <= twiddle_rsc_0_4_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_5_i_q_d <= twiddle_rsc_0_5_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_6_i_q_d <= twiddle_rsc_0_6_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_7_i_q_d <= twiddle_rsc_0_7_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_8_i_q_d <= twiddle_rsc_0_8_i_q_d;
  twiddle_rsc_0_8_i_radr_d <= inPlaceNTT_DIF_core_inst_twiddle_rsc_0_8_i_radr_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_9_i_q_d <= twiddle_rsc_0_9_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_10_i_q_d <= twiddle_rsc_0_10_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_11_i_q_d <= twiddle_rsc_0_11_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_12_i_q_d <= twiddle_rsc_0_12_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_13_i_q_d <= twiddle_rsc_0_13_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_14_i_q_d <= twiddle_rsc_0_14_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_15_i_q_d <= twiddle_rsc_0_15_i_q_d;
  vec_rsc_0_0_i_d_d_iff <= inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_d_d_pff;
  vec_rsc_0_0_i_radr_d_iff <= inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_radr_d_pff;
  vec_rsc_0_0_i_wadr_d_iff <= inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_wadr_d_pff;
  twiddle_rsc_0_1_i_radr_d_iff <= inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_radr_d_pff;
  twiddle_rsc_0_2_i_radr_d_iff <= inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_radr_d_pff;
  twiddle_rsc_0_4_i_radr_d_iff <= inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_radr_d_pff;

END v7;



