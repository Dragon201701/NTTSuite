
--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_pkg_v1 IS

COMPONENT ccs_in_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    dat    : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_in_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    dat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_in_v1;

ARCHITECTURE beh OF ccs_in_v1 IS
BEGIN

  idat <= dat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/src/funcs.vhd 

-- a package of attributes that give verification tools a hint about
-- the function being implemented
PACKAGE attributes IS
  ATTRIBUTE CALYPTO_FUNC : string;
  ATTRIBUTE CALYPTO_DATA_ORDER : string;
end attributes;

-----------------------------------------------------------------------
-- Package that declares synthesizable functions needed for RTL output
-----------------------------------------------------------------------

LIBRARY ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

PACKAGE funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

   FUNCTION maximum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION minimum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2 : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;
   
-----------------------------------------------------------------
-- logic functions
-----------------------------------------------------------------

   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION or_v (inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- mux functions
-----------------------------------------------------------------

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC_VECTOR;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- latch functions
-----------------------------------------------------------------
   FUNCTION lat_s(dinput: STD_LOGIC       ; clk: STD_LOGIC; doutput: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- tristate functions
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC       ; control: STD_LOGIC) RETURN STD_LOGIC;
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: SIGNED  ) RETURN STD_LOGIC;

   -- RETURN 2 bits (left => lt, right => eq)
   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED;
 
   FUNCTION fabs(arg1: SIGNED  ) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "**" (l, r: UNSIGNED) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "**" (l, r: SIGNED  ) RETURN SIGNED  ;

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-- *_stdar functions use shift functions from std_logic_arith
-----------------------------------------------------------------

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;

   -----------------------------------------------------------------
   -- *_stdar functions use shift functions from std_logic_arith
   -----------------------------------------------------------------
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC;
   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE;
   --FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR ;

   FUNCTION ceil_log2(size : NATURAL) return NATURAL;
   FUNCTION bits(size : NATURAL) return NATURAL;    

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   
END funcs;


--------------------------- B O D Y ----------------------------


PACKAGE BODY funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC IS
     BEGIN IF arg1 THEN RETURN '1'; ELSE RETURN '0'; END IF; END;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
--     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;

   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
     VARIABLE result: STD_LOGIC_VECTOR(0 DOWNTO 0);
   BEGIN
     result := (0 => arg1);
     RETURN result;
   END;

   FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 > arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION minimum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 < arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;

   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := input1'LENGTH;
     ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
     ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     --synopsys translate_off
     FOR i IN len-1 DOWNTO 0 LOOP
       result(i) := resolved(input1a(i) & input2a(i));
     END LOOP;
     --synopsys translate_on
     RETURN result;
   END;

   FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED) RETURN UNSIGNED IS
   BEGIN RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

   FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED) RETURN SIGNED IS
   BEGIN RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

-----------------------------------------------------------------
-- Logic Functions
-----------------------------------------------------------------

   FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;
   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(and_v(inputs, 1)); END;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(or_v(inputs, 1)); END;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(xor_v(inputs, 1)); END;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result AND inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

   FUNCTION or_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     -- this if is added as a quick fix for a bug in catapult evaluating the loop even if inputs'LENGTH==1
     -- see dts0100971279
     IF icnt2 > 1 THEN
       FOR i IN icnt2-1 DOWNTO 1 LOOP
         inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
         result := result OR inputsx(olenM1 DOWNTO 0);
       END LOOP;
     END IF;
     RETURN result;
   END;

   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result XOR inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

-----------------------------------------------------------------
-- Muxes
-----------------------------------------------------------------
   
   FUNCTION mux_sel2_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(1 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 4;
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector( size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "01" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "10" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "11" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel3_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(2 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 8;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "001" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "010" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "011" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN "100" =>
       result := inputs0(5*size-1 DOWNTO 4*size);
     WHEN "101" =>
       result := inputs0(6*size-1 DOWNTO 5*size);
     WHEN "110" =>
       result := inputs0(7*size-1 DOWNTO 6*size);
     WHEN "111" =>
       result := inputs0(8*size-1 DOWNTO 7*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel4_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(3 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 16;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "0000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "0001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "0010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "0011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "0100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "0101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "0110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "0111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "1000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "1001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "1010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "1011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "1100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "1101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "1110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "1111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel5_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(4 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 32;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0 );
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "00001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "00010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "00011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "00100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "00101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "00110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "00111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "01000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "01001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "01010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "01011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "01100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "01101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "01110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "01111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "10000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "10001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "10010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "10011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "10100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "10101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "10110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "10111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "11000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "11001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "11010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "11011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "11100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "11101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "11110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "11111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel6_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(5 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 64;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "000001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "000010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "000011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "000100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "000101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "000110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "000111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "001000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "001001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "001010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "001011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "001100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "001101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "001110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "001111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "010000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "010001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "010010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "010011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "010100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "010101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "010110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "010111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "011000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "011001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "011010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "011011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "011100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "011101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "011110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "011111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN "100000" =>
       result := inputs0( 33*size-1 DOWNTO 32*size);
     WHEN "100001" =>
       result := inputs0( 34*size-1 DOWNTO 33*size);
     WHEN "100010" =>
       result := inputs0( 35*size-1 DOWNTO 34*size);
     WHEN "100011" =>
       result := inputs0( 36*size-1 DOWNTO 35*size);
     WHEN "100100" =>
       result := inputs0( 37*size-1 DOWNTO 36*size);
     WHEN "100101" =>
       result := inputs0( 38*size-1 DOWNTO 37*size);
     WHEN "100110" =>
       result := inputs0( 39*size-1 DOWNTO 38*size);
     WHEN "100111" =>
       result := inputs0( 40*size-1 DOWNTO 39*size);
     WHEN "101000" =>
       result := inputs0( 41*size-1 DOWNTO 40*size);
     WHEN "101001" =>
       result := inputs0( 42*size-1 DOWNTO 41*size);
     WHEN "101010" =>
       result := inputs0( 43*size-1 DOWNTO 42*size);
     WHEN "101011" =>
       result := inputs0( 44*size-1 DOWNTO 43*size);
     WHEN "101100" =>
       result := inputs0( 45*size-1 DOWNTO 44*size);
     WHEN "101101" =>
       result := inputs0( 46*size-1 DOWNTO 45*size);
     WHEN "101110" =>
       result := inputs0( 47*size-1 DOWNTO 46*size);
     WHEN "101111" =>
       result := inputs0( 48*size-1 DOWNTO 47*size);
     WHEN "110000" =>
       result := inputs0( 49*size-1 DOWNTO 48*size);
     WHEN "110001" =>
       result := inputs0( 50*size-1 DOWNTO 49*size);
     WHEN "110010" =>
       result := inputs0( 51*size-1 DOWNTO 50*size);
     WHEN "110011" =>
       result := inputs0( 52*size-1 DOWNTO 51*size);
     WHEN "110100" =>
       result := inputs0( 53*size-1 DOWNTO 52*size);
     WHEN "110101" =>
       result := inputs0( 54*size-1 DOWNTO 53*size);
     WHEN "110110" =>
       result := inputs0( 55*size-1 DOWNTO 54*size);
     WHEN "110111" =>
       result := inputs0( 56*size-1 DOWNTO 55*size);
     WHEN "111000" =>
       result := inputs0( 57*size-1 DOWNTO 56*size);
     WHEN "111001" =>
       result := inputs0( 58*size-1 DOWNTO 57*size);
     WHEN "111010" =>
       result := inputs0( 59*size-1 DOWNTO 58*size);
     WHEN "111011" =>
       result := inputs0( 60*size-1 DOWNTO 59*size);
     WHEN "111100" =>
       result := inputs0( 61*size-1 DOWNTO 60*size);
     WHEN "111101" =>
       result := inputs0( 62*size-1 DOWNTO 61*size);
     WHEN "111110" =>
       result := inputs0( 63*size-1 DOWNTO 62*size);
     WHEN "111111" =>
       result := inputs0( 64*size-1 DOWNTO 63*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS  --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2 SEVERITY FAILURE;
     --synopsys translate_on
       CASE sel IS
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0( size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1  DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0(size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
       RETURN result;
   END;
--   BEGIN RETURN mux_v(inputs, TO_STDLOGICVECTOR(sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     ALIAS    sel0   : STD_LOGIC_VECTOR( sel'LENGTH-1 DOWNTO 0 ) IS sel;

     VARIABLE sellen : INTEGER RANGE 2-sel'LENGTH TO sel'LENGTH;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2**sel'LENGTH;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
     TYPE inputs_array_type is array(natural range <>) of std_logic_vector( olen - 1 DOWNTO 0);
     VARIABLE inputs_array : inputs_array_type( 2**sel'LENGTH - 1 DOWNTO 0);
   BEGIN
     sellen := sel'LENGTH;
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2**sellen SEVERITY FAILURE;
     sellen := 2-sellen;
     --synopsys translate_on
     CASE sellen IS
     WHEN 1 =>
       CASE sel0(0) IS

       WHEN '1' 
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0(  size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1 DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0( size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
     WHEN 2 =>
       result := mux_sel2_v(inputs, not sel);
     WHEN 3 =>
       result := mux_sel3_v(inputs, not sel);
     WHEN 4 =>
       result := mux_sel4_v(inputs, not sel);
     WHEN 5 =>
       result := mux_sel5_v(inputs, not sel);
     WHEN 6 =>
       result := mux_sel6_v(inputs, not sel);
     WHEN others =>
       -- synopsys translate_off
       IF(Is_X(sel0)) THEN
         result := (others => 'X');
       ELSE
       -- synopsys translate_on
         FOR i in 0 to 2**sel'LENGTH - 1 LOOP
           inputs_array(i) := inputs0( ((i + 1) * olen) - 1  DOWNTO i*olen);
         END LOOP;
         result := inputs_array(CONV_INTEGER( (UNSIGNED(NOT sel0)) ));
       -- synopsys translate_off
       END IF;
       -- synopsys translate_on
     END CASE;
     RETURN result;
   END;

 
-----------------------------------------------------------------
-- Latches
-----------------------------------------------------------------

   FUNCTION lat_s(dinput: STD_LOGIC; clk: STD_LOGIC; doutput: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN mux_s(STD_LOGIC_VECTOR'(doutput & dinput), clk); END;

   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR ; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR ) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     --synopsys translate_off
     ASSERT dinput'LENGTH = doutput'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN mux_v(doutput & dinput, clk);
   END;

-----------------------------------------------------------------
-- Tri-States
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC; control: STD_LOGIC) RETURN STD_LOGIC IS
--   BEGIN RETURN TO_STDLOGIC(tri_v(TO_STDLOGICVECTOR(dinput), control)); END;
--
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR ; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
--     VARIABLE result: STD_LOGIC_VECTOR(dinput'range);
--   BEGIN
--     CASE control IS
--     WHEN '0' | 'L' =>
--       result := (others => 'Z');
--     WHEN '1' | 'H' =>
--       FOR i IN dinput'range LOOP
--         result(i) := to_UX01(dinput(i));
--       END LOOP;
--     WHEN others =>
--       -- synopsys translate_off
--       result := (others => 'X');
--       -- synopsys translate_on
--     END CASE;
--     RETURN result;
--   END;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;

   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     VARIABLE diff: UNSIGNED(l'LENGTH DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     diff := ('0'&l) - ('0'&r);
     RETURN diff(l'LENGTH);
   END;
   FUNCTION "<"(l, r: SIGNED  ) RETURN STD_LOGIC IS
   BEGIN
     RETURN (UNSIGNED(l) < UNSIGNED(r)) xor (l(l'LEFT) xor r(r'LEFT));
   END;

   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION "<=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">"(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;
   FUNCTION ">=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;

   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN not or_s(l xor r);
   END;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   --some functions to placate spyglass
   FUNCTION mult_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a*b;
   END mult_natural;

   FUNCTION div_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a/b;
   END div_natural;

   FUNCTION mod_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a mod b;
   END mod_natural;

   FUNCTION add_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a+b;
   END add_unsigned;

   FUNCTION sub_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a-b;
   END sub_unsigned;

   FUNCTION sub_int(a,b : INTEGER) RETURN INTEGER IS
   BEGIN
     return a-b;
   END sub_int;

   FUNCTION concat_0(b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return '0' & b;
   END concat_0;

   FUNCTION concat_uns(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a&b;
   END concat_uns;

   FUNCTION concat_vect(a,b : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     return a&b;
   END concat_vect;





   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED IS
     CONSTANT ninps : NATURAL := arg'LENGTH / width;
     ALIAS    arg0  : UNSIGNED(arg'LENGTH-1 DOWNTO 0) IS arg;
     VARIABLE result: UNSIGNED(width-1 DOWNTO 0);
     VARIABLE from  : INTEGER;
     VARIABLE dto   : INTEGER;
   BEGIN
     --synopsys translate_off
     ASSERT arg'LENGTH = width * ninps SEVERITY FAILURE;
     --synopsys translate_on
     result := (OTHERS => '0');
     FOR i IN ninps-1 DOWNTO 0 LOOP
       --result := result + arg0((i+1)*width-1 DOWNTO i*width);
       from := mult_natural((i+1), width)-1; --2.1.6.3
       dto  := mult_natural(i,width); --2.1.6.3
       result := add_unsigned(result , arg0(from DOWNTO dto) );
     END LOOP;
     RETURN result;
   END faccu;

   FUNCTION  fabs (arg1: SIGNED) RETURN UNSIGNED IS
   BEGIN
     CASE arg1(arg1'LEFT) IS
     WHEN '1'
     --synopsys translate_off
          | 'H'
     --synopsys translate_on
       =>
       RETURN UNSIGNED'("0") - UNSIGNED(arg1);
     WHEN '0'
     --synopsys translate_off
          | 'L'
     --synopsys translate_on
       =>
       RETURN UNSIGNED(arg1);
     WHEN others =>
       RETURN resolve_unsigned(UNSIGNED(arg1), UNSIGNED'("0") - UNSIGNED(arg1));
     END CASE;
   END;

   PROCEDURE divmod(l, r: UNSIGNED; rdiv, rmod: OUT UNSIGNED) IS
     CONSTANT llen: INTEGER := l'LENGTH;
     CONSTANT rlen: INTEGER := r'LENGTH;
     CONSTANT llen_plus_rlen: INTEGER := llen + rlen;
     VARIABLE lbuf: UNSIGNED(llen+rlen-1 DOWNTO 0);
     VARIABLE diff: UNSIGNED(rlen DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT rdiv'LENGTH = llen AND rmod'LENGTH = rlen SEVERITY FAILURE;
     --synopsys translate_on
     lbuf := (others => '0');
     lbuf(llen-1 DOWNTO 0) := l;
     FOR i IN rdiv'range LOOP
       diff := sub_unsigned(lbuf(llen_plus_rlen-1 DOWNTO llen-1) ,(concat_0(r)));
       rdiv(i) := not diff(rlen);
       IF diff(rlen) = '0' THEN
         lbuf(llen_plus_rlen-1 DOWNTO llen-1) := diff;
       END IF;
       lbuf(llen_plus_rlen-1 DOWNTO 1) := lbuf(llen_plus_rlen-2 DOWNTO 0);
     END LOOP;
     rmod := lbuf(llen_plus_rlen-1 DOWNTO llen);
   END divmod;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rdiv;
   END "/";

   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rmod;
   END;

   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN l MOD r; END;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rdiv := UNSIGNED'("0") - rdiv;
     END IF;
     RETURN SIGNED(rdiv); -- overflow problem "1000" / "11"
   END "/";

   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
     CONSTANT rnul: UNSIGNED(r'LENGTH-1 DOWNTO 0) := (others => '0');
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     IF rmod /= rnul AND to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rmod := UNSIGNED(r) + rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "MOD";

   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "REM";

   FUNCTION mult_unsigned(l,r : UNSIGNED) return UNSIGNED is
   BEGIN
     return l*r; 
   END mult_unsigned;

   FUNCTION "**" (l, r : UNSIGNED) RETURN UNSIGNED IS
     CONSTANT llen  : NATURAL := l'LENGTH;
     VARIABLE result: UNSIGNED(llen-1 DOWNTO 0);
     VARIABLE fak   : UNSIGNED(llen-1 DOWNTO 0);
   BEGIN
     fak := l;
     result := (others => '0'); result(0) := '1';
     FOR i IN r'reverse_range LOOP
       --was:result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(result & (result*fak)), r(i)));
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR( concat_uns(result , mult_unsigned(result,fak) )), r(i)));

       fak := mult_unsigned(fak , fak);
     END LOOP;
     RETURN result;
   END "**";

   FUNCTION "**" (l, r : SIGNED) RETURN SIGNED IS
     CONSTANT rlen  : NATURAL := r'LENGTH;
     ALIAS    r0    : SIGNED(0 TO r'LENGTH-1) IS r;
     VARIABLE result: SIGNED(l'range);
   BEGIN
     CASE r(r'LEFT) IS
     WHEN '0'
   --synopsys translate_off
          | 'L'
   --synopsys translate_on
     =>
       result := SIGNED(UNSIGNED(l) ** UNSIGNED(r0(1 TO r'LENGTH-1)));
     WHEN '1'
   --synopsys translate_off
          | 'H'
   --synopsys translate_on
     =>
       result := (others => '0');
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END "**";

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-----------------------------------------------------------------

   FUNCTION add_nat(arg1 : NATURAL; arg2 : NATURAL ) RETURN NATURAL IS
   BEGIN
     return (arg1 + arg2);
   END;
   
--   FUNCTION UNSIGNED_2_BIT_VECTOR(arg1 : NATURAL; arg2 : NATURAL ) RETURN BIT_VECTOR IS
--   BEGIN
--     return (arg1 + arg2);
--   END;
   
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(SIGNED(result), arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
        =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
        =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;


   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     --SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: NATURAL range 1 TO len;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => '0');
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         --was:temp(i2+sw) := result(i2);
         temp_idx := add_nat(i2,sw);
         temp(temp_idx) := result(i2);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: sw_range;
     VARIABLE result_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => sbit);
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         -- was: temp(i2) := result(i2+sw);
         result_idx := add_nat(i2,sw);
         temp(i2) := result(result_idx);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;


   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := arg1'LENGTH;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     VARIABLE temp: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     SUBTYPE sw_range IS NATURAL range 0 TO len-1;
     VARIABLE sw: sw_range;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     result := (others=>'0');
     result := arg1;
     sw := sdir MOD len;
     FOR i IN arg2'reverse_range LOOP
       EXIT WHEN sw = 0;
       IF signd2 AND i = arg2'LEFT THEN 
         sw := sub_int(len,sw); 
       END IF;
       -- temp := result(len-sw-1 DOWNTO 0) & result(len-1 DOWNTO len-sw)
       FOR i2 IN len-1 DOWNTO 0 LOOP
         --was: temp((i2+sw) MOD len) := result(i2);
         temp_idx := add_nat(i2,sw) MOD len;
         temp(temp_idx) := result(i2);
       END LOOP;
       result := mux_v(STD_LOGIC_VECTOR(concat_vect(result,temp)), arg2(i));
       sw := mod_natural(mult_natural(sw,2), len);
     END LOOP;
     RETURN result;
   END frot;

   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, -1); END;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, -1); END;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC IS
     CONSTANT len : INTEGER := vec'LENGTH;
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
   BEGIN
     IF index >= len OR index < 0 THEN
       RETURN 'X';
     END IF;
     RETURN vec0(index);
   END;

   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     CONSTANT indexPwidthM1 : INTEGER := index+width-1; --2.1.6.3
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
     CONSTANT xxx : STD_LOGIC_VECTOR(width-1 DOWNTO 0) := (others => 'X');
   BEGIN
     IF index+width > len OR index < 0 THEN
       RETURN xxx;
     END IF;
     RETURN vec0(indexPwidthM1 DOWNTO index);
   END;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     VARIABLE vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     CONSTANT xxx : STD_LOGIC_VECTOR(len-1 DOWNTO 0) := (others => 'X');
   BEGIN
     vec0 := vec;
     IF index >= len OR index < 0 THEN
       RETURN xxx;
     END IF;
     vec0(index) := dinput;
     RETURN vec0;
   END;

   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE IS
     VARIABLE n_b : POSITIVE;
     VARIABLE p_v : NATURAL;
   BEGIN
     p_v := p;
     FOR i IN 1 TO 32 LOOP
       p_v := div_natural(p_v,2);
       n_b := i;
       EXIT WHEN (p_v = 0);
     END LOOP;
     RETURN n_b;
   END;


--   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
--
--     CONSTANT vlen: INTEGER := vec'LENGTH;
--     CONSTANT ilen: INTEGER := dinput'LENGTH;
--     CONSTANT max_shift: INTEGER := vlen-ilen;
--     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
--     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
--     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
--     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
--     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
--     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
--   BEGIN
--     inp := (others => '0');
--     mask := (others => '0');
--
--     IF index > max_shift OR index < 0 THEN
--       RETURN xxx;
--     END IF;
--
--     shift := CONV_UNSIGNED(index, shift'LENGTH);
--     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
--     mask(ilen-1 DOWNTO 0) := ones;
--     inp := fshl(inp, shift, vlen);
--     mask := fshl(mask, shift, vlen);
--     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
--     RETURN vec0;
--   END;

   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR IS

     type enable_matrix is array (0 to enable'LENGTH-1 ) of std_logic_vector(byte_width-1 downto 0);
     CONSTANT vlen: INTEGER := vec'LENGTH;
     CONSTANT ilen: INTEGER := dinput'LENGTH;
     CONSTANT max_shift: INTEGER := vlen-ilen;
     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask2: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE enables: enable_matrix;
     VARIABLE cat_enables: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0 );
     VARIABLE lsbi : INTEGER;
     VARIABLE msbi : INTEGER;

   BEGIN
     cat_enables := (others => '0');
     lsbi := 0;
     msbi := byte_width-1;
     inp := (others => '0');
     mask := (others => '0');

     IF index > max_shift OR index < 0 THEN
       RETURN xxx;
     END IF;

     --initialize enables
     for i in 0 TO (enable'LENGTH-1) loop
       enables(i)  := (others => enable(i));
       cat_enables(msbi downto lsbi) := enables(i) ;
       lsbi := msbi+1;
       msbi := msbi+byte_width;
     end loop;


     shift := CONV_UNSIGNED(index, shift'LENGTH);
     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
     mask(ilen-1 DOWNTO 0) := UNSIGNED((STD_LOGIC_VECTOR(ones) AND cat_enables));
     inp := fshl(inp, shift, vlen);
     mask := fshl(mask, shift, vlen);
     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
     RETURN vec0;
   END;


   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;
   
   FUNCTION bits(size : NATURAL) return NATURAL is
   begin
     return ceil_log2(size);
   END;

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH) xor conv_std_logic_vector(c, s'LENGTH);
     cout := ( (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH)) or (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) or (conv_std_logic_vector(b, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) );
   END PROCEDURE csa;

   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH);
     cout := (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH));
   END PROCEDURE csha;

END funcs;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_comps.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_comps IS
 
FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
FUNCTION ceil_log2(size : NATURAL) return NATURAL;
 

COMPONENT mgc_not
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_and
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nand
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_or
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xnor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux
  GENERIC (
    width  :  NATURAL;
    ctrlw  :  NATURAL;
    p2ctrlw : NATURAL := 0
  );
  PORT (
    a: in  std_logic_vector(width*(2**ctrlw) - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw            - 1 DOWNTO 0);
    z: out std_logic_vector(width            - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux1hot
  GENERIC (
    width  : NATURAL;
    ctrlw  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ctrlw - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw       - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_reg_pos
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;  -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL  -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_reg_neg
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;   -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_generic_reg
  GENERIC(
   width: natural := 8;
   ph_clk: integer range 0 to 1 := 1; -- clock polarity, 1=rising_edge
   ph_en: integer range 0 to 1 := 1;
   ph_a_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   ph_s_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   a_rst_used: integer range 0 to 1 := 1;
   s_rst_used: integer range 0 to 1 := 0;
   en_used: integer range 0 to 1 := 1
  );
  PORT(
   d: std_logic_vector(width-1 downto 0);
   clk: in std_logic;
   en: in std_logic;
   a_rst: in std_logic;
   s_rst: in std_logic;
   q: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_equal
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a : in  std_logic_vector(width-1 DOWNTO 0);
    b : in  std_logic_vector(width-1 DOWNTO 0);
    eq: out std_logic;
    ne: out std_logic
  );
END COMPONENT;

COMPONENT mgc_shift_l
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rot
  GENERIC (
    width  : NATURAL;
    width_s: NATURAL;
    signd_s: NATURAL;      -- 0:unsigned 1:signed
    sleft  : NATURAL;      -- 0:right 1:left;
    log2w  : NATURAL := 0; -- LOG2(width)
    l2wp2  : NATURAL := 0  --2**LOG2(width)
  );
  PORT (
    a : in  std_logic_vector(width  -1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width  -1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_sub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_ci
  GENERIC (
    width_a : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width_a, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width_a, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width_a,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width_a,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_addc
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add3
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_c : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_c : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(ifeqsel(width_c,0,width,width_c)-1 DOWNTO 0);
    d: in  std_logic_vector(0 DOWNTO 0);
    e: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_sub_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addc_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     c: in std_logic_vector(0 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addsub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    add: in  std_logic;
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_accu
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_abs
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_fast
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_pipe
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2  : NATURAL;
    add_d2  : NATURAL
  );
  PORT (
    a   : in  std_logic_vector(width_a-1 DOWNTO 0);
    b   : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2  : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c   : in  std_logic_vector(width_c-1 DOWNTO 0);
    d   : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2  : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst : in  std_logic_vector(width_e-1 DOWNTO 0);
    z   : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1_pipe
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2   : NATURAL;
    add_d2   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2     : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2     : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_e-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL
  );
  PORT (
    a:   in  std_logic_vector(width_a-1 DOWNTO 0);
    b:   in  std_logic_vector(width_b-1 DOWNTO 0);
    c:   in  std_logic_vector(width_c-1 DOWNTO 0);
    cst: in  std_logic_vector(width_cst-1 DOWNTO 0);
    d:   in  std_logic_vector(width_d-1 DOWNTO 0);
    z:   out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1_pipe
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_cst-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mulacc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2acc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    add_cxd : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    d         : in  std_logic_vector(width_d-1 DOWNTO 0);
    e         : in  std_logic_vector(width_e-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_div
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mod
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rem
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_csa
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     c: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_csha
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_rom
    GENERIC (
      rom_id : natural := 1;
      size : natural := 33;
      width : natural := 32
      );
    PORT (
      data_in : std_logic_vector((size*width)-1 downto 0);
      addr : std_logic_vector(ceil_log2(size)-1 downto 0);
      data_out : out std_logic_vector(width-1 downto 0)
    );
END COMPONENT;

END mgc_comps;

PACKAGE BODY mgc_comps IS
 
   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;
 
END mgc_comps;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_mul_pipe IS
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_mul_pipe;

LIBRARY IEEE;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_mul_pipe IS
  TYPE reg_array_type is array(natural range<>) of std_logic_vector(width_z-1 DOWNTO 0); 
  SIGNAL xz : std_logic_vector(width_a+width_b DOWNTO 0);

--MF Added pipelined input
    signal a_f     : STD_LOGIC_VECTOR(width_a-1 downto 0); 
    signal b_f     : STD_LOGIC_VECTOR(width_b-1 downto 0);
   type a_array is array (natural range <>) of STD_LOGIC_VECTOR(width_a-1 downto 0);
   type b_array is array (natural range <>) of STD_LOGIC_VECTOR(width_b-1 downto 0);
BEGIN
  n_inreg_gt_0: if n_inreg > 0 generate
    GENPOS_INREG: IF clock_edge = 1 GENERATE
     I0: process(clk)
        variable a_in_reg: a_array(n_inreg-1 downto 0);
        variable b_in_reg: b_array(n_inreg-1 downto 0);
      begin
        if (clk'event and clk = '1' ) then
          if (conv_integer(en) = enable_active) then
            for i in n_inreg - 2 downto 0 loop
              a_in_reg(i+1) := a_in_reg(i);
              b_in_reg(i+1) := b_in_reg(i);
            end loop;                                                                                                                             
            a_in_reg(0) := a;
            b_in_reg(0) := b;

            a_f <= a_in_reg(n_inreg-1);             
            b_f <= b_in_reg(n_inreg-1);    
                                                   
          end if;
        end if;
      end process;
    END GENERATE;
  
   GENNEG_INREG: IF clock_edge = 0 GENERATE
     I0: process(clk)
        variable a_in_reg: a_array(n_inreg-1 downto 0);
        variable b_in_reg: b_array(n_inreg-1 downto 0);
      begin
        if (clk'event and clk = '0' ) then
          if (conv_integer(en) = enable_active) then
            for i in n_inreg - 2 downto 0 loop
              a_in_reg(i+1) := a_in_reg(i);
              b_in_reg(i+1) := b_in_reg(i);
            end loop;                                                                                                                             
            a_in_reg(0) := a;
            b_in_reg(0) := b;            
                                 
            a_f <= a_in_reg(n_inreg-1);             
            b_f <= b_in_reg(n_inreg-1);
                                                        
          end if;
        end if;
      end process;
    END GENERATE;
  END GENERATE;

  n_inreg_eq_0: if n_inreg = 0 generate
    a_f <= a;
    b_f <= b;
  end generate n_inreg_eq_0;

  xz <= '0'&(unsigned(a_f) * unsigned(b_f)) WHEN signd_a = 0 AND signd_b = 0 ELSE
            (  signed(a_f) * unsigned(b_f)) WHEN signd_a = 1 AND signd_b = 0 ELSE
            (unsigned(a_f) *   signed(b_f)) WHEN signd_a = 0 AND signd_b = 1 ELSE
        '0'&(  signed(a_f) *   signed(b_f));

  GENPOS: IF clock_edge = 1 GENERATE
    PROCESS (clk)
    VARIABLE reg_array: reg_array_type(stages-2 DOWNTO 0);
    BEGIN
      IF ( clk'EVENT AND clk = '1') THEN
        IF ( conv_integer(en) = enable_active) THEN
          FOR I IN stages-2 DOWNTO 1 LOOP
            reg_array(I) := reg_array(I-1);
          END LOOP;
          reg_array(0) := xz(width_z-1 DOWNTO 0);
          z <= reg_array(stages-2);
        END IF;
      END IF;
    END PROCESS;
  END GENERATE;

  GENNEG: IF clock_edge = 0 GENERATE
    PROCESS (clk)
    VARIABLE reg_array: reg_array_type(stages-2 DOWNTO 0);
    BEGIN
      IF ( clk'EVENT AND clk = '0') THEN
        IF ( conv_integer(en) = enable_active) THEN
          FOR I IN stages-2 DOWNTO 1 LOOP
            reg_array(I) := reg_array(I-1);
          END LOOP;
          reg_array(0) := xz(width_z-1 DOWNTO 0);
          z <= reg_array(stages-2);
        END IF;
      END IF;
    END PROCESS;
  END GENERATE;
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_comps_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_shift_comps_v5 IS

COMPONENT mgc_shift_l_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_shift_comps_v5;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_bl_beh_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_shift_bl_v5 IS
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_shift_bl_v5;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_shift_bl_v5 IS

  FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
    CONSTANT len: INTEGER := input1'LENGTH;
    ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
    ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
    VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
  BEGIN
    result := (others => '0');
    --synopsys translate_off
    FOR i IN len-1 DOWNTO 0 LOOP
      result(i) := resolved(input1a(i) & input2a(i));
    END LOOP;
    --synopsys translate_on
    RETURN result;
  END;

  FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED)
  RETURN UNSIGNED IS
  BEGIN
    RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1),
                                             STD_LOGIC_VECTOR(input2)));
  END;

  FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED)
  RETURN SIGNED IS
  BEGIN
    RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1),
                                           STD_LOGIC_VECTOR(input2)));
  END;

  FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
    BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;

  FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1 > arg2) THEN
      RETURN(arg1) ;
    ELSE
      RETURN(arg2) ;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shr(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(SIGNED(result), arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shr(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

 FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
    ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
    CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
    ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
    VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
    VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
  BEGIN
    result := (others=>'0');
    arg1x_pad(arg1l+1) := sbit;
    arg1x_pad(arg1l downto 0) := arg1x;
    IF arg2l = 0 THEN
      RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
    -- ELSIF arg1l = 0 THEN
    --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
    ELSE
      CASE arg2x(arg2l) IS
      WHEN '0'
    --synopsys translate_off
           | 'L'
    --synopsys translate_on
      =>
        RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
      WHEN '1'
    --synopsys translate_off
           | 'H'
    --synopsys translate_on
      =>
        RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
      WHEN others =>
        --synopsys translate_off
        result := resolve_unsigned(
          fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
          fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
        );
        --synopsys translate_on
        RETURN result;
      END CASE;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
    ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
    CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
    ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
    VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
    VARIABLE result: SIGNED(olen-1 DOWNTO 0);
  BEGIN
    result := (others=>'0');
    arg1x_pad(arg1l+1) := sbit;
    arg1x_pad(arg1l downto 0) := arg1x;
    IF arg2l = 0 THEN
      RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
    -- ELSIF arg1l = 0 THEN
    --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
    ELSE
      CASE arg2x(arg2l) IS
      WHEN '0'
      --synopsys translate_off
           | 'L'
      --synopsys translate_on
      =>
        RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
      WHEN '1'
      --synopsys translate_off
           | 'H'
      --synopsys translate_on
      =>
        RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
      WHEN others =>
        --synopsys translate_off
        result := resolve_signed(
          fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
          fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
        );
        --synopsys translate_on
        RETURN result;
      END CASE;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE)
  RETURN UNSIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, '0', olen);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE)
  RETURN SIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen);
  END;

BEGIN
UNSGNED:  IF signd_a = 0 GENERATE
    z <= std_logic_vector(fshl_stdar(unsigned(a), signed(s), width_z));
  END GENERATE;
SGNED:  IF signd_a /= 0 GENERATE
    z <= std_logic_vector(fshl_stdar(  signed(a), signed(s), width_z));
  END GENERATE;
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_shift_l_v5 IS
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_shift_l_v5;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_shift_l_v5 IS

  FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1 > arg2) THEN
      RETURN(arg1) ;
    ELSE
      RETURN(arg2) ;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(SIGNED(result), arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE)
  RETURN UNSIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, '0', olen);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE)
  RETURN SIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen);
  END;

BEGIN
UNSGNED:  IF signd_a = 0 GENERATE
    z <= std_logic_vector(fshl_stdar(unsigned(a), unsigned(s), width_z));
  END GENERATE;
SGNED:  IF signd_a /= 0 GENERATE
    z <= std_logic_vector(fshl_stdar(  signed(a), unsigned(s), width_z));
  END GENERATE;
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_DPRAM_RBW_DUAL.vhd 
-- Memory Type:            BLOCK
-- Operating Mode:         True Dual Port (2-Port)
-- Clock Mode:             Dual Clock
-- 
-- RTL Code RW Resolution: RBW
-- Catapult RW Resolution: RBW
-- 
-- HDL Work Library:       Xilinx_RAMS_lib
-- Component Name:         BLOCK_DPRAM_RBW_DUAL
-- Latency = 1:            RAM with no registers on inputs or outputs
--         = 2:            adds embedded register on RAM output
--         = 3:            adds fabric registers to non-clock input RAM pins
--         = 4:            adds fabric register to output (driven by embedded register from latency=2)

LIBRARY ieee;

  USE ieee.std_logic_1164.all;
  USE ieee.numeric_std.all;
PACKAGE BLOCK_DPRAM_RBW_DUAL_pkg IS
  COMPONENT BLOCK_DPRAM_RBW_DUAL IS
  GENERIC (
    addr_width : integer := 8 ;
    data_width : integer := 7 ;
    depth : integer := 256 ;
    latency : integer := 1 
    
  );
  PORT (
    adra : in std_logic_vector(addr_width-1 downto 0) ;
    adrb : in std_logic_vector(addr_width-1 downto 0) ;
    clka : in std_logic ;
    clka_en : in std_logic ;
    clkb : in std_logic ;
    clkb_en : in std_logic ;
    da : in std_logic_vector(data_width-1 downto 0) ;
    db : in std_logic_vector(data_width-1 downto 0) ;
    qa : out std_logic_vector(data_width-1 downto 0) ;
    qb : out std_logic_vector(data_width-1 downto 0) ;
    wea : in std_logic ;
    web : in std_logic 
    
  );
  END COMPONENT;
END BLOCK_DPRAM_RBW_DUAL_pkg;
LIBRARY ieee;

  USE ieee.std_logic_1164.all;
  USE ieee.numeric_std.all;
ENTITY BLOCK_DPRAM_RBW_DUAL IS
  GENERIC (
    addr_width : integer := 8 ;
    data_width : integer := 7 ;
    depth : integer := 256 ;
    latency : integer := 1 
    
  );
  PORT (
    adra : in std_logic_vector(addr_width-1 downto 0) ;
    adrb : in std_logic_vector(addr_width-1 downto 0) ;
    clka : in std_logic ;
    clka_en : in std_logic ;
    clkb : in std_logic ;
    clkb_en : in std_logic ;
    da : in std_logic_vector(data_width-1 downto 0) ;
    db : in std_logic_vector(data_width-1 downto 0) ;
    qa : out std_logic_vector(data_width-1 downto 0) ;
    qb : out std_logic_vector(data_width-1 downto 0) ;
    wea : in std_logic ;
    web : in std_logic 
    
  );
 END BLOCK_DPRAM_RBW_DUAL;
ARCHITECTURE rtl OF BLOCK_DPRAM_RBW_DUAL IS
  TYPE ram_t IS ARRAY (depth-1 DOWNTO 0) OF std_logic_vector(data_width-1 DOWNTO 0);
  SHARED VARIABLE mem : ram_t := (OTHERS => (OTHERS => '0'));
  ATTRIBUTE ram_style: STRING;
  ATTRIBUTE ram_style OF mem : VARIABLE IS "block";
  ATTRIBUTE syn_ramstyle: STRING;
  ATTRIBUTE syn_ramstyle OF mem : VARIABLE IS "block";
  
  SIGNAL ramqa : std_logic_vector(data_width-1 downto 0);
  SIGNAL ramqb : std_logic_vector(data_width-1 downto 0);
  
BEGIN
-- Port Map
-- rwA :: ADDRESS adra CLOCK clka ENABLE clka_en DATA_IN da DATA_OUT qa WRITE_ENABLE wea
-- rwB :: ADDRESS adrb CLOCK clkb ENABLE clkb_en DATA_IN db DATA_OUT qb WRITE_ENABLE web

-- Access memory with non-registered inputs (latency = 1||2)
  IN_PIN :  IF latency < 3 GENERATE
  BEGIN
    PROCESS (clka)
    BEGIN
      IF (rising_edge(clka)) THEN
         IF (clka_en = '1') THEN
          -- workaround for simulation when read address out-of-range during inactive cycle
          --pragma translate_off
          IF (to_integer(unsigned(adra)) < depth) THEN
          --pragma translate_on
          ramqa <= mem(to_integer(unsigned(adra)));
          --pragma translate_off
          END IF;
          --pragma translate_on
          IF (wea = '1') THEN
            mem(to_integer(unsigned(adra))) := da;
          END IF;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clka)
    BEGIN
      IF (rising_edge(clka)) THEN
         IF (clka_en = '1') THEN
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkb)
    BEGIN
      IF (rising_edge(clkb)) THEN
         IF (clkb_en = '1') THEN
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkb)
    BEGIN
      IF (rising_edge(clkb)) THEN
         IF (clkb_en = '1') THEN
          -- workaround for simulation when read address out-of-range during inactive cycle
          --pragma translate_off
          IF (to_integer(unsigned(adrb)) < depth) THEN
          --pragma translate_on
          ramqb <= mem(to_integer(unsigned(adrb)));
          --pragma translate_off
          END IF;
          --pragma translate_on
          IF (web = '1') THEN
            mem(to_integer(unsigned(adrb))) := db;
          END IF;
        END IF;
      END IF;
    END PROCESS;
    
  END GENERATE IN_PIN; 

-- Register all non-clock inputs (latency = 3||4)
  IN_REG :  IF latency > 2 GENERATE
    SIGNAL adra_reg : std_logic_vector(addr_width-1 downto 0);
    SIGNAL da_reg : std_logic_vector(data_width-1 downto 0);
    SIGNAL wea_reg : std_logic;
    SIGNAL adrb_reg : std_logic_vector(addr_width-1 downto 0);
    SIGNAL db_reg : std_logic_vector(data_width-1 downto 0);
    SIGNAL web_reg : std_logic;
    
  BEGIN
    PROCESS (clka)
    BEGIN
      IF (rising_edge(clka)) THEN
        IF (clka_en = '1') THEN
          adra_reg <= adra;
          da_reg <= da;
          wea_reg <= wea;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkb)
    BEGIN
      IF (rising_edge(clkb)) THEN
        IF (clkb_en = '1') THEN
          adrb_reg <= adrb;
          db_reg <= db;
          web_reg <= web;
        END IF;
      END IF;
    END PROCESS;
    
    PROCESS (clka)
    BEGIN
      IF (rising_edge(clka)) THEN
         IF (clka_en = '1') THEN
          -- workaround for simulation when read address out-of-range during inactive cycle
          --pragma translate_off
          IF (to_integer(unsigned(adra_reg)) < depth) THEN
          --pragma translate_on
          ramqa <= mem(to_integer(unsigned(adra_reg)));
          --pragma translate_off
          END IF;
          --pragma translate_on
          IF (wea_reg = '1') THEN
            mem(to_integer(unsigned(adra_reg))) := da_reg;
          END IF;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clka)
    BEGIN
      IF (rising_edge(clka)) THEN
         IF (clka_en = '1') THEN
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkb)
    BEGIN
      IF (rising_edge(clkb)) THEN
         IF (clkb_en = '1') THEN
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkb)
    BEGIN
      IF (rising_edge(clkb)) THEN
         IF (clkb_en = '1') THEN
          -- workaround for simulation when read address out-of-range during inactive cycle
          --pragma translate_off
          IF (to_integer(unsigned(adrb_reg)) < depth) THEN
          --pragma translate_on
          ramqb <= mem(to_integer(unsigned(adrb_reg)));
          --pragma translate_off
          END IF;
          --pragma translate_on
          IF (web_reg = '1') THEN
            mem(to_integer(unsigned(adrb_reg))) := db_reg;
          END IF;
        END IF;
      END IF;
    END PROCESS;
    
  END GENERATE IN_REG;

  out_ram : IF latency = 1 GENERATE
  BEGIN
    qa <= ramqa;
    qb <= ramqb;
    
  END GENERATE out_ram;

  out_reg1 : IF ((latency = 2) OR (latency = 3)) GENERATE
    SIGNAL tmpqa : std_logic_vector(data_width-1 downto 0);
    SIGNAL tmpqb : std_logic_vector(data_width-1 downto 0);
    
  BEGIN
    PROCESS (clka)
    BEGIN
      IF (rising_edge(clka)) THEN
        IF (clka_en = '1') THEN
          tmpqa <= ramqa;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkb)
    BEGIN
      IF (rising_edge(clkb)) THEN
        IF (clkb_en = '1') THEN
          tmpqb <= ramqb;
        END IF;
      END IF;
    END PROCESS;
    
    qa <= tmpqa;
    qb <= tmpqb;
    
  END GENERATE out_reg1;

  out_reg2 : IF latency = 4 GENERATE
    SIGNAL tmp1qa : std_logic_vector(data_width-1 downto 0);
    SIGNAL tmp1qb : std_logic_vector(data_width-1 downto 0);
    
    SIGNAL tmp2qa : std_logic_vector(data_width-1 downto 0);
    SIGNAL tmp2qb : std_logic_vector(data_width-1 downto 0);
    
  BEGIN
    PROCESS (clka)
    BEGIN
      IF (rising_edge(clka)) THEN
        IF (clka_en = '1') THEN
          tmp1qa <= ramqa;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkb)
    BEGIN
      IF (rising_edge(clkb)) THEN
        IF (clkb_en = '1') THEN
          tmp1qb <= ramqb;
        END IF;
      END IF;
    END PROCESS;
    
    PROCESS (clka)
    BEGIN
      IF (rising_edge(clka)) THEN
        IF (clka_en = '1') THEN
          tmp2qa <= tmp1qa;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkb)
    BEGIN
      IF (rising_edge(clkb)) THEN
        IF (clkb_en = '1') THEN
          tmp2qb <= tmp1qb;
        END IF;
      END IF;
    END PROCESS;
    
    qa <= tmp2qa;
    qb <= tmp2qb;
    
  END GENERATE out_reg2;


END rtl;

--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Tue Sep 14 21:33:02 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_102_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_102_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_102_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_102_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_101_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_101_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_101_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_101_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_100_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_100_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_100_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_100_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_99_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_99_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_99_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_99_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_98_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_98_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_98_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_98_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_97_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_97_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_97_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_97_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_96_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_96_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_96_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_96_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_95_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_95_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_95_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_95_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_94_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_94_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_94_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_94_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_93_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_93_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_93_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_93_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_92_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_92_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_92_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_92_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_91_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_91_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_91_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_91_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_90_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_90_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_90_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_90_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_89_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_89_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_89_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_89_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_88_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_88_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_88_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_88_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_87_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_87_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_87_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_87_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_86_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_86_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_86_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_86_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_85_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_85_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_85_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_85_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_84_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_84_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_84_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_84_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_83_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_83_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_83_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_83_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_82_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_82_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_82_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_82_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_81_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_81_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_81_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_81_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_80_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_80_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_80_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_80_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_79_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_79_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_79_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_79_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_78_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_78_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_78_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_78_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_77_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_77_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_77_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_77_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_76_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_76_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_76_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_76_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_75_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_75_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_75_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_75_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_74_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_74_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_74_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_74_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_73_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_73_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_73_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_73_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_72_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_72_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_72_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_72_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_71_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_71_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_71_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_71_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_70_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_70_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_70_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_70_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_69_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_69_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_69_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_69_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_68_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_68_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_68_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_68_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_67_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_67_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_67_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_67_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_66_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_66_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_66_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_66_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_65_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_65_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_65_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_65_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_64_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_64_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_64_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_64_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_63_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_63_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_63_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_63_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_62_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_62_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_62_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_62_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_61_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_61_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_61_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_61_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_60_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_60_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_60_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_60_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_59_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_59_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_59_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_59_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_58_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_58_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_58_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_58_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_57_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_57_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_57_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_57_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_56_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_56_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_56_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_56_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_55_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_55_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_55_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_55_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_54_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_54_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_54_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_54_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_53_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_53_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_53_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_53_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_52_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_52_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_52_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_52_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_51_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_51_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_51_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_51_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_50_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_50_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_50_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_50_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_49_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_49_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_49_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_49_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_48_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_48_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_48_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_48_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_47_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_47_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_47_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_47_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_46_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_46_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_46_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_46_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_45_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_45_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_45_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_45_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_44_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_44_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_44_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_44_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_43_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_43_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_43_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_43_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_42_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_42_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_42_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_42_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_41_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_41_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_41_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_41_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_40_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_40_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_40_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_40_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_39_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_39_8_32_256_256_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_39_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_39_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_38_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_38_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_38_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_38_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_37_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_37_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_37_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_37_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_36_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_36_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_36_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_36_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_35_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_35_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_35_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_35_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_34_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_34_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_34_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_34_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_33_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_33_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_33_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_33_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_32_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_32_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_32_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_32_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_31_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_31_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_31_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_31_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_30_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_30_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_30_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_30_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_29_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_29_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_29_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_29_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_28_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_28_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_28_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_28_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_27_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_27_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_27_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_27_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_26_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_26_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_26_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_26_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_25_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_25_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_25_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_25_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_24_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_24_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_24_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_24_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_23_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_23_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_23_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_23_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_22_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_22_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_22_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_22_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_21_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_21_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_21_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_21_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_20_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_20_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_20_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_20_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_19_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_19_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_19_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_19_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_18_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_18_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_18_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_18_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_17_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_17_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_17_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_17_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_16_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_16_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_16_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_16_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_15_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_15_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_15_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_15_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_14_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_14_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_14_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_14_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_13_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_13_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_13_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_13_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_12_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_12_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_12_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_12_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_11_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_11_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_11_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_11_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_10_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_10_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_10_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_10_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_9_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_9_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_9_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_9_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_8_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_8_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_8_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_8_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_7_8_32_256_256_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_7_8_32_256_256_32_1_gen
    IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_7_8_32_256_256_32_1_gen;

ARCHITECTURE v11 OF peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_7_8_32_256_256_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(15 DOWNTO 8));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(7 DOWNTO 0));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    INNER_LOOP1_C_0_tr0 : IN STD_LOGIC;
    INNER_LOOP2_C_0_tr0 : IN STD_LOGIC;
    STAGE_LOOP_C_2_tr0 : IN STD_LOGIC;
    INNER_LOOP3_C_0_tr0 : IN STD_LOGIC;
    INNER_LOOP4_C_0_tr0 : IN STD_LOGIC;
    INNER_LOOP4_C_0_tr1 : IN STD_LOGIC
  );
END peaseNTT_core_core_fsm;

ARCHITECTURE v11 OF peaseNTT_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for peaseNTT_core_core_fsm_1
  TYPE peaseNTT_core_core_fsm_1_ST IS (main_C_0, STAGE_LOOP_C_0, INNER_LOOP1_C_0,
      STAGE_LOOP_C_1, INNER_LOOP2_C_0, STAGE_LOOP_C_2, STAGE_LOOP1_C_0, INNER_LOOP3_C_0,
      STAGE_LOOP1_C_1, INNER_LOOP4_C_0, main_C_1);

  SIGNAL state_var : peaseNTT_core_core_fsm_1_ST;
  SIGNAL state_var_NS : peaseNTT_core_core_fsm_1_ST;

BEGIN
  peaseNTT_core_core_fsm_1 : PROCESS (INNER_LOOP1_C_0_tr0, INNER_LOOP2_C_0_tr0, STAGE_LOOP_C_2_tr0,
      INNER_LOOP3_C_0_tr0, INNER_LOOP4_C_0_tr0, INNER_LOOP4_C_0_tr1, state_var)
  BEGIN
    CASE state_var IS
      WHEN STAGE_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000010");
        state_var_NS <= INNER_LOOP1_C_0;
      WHEN INNER_LOOP1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000100");
        IF ( INNER_LOOP1_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP_C_1;
        ELSE
          state_var_NS <= INNER_LOOP1_C_0;
        END IF;
      WHEN STAGE_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001000");
        state_var_NS <= INNER_LOOP2_C_0;
      WHEN INNER_LOOP2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010000");
        IF ( INNER_LOOP2_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP_C_2;
        ELSE
          state_var_NS <= INNER_LOOP2_C_0;
        END IF;
      WHEN STAGE_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100000");
        IF ( STAGE_LOOP_C_2_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP1_C_0;
        ELSE
          state_var_NS <= STAGE_LOOP_C_0;
        END IF;
      WHEN STAGE_LOOP1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000000");
        state_var_NS <= INNER_LOOP3_C_0;
      WHEN INNER_LOOP3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000000");
        IF ( INNER_LOOP3_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP1_C_1;
        ELSE
          state_var_NS <= INNER_LOOP3_C_0;
        END IF;
      WHEN STAGE_LOOP1_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000000");
        state_var_NS <= INNER_LOOP4_C_0;
      WHEN INNER_LOOP4_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000000");
        IF ( INNER_LOOP4_C_0_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSIF ( INNER_LOOP4_C_0_tr1 = '1' ) THEN
          state_var_NS <= INNER_LOOP4_C_0;
        ELSE
          state_var_NS <= STAGE_LOOP1_C_0;
        END IF;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000000");
        state_var_NS <= main_C_0;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000001");
        state_var_NS <= STAGE_LOOP_C_0;
    END CASE;
  END PROCESS peaseNTT_core_core_fsm_1;

  peaseNTT_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        state_var <= state_var_NS;
      END IF;
    END IF;
  END PROCESS peaseNTT_core_core_fsm_1_REG;

END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_core_wait_dp IS
  PORT(
    yt_rsc_0_0_cgo_iro : IN STD_LOGIC;
    yt_rsc_0_0_i_clka_en_d : OUT STD_LOGIC;
    yt_rsc_0_16_cgo_iro : IN STD_LOGIC;
    yt_rsc_0_16_i_clka_en_d : OUT STD_LOGIC;
    ensig_cgo_iro : IN STD_LOGIC;
    ensig_cgo_iro_17 : IN STD_LOGIC;
    yt_rsc_0_0_cgo : IN STD_LOGIC;
    yt_rsc_0_16_cgo : IN STD_LOGIC;
    ensig_cgo : IN STD_LOGIC;
    mult_t_mul_cmp_en : OUT STD_LOGIC;
    ensig_cgo_17 : IN STD_LOGIC;
    mult_z_mul_cmp_1_en : OUT STD_LOGIC
  );
END peaseNTT_core_wait_dp;

ARCHITECTURE v11 OF peaseNTT_core_wait_dp IS
  -- Default Constants

BEGIN
  yt_rsc_0_0_i_clka_en_d <= yt_rsc_0_0_cgo OR yt_rsc_0_0_cgo_iro;
  yt_rsc_0_16_i_clka_en_d <= yt_rsc_0_16_cgo OR yt_rsc_0_16_cgo_iro;
  mult_t_mul_cmp_en <= ensig_cgo OR ensig_cgo_iro;
  mult_z_mul_cmp_1_en <= ensig_cgo_17 OR ensig_cgo_iro_17;
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_16_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_17_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_18_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_19_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_20_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_21_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_22_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_23_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_24_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_25_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_26_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_27_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_28_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_29_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_30_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_31_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    yt_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_0_i_clka_en_d : OUT STD_LOGIC;
    yt_rsc_0_0_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_1_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_1_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_2_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_2_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_3_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_3_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_4_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_4_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_5_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_5_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_6_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_6_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_7_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_7_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_8_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_8_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_9_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_9_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_10_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_10_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_11_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_11_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_12_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_12_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_13_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_13_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_14_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_14_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_15_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_15_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_16_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_16_i_clka_en_d : OUT STD_LOGIC;
    yt_rsc_0_16_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_16_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_17_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_17_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_17_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_18_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_18_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_18_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_19_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_19_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_19_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_20_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_20_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_20_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_21_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_21_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_21_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_22_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_22_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_22_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_23_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_23_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_23_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_24_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_24_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_24_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_25_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_25_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_25_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_26_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_26_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_26_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_27_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_27_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_27_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_28_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_28_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_28_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_29_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_29_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_29_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_30_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_30_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_30_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yt_rsc_0_31_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    yt_rsc_0_31_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_31_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_0_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_1_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_1_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_2_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_2_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_3_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_3_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_4_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_4_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_5_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_5_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_6_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_6_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_7_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_7_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_8_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_8_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_9_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_9_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_10_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_10_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_11_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_11_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_12_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_12_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_13_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_13_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_14_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_14_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_15_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_15_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_16_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_16_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_16_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_17_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_17_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_17_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_18_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_18_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_18_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_19_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_19_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_19_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_20_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_20_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_20_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_21_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_21_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_21_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_22_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_22_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_22_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_23_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_23_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_23_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_24_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_24_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_24_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_25_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_25_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_25_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_26_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_26_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_26_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_27_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_27_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_27_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_28_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_28_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_28_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_29_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_29_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_29_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_30_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_30_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_30_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xt_rsc_0_31_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    xt_rsc_0_31_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_31_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    twiddle_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_1_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_2_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_3_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_4_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_5_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_6_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_7_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_8_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_9_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_10_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_11_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_12_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_13_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_14_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_rsc_0_15_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_1_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_2_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_3_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_4_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_5_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_6_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_7_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_8_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_9_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
        DOWNTO 0);
    twiddle_h_rsc_0_10_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    twiddle_h_rsc_0_11_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    twiddle_h_rsc_0_12_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    twiddle_h_rsc_0_13_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    twiddle_h_rsc_0_14_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    twiddle_h_rsc_0_15_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    yt_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yt_rsc_0_16_i_wea_d_pff : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xt_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xt_rsc_0_16_i_wea_d_pff : OUT STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END peaseNTT_core;

ARCHITECTURE v11 OF peaseNTT_core IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL p_rsci_idat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_en : STD_LOGIC;
  SIGNAL mult_t_mul_cmp_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_1_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_2_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_3_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_4_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_5_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_6_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_7_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_8_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_9_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_10_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_11_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_12_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_13_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_14_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_15_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_1_en : STD_LOGIC;
  SIGNAL mult_z_mul_cmp_1_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_2_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_3_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_4_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_5_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_6_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_7_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_8_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_9_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_10_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_11_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_12_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_13_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_14_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_15_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_16_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_17_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_18_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_19_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_20_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_21_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_22_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_23_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_24_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_25_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_26_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_27_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_28_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_29_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_30_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_31_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL fsm_output : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL INNER_LOOP4_nor_tmp : STD_LOGIC;
  SIGNAL or_dcpl_13 : STD_LOGIC;
  SIGNAL or_dcpl_22 : STD_LOGIC;
  SIGNAL or_dcpl_45 : STD_LOGIC;
  SIGNAL or_dcpl_65 : STD_LOGIC;
  SIGNAL or_dcpl_101 : STD_LOGIC;
  SIGNAL or_dcpl_121 : STD_LOGIC;
  SIGNAL and_dcpl_51 : STD_LOGIC;
  SIGNAL and_dcpl_56 : STD_LOGIC;
  SIGNAL and_dcpl_57 : STD_LOGIC;
  SIGNAL or_dcpl_194 : STD_LOGIC;
  SIGNAL and_dcpl_58 : STD_LOGIC;
  SIGNAL and_dcpl_59 : STD_LOGIC;
  SIGNAL or_dcpl_197 : STD_LOGIC;
  SIGNAL or_dcpl_198 : STD_LOGIC;
  SIGNAL or_dcpl_199 : STD_LOGIC;
  SIGNAL or_dcpl_200 : STD_LOGIC;
  SIGNAL and_dcpl_67 : STD_LOGIC;
  SIGNAL and_dcpl_68 : STD_LOGIC;
  SIGNAL and_dcpl_69 : STD_LOGIC;
  SIGNAL and_dcpl_70 : STD_LOGIC;
  SIGNAL or_dcpl_205 : STD_LOGIC;
  SIGNAL or_dcpl_206 : STD_LOGIC;
  SIGNAL or_dcpl_207 : STD_LOGIC;
  SIGNAL or_dcpl_208 : STD_LOGIC;
  SIGNAL or_dcpl_210 : STD_LOGIC;
  SIGNAL or_dcpl_212 : STD_LOGIC;
  SIGNAL or_dcpl_214 : STD_LOGIC;
  SIGNAL and_dcpl_79 : STD_LOGIC;
  SIGNAL and_dcpl_81 : STD_LOGIC;
  SIGNAL and_dcpl_82 : STD_LOGIC;
  SIGNAL or_dcpl_217 : STD_LOGIC;
  SIGNAL or_dcpl_218 : STD_LOGIC;
  SIGNAL and_dcpl_90 : STD_LOGIC;
  SIGNAL or_dcpl_233 : STD_LOGIC;
  SIGNAL or_tmp_21 : STD_LOGIC;
  SIGNAL or_tmp_22 : STD_LOGIC;
  SIGNAL or_tmp_25 : STD_LOGIC;
  SIGNAL or_tmp_26 : STD_LOGIC;
  SIGNAL or_tmp_203 : STD_LOGIC;
  SIGNAL or_tmp_204 : STD_LOGIC;
  SIGNAL or_tmp_207 : STD_LOGIC;
  SIGNAL or_tmp_208 : STD_LOGIC;
  SIGNAL or_tmp_771 : STD_LOGIC;
  SIGNAL or_tmp_779 : STD_LOGIC;
  SIGNAL or_tmp_782 : STD_LOGIC;
  SIGNAL or_tmp_790 : STD_LOGIC;
  SIGNAL or_tmp_792 : STD_LOGIC;
  SIGNAL or_tmp_809 : STD_LOGIC;
  SIGNAL or_tmp_819 : STD_LOGIC;
  SIGNAL or_tmp_885 : STD_LOGIC;
  SIGNAL or_tmp_894 : STD_LOGIC;
  SIGNAL or_tmp_1134 : STD_LOGIC;
  SIGNAL or_tmp_1138 : STD_LOGIC;
  SIGNAL or_tmp_1189 : STD_LOGIC;
  SIGNAL and_167_cse : STD_LOGIC;
  SIGNAL and_192_cse : STD_LOGIC;
  SIGNAL and_1445_cse : STD_LOGIC;
  SIGNAL and_1454_cse : STD_LOGIC;
  SIGNAL and_1463_cse : STD_LOGIC;
  SIGNAL and_1700_cse : STD_LOGIC;
  SIGNAL and_1719_cse : STD_LOGIC;
  SIGNAL and_1725_cse : STD_LOGIC;
  SIGNAL and_1763_cse : STD_LOGIC;
  SIGNAL and_1783_cse : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_11_4_sva_6_0 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL INNER_LOOP3_r_11_4_sva_6_0 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL INNER_LOOP2_r_11_4_sva_6_0 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_11_4_sva_6_0 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly2_11_tw_h_slc_operator_33_true_2_lshift_psp_2_0_1_0_itm : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL c_1_sva : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_10 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_9 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_11 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 : STD_LOGIC;
  SIGNAL operator_20_false_acc_cse_sva : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL operator_33_true_3_lshift_psp_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL INNER_LOOP1_stage_0_4 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_2 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_3 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_6 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_7 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_5 : STD_LOGIC;
  SIGNAL p_sva : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_yt_rsc_0_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_0_16_cgo_cse : STD_LOGIC;
  SIGNAL reg_xt_rsc_triosy_0_31_obj_ld_cse : STD_LOGIC;
  SIGNAL reg_ensig_cgo_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_49_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_51_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_53_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_55_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_44_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_45_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_46_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_47_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_48_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_50_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_52_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_54_cse : STD_LOGIC;
  SIGNAL reg_ensig_cgo_17_cse : STD_LOGIC;
  SIGNAL butterFly1_or_5_cse : STD_LOGIC;
  SIGNAL butterFly1_or_1_cse : STD_LOGIC;
  SIGNAL butterFly1_mux_17_cse : STD_LOGIC;
  SIGNAL butterFly1_or_4_cse : STD_LOGIC;
  SIGNAL butterFly1_or_cse : STD_LOGIC;
  SIGNAL mult_15_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_14_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_13_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_11_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_9_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_8_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_7_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_6_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_5_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_4_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_3_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_2_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly2_7_tw_nor_cse : STD_LOGIC;
  SIGNAL butterFly2_7_tw_nor_1_cse : STD_LOGIC;
  SIGNAL butterFly2_7_tw_nor_2_cse : STD_LOGIC;
  SIGNAL mult_15_t_or_9_cse : STD_LOGIC;
  SIGNAL mult_15_t_or_10_cse : STD_LOGIC;
  SIGNAL mult_15_t_or_11_cse : STD_LOGIC;
  SIGNAL mult_15_t_or_12_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_41_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_42_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_43_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_37_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_38_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_39_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_30_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_31_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_32_cse : STD_LOGIC;
  SIGNAL mult_15_t_or_3_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_40_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_36_cse : STD_LOGIC;
  SIGNAL mult_15_t_and_29_cse : STD_LOGIC;
  SIGNAL nor_7_cse : STD_LOGIC;
  SIGNAL mult_15_t_or_1_cse : STD_LOGIC;
  SIGNAL mult_15_t_or_cse : STD_LOGIC;
  SIGNAL reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_570_itm_8_cse : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_602_itm_9_cse : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_633_itm_8_cse : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_114_itm_9_cse : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_129_itm_8_cse : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_161_itm_9_cse : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_192_itm_8_cse : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_224_itm_9_cse : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_255_itm_8_cse : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_287_itm_9_cse : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_318_itm_8_cse : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_350_itm_9_cse : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_381_itm_8_cse : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL or_261_rmff : STD_LOGIC;
  SIGNAL butterFly1_nor_7_rmff : STD_LOGIC;
  SIGNAL butterFly1_butterFly1_or_1_rmff : STD_LOGIC;
  SIGNAL butterFly1_butterFly1_mux_3_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_butterFly1_and_17_rmff : STD_LOGIC;
  SIGNAL butterFly1_mux1h_15_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL and_202_rmff : STD_LOGIC;
  SIGNAL butterFly1_1_butterFly1_1_mux_3_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_1_mux1h_11_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_2_butterFly1_2_mux_3_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_2_mux1h_11_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_3_butterFly1_3_mux_3_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_3_mux1h_11_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_4_butterFly1_4_mux_3_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_4_mux1h_11_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_7_butterFly1_7_mux_3_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_8_butterFly1_8_mux_3_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_8_mux1h_11_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL or_443_rmff : STD_LOGIC;
  SIGNAL butterFly1_nor_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_butterFly1_or_rmff : STD_LOGIC;
  SIGNAL butterFly1_butterFly1_mux_4_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_butterFly1_and_15_rmff : STD_LOGIC;
  SIGNAL butterFly1_mux1h_13_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_1_butterFly1_1_mux_4_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_1_mux1h_9_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_2_butterFly1_2_mux_4_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_2_mux1h_9_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_3_butterFly1_3_mux_4_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_3_mux1h_9_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_4_butterFly1_4_mux_4_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_4_mux1h_9_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_7_butterFly1_7_mux_4_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_8_butterFly1_8_mux_4_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_8_mux1h_9_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_15_f2_mux1h_65_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_f1_butterFly1_f1_mux_2_rmff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_f1_butterFly1_f1_mux_3_rmff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_f1_butterFly1_f1_butterFly1_f1_butterFly1_f1_nor_rmff : STD_LOGIC;
  SIGNAL and_921_rmff : STD_LOGIC;
  SIGNAL butterFly1_15_f2_mux1h_64_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_f2_butterFly1_f2_mux_2_rmff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_f2_butterFly1_f2_mux_3_rmff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_15_f2_mux1h_63_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_1_f1_butterFly1_1_f1_mux_2_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_1_f1_butterFly1_1_f1_mux_3_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_15_f2_mux1h_62_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_1_f2_butterFly1_1_f2_mux_2_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_1_f2_butterFly1_1_f2_mux_3_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_15_f2_mux1h_61_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_2_f1_butterFly1_2_f1_mux_2_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_2_f1_butterFly1_2_f1_mux_3_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_15_f2_mux1h_60_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_2_f2_butterFly1_2_f2_mux_2_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_2_f2_butterFly1_2_f2_mux_3_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_15_f2_mux1h_59_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_3_f1_butterFly1_3_f1_mux_2_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_3_f1_butterFly1_3_f1_mux_3_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_15_f2_mux1h_58_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_3_f2_butterFly1_3_f2_mux_2_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_3_f2_butterFly1_3_f2_mux_3_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_15_f2_mux1h_57_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_4_f1_butterFly1_4_f1_mux_2_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_4_f1_butterFly1_4_f1_mux_3_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_15_f2_mux1h_56_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_4_f2_butterFly1_4_f2_mux_2_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_4_f2_butterFly1_4_f2_mux_3_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_15_f2_mux1h_55_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_5_f1_butterFly1_5_f1_mux_2_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_5_f1_butterFly1_5_f1_mux_3_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_15_f2_mux1h_54_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_5_f2_butterFly1_5_f2_mux_2_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_5_f2_butterFly1_5_f2_mux_3_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_15_f2_mux1h_53_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_6_f1_butterFly1_6_f1_mux_2_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_6_f1_butterFly1_6_f1_mux_3_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_15_f2_mux1h_52_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_6_f2_butterFly1_6_f2_mux_2_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_6_f2_butterFly1_6_f2_mux_3_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_15_f2_mux1h_51_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_7_f1_butterFly1_7_f1_mux_2_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_7_f1_butterFly1_7_f1_mux_3_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_15_f2_mux1h_50_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL butterFly1_7_f2_butterFly1_7_f2_mux_2_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_7_f2_butterFly1_7_f2_mux_3_rmff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL butterFly1_f1_butterFly1_f1_butterFly1_f1_butterFly1_8_f1_nor_rmff : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_mux1h_4_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL and_1435_rmff : STD_LOGIC;
  SIGNAL butterFly2_1_tw_butterFly2_1_tw_mux_rmff : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL or_896_rmff : STD_LOGIC;
  SIGNAL or_900_rmff : STD_LOGIC;
  SIGNAL or_904_rmff : STD_LOGIC;
  SIGNAL or_908_rmff : STD_LOGIC;
  SIGNAL or_912_rmff : STD_LOGIC;
  SIGNAL or_916_rmff : STD_LOGIC;
  SIGNAL or_920_rmff : STD_LOGIC;
  SIGNAL and_1506_rmff : STD_LOGIC;
  SIGNAL or_997_rmff : STD_LOGIC;
  SIGNAL or_1156_rmff : STD_LOGIC;
  SIGNAL mult_4_t_mux1h_1_rmff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_da_d_mx0w0_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_da_d_mx0w2_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_15_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_31_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_da_d_mx0w0_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_da_d_mx0w2_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_14_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_30_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_da_d_mx0w0_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_da_d_mx0w2_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_13_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_29_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_da_d_mx0w0_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_da_d_mx0w2_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_12_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_28_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_da_d_mx0w0_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_da_d_mx0w2_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_11_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_27_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_da_d_mx0w0_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_da_d_mx0w2_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_10_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_26_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_da_d_mx0w0_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_da_d_mx0w2_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_25_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_da_d_mx0w0_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_da_d_mx0w2_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_24_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_da_d_mx0w0_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_23_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_9 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_da_d_mx0w0_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_da_d_mx0w2_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_1_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_9 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_da_d_mx0w2_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_da_d_mx0w0_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_da_d_mx0w2_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_da_d_mx0w0_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_da_d_mx0w2_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_da_d_mx0w0_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_da_d_mx0w2_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_da_d_mx0w0_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_da_d_mx0w2_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_da_d_mx0w0_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_da_d_mx0w2_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_8 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_8 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_wea_d_mx0c2 : STD_LOGIC;
  SIGNAL yt_rsc_0_0_i_wea_d_mx0c0 : STD_LOGIC;
  SIGNAL yt_rsc_0_16_i_wea_d_mx0c2 : STD_LOGIC;
  SIGNAL yt_rsc_0_16_i_wea_d_mx0c0 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_8 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_9 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL z_out : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL z_out_1 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL z_out_2 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL z_out_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_9 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_10 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_12 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_13 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_14 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_16 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_17 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_18 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_20 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_21 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_22 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_24 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_25 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_26 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_28 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_29 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_31 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_34 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_36 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_37 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_39 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_41 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_42 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_44 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_46 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_47 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_49 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_51 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_52 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_53 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_54 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_55 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_56 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_57 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_58 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_59 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_60 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_61 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_62 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_63 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_64 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_65 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_66 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_67 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_68 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_69 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_70 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_71 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_72 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_73 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_74 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_75 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_76 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_77 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_78 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_79 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_80 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_81 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_82 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL operator_33_true_1_lshift_psp_9_4_sva : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL INNER_LOOP1_stage_0_8 : STD_LOGIC;
  SIGNAL mult_res_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_res_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_2_res_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_3_res_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_4_res_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_5_res_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_6_res_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_7_res_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_8_res_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_9_res_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_res_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_11_res_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_res_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_13_res_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_14_res_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_15_res_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_8 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_8 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL mult_10_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_8 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL mult_11_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_11_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_11_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_8 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL mult_12_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_8 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL mult_13_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_13_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_13_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_8 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL mult_14_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_14_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_14_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_8 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL mult_15_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_15_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_15_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_8 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 : STD_LOGIC;
  SIGNAL tmp_10_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_16_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_17_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_18_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_19_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_20_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_21_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_22_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_23_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_23_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_23_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_24_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_24_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_24_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_25_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_25_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_25_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_26_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_26_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_27_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_27_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_28_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_28_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_29_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_29_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_8 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL mult_30_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_30_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_1 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_2 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_3 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_4 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_5 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_6 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_7 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_8 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_9 : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL mult_31_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_31_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly2_15_tw_equal_tmp_1 : STD_LOGIC;
  SIGNAL butterFly2_15_tw_equal_tmp_3_1 : STD_LOGIC;
  SIGNAL butterFly2_15_tw_equal_tmp_5_1 : STD_LOGIC;
  SIGNAL butterFly2_15_tw_equal_tmp_6_1 : STD_LOGIC;
  SIGNAL butterFly2_15_tw_equal_tmp_7_1 : STD_LOGIC;
  SIGNAL tmp_60_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL operator_33_true_3_lshift_psp_1_0_sva_mx0w3 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL mult_15_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_14_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_13_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_11_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_9_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_8_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_7_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_6_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_5_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_4_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_3_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_2_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_res_lpi_3_dfm_1_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_31_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_31_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_30_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_30_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_29_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_29_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_28_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_28_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_27_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_27_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_26_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_26_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_25_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_25_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_24_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_24_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_23_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_23_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_22_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_22_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_21_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_21_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_20_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_20_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_19_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_19_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_18_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_18_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_17_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_17_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_16_qelse_and_ssc : STD_LOGIC;
  SIGNAL modulo_sub_16_qelse_and_ssc_1 : STD_LOGIC;
  SIGNAL reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd : STD_LOGIC;
  SIGNAL reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd_1 : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_add_1_qelse_or_m1c : STD_LOGIC;
  SIGNAL reg_mult_17_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_25_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_28_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_20_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_22_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_30_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_26_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_18_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_19_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_23_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_27_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_31_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_29_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_24_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_21_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_16_res_lpi_3_dfm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL or_12_cse : STD_LOGIC;
  SIGNAL or_44_cse : STD_LOGIC;
  SIGNAL or_64_cse : STD_LOGIC;
  SIGNAL or_84_cse : STD_LOGIC;
  SIGNAL or_103_cse : STD_LOGIC;
  SIGNAL or_123_cse : STD_LOGIC;
  SIGNAL or_143_cse : STD_LOGIC;
  SIGNAL or_142_cse : STD_LOGIC;
  SIGNAL modulo_sub_5_qelse_mux_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_83_32 : STD_LOGIC;
  SIGNAL z_out_84_32 : STD_LOGIC;
  SIGNAL z_out_85_32 : STD_LOGIC;
  SIGNAL z_out_86_32 : STD_LOGIC;
  SIGNAL z_out_87_32 : STD_LOGIC;
  SIGNAL z_out_88_32 : STD_LOGIC;
  SIGNAL z_out_89_32 : STD_LOGIC;
  SIGNAL z_out_90_32 : STD_LOGIC;
  SIGNAL z_out_91_32 : STD_LOGIC;
  SIGNAL z_out_92_32 : STD_LOGIC;
  SIGNAL z_out_93_32 : STD_LOGIC;
  SIGNAL z_out_94_32 : STD_LOGIC;
  SIGNAL z_out_95_32 : STD_LOGIC;
  SIGNAL z_out_96_32 : STD_LOGIC;
  SIGNAL z_out_97_32 : STD_LOGIC;
  SIGNAL z_out_98_32 : STD_LOGIC;

  SIGNAL c_mux_nl : STD_LOGIC;
  SIGNAL butterFly2_21_tw_butterFly2_21_tw_or_nl : STD_LOGIC;
  SIGNAL STAGE_LOOP_mux1h_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL STAGE_LOOP_and_nl : STD_LOGIC;
  SIGNAL nor_4_nl : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_mux_44_nl : STD_LOGIC;
  SIGNAL acc_2_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_1_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_1_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_1_qelse_or_1_nl : STD_LOGIC;
  SIGNAL modulo_add_1_qelse_and_4_nl : STD_LOGIC;
  SIGNAL modulo_add_1_qelse_and_5_nl : STD_LOGIC;
  SIGNAL acc_6_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_10_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_10_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_10_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_10_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_10_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_10_qelse_and_7_nl : STD_LOGIC;
  SIGNAL acc_10_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_11_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_11_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_11_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_11_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_11_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_11_qelse_and_7_nl : STD_LOGIC;
  SIGNAL acc_14_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_12_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_12_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_12_qelse_or_1_nl : STD_LOGIC;
  SIGNAL modulo_add_12_qelse_and_4_nl : STD_LOGIC;
  SIGNAL modulo_add_12_qelse_and_5_nl : STD_LOGIC;
  SIGNAL acc_18_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_13_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_13_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_13_qelse_or_1_nl : STD_LOGIC;
  SIGNAL modulo_add_13_qelse_and_4_nl : STD_LOGIC;
  SIGNAL modulo_add_13_qelse_and_5_nl : STD_LOGIC;
  SIGNAL acc_22_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_14_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_14_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_14_qelse_or_1_nl : STD_LOGIC;
  SIGNAL modulo_add_14_qelse_and_4_nl : STD_LOGIC;
  SIGNAL modulo_add_14_qelse_and_5_nl : STD_LOGIC;
  SIGNAL acc_26_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_15_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_15_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_15_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_15_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_15_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_15_qelse_and_7_nl : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_mux_45_nl : STD_LOGIC;
  SIGNAL INNER_LOOP1_mux_nl : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_mux1h_46_nl : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_INNER_LOOP1_r_and_1_nl : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_INNER_LOOP1_r_and_3_nl : STD_LOGIC;
  SIGNAL or_1465_nl : STD_LOGIC;
  SIGNAL INNER_LOOP1_mux_11_nl : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_INNER_LOOP1_r_and_2_nl : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_INNER_LOOP1_r_and_nl : STD_LOGIC;
  SIGNAL STAGE_LOOP_base_STAGE_LOOP_base_mux_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL INNER_LOOP2_r_or_nl : STD_LOGIC;
  SIGNAL acc_29_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_2_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_23_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_23_qelse_or_1_nl : STD_LOGIC;
  SIGNAL modulo_add_23_qelse_and_4_nl : STD_LOGIC;
  SIGNAL modulo_add_23_qelse_and_5_nl : STD_LOGIC;
  SIGNAL acc_32_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_3_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_24_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_24_qelse_or_1_nl : STD_LOGIC;
  SIGNAL modulo_add_24_qelse_and_4_nl : STD_LOGIC;
  SIGNAL modulo_add_24_qelse_and_5_nl : STD_LOGIC;
  SIGNAL acc_34_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_4_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_25_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_25_qelse_or_1_nl : STD_LOGIC;
  SIGNAL modulo_add_25_qelse_and_4_nl : STD_LOGIC;
  SIGNAL modulo_add_25_qelse_and_5_nl : STD_LOGIC;
  SIGNAL acc_37_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_5_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_26_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_26_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_26_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_26_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_26_qelse_and_7_nl : STD_LOGIC;
  SIGNAL acc_39_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_6_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_27_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_27_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_27_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_27_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_27_qelse_and_7_nl : STD_LOGIC;
  SIGNAL acc_42_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_7_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_28_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_28_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_28_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_28_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_28_qelse_and_7_nl : STD_LOGIC;
  SIGNAL acc_44_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_8_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_29_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_29_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_29_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_29_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_29_qelse_and_7_nl : STD_LOGIC;
  SIGNAL acc_47_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_9_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_30_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_30_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_30_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_30_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_30_qelse_and_7_nl : STD_LOGIC;
  SIGNAL acc_49_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_31_qelse_and_nl : STD_LOGIC;
  SIGNAL modulo_add_31_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_add_31_qelse_and_5_nl : STD_LOGIC;
  SIGNAL modulo_add_31_qelse_and_6_nl : STD_LOGIC;
  SIGNAL modulo_add_31_qelse_and_7_nl : STD_LOGIC;
  SIGNAL modulo_sub_16_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_17_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_18_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_19_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_20_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_21_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_22_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_23_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_24_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_25_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_26_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_27_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_28_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_29_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_30_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_31_qelse_or_nl : STD_LOGIC;
  SIGNAL modulo_sub_5_qif_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_15_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_31_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_14_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_30_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_13_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_29_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_12_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_28_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_11_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_27_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_10_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_26_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_9_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_25_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_8_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_24_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_7_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_23_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_6_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_22_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_5_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_21_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_4_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_20_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_3_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_19_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_2_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_18_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_1_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_17_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_16_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL INNER_LOOP1_tw_and_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL INNER_LOOP2_tw_and_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_butterFly1_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_butterFly1_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_butterFly1_nor_2_nl : STD_LOGIC;
  SIGNAL butterFly1_butterFly1_nor_3_nl : STD_LOGIC;
  SIGNAL butterFly1_mux_15_nl : STD_LOGIC;
  SIGNAL butterFly1_1_butterFly1_1_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_1_butterFly1_1_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_2_butterFly1_2_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_2_butterFly1_2_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_3_butterFly1_3_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_3_butterFly1_3_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_4_butterFly1_4_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_4_butterFly1_4_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_5_butterFly1_5_mux_3_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_5_mux1h_11_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_5_butterFly1_5_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_5_butterFly1_5_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_6_butterFly1_6_mux_3_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_6_mux1h_11_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_6_butterFly1_6_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_6_butterFly1_6_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_7_mux1h_11_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_7_butterFly1_7_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_7_butterFly1_7_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_8_butterFly1_8_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_8_butterFly1_8_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_9_butterFly1_9_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_9_butterFly1_9_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_10_butterFly1_10_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_10_butterFly1_10_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_11_butterFly1_11_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_11_butterFly1_11_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_12_butterFly1_12_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_12_butterFly1_12_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_13_butterFly1_13_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_13_butterFly1_13_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_14_mux1h_11_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_14_butterFly1_14_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_14_butterFly1_14_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_15_butterFly1_15_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_15_butterFly1_15_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_butterFly1_mux_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_butterFly1_mux_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_butterFly1_nor_nl : STD_LOGIC;
  SIGNAL butterFly1_butterFly1_nor_1_nl : STD_LOGIC;
  SIGNAL butterFly1_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_1_butterFly1_1_mux_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_1_butterFly1_1_mux_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_2_butterFly1_2_mux_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_2_butterFly1_2_mux_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_3_butterFly1_3_mux_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_3_butterFly1_3_mux_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_4_butterFly1_4_mux_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_4_butterFly1_4_mux_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_5_butterFly1_5_mux_4_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_5_mux1h_9_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_5_butterFly1_5_mux_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_5_butterFly1_5_mux_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_6_butterFly1_6_mux_4_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_6_mux1h_9_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_6_butterFly1_6_mux_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_6_butterFly1_6_mux_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_7_mux1h_9_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_7_butterFly1_7_mux_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_7_butterFly1_7_mux_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_8_butterFly1_8_mux_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_8_butterFly1_8_mux_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_9_butterFly1_9_mux_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_9_butterFly1_9_mux_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_10_butterFly1_10_mux_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_10_butterFly1_10_mux_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_11_butterFly1_11_mux_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_11_butterFly1_11_mux_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_12_butterFly1_12_mux_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_12_butterFly1_12_mux_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_13_butterFly1_13_mux_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_13_butterFly1_13_mux_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_14_mux1h_9_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL butterFly1_14_butterFly1_14_mux_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_14_butterFly1_14_mux_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_15_butterFly1_15_mux_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_15_butterFly1_15_mux_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL operator_20_false_mux_2_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL operator_20_false_mux1h_2_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL modulo_sub_6_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_37_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_36_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_4_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_35_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_3_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_34_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_2_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_33_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_1_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_32_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_31_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_13_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_30_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_45_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_29_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_15_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_28_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_27_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_26_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_25_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_24_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_23_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_22_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_21_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_20_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_19_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_18_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_17_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_16_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL acc_50_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_mux1h_17_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_51_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_1_mux1h_13_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_52_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_2_mux1h_13_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_53_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_3_mux1h_13_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_54_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_4_mux1h_13_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_55_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_5_mux1h_13_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_56_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_6_mux1h_13_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_57_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_7_mux1h_13_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_58_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_8_mux1h_13_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_59_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_9_mux1h_13_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_60_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_10_mux1h_13_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_61_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_11_mux1h_13_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_62_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_12_mux1h_13_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_63_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_13_mux1h_13_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_64_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_14_mux1h_13_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_65_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_15_mux1h_13_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_15_mux1h_14_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_14_mux1h_14_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_13_mux1h_14_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_12_mux1h_14_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_11_mux1h_14_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_10_mux1h_14_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_9_mux1h_14_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_8_mux1h_14_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_7_mux1h_14_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_6_mux1h_14_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_5_mux1h_14_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_4_mux1h_14_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_3_mux1h_14_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_2_mux1h_14_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_1_mux1h_14_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_mux1h_18_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_82_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_1_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_83_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_10_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_84_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_54_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_85_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_48_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_86_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_33_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_87_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_34_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_88_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_6_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_89_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_50_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_90_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_51_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_91_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_14_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_92_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_36_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_93_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_52_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_94_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_41_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_95_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_2_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_96_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_53_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_97_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_55_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL p_rsci_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL p_rsci_idat_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_1_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_1_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_1_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_2_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_2_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_2_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_3_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_3_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_3_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_4_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_4_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_4_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_5_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_5_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_5_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_6_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_6_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_6_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_7_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_7_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_7_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_8_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_8_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_8_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_9_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_9_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_9_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_10_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_10_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_10_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_11_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_11_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_11_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_12_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_12_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_12_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_13_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_13_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_13_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_14_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_14_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_14_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_15_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_15_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_15_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_1_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_1_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_1_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_2_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_2_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_2_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_3_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_3_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_3_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_4_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_4_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_4_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_5_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_5_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_5_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_6_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_6_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_6_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_7_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_7_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_7_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_8_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_8_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_8_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_9_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_9_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_9_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_10_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_10_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_10_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_11_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_11_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_11_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_12_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_12_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_12_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_13_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_13_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_13_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_14_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_14_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_14_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_15_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_15_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_15_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_16_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_16_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_16_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_17_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_17_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_17_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_18_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_18_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_18_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_19_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_19_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_19_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_20_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_20_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_20_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_21_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_21_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_21_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_22_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_22_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_22_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_23_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_23_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_23_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_24_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_24_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_24_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_25_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_25_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_25_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_26_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_26_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_26_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_27_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_27_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_27_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_28_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_28_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_28_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_29_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_29_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_29_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_30_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_30_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_30_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_31_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_31_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_31_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL operator_33_true_3_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL operator_33_true_3_lshift_rg_s : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL operator_33_true_3_lshift_rg_z : STD_LOGIC_VECTOR (1 DOWNTO 0);

  SIGNAL operator_33_true_1_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL operator_33_true_1_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL operator_33_true_1_lshift_rg_z : STD_LOGIC_VECTOR (10 DOWNTO 0);

  COMPONENT peaseNTT_core_wait_dp
    PORT(
      yt_rsc_0_0_cgo_iro : IN STD_LOGIC;
      yt_rsc_0_0_i_clka_en_d : OUT STD_LOGIC;
      yt_rsc_0_16_cgo_iro : IN STD_LOGIC;
      yt_rsc_0_16_i_clka_en_d : OUT STD_LOGIC;
      ensig_cgo_iro : IN STD_LOGIC;
      ensig_cgo_iro_17 : IN STD_LOGIC;
      yt_rsc_0_0_cgo : IN STD_LOGIC;
      yt_rsc_0_16_cgo : IN STD_LOGIC;
      ensig_cgo : IN STD_LOGIC;
      mult_t_mul_cmp_en : OUT STD_LOGIC;
      ensig_cgo_17 : IN STD_LOGIC;
      mult_z_mul_cmp_1_en : OUT STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      INNER_LOOP1_C_0_tr0 : IN STD_LOGIC;
      INNER_LOOP2_C_0_tr0 : IN STD_LOGIC;
      STAGE_LOOP_C_2_tr0 : IN STD_LOGIC;
      INNER_LOOP3_C_0_tr0 : IN STD_LOGIC;
      INNER_LOOP4_C_0_tr0 : IN STD_LOGIC;
      INNER_LOOP4_C_0_tr1 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL peaseNTT_core_core_fsm_inst_INNER_LOOP1_C_0_tr0 : STD_LOGIC;
  SIGNAL peaseNTT_core_core_fsm_inst_STAGE_LOOP_C_2_tr0 : STD_LOGIC;
  SIGNAL peaseNTT_core_core_fsm_inst_INNER_LOOP4_C_0_tr1 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_s_1_4_2(input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_2_5_2(input_4 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_31_3_2(input_2 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(30 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(30 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_12_2(input_11 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(11 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_3_2(input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_4_2(input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_5_2(input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_6_2(input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_8_2(input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(7 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_9_2(input_8 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(8 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_3_2(input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_3_2(input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_4_2(input_3 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_7_4_2(input_3 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_2_2_2(input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_31_2_2(input_0 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(30 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_3_2_2(input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_6_2_2(input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_7_2_2(input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  p_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 2,
      width => 32
      )
    PORT MAP(
      dat => p_rsci_dat,
      idat => p_rsci_idat_1
    );
  p_rsci_dat <= p_rsc_dat;
  p_rsci_idat <= p_rsci_idat_1;

  xt_rsc_triosy_0_31_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_31_lz
    );
  xt_rsc_triosy_0_30_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_30_lz
    );
  xt_rsc_triosy_0_29_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_29_lz
    );
  xt_rsc_triosy_0_28_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_28_lz
    );
  xt_rsc_triosy_0_27_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_27_lz
    );
  xt_rsc_triosy_0_26_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_26_lz
    );
  xt_rsc_triosy_0_25_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_25_lz
    );
  xt_rsc_triosy_0_24_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_24_lz
    );
  xt_rsc_triosy_0_23_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_23_lz
    );
  xt_rsc_triosy_0_22_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_22_lz
    );
  xt_rsc_triosy_0_21_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_21_lz
    );
  xt_rsc_triosy_0_20_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_20_lz
    );
  xt_rsc_triosy_0_19_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_19_lz
    );
  xt_rsc_triosy_0_18_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_18_lz
    );
  xt_rsc_triosy_0_17_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_17_lz
    );
  xt_rsc_triosy_0_16_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_16_lz
    );
  xt_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_15_lz
    );
  xt_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_14_lz
    );
  xt_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_13_lz
    );
  xt_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_12_lz
    );
  xt_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_11_lz
    );
  xt_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_10_lz
    );
  xt_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_9_lz
    );
  xt_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_8_lz
    );
  xt_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_7_lz
    );
  xt_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_6_lz
    );
  xt_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_5_lz
    );
  xt_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_4_lz
    );
  xt_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_3_lz
    );
  xt_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_2_lz
    );
  xt_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_1_lz
    );
  xt_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => xt_rsc_triosy_0_0_lz
    );
  p_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => p_rsc_triosy_lz
    );
  r_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => r_rsc_triosy_lz
    );
  twiddle_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_15_lz
    );
  twiddle_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_14_lz
    );
  twiddle_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_13_lz
    );
  twiddle_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_12_lz
    );
  twiddle_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_11_lz
    );
  twiddle_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_10_lz
    );
  twiddle_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_9_lz
    );
  twiddle_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_8_lz
    );
  twiddle_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_7_lz
    );
  twiddle_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_6_lz
    );
  twiddle_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_5_lz
    );
  twiddle_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_4_lz
    );
  twiddle_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_3_lz
    );
  twiddle_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_2_lz
    );
  twiddle_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_1_lz
    );
  twiddle_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_0_lz
    );
  twiddle_h_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_15_lz
    );
  twiddle_h_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_14_lz
    );
  twiddle_h_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_13_lz
    );
  twiddle_h_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_12_lz
    );
  twiddle_h_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_11_lz
    );
  twiddle_h_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_10_lz
    );
  twiddle_h_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_9_lz
    );
  twiddle_h_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_8_lz
    );
  twiddle_h_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_7_lz
    );
  twiddle_h_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_6_lz
    );
  twiddle_h_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_5_lz
    );
  twiddle_h_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_4_lz
    );
  twiddle_h_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_3_lz
    );
  twiddle_h_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_2_lz
    );
  twiddle_h_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_1_lz
    );
  twiddle_h_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_xt_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_h_rsc_triosy_0_0_lz
    );
  mult_t_mul_cmp : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_a,
      b => mult_t_mul_cmp_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_z_1
    );
  mult_t_mul_cmp_a <= MUX1HOT_v_32_4_2((xt_rsc_0_1_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_1_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_31_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_31_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_b <= MUX1HOT_v_32_9_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_8_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_9_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_10_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_11_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_12_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_13_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_14_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_15_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & mult_15_t_and_44_cse & mult_15_t_and_45_cse & mult_15_t_and_46_cse & mult_15_t_and_47_cse
      & mult_15_t_or_9_cse & mult_15_t_or_10_cse & mult_15_t_or_11_cse & mult_15_t_or_12_cse));
  mult_t_mul_cmp_z <= mult_t_mul_cmp_z_1;

  mult_t_mul_cmp_1 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_1_a,
      b => mult_t_mul_cmp_1_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_1_z_1
    );
  mult_t_mul_cmp_1_a <= MUX1HOT_v_32_4_2((xt_rsc_0_31_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_31_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_29_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_1_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_1_b <= MUX1HOT_v_32_5_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_10_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_12_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_14_i_qa_d(31
      DOWNTO 0)), STD_LOGIC_VECTOR'( or_tmp_771 & mult_15_t_and_40_cse & mult_15_t_and_41_cse
      & mult_15_t_and_42_cse & mult_15_t_and_43_cse));
  mult_t_mul_cmp_1_z <= mult_t_mul_cmp_1_z_1;

  mult_t_mul_cmp_2 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_2_a,
      b => mult_t_mul_cmp_2_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_2_z_1
    );
  mult_t_mul_cmp_2_a <= MUX1HOT_v_32_4_2((xt_rsc_0_29_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_29_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_27_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_3_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_2_b <= MUX1HOT_v_32_6_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_9_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_12_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_13_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_1_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( or_tmp_779
      & mult_15_t_and_36_cse & mult_15_t_and_37_cse & mult_15_t_and_38_cse & mult_15_t_and_39_cse
      & or_tmp_782));
  mult_t_mul_cmp_2_z <= mult_t_mul_cmp_2_z_1;

  mult_t_mul_cmp_3 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_3_a,
      b => mult_t_mul_cmp_3_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_3_z_1
    );
  mult_t_mul_cmp_3_a <= MUX1HOT_v_32_4_2((xt_rsc_0_27_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_27_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_25_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_5_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_3_b <= MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_12_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_2_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( (and_1719_cse
      OR modulo_add_1_qelse_or_m1c) & or_tmp_790 & and_1725_cse & or_tmp_792));
  mult_t_mul_cmp_3_z <= mult_t_mul_cmp_3_z_1;

  mult_t_mul_cmp_4 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_4_a,
      b => mult_t_mul_cmp_4_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_4_z_1
    );
  mult_t_mul_cmp_4_a <= MUX1HOT_v_32_4_2((xt_rsc_0_25_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_25_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_23_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_7_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_4_b <= MUX1HOT_v_32_8_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_9_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_10_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_11_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_1_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_2_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_3_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( (modulo_add_1_qelse_or_m1c
      OR mult_15_t_and_49_cse) & mult_15_t_and_29_cse & mult_15_t_and_30_cse & mult_15_t_and_31_cse
      & mult_15_t_and_32_cse & mult_15_t_and_51_cse & mult_15_t_and_53_cse & mult_15_t_and_55_cse));
  mult_t_mul_cmp_4_z <= mult_t_mul_cmp_4_z_1;

  mult_t_mul_cmp_5 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_5_a,
      b => mult_t_mul_cmp_5_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_5_z_1
    );
  mult_t_mul_cmp_5_a <= MUX1HOT_v_32_4_2((xt_rsc_0_23_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_23_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_21_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_9_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_5_b <= MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_10_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_4_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & or_tmp_809 & and_1763_cse & (fsm_output(9))));
  mult_t_mul_cmp_5_z <= mult_t_mul_cmp_5_z_1;

  mult_t_mul_cmp_6 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_6_a,
      b => mult_t_mul_cmp_6_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_6_z_1
    );
  mult_t_mul_cmp_6_a <= MUX1HOT_v_32_4_2((xt_rsc_0_21_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_21_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_19_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_11_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_6_b <= MUX1HOT_v_32_5_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_9_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_5_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_4_i_qa_d(31
      DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & or_tmp_819 & and_1783_cse
      & or_tmp_782 & and_1700_cse));
  mult_t_mul_cmp_6_z <= mult_t_mul_cmp_6_z_1;

  mult_t_mul_cmp_7 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_7_a,
      b => mult_t_mul_cmp_7_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_7_z_1
    );
  mult_t_mul_cmp_7_a <= MUX1HOT_v_32_4_2((xt_rsc_0_19_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_19_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_17_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_13_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_7_b <= MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_6_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_4_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & or_tmp_792 & and_1719_cse));
  mult_t_mul_cmp_7_z <= mult_t_mul_cmp_7_z_1;

  mult_t_mul_cmp_8 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_8_a,
      b => mult_t_mul_cmp_8_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_8_z_1
    );
  mult_t_mul_cmp_8_a <= MUX1HOT_v_32_4_2((xt_rsc_0_17_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_17_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_15_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_15_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_8_b <= MUX1HOT_v_32_8_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_1_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_2_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_3_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_4_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_5_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_6_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_7_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( mult_15_t_or_3_cse
      & mult_15_t_and_45_cse & mult_15_t_and_46_cse & mult_15_t_and_47_cse & mult_15_t_or_9_cse
      & mult_15_t_or_10_cse & mult_15_t_or_11_cse & mult_15_t_or_12_cse));
  mult_t_mul_cmp_8_z <= mult_t_mul_cmp_8_z_1;

  mult_t_mul_cmp_9 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_9_a,
      b => mult_t_mul_cmp_9_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_9_z_1
    );
  mult_t_mul_cmp_9_a <= MUX1HOT_v_32_4_2((xt_rsc_0_15_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_15_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_13_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_17_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_9_b <= MUX1HOT_v_32_5_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_2_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_4_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_6_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_8_i_qa_d(31
      DOWNTO 0)), STD_LOGIC_VECTOR'( (modulo_add_1_qelse_or_m1c OR mult_15_t_and_40_cse)
      & mult_15_t_and_41_cse & mult_15_t_and_42_cse & mult_15_t_and_43_cse & (fsm_output(9))));
  mult_t_mul_cmp_9_z <= mult_t_mul_cmp_9_z_1;

  mult_t_mul_cmp_10 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_10_a,
      b => mult_t_mul_cmp_10_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_10_z_1
    );
  mult_t_mul_cmp_10_a <= MUX1HOT_v_32_4_2((xt_rsc_0_13_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_13_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_11_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_19_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_10_b <= MUX1HOT_v_32_6_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_1_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_4_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_5_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_9_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( mult_15_t_or_1_cse
      & mult_15_t_and_37_cse & mult_15_t_and_38_cse & mult_15_t_and_39_cse & or_tmp_782
      & and_1700_cse));
  mult_t_mul_cmp_10_z <= mult_t_mul_cmp_10_z_1;

  mult_t_mul_cmp_11 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_11_a,
      b => mult_t_mul_cmp_11_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_11_z_1
    );
  mult_t_mul_cmp_11_a <= MUX1HOT_v_32_4_2((xt_rsc_0_11_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_11_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_9_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_21_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_11_b <= MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_4_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_10_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_8_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( (and_1725_cse
      OR modulo_add_1_qelse_or_m1c) & or_tmp_790 & or_tmp_792 & and_1719_cse));
  mult_t_mul_cmp_11_z <= mult_t_mul_cmp_11_z_1;

  mult_t_mul_cmp_12 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_12_a,
      b => mult_t_mul_cmp_12_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_12_z_1
    );
  mult_t_mul_cmp_12_a <= mult_4_t_mux1h_1_rmff;
  mult_t_mul_cmp_12_b <= MUX1HOT_v_32_8_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_1_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_2_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_3_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_8_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_9_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_10_i_qa_d(31
      DOWNTO 0)), (twiddle_h_rsc_0_11_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( mult_15_t_or_cse
      & mult_15_t_and_30_cse & mult_15_t_and_31_cse & mult_15_t_and_32_cse & mult_15_t_and_49_cse
      & mult_15_t_and_51_cse & mult_15_t_and_53_cse & mult_15_t_and_55_cse));
  mult_t_mul_cmp_12_z <= mult_t_mul_cmp_12_z_1;

  mult_t_mul_cmp_13 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_13_a,
      b => mult_t_mul_cmp_13_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_13_z_1
    );
  mult_t_mul_cmp_13_a <= MUX1HOT_v_32_4_2((xt_rsc_0_7_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_7_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_5_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_25_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_13_b <= MUX1HOT_v_32_3_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_2_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_12_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( or_tmp_885 & or_tmp_809 & (fsm_output(9))));
  mult_t_mul_cmp_13_z <= mult_t_mul_cmp_13_z_1;

  mult_t_mul_cmp_14 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_14_a,
      b => mult_t_mul_cmp_14_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_14_z_1
    );
  mult_t_mul_cmp_14_a <= MUX1HOT_v_32_4_2((xt_rsc_0_5_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_5_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_3_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_27_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_14_b <= MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_1_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_13_i_qa_d(31 DOWNTO
      0)), (twiddle_h_rsc_0_12_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( or_tmp_894
      & or_tmp_819 & or_tmp_782 & and_1700_cse));
  mult_t_mul_cmp_14_z <= mult_t_mul_cmp_14_z_1;

  mult_t_mul_cmp_15 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_t_mul_cmp_15_a,
      b => mult_t_mul_cmp_15_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_15_z_1
    );
  mult_t_mul_cmp_15_a <= MUX1HOT_v_32_4_2((xt_rsc_0_3_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_3_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_1_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_29_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_t_mul_cmp_15_b <= MUX1HOT_v_32_3_2((twiddle_h_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_h_rsc_0_14_i_qa_d(31 DOWNTO 0)), (twiddle_h_rsc_0_12_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (modulo_add_1_qelse_or_m1c OR (fsm_output(7))) & or_tmp_792
      & and_1719_cse));
  mult_t_mul_cmp_15_z <= mult_t_mul_cmp_15_z_1;

  mult_z_mul_cmp : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_a,
      b => mult_z_mul_cmp_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_z_1
    );
  mult_z_mul_cmp_a <= MUX1HOT_v_32_3_2((xt_rsc_0_1_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_1_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_31_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( (fsm_output(2))
      & or_dcpl_194 & (fsm_output(7))));
  mult_z_mul_cmp_b <= MUX1HOT_v_32_9_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_8_i_qa_d(31
      DOWNTO 0)), (twiddle_rsc_0_9_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_10_i_qa_d(31
      DOWNTO 0)), (twiddle_rsc_0_11_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_12_i_qa_d(31
      DOWNTO 0)), (twiddle_rsc_0_13_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_14_i_qa_d(31
      DOWNTO 0)), (twiddle_rsc_0_15_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( or_tmp_771
      & mult_15_t_and_44_cse & mult_15_t_and_45_cse & mult_15_t_and_46_cse & mult_15_t_and_47_cse
      & mult_15_t_and_48_cse & mult_15_t_and_50_cse & mult_15_t_and_52_cse & mult_15_t_and_54_cse));
  mult_z_mul_cmp_z <= mult_z_mul_cmp_z_1;

  mult_z_mul_cmp_1 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_1_a,
      b => mult_z_mul_cmp_1_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_1_z_1
    );
  mult_z_mul_cmp_1_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_1_z(63 DOWNTO 32)), (mult_t_mul_cmp_11_z(63
      DOWNTO 32)), (mult_t_mul_cmp_12_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_1_b <= p_sva;
  mult_z_mul_cmp_1_z <= mult_z_mul_cmp_1_z_1;

  mult_z_mul_cmp_2 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_2_a,
      b => mult_z_mul_cmp_2_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_2_z_1
    );
  mult_z_mul_cmp_2_a <= MUX1HOT_v_32_4_2((xt_rsc_0_31_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_31_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_1_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_17_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_z_mul_cmp_2_b <= MUX_v_32_2_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_8_i_qa_d(31
      DOWNTO 0)), fsm_output(9));
  mult_z_mul_cmp_2_z <= mult_z_mul_cmp_2_z_1;

  mult_z_mul_cmp_3 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_3_a,
      b => mult_z_mul_cmp_3_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_3_z_1
    );
  mult_z_mul_cmp_3_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_2_z(63 DOWNTO 32)), (mult_t_mul_cmp_5_z(63
      DOWNTO 32)), (mult_t_mul_cmp_6_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_3_b <= p_sva;
  mult_z_mul_cmp_3_z <= mult_z_mul_cmp_3_z_1;

  mult_z_mul_cmp_4 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_4_a,
      b => mult_z_mul_cmp_4_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_4_z_1
    );
  mult_z_mul_cmp_4_a <= MUX1HOT_v_32_3_2((xt_rsc_0_29_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_29_i_qa_d(31
      DOWNTO 0)), (yt_rsc_0_9_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( or_dcpl_210
      & (fsm_output(4)) & (fsm_output(9))));
  mult_z_mul_cmp_4_b <= MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_8_i_qa_d(31
      DOWNTO 0)), (twiddle_rsc_0_10_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_12_i_qa_d(31
      DOWNTO 0)), (twiddle_rsc_0_14_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_4_i_qa_d(31
      DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & mult_15_t_and_40_cse
      & mult_15_t_and_41_cse & mult_15_t_and_42_cse & mult_15_t_and_43_cse & (fsm_output(9))));
  mult_z_mul_cmp_4_z <= mult_z_mul_cmp_4_z_1;

  mult_z_mul_cmp_5 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_5_a,
      b => mult_z_mul_cmp_5_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_5_z_1
    );
  mult_z_mul_cmp_5_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_3_z(63 DOWNTO 32)), (mult_t_mul_cmp_12_z(63
      DOWNTO 32)), (mult_t_mul_cmp_13_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_5_b <= p_sva;
  mult_z_mul_cmp_5_z <= mult_z_mul_cmp_5_z_1;

  mult_z_mul_cmp_6 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_6_a,
      b => mult_z_mul_cmp_6_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_6_z_1
    );
  mult_z_mul_cmp_6_a <= MUX1HOT_v_32_4_2((xt_rsc_0_27_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_27_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_15_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_31_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_z_mul_cmp_6_b <= MUX1HOT_v_32_12_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_1_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_2_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_3_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_4_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_5_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_6_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_7_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_12_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_13_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_14_i_qa_d(31 DOWNTO
      0)), (twiddle_rsc_0_15_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( mult_15_t_or_3_cse
      & mult_15_t_and_45_cse & mult_15_t_and_46_cse & mult_15_t_and_47_cse & mult_15_t_and_48_cse
      & mult_15_t_and_50_cse & mult_15_t_and_52_cse & mult_15_t_and_54_cse & mult_15_t_and_49_cse
      & mult_15_t_and_51_cse & mult_15_t_and_53_cse & mult_15_t_and_55_cse));
  mult_z_mul_cmp_6_z <= mult_z_mul_cmp_6_z_1;

  mult_z_mul_cmp_7 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_7_a,
      b => mult_z_mul_cmp_7_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_7_z_1
    );
  mult_z_mul_cmp_7_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_4_z(63 DOWNTO 32)), (mult_t_mul_cmp_2_z(63
      DOWNTO 32)), (mult_t_mul_cmp_3_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_7_b <= p_sva;
  mult_z_mul_cmp_7_z <= mult_z_mul_cmp_7_z_1;

  mult_z_mul_cmp_8 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_8_a,
      b => mult_z_mul_cmp_8_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_8_z_1
    );
  mult_z_mul_cmp_8_a <= MUX1HOT_v_32_4_2((xt_rsc_0_25_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_25_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_3_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_19_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_z_mul_cmp_8_b <= MUX1HOT_v_32_4_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_1_i_qa_d(31
      DOWNTO 0)), (twiddle_rsc_0_9_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_8_i_qa_d(31
      DOWNTO 0)), STD_LOGIC_VECTOR'( or_tmp_894 & or_tmp_819 & or_tmp_782 & and_1700_cse));
  mult_z_mul_cmp_8_z <= mult_z_mul_cmp_8_z_1;

  mult_z_mul_cmp_9 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_9_a,
      b => mult_z_mul_cmp_9_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_9_z_1
    );
  mult_z_mul_cmp_9_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_5_z(63 DOWNTO 32)), (mult_t_mul_cmp_10_z(63
      DOWNTO 32)), (mult_t_mul_cmp_11_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_9_b <= p_sva;
  mult_z_mul_cmp_9_z <= mult_z_mul_cmp_9_z_1;

  mult_z_mul_cmp_10 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_10_a,
      b => mult_z_mul_cmp_10_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_10_z_1
    );
  mult_z_mul_cmp_10_a <= MUX1HOT_v_32_4_2((xt_rsc_0_23_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_23_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_17_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_15_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_z_mul_cmp_10_b <= MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_8_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_4_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_5_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_6_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_7_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & mult_15_t_and_49_cse & mult_15_t_and_51_cse & mult_15_t_and_53_cse
      & mult_15_t_and_55_cse));
  mult_z_mul_cmp_10_z <= mult_z_mul_cmp_10_z_1;

  mult_z_mul_cmp_11 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_11_a,
      b => mult_z_mul_cmp_11_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_11_z_1
    );
  mult_z_mul_cmp_11_a <= MUX_v_32_2_2((mult_t_mul_cmp_6_z(63 DOWNTO 32)), (mult_t_mul_cmp_7_z(63
      DOWNTO 32)), fsm_output(9));
  mult_z_mul_cmp_11_b <= p_sva;
  mult_z_mul_cmp_11_z <= mult_z_mul_cmp_11_z_1;

  mult_z_mul_cmp_12 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_12_a,
      b => mult_z_mul_cmp_12_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_12_z_1
    );
  mult_z_mul_cmp_12_a <= MUX1HOT_v_32_4_2((xt_rsc_0_21_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_21_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_5_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_7_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_z_mul_cmp_12_b <= MUX1HOT_v_32_4_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_2_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_1_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_3_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( (or_tmp_885 OR mult_15_t_and_49_cse)
      & (or_tmp_809 OR mult_15_t_and_53_cse) & mult_15_t_and_51_cse & mult_15_t_and_55_cse));
  mult_z_mul_cmp_12_z <= mult_z_mul_cmp_12_z_1;

  mult_z_mul_cmp_13 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_13_a,
      b => mult_z_mul_cmp_13_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_13_z_1
    );
  mult_z_mul_cmp_13_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_7_z(63 DOWNTO 32)), (mult_t_mul_cmp_1_z(63
      DOWNTO 32)), (mult_t_mul_cmp_2_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_13_b <= p_sva;
  mult_z_mul_cmp_13_z <= mult_z_mul_cmp_13_z_1;

  mult_z_mul_cmp_14 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_14_a,
      b => mult_z_mul_cmp_14_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_14_z_1
    );
  mult_z_mul_cmp_14_a <= MUX1HOT_v_32_4_2((xt_rsc_0_19_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_19_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_27_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_29_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_z_mul_cmp_14_b <= MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_8_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_9_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_12_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_13_i_qa_d(31 DOWNTO
      0)), (twiddle_rsc_0_14_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & mult_15_t_and_36_cse & mult_15_t_and_37_cse & (mult_15_t_and_38_cse OR and_1719_cse)
      & mult_15_t_and_39_cse & or_tmp_792));
  mult_z_mul_cmp_14_z <= mult_z_mul_cmp_14_z_1;

  mult_z_mul_cmp_15 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_15_a,
      b => mult_z_mul_cmp_15_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_15_z_1
    );
  mult_z_mul_cmp_15_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_8_z(63 DOWNTO 32)), (mult_t_mul_cmp_13_z(63
      DOWNTO 32)), (mult_t_mul_cmp_14_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_15_b <= p_sva;
  mult_z_mul_cmp_15_z <= mult_z_mul_cmp_15_z_1;

  mult_z_mul_cmp_16 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_16_a,
      b => mult_z_mul_cmp_16_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_16_z_1
    );
  mult_z_mul_cmp_16_a <= MUX1HOT_v_32_4_2((xt_rsc_0_17_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_17_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_13_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_3_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_z_mul_cmp_16_b <= MUX1HOT_v_32_5_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_2_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_4_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_6_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_1_i_qa_d(31 DOWNTO 0)),
      STD_LOGIC_VECTOR'( (or_tmp_779 OR mult_15_t_and_40_cse) & mult_15_t_and_41_cse
      & mult_15_t_and_42_cse & mult_15_t_and_43_cse & or_tmp_782));
  mult_z_mul_cmp_16_z <= mult_z_mul_cmp_16_z_1;

  mult_z_mul_cmp_17 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_17_a,
      b => mult_z_mul_cmp_17_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_17_z_1
    );
  mult_z_mul_cmp_17_a <= MUX_v_32_2_2((mult_t_mul_cmp_9_z(63 DOWNTO 32)), (mult_t_mul_cmp_10_z(63
      DOWNTO 32)), fsm_output(9));
  mult_z_mul_cmp_17_b <= p_sva;
  mult_z_mul_cmp_17_z <= mult_z_mul_cmp_17_z_1;

  mult_z_mul_cmp_18 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_18_a,
      b => mult_z_mul_cmp_18_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_18_z_1
    );
  mult_z_mul_cmp_18_a <= MUX1HOT_v_32_4_2((xt_rsc_0_15_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_15_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_19_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_21_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_z_mul_cmp_18_b <= MUX1HOT_v_32_4_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_9_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_8_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_10_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & or_tmp_819 & (and_1783_cse OR and_1719_cse) & or_tmp_792));
  mult_z_mul_cmp_18_z <= mult_z_mul_cmp_18_z_1;

  mult_z_mul_cmp_19 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_19_a,
      b => mult_z_mul_cmp_19_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_19_z_1
    );
  mult_z_mul_cmp_19_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_10_z(63 DOWNTO 32)), (mult_t_mul_cmp_4_z(63
      DOWNTO 32)), (mult_t_mul_cmp_5_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_19_b <= p_sva;
  mult_z_mul_cmp_19_z <= mult_z_mul_cmp_19_z_1;

  mult_z_mul_cmp_20 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_20_a,
      b => mult_z_mul_cmp_20_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_20_z_1
    );
  mult_z_mul_cmp_20_a <= MUX1HOT_v_32_4_2((xt_rsc_0_13_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_13_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_25_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_11_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_z_mul_cmp_20_b <= MUX1HOT_v_32_5_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_12_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_8_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_5_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_4_i_qa_d(31 DOWNTO 0)),
      STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & or_tmp_790 & and_1725_cse &
      or_tmp_782 & and_1700_cse));
  mult_z_mul_cmp_20_z <= mult_z_mul_cmp_20_z_1;

  mult_z_mul_cmp_21 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_21_a,
      b => mult_z_mul_cmp_21_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_21_z_1
    );
  mult_z_mul_cmp_21_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_11_z(63 DOWNTO 32)), (mult_t_mul_cmp_14_z(63
      DOWNTO 32)), (mult_t_mul_cmp_15_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_21_b <= p_sva;
  mult_z_mul_cmp_21_z <= mult_z_mul_cmp_21_z_1;

  mult_z_mul_cmp_22 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_22_a,
      b => mult_z_mul_cmp_22_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_22_z_1
    );
  mult_z_mul_cmp_22_a <= MUX1HOT_v_32_3_2((xt_rsc_0_11_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_11_i_qa_d(31
      DOWNTO 0)), (yt_rsc_0_27_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( or_dcpl_210
      & (fsm_output(4)) & (fsm_output(9))));
  mult_z_mul_cmp_22_b <= MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_1_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_4_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_5_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_13_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_12_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( mult_15_t_or_1_cse
      & mult_15_t_and_37_cse & mult_15_t_and_38_cse & mult_15_t_and_39_cse & or_tmp_782
      & and_1700_cse));
  mult_z_mul_cmp_22_z <= mult_z_mul_cmp_22_z_1;

  mult_z_mul_cmp_23 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_23_a,
      b => mult_z_mul_cmp_23_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_23_z_1
    );
  mult_z_mul_cmp_23_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_12_z(63 DOWNTO 32)), (mult_t_mul_cmp_3_z(63
      DOWNTO 32)), (mult_t_mul_cmp_4_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_23_b <= p_sva;
  mult_z_mul_cmp_23_z <= mult_z_mul_cmp_23_z_1;

  mult_z_mul_cmp_24 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_24_a,
      b => mult_z_mul_cmp_24_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_24_z_1
    );
  mult_z_mul_cmp_24_a <= mult_4_t_mux1h_1_rmff;
  mult_z_mul_cmp_24_b <= MUX1HOT_v_32_8_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_1_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_2_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_3_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_8_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_9_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_10_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_11_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( mult_15_t_or_cse
      & mult_15_t_and_30_cse & mult_15_t_and_31_cse & mult_15_t_and_32_cse & mult_15_t_and_49_cse
      & mult_15_t_and_51_cse & mult_15_t_and_53_cse & mult_15_t_and_55_cse));
  mult_z_mul_cmp_24_z <= mult_z_mul_cmp_24_z_1;

  mult_z_mul_cmp_25 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_25_a,
      b => mult_z_mul_cmp_25_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_25_z_1
    );
  mult_z_mul_cmp_25_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_13_z(63 DOWNTO 32)), (mult_t_mul_cmp_8_z(63
      DOWNTO 32)), (mult_t_mul_cmp_9_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_25_b <= p_sva;
  mult_z_mul_cmp_25_z <= mult_z_mul_cmp_25_z_1;

  mult_z_mul_cmp_26 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_26_a,
      b => mult_z_mul_cmp_26_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_26_z_1
    );
  mult_z_mul_cmp_26_a <= MUX1HOT_v_32_4_2((xt_rsc_0_7_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_7_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_21_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_13_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_z_mul_cmp_26_b <= MUX1HOT_v_32_5_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_10_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_8_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_6_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_4_i_qa_d(31 DOWNTO 0)),
      STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & or_tmp_809 & and_1763_cse &
      or_tmp_792 & and_1719_cse));
  mult_z_mul_cmp_26_z <= mult_z_mul_cmp_26_z_1;

  mult_z_mul_cmp_27 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_27_a,
      b => mult_z_mul_cmp_27_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_27_z_1
    );
  mult_z_mul_cmp_27_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_14_z(63 DOWNTO 32)), (mult_t_mul_cmp_7_z(63
      DOWNTO 32)), (mult_t_mul_cmp_8_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_27_b <= p_sva;
  mult_z_mul_cmp_27_z <= mult_z_mul_cmp_27_z_1;

  mult_z_mul_cmp_28 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_28_a,
      b => mult_z_mul_cmp_28_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_28_z_1
    );
  mult_z_mul_cmp_28_a <= MUX1HOT_v_32_3_2((xt_rsc_0_5_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_5_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_9_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( (fsm_output(2))
      & or_dcpl_194 & (fsm_output(7))));
  mult_z_mul_cmp_28_b <= MUX1HOT_v_32_3_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_4_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_2_i_qa_d(31 DOWNTO 0)),
      STD_LOGIC_VECTOR'( (and_1725_cse OR and_1719_cse OR modulo_add_1_qelse_or_m1c)
      & or_tmp_790 & or_tmp_792));
  mult_z_mul_cmp_28_z <= mult_z_mul_cmp_28_z_1;

  mult_z_mul_cmp_29 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_29_a,
      b => mult_z_mul_cmp_29_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_29_z_1
    );
  mult_z_mul_cmp_29_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_15_z(63 DOWNTO 32)), (mult_t_mul_cmp_z(63
      DOWNTO 32)), (mult_t_mul_cmp_1_z(63 DOWNTO 32)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & (fsm_output(7)) & (fsm_output(9))));
  mult_z_mul_cmp_29_b <= p_sva;
  mult_z_mul_cmp_29_z <= mult_z_mul_cmp_29_z_1;

  mult_z_mul_cmp_30 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_30_a,
      b => mult_z_mul_cmp_30_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_30_z_1
    );
  mult_z_mul_cmp_30_a <= MUX1HOT_v_32_4_2((xt_rsc_0_3_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_3_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_23_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_25_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_z_mul_cmp_30_b <= MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_8_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_9_i_qa_d(31 DOWNTO 0)),
      (twiddle_rsc_0_10_i_qa_d(31 DOWNTO 0)), (twiddle_rsc_0_11_i_qa_d(31 DOWNTO
      0)), (twiddle_rsc_0_12_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c
      & mult_15_t_and_29_cse & mult_15_t_and_30_cse & mult_15_t_and_31_cse & mult_15_t_and_32_cse
      & (fsm_output(9))));
  mult_z_mul_cmp_30_z <= mult_z_mul_cmp_30_z_1;

  mult_z_mul_cmp_31 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 3,
      n_inreg => 1
      )
    PORT MAP(
      a => mult_z_mul_cmp_31_a,
      b => mult_z_mul_cmp_31_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_31_z_1
    );
  mult_z_mul_cmp_31_a <= MUX_v_32_2_2((mult_t_mul_cmp_z(63 DOWNTO 32)), (mult_t_mul_cmp_15_z(63
      DOWNTO 32)), fsm_output(7));
  mult_z_mul_cmp_31_b <= p_sva;
  mult_z_mul_cmp_31_z <= mult_z_mul_cmp_31_z_1;

  operator_33_true_3_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_bl_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 1,
      width_s => 3,
      width_z => 2
      )
    PORT MAP(
      a => operator_33_true_3_lshift_rg_a,
      s => operator_33_true_3_lshift_rg_s,
      z => operator_33_true_3_lshift_rg_z
    );
  operator_33_true_3_lshift_rg_a(0) <= '1';
  operator_33_true_3_lshift_rg_s <= STD_LOGIC_VECTOR'( '0' & (NOT c_1_sva) & '0');
  operator_33_true_3_lshift_psp_1_0_sva_mx0w3 <= operator_33_true_3_lshift_rg_z;

  operator_33_true_1_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_l_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 1,
      width_s => 4,
      width_z => 11
      )
    PORT MAP(
      a => operator_33_true_1_lshift_rg_a,
      s => operator_33_true_1_lshift_rg_s,
      z => operator_33_true_1_lshift_rg_z
    );
  operator_33_true_1_lshift_rg_a(0) <= '1';
  operator_33_true_1_lshift_rg_s <= (MUX1HOT_v_3_3_2(z_out_1, operator_20_false_acc_cse_sva,
      (STD_LOGIC_VECTOR'( "00") & (NOT c_1_sva)), STD_LOGIC_VECTOR'( (fsm_output(1))
      & (fsm_output(3)) & (fsm_output(6))))) & ((NOT (fsm_output(3))) OR (fsm_output(1))
      OR (fsm_output(6)));
  z_out <= operator_33_true_1_lshift_rg_z;

  peaseNTT_core_wait_dp_inst : peaseNTT_core_wait_dp
    PORT MAP(
      yt_rsc_0_0_cgo_iro => or_261_rmff,
      yt_rsc_0_0_i_clka_en_d => yt_rsc_0_0_i_clka_en_d,
      yt_rsc_0_16_cgo_iro => or_443_rmff,
      yt_rsc_0_16_i_clka_en_d => yt_rsc_0_16_i_clka_en_d,
      ensig_cgo_iro => or_997_rmff,
      ensig_cgo_iro_17 => or_1156_rmff,
      yt_rsc_0_0_cgo => reg_yt_rsc_0_0_cgo_cse,
      yt_rsc_0_16_cgo => reg_yt_rsc_0_16_cgo_cse,
      ensig_cgo => reg_ensig_cgo_cse,
      mult_t_mul_cmp_en => mult_t_mul_cmp_en,
      ensig_cgo_17 => reg_ensig_cgo_17_cse,
      mult_z_mul_cmp_1_en => mult_z_mul_cmp_1_en
    );
  peaseNTT_core_core_fsm_inst : peaseNTT_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      fsm_output => peaseNTT_core_core_fsm_inst_fsm_output,
      INNER_LOOP1_C_0_tr0 => peaseNTT_core_core_fsm_inst_INNER_LOOP1_C_0_tr0,
      INNER_LOOP2_C_0_tr0 => INNER_LOOP4_nor_tmp,
      STAGE_LOOP_C_2_tr0 => peaseNTT_core_core_fsm_inst_STAGE_LOOP_C_2_tr0,
      INNER_LOOP3_C_0_tr0 => INNER_LOOP4_nor_tmp,
      INNER_LOOP4_C_0_tr0 => and_dcpl_51,
      INNER_LOOP4_C_0_tr1 => peaseNTT_core_core_fsm_inst_INNER_LOOP4_C_0_tr1
    );
  fsm_output <= peaseNTT_core_core_fsm_inst_fsm_output;
  peaseNTT_core_core_fsm_inst_INNER_LOOP1_C_0_tr0 <= NOT(INNER_LOOP1_stage_0 OR INNER_LOOP1_stage_0_2
      OR INNER_LOOP1_stage_0_3 OR INNER_LOOP1_stage_0_4 OR INNER_LOOP1_stage_0_5
      OR INNER_LOOP1_stage_0_6 OR INNER_LOOP1_stage_0_7 OR INNER_LOOP1_stage_0_8
      OR INNER_LOOP1_stage_0_9 OR INNER_LOOP1_stage_0_10);
  peaseNTT_core_core_fsm_inst_STAGE_LOOP_C_2_tr0 <= z_out_1(2);
  peaseNTT_core_core_fsm_inst_INNER_LOOP4_C_0_tr1 <= NOT INNER_LOOP4_nor_tmp;

  or_261_rmff <= ((and_dcpl_57 OR and_dcpl_56 OR ((NOT INNER_LOOP1_stage_0_10) AND
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8)) AND (fsm_output(7))) OR
      and_167_cse OR (((INNER_LOOP1_stage_0_11 AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10))
      OR and_dcpl_59 OR and_dcpl_58) AND (fsm_output(2)));
  and_202_rmff <= INNER_LOOP1_stage_0 AND or_dcpl_194;
  or_443_rmff <= ((and_dcpl_68 OR and_dcpl_67 OR (INNER_LOOP1_stage_0_10 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8))
      AND (fsm_output(7))) OR and_167_cse OR (((INNER_LOOP1_stage_0_11 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10)
      OR and_dcpl_70 OR and_dcpl_69) AND (fsm_output(2)));
  and_921_rmff <= INNER_LOOP1_stage_0 AND or_dcpl_210;
  and_1435_rmff <= INNER_LOOP1_stage_0 AND or_dcpl_214;
  butterFly2_1_tw_butterFly2_1_tw_mux_rmff <= MUX_v_7_2_2(INNER_LOOP3_r_11_4_sva_6_0,
      INNER_LOOP4_r_11_4_sva_6_0, fsm_output(9));
  or_896_rmff <= (and_dcpl_79 AND (fsm_output(7))) OR and_1445_cse;
  or_900_rmff <= (and_dcpl_81 AND (fsm_output(7))) OR and_1454_cse;
  or_904_rmff <= (and_dcpl_79 AND (operator_20_false_acc_cse_sva(1)) AND (fsm_output(7)))
      OR and_1463_cse;
  or_908_rmff <= (INNER_LOOP1_stage_0 AND (operator_20_false_acc_cse_sva(2)) AND
      (fsm_output(7))) OR (INNER_LOOP1_stage_0 AND (fsm_output(9)));
  or_912_rmff <= (and_dcpl_79 AND (operator_20_false_acc_cse_sva(2)) AND (fsm_output(7)))
      OR and_1445_cse;
  or_916_rmff <= (and_dcpl_81 AND (operator_20_false_acc_cse_sva(2)) AND (fsm_output(7)))
      OR and_1454_cse;
  or_920_rmff <= (and_dcpl_79 AND CONV_SL_1_1(operator_20_false_acc_cse_sva(2 DOWNTO
      1)=STD_LOGIC_VECTOR'("11")) AND (fsm_output(7))) OR and_1463_cse;
  and_1506_rmff <= INNER_LOOP1_stage_0 AND or_dcpl_212;
  or_997_rmff <= ((INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2
      OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1) AND or_dcpl_218) OR ((INNER_LOOP1_stage_0_4
      OR INNER_LOOP1_stage_0_2 OR INNER_LOOP1_stage_0_3) AND (fsm_output(2)));
  mult_15_t_and_49_cse <= CONV_SL_1_1(operator_33_true_3_lshift_psp_1_0_sva=STD_LOGIC_VECTOR'("00"))
      AND (fsm_output(9));
  mult_15_t_and_51_cse <= CONV_SL_1_1(operator_33_true_3_lshift_psp_1_0_sva=STD_LOGIC_VECTOR'("01"))
      AND (fsm_output(9));
  mult_15_t_and_53_cse <= CONV_SL_1_1(operator_33_true_3_lshift_psp_1_0_sva=STD_LOGIC_VECTOR'("10"))
      AND (fsm_output(9));
  mult_15_t_and_55_cse <= CONV_SL_1_1(operator_33_true_3_lshift_psp_1_0_sva=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(9));
  mult_15_t_and_44_cse <= butterFly2_15_tw_equal_tmp_1 AND (fsm_output(7));
  butterFly2_7_tw_nor_cse <= NOT(CONV_SL_1_1(operator_20_false_acc_cse_sva(2 DOWNTO
      1)/=STD_LOGIC_VECTOR'("00")));
  mult_15_t_and_45_cse <= (operator_20_false_acc_cse_sva(0)) AND butterFly2_7_tw_nor_cse
      AND (fsm_output(7));
  butterFly2_7_tw_nor_1_cse <= NOT((operator_20_false_acc_cse_sva(2)) OR (operator_20_false_acc_cse_sva(0)));
  mult_15_t_and_46_cse <= (operator_20_false_acc_cse_sva(1)) AND butterFly2_7_tw_nor_1_cse
      AND (fsm_output(7));
  mult_15_t_and_47_cse <= butterFly2_15_tw_equal_tmp_3_1 AND (fsm_output(7));
  butterFly2_7_tw_nor_2_cse <= NOT(CONV_SL_1_1(operator_20_false_acc_cse_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("00")));
  mult_15_t_and_48_cse <= (operator_20_false_acc_cse_sva(2)) AND butterFly2_7_tw_nor_2_cse
      AND (fsm_output(7));
  mult_15_t_and_50_cse <= butterFly2_15_tw_equal_tmp_5_1 AND (fsm_output(7));
  mult_15_t_and_52_cse <= butterFly2_15_tw_equal_tmp_6_1 AND (fsm_output(7));
  mult_15_t_and_54_cse <= butterFly2_15_tw_equal_tmp_7_1 AND (fsm_output(7));
  mult_15_t_or_9_cse <= mult_15_t_and_48_cse OR mult_15_t_and_49_cse;
  mult_15_t_or_10_cse <= mult_15_t_and_50_cse OR mult_15_t_and_51_cse;
  mult_15_t_or_11_cse <= mult_15_t_and_52_cse OR mult_15_t_and_53_cse;
  mult_15_t_or_12_cse <= mult_15_t_and_54_cse OR mult_15_t_and_55_cse;
  mult_15_t_and_41_cse <= CONV_SL_1_1(operator_20_false_acc_cse_sva(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"))
      AND (fsm_output(7));
  mult_15_t_and_42_cse <= CONV_SL_1_1(operator_20_false_acc_cse_sva(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10"))
      AND (fsm_output(7));
  mult_15_t_and_43_cse <= CONV_SL_1_1(operator_20_false_acc_cse_sva(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(7));
  mult_15_t_and_40_cse <= butterFly2_7_tw_nor_cse AND (fsm_output(7));
  mult_15_t_and_37_cse <= (operator_20_false_acc_cse_sva(0)) AND (NOT (operator_20_false_acc_cse_sva(2)))
      AND (fsm_output(7));
  mult_15_t_and_38_cse <= (operator_20_false_acc_cse_sva(2)) AND (NOT (operator_20_false_acc_cse_sva(0)))
      AND (fsm_output(7));
  mult_15_t_and_39_cse <= (operator_20_false_acc_cse_sva(2)) AND (operator_20_false_acc_cse_sva(0))
      AND (fsm_output(7));
  mult_15_t_and_36_cse <= butterFly2_7_tw_nor_1_cse AND (fsm_output(7));
  mult_15_t_and_30_cse <= CONV_SL_1_1(operator_20_false_acc_cse_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND (fsm_output(7));
  mult_15_t_and_31_cse <= CONV_SL_1_1(operator_20_false_acc_cse_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND (fsm_output(7));
  mult_15_t_and_32_cse <= CONV_SL_1_1(operator_20_false_acc_cse_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(7));
  mult_15_t_and_29_cse <= butterFly2_7_tw_nor_2_cse AND (fsm_output(7));
  mult_15_t_or_3_cse <= modulo_add_1_qelse_or_m1c OR mult_15_t_and_44_cse;
  mult_15_t_or_1_cse <= modulo_add_1_qelse_or_m1c OR mult_15_t_and_36_cse;
  mult_4_t_mux1h_1_rmff <= MUX1HOT_v_32_4_2((xt_rsc_0_9_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_9_i_qa_d(31
      DOWNTO 0)), (xt_rsc_0_7_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_23_i_qa_d(31 DOWNTO
      0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  mult_15_t_or_cse <= modulo_add_1_qelse_or_m1c OR mult_15_t_and_29_cse;
  or_1156_rmff <= ((INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4
      OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3) AND or_dcpl_218) OR ((INNER_LOOP1_stage_0_6
      OR INNER_LOOP1_stage_0_7 OR INNER_LOOP1_stage_0_5) AND (fsm_output(2)));
  modulo_add_1_qelse_or_m1c <= (fsm_output(2)) OR (fsm_output(4));
  or_12_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 OR INNER_LOOP1_stage_0_9;
  or_44_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 OR INNER_LOOP1_stage_0_8;
  or_64_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 OR INNER_LOOP1_stage_0_7;
  or_84_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 OR INNER_LOOP1_stage_0_6;
  or_103_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 OR INNER_LOOP1_stage_0_5;
  or_123_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 OR INNER_LOOP1_stage_0_4;
  or_142_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm OR INNER_LOOP1_stage_0_3;
  or_143_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm OR INNER_LOOP1_stage_0_2;
  modulo_sub_16_qelse_and_ssc <= NOT((z_out_66(31)) OR (fsm_output(9)));
  modulo_sub_16_qelse_and_ssc_1 <= (NOT (z_out_51(31))) AND (fsm_output(9));
  modulo_sub_17_qelse_and_ssc <= NOT((z_out_56(31)) OR (fsm_output(9)));
  modulo_sub_17_qelse_and_ssc_1 <= (NOT (z_out_52(31))) AND (fsm_output(9));
  modulo_sub_18_qelse_and_ssc <= NOT((z_out_63(31)) OR (fsm_output(9)));
  modulo_sub_18_qelse_and_ssc_1 <= (NOT (z_out_53(31))) AND (fsm_output(9));
  modulo_sub_19_qelse_and_ssc <= NOT((z_out_64(31)) OR (fsm_output(9)));
  modulo_sub_19_qelse_and_ssc_1 <= (NOT (z_out_54(31))) AND (fsm_output(9));
  modulo_sub_20_qelse_and_ssc <= NOT((z_out_65(31)) OR (fsm_output(9)));
  modulo_sub_20_qelse_and_ssc_1 <= (NOT (z_out_55(31))) AND (fsm_output(9));
  modulo_sub_21_qelse_and_ssc <= NOT((z_out_51(31)) OR (fsm_output(9)));
  modulo_sub_21_qelse_and_ssc_1 <= (NOT (z_out_56(31))) AND (fsm_output(9));
  modulo_sub_22_qelse_and_ssc <= NOT((z_out_52(31)) OR (fsm_output(9)));
  modulo_sub_22_qelse_and_ssc_1 <= (NOT (z_out_57(31))) AND (fsm_output(9));
  modulo_sub_23_qelse_and_ssc <= NOT((z_out_53(31)) OR (fsm_output(9)));
  modulo_sub_23_qelse_and_ssc_1 <= (NOT (z_out_58(31))) AND (fsm_output(9));
  modulo_sub_24_qelse_and_ssc <= NOT((z_out_54(31)) OR (fsm_output(9)));
  modulo_sub_24_qelse_and_ssc_1 <= (NOT (z_out_59(31))) AND (fsm_output(9));
  modulo_sub_25_qelse_and_ssc <= NOT((z_out_55(31)) OR (fsm_output(9)));
  modulo_sub_25_qelse_and_ssc_1 <= (NOT (z_out_60(31))) AND (fsm_output(9));
  modulo_sub_26_qelse_and_ssc <= NOT((z_out_57(31)) OR (fsm_output(9)));
  modulo_sub_26_qelse_and_ssc_1 <= (NOT (z_out_61(31))) AND (fsm_output(9));
  modulo_sub_27_qelse_and_ssc <= NOT((z_out_58(31)) OR (fsm_output(9)));
  modulo_sub_27_qelse_and_ssc_1 <= (NOT (z_out_62(31))) AND (fsm_output(9));
  modulo_sub_28_qelse_and_ssc <= NOT((z_out_59(31)) OR (fsm_output(9)));
  modulo_sub_28_qelse_and_ssc_1 <= (NOT (z_out_63(31))) AND (fsm_output(9));
  modulo_sub_29_qelse_and_ssc <= NOT((z_out_60(31)) OR (fsm_output(9)));
  modulo_sub_29_qelse_and_ssc_1 <= (NOT (z_out_64(31))) AND (fsm_output(9));
  modulo_sub_30_qelse_and_ssc <= NOT((z_out_61(31)) OR (fsm_output(9)));
  modulo_sub_30_qelse_and_ssc_1 <= (NOT (z_out_65(31))) AND (fsm_output(9));
  modulo_sub_31_qelse_and_ssc <= NOT((z_out_62(31)) OR (fsm_output(9)));
  modulo_sub_31_qelse_and_ssc_1 <= (NOT (z_out_66(31))) AND (fsm_output(9));
  yt_rsc_0_0_i_da_d_mx0w0_63_32 <= MUX_v_32_2_2(('0' & (z_out_51(30 DOWNTO 0))),
      z_out_20, z_out_51(31));
  yt_rsc_0_0_i_da_d_mx0w2_63_32 <= MUX_v_32_2_2(('0' & (z_out_65(30 DOWNTO 0))),
      z_out_18, z_out_65(31));
  yt_rsc_0_1_i_da_d_mx0w0_63_32 <= MUX_v_32_2_2(('0' & (z_out_52(30 DOWNTO 0))),
      z_out_17, z_out_52(31));
  yt_rsc_0_1_i_da_d_mx0w2_63_32 <= MUX_v_32_2_2(('0' & (z_out_66(30 DOWNTO 0))),
      z_out_16, z_out_66(31));
  yt_rsc_0_2_i_da_d_mx0w0_63_32 <= MUX_v_32_2_2(('0' & (z_out_53(30 DOWNTO 0))),
      z_out_14, z_out_53(31));
  yt_rsc_0_2_i_da_d_mx0w2_63_32 <= MUX_v_32_2_2(('0' & (z_out_51(30 DOWNTO 0))),
      z_out_13, z_out_51(31));
  yt_rsc_0_3_i_da_d_mx0w0_63_32 <= MUX_v_32_2_2(('0' & (z_out_54(30 DOWNTO 0))),
      z_out_12, z_out_54(31));
  yt_rsc_0_3_i_da_d_mx0w2_63_32 <= MUX_v_32_2_2(('0' & (z_out_52(30 DOWNTO 0))),
      z_out_10, z_out_52(31));
  yt_rsc_0_4_i_da_d_mx0w0_63_32 <= MUX_v_32_2_2(('0' & (z_out_55(30 DOWNTO 0))),
      z_out_9, z_out_55(31));
  yt_rsc_0_4_i_da_d_mx0w2_63_32 <= MUX_v_32_2_2(('0' & (z_out_53(30 DOWNTO 0))),
      z_out_8, z_out_53(31));
  modulo_sub_5_qif_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & (z_out_56(30
      DOWNTO 0))) + UNSIGNED(p_sva), 32));
  modulo_sub_5_qelse_mux_cse <= MUX_v_32_2_2(('0' & (z_out_56(30 DOWNTO 0))), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_sub_5_qif_acc_nl),
      32)), z_out_56(31));
  yt_rsc_0_5_i_da_d_mx0w2_63_32 <= MUX_v_32_2_2(('0' & (z_out_54(30 DOWNTO 0))),
      z_out_5, z_out_54(31));
  yt_rsc_0_6_i_da_d_mx0w0_63_32 <= MUX_v_32_2_2(('0' & (z_out_57(30 DOWNTO 0))),
      z_out_4, z_out_57(31));
  yt_rsc_0_6_i_da_d_mx0w2_63_32 <= MUX_v_32_2_2(('0' & (z_out_55(30 DOWNTO 0))),
      z_out_4, z_out_55(31));
  yt_rsc_0_7_i_da_d_mx0w0_63_32 <= MUX_v_32_2_2(('0' & (z_out_58(30 DOWNTO 0))),
      z_out_5, z_out_58(31));
  yt_rsc_0_8_i_da_d_mx0w0_63_32 <= MUX_v_32_2_2(('0' & (z_out_59(30 DOWNTO 0))),
      z_out_8, z_out_59(31));
  yt_rsc_0_8_i_da_d_mx0w2_63_32 <= MUX_v_32_2_2(('0' & (z_out_57(30 DOWNTO 0))),
      z_out_9, z_out_57(31));
  yt_rsc_0_9_i_da_d_mx0w0_63_32 <= MUX_v_32_2_2(('0' & (z_out_60(30 DOWNTO 0))),
      z_out_10, z_out_60(31));
  yt_rsc_0_9_i_da_d_mx0w2_63_32 <= MUX_v_32_2_2(('0' & (z_out_58(30 DOWNTO 0))),
      z_out_12, z_out_58(31));
  yt_rsc_0_10_i_da_d_mx0w0_63_32 <= MUX_v_32_2_2(('0' & (z_out_61(30 DOWNTO 0))),
      z_out_13, z_out_61(31));
  yt_rsc_0_10_i_da_d_mx0w2_63_32 <= MUX_v_32_2_2(('0' & (z_out_59(30 DOWNTO 0))),
      z_out_14, z_out_59(31));
  yt_rsc_0_11_i_da_d_mx0w0_63_32 <= MUX_v_32_2_2(('0' & (z_out_62(30 DOWNTO 0))),
      z_out_16, z_out_62(31));
  yt_rsc_0_11_i_da_d_mx0w2_63_32 <= MUX_v_32_2_2(('0' & (z_out_60(30 DOWNTO 0))),
      z_out_17, z_out_60(31));
  yt_rsc_0_12_i_da_d_mx0w0_63_32 <= MUX_v_32_2_2(('0' & (z_out_63(30 DOWNTO 0))),
      z_out_18, z_out_63(31));
  yt_rsc_0_12_i_da_d_mx0w2_63_32 <= MUX_v_32_2_2(('0' & (z_out_61(30 DOWNTO 0))),
      z_out_20, z_out_61(31));
  yt_rsc_0_13_i_da_d_mx0w0_63_32 <= MUX_v_32_2_2(('0' & (z_out_64(30 DOWNTO 0))),
      z_out_22, z_out_64(31));
  yt_rsc_0_13_i_da_d_mx0w2_63_32 <= MUX_v_32_2_2(('0' & (z_out_62(30 DOWNTO 0))),
      z_out_25, z_out_62(31));
  yt_rsc_0_14_i_da_d_mx0w0_63_32 <= MUX_v_32_2_2(('0' & (z_out_65(30 DOWNTO 0))),
      z_out_25, z_out_65(31));
  yt_rsc_0_14_i_da_d_mx0w2_63_32 <= MUX_v_32_2_2(('0' & (z_out_63(30 DOWNTO 0))),
      z_out_22, z_out_63(31));
  yt_rsc_0_15_i_da_d_mx0w0_63_32 <= MUX_v_32_2_2(('0' & (z_out_66(30 DOWNTO 0))),
      z_out_28, z_out_66(31));
  yt_rsc_0_15_i_da_d_mx0w2_63_32 <= MUX_v_32_2_2(('0' & (z_out_64(30 DOWNTO 0))),
      z_out_28, z_out_64(31));
  mult_15_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_15_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_31_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_15_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_15_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_15_if_acc_nl),
      32)), mult_15_res_sva_1, mult_31_acc_1_nl(32));
  mult_14_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_14_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_30_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_14_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_14_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_14_if_acc_nl),
      32)), mult_14_res_sva_1, mult_30_acc_1_nl(32));
  mult_13_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_13_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_29_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_13_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_13_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_13_if_acc_nl),
      32)), mult_13_res_sva_1, mult_29_acc_1_nl(32));
  mult_12_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_12_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_28_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_12_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_12_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_12_if_acc_nl),
      32)), mult_12_res_sva_1, mult_28_acc_1_nl(32));
  mult_11_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_11_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_27_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_11_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_11_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_11_if_acc_nl),
      32)), mult_11_res_sva_1, mult_27_acc_1_nl(32));
  mult_10_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_10_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_26_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_10_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_10_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_10_if_acc_nl),
      32)), mult_10_res_sva_1, mult_26_acc_1_nl(32));
  mult_9_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_9_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_25_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_9_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_9_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_9_if_acc_nl),
      32)), mult_9_res_sva_1, mult_25_acc_1_nl(32));
  mult_8_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_8_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_24_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_8_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_8_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_8_if_acc_nl),
      32)), mult_8_res_sva_1, mult_24_acc_1_nl(32));
  mult_7_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_7_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_23_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_7_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_7_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_7_if_acc_nl),
      32)), mult_7_res_sva_1, mult_23_acc_1_nl(32));
  mult_6_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_6_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_22_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_6_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_6_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_6_if_acc_nl),
      32)), mult_6_res_sva_1, mult_22_acc_1_nl(32));
  mult_5_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_5_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_21_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_5_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_5_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_5_if_acc_nl),
      32)), mult_5_res_sva_1, mult_21_acc_1_nl(32));
  mult_4_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_4_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_20_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_4_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_4_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_4_if_acc_nl),
      32)), mult_4_res_sva_1, mult_20_acc_1_nl(32));
  mult_3_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_3_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_19_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_3_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_3_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_3_if_acc_nl),
      32)), mult_3_res_sva_1, mult_19_acc_1_nl(32));
  mult_2_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_2_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_18_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_2_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_2_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_2_if_acc_nl),
      32)), mult_2_res_sva_1, mult_18_acc_1_nl(32));
  mult_1_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_1_res_sva_1) -
      UNSIGNED(p_sva), 32));
  mult_17_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_1_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_1_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_1_if_acc_nl),
      32)), mult_1_res_sva_1, mult_17_acc_1_nl(32));
  mult_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_res_sva_1) - UNSIGNED(p_sva),
      32));
  mult_16_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_res_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_res_lpi_3_dfm_1_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_if_acc_nl),
      32)), mult_res_sva_1, mult_16_acc_1_nl(32));
  mult_15_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_15_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_1_z), 32));
  mult_14_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_14_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_3_z), 32));
  mult_13_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_13_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_5_z), 32));
  mult_12_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_12_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_7_z), 32));
  mult_11_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_11_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_9_z), 32));
  mult_10_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_10_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_11_z), 32));
  mult_9_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_25_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_13_z), 32));
  mult_8_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_24_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_15_z), 32));
  mult_7_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_23_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_17_z), 32));
  mult_6_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_22_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_19_z), 32));
  mult_5_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_21_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_21_z), 32));
  mult_4_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_20_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_23_z), 32));
  mult_3_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_19_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_25_z), 32));
  mult_2_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_18_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_27_z), 32));
  mult_1_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_17_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_29_z), 32));
  mult_res_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_16_z_asn_itm_3)
      - UNSIGNED(mult_z_mul_cmp_31_z), 32));
  INNER_LOOP4_nor_tmp <= NOT(INNER_LOOP1_stage_0 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm
      OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2
      OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4
      OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6
      OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10);
  or_dcpl_13 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 OR INNER_LOOP1_stage_0_8;
  or_dcpl_22 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 OR INNER_LOOP1_stage_0_7;
  or_dcpl_45 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 OR INNER_LOOP1_stage_0_6;
  or_dcpl_65 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 OR INNER_LOOP1_stage_0_5;
  or_dcpl_101 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 OR INNER_LOOP1_stage_0_4;
  or_dcpl_121 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 OR INNER_LOOP1_stage_0_3;
  and_dcpl_51 <= INNER_LOOP4_nor_tmp AND c_1_sva;
  and_dcpl_56 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 AND (NOT INNER_LOOP1_stage_0_9);
  and_dcpl_57 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10 AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9);
  or_dcpl_194 <= (fsm_output(4)) OR (fsm_output(9));
  and_dcpl_58 <= INNER_LOOP1_stage_0_9 AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8);
  and_dcpl_59 <= (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9) AND INNER_LOOP1_stage_0_10;
  or_dcpl_197 <= (NOT INNER_LOOP1_stage_0_9) OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8;
  or_dcpl_198 <= (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7) OR INNER_LOOP1_stage_0_9;
  or_dcpl_199 <= (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10) OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9;
  or_dcpl_200 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9 OR (NOT INNER_LOOP1_stage_0_10);
  and_dcpl_67 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 AND INNER_LOOP1_stage_0_9;
  and_dcpl_68 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9;
  and_dcpl_69 <= INNER_LOOP1_stage_0_9 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8;
  and_dcpl_70 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9 AND INNER_LOOP1_stage_0_10;
  or_dcpl_205 <= NOT(INNER_LOOP1_stage_0_9 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8);
  or_dcpl_206 <= NOT(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 AND INNER_LOOP1_stage_0_9);
  or_dcpl_207 <= NOT(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9);
  or_dcpl_208 <= NOT(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9 AND INNER_LOOP1_stage_0_10);
  or_dcpl_210 <= (fsm_output(2)) OR (fsm_output(7));
  or_dcpl_212 <= (fsm_output(7)) OR (fsm_output(9));
  or_dcpl_214 <= modulo_add_1_qelse_or_m1c OR or_dcpl_212;
  and_dcpl_79 <= INNER_LOOP1_stage_0 AND (operator_20_false_acc_cse_sva(0));
  and_dcpl_81 <= INNER_LOOP1_stage_0 AND (operator_20_false_acc_cse_sva(1));
  and_dcpl_82 <= INNER_LOOP1_stage_0 AND (operator_33_true_3_lshift_psp_1_0_sva(1));
  or_dcpl_217 <= (fsm_output(4)) OR (fsm_output(7));
  or_dcpl_218 <= or_dcpl_217 OR (fsm_output(9));
  and_dcpl_90 <= NOT((fsm_output(7)) OR (fsm_output(9)));
  or_dcpl_233 <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"));
  and_167_cse <= (INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm OR INNER_LOOP1_stage_0)
      AND or_dcpl_194;
  or_tmp_21 <= and_dcpl_58 AND (fsm_output(2));
  or_tmp_22 <= or_dcpl_197 AND (fsm_output(2));
  or_tmp_25 <= and_dcpl_56 AND (fsm_output(7));
  or_tmp_26 <= or_dcpl_198 AND (fsm_output(7));
  and_192_cse <= NOT((fsm_output(2)) OR (fsm_output(7)));
  or_tmp_203 <= and_dcpl_69 AND (fsm_output(2));
  or_tmp_204 <= or_dcpl_205 AND (fsm_output(2));
  or_tmp_207 <= and_dcpl_67 AND (fsm_output(7));
  or_tmp_208 <= or_dcpl_206 AND (fsm_output(7));
  nor_7_cse <= NOT((fsm_output(4)) OR (fsm_output(9)));
  and_1445_cse <= INNER_LOOP1_stage_0 AND (operator_33_true_3_lshift_psp_1_0_sva(0))
      AND (fsm_output(9));
  and_1454_cse <= and_dcpl_82 AND (fsm_output(9));
  and_1463_cse <= and_dcpl_82 AND (operator_33_true_3_lshift_psp_1_0_sva(0)) AND
      (fsm_output(9));
  or_tmp_771 <= modulo_add_1_qelse_or_m1c OR (fsm_output(9));
  and_1700_cse <= (NOT (operator_33_true_3_lshift_psp_1_0_sva(0))) AND (fsm_output(9));
  or_tmp_779 <= and_1700_cse OR modulo_add_1_qelse_or_m1c;
  or_tmp_782 <= (operator_33_true_3_lshift_psp_1_0_sva(0)) AND (fsm_output(9));
  and_1719_cse <= (NOT (operator_33_true_3_lshift_psp_1_0_sva(1))) AND (fsm_output(9));
  or_tmp_790 <= (operator_20_false_acc_cse_sva(2)) AND (fsm_output(7));
  and_1725_cse <= (NOT (operator_20_false_acc_cse_sva(2))) AND (fsm_output(7));
  or_tmp_792 <= (operator_33_true_3_lshift_psp_1_0_sva(1)) AND (fsm_output(9));
  or_tmp_809 <= (operator_20_false_acc_cse_sva(1)) AND (fsm_output(7));
  and_1763_cse <= (NOT (operator_20_false_acc_cse_sva(1))) AND (fsm_output(7));
  or_tmp_819 <= (operator_20_false_acc_cse_sva(0)) AND (fsm_output(7));
  and_1783_cse <= (NOT (operator_20_false_acc_cse_sva(0))) AND (fsm_output(7));
  or_tmp_885 <= and_1763_cse OR modulo_add_1_qelse_or_m1c;
  or_tmp_894 <= and_1783_cse OR modulo_add_1_qelse_or_m1c;
  or_tmp_1134 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  or_tmp_1138 <= (NOT (fsm_output(4))) AND (NOT (fsm_output(2))) AND and_dcpl_90;
  or_tmp_1189 <= (fsm_output(2)) OR (fsm_output(9));
  yt_rsc_0_0_i_wea_d_mx0c0 <= (or_dcpl_199 AND or_dcpl_198 AND (fsm_output(7))) OR
      and_192_cse OR (or_dcpl_200 AND or_dcpl_197 AND (fsm_output(2)));
  yt_rsc_0_0_i_wea_d_mx0c2 <= (and_dcpl_57 AND or_dcpl_198 AND (fsm_output(7))) OR
      (and_dcpl_59 AND or_dcpl_197 AND (fsm_output(2)));
  yt_rsc_0_16_i_wea_d_mx0c0 <= (or_dcpl_207 AND or_dcpl_206 AND (fsm_output(7)))
      OR and_192_cse OR (or_dcpl_208 AND or_dcpl_205 AND (fsm_output(2)));
  yt_rsc_0_16_i_wea_d_mx0c2 <= (and_dcpl_68 AND or_dcpl_206 AND (fsm_output(7)))
      OR (and_dcpl_70 AND or_dcpl_205 AND (fsm_output(2)));
  butterFly1_nor_7_rmff <= NOT(or_tmp_21 OR or_tmp_25);
  butterFly1_mux_17_cse <= MUX_s_1_2_2((INNER_LOOP2_r_11_4_sva_6_0(6)), (INNER_LOOP4_r_11_4_sva_6_0(6)),
      fsm_output(9));
  butterFly1_butterFly1_and_17_rmff <= butterFly1_mux_17_cse AND (NOT(or_tmp_21 OR
      or_tmp_22 OR or_tmp_25 OR or_tmp_26));
  butterFly1_or_5_cse <= or_tmp_25 OR or_tmp_26;
  butterFly1_or_1_cse <= or_tmp_21 OR or_tmp_22;
  butterFly1_mux1h_15_rmff <= MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_114_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_1_cse
      & (fsm_output(4)) & butterFly1_or_5_cse & (fsm_output(9))));
  butterFly1_1_mux1h_11_rmff <= MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_161_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_1_cse
      & (fsm_output(4)) & butterFly1_or_5_cse & (fsm_output(9))));
  butterFly1_2_mux1h_11_rmff <= MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_224_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_1_cse
      & (fsm_output(4)) & butterFly1_or_5_cse & (fsm_output(9))));
  butterFly1_3_mux1h_11_rmff <= MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_287_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_1_cse
      & (fsm_output(4)) & butterFly1_or_5_cse & (fsm_output(9))));
  butterFly1_4_mux1h_11_rmff <= MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_350_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_1_cse
      & (fsm_output(4)) & butterFly1_or_5_cse & (fsm_output(9))));
  butterFly1_8_mux1h_11_rmff <= MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_602_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_1_cse
      & (fsm_output(4)) & butterFly1_or_5_cse & (fsm_output(9))));
  butterFly1_nor_4_rmff <= NOT(or_tmp_203 OR or_tmp_207);
  butterFly1_butterFly1_and_15_rmff <= butterFly1_mux_17_cse AND (NOT(or_tmp_203
      OR or_tmp_204 OR or_tmp_207 OR or_tmp_208));
  butterFly1_or_4_cse <= or_tmp_207 OR or_tmp_208;
  butterFly1_or_cse <= or_tmp_203 OR or_tmp_204;
  butterFly1_mux1h_13_rmff <= MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_114_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_cse
      & (fsm_output(4)) & butterFly1_or_4_cse & (fsm_output(9))));
  butterFly1_1_mux1h_9_rmff <= MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_161_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_cse
      & (fsm_output(4)) & butterFly1_or_4_cse & (fsm_output(9))));
  butterFly1_2_mux1h_9_rmff <= MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_224_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_cse
      & (fsm_output(4)) & butterFly1_or_4_cse & (fsm_output(9))));
  butterFly1_3_mux1h_9_rmff <= MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_287_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_cse
      & (fsm_output(4)) & butterFly1_or_4_cse & (fsm_output(9))));
  butterFly1_4_mux1h_9_rmff <= MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_350_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_cse
      & (fsm_output(4)) & butterFly1_or_4_cse & (fsm_output(9))));
  butterFly1_8_mux1h_9_rmff <= MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_602_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_cse
      & (fsm_output(4)) & butterFly1_or_4_cse & (fsm_output(9))));
  butterFly1_15_f2_mux1h_65_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, ('0'
      & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_2), INNER_LOOP3_r_11_4_sva_6_0,
      ('1' & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_3), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_f1_butterFly1_f1_mux_2_rmff <= MUX_v_32_2_2((reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd
      & reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd_1), modulo_add_10_qr_lpi_3_dfm_1, fsm_output(9));
  butterFly1_f1_butterFly1_f1_mux_3_rmff <= MUX_v_32_2_2(modulo_add_10_qr_lpi_3_dfm_1,
      (reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd_1),
      fsm_output(9));
  butterFly1_15_f2_mux1h_64_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, ('0'
      & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_3), INNER_LOOP3_r_11_4_sva_6_0,
      ('1' & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_4), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_f2_butterFly1_f2_mux_2_rmff <= MUX_v_32_2_2((reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd
      & reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd_1), modulo_add_11_qr_lpi_3_dfm_1, fsm_output(9));
  butterFly1_f2_butterFly1_f2_mux_3_rmff <= MUX_v_32_2_2(modulo_add_11_qr_lpi_3_dfm_1,
      (reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd_1),
      fsm_output(9));
  butterFly1_15_f2_mux1h_63_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, ('0'
      & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_4), INNER_LOOP3_r_11_4_sva_6_0,
      ('1' & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_5), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_1_f1_butterFly1_1_f1_mux_2_rmff <= MUX_v_32_2_2((reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd
      & reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd_1), modulo_add_12_qr_lpi_3_dfm_1, fsm_output(9));
  butterFly1_1_f1_butterFly1_1_f1_mux_3_rmff <= MUX_v_32_2_2(modulo_add_12_qr_lpi_3_dfm_1,
      (reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd_1),
      fsm_output(9));
  butterFly1_15_f2_mux1h_62_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, ('0'
      & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_5), INNER_LOOP3_r_11_4_sva_6_0,
      ('1' & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_6), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_1_f2_butterFly1_1_f2_mux_2_rmff <= MUX_v_32_2_2((reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd
      & reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd_1), modulo_add_13_qr_lpi_3_dfm_1, fsm_output(9));
  butterFly1_1_f2_butterFly1_1_f2_mux_3_rmff <= MUX_v_32_2_2(modulo_add_13_qr_lpi_3_dfm_1,
      (reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd_1),
      fsm_output(9));
  butterFly1_15_f2_mux1h_61_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, ('0'
      & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_6), INNER_LOOP3_r_11_4_sva_6_0,
      ('1' & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_7), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_2_f1_butterFly1_2_f1_mux_2_rmff <= MUX_v_32_2_2((reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd
      & reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd_1), modulo_add_14_qr_lpi_3_dfm_1, fsm_output(9));
  butterFly1_2_f1_butterFly1_2_f1_mux_3_rmff <= MUX_v_32_2_2(modulo_add_14_qr_lpi_3_dfm_1,
      (reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd_1),
      fsm_output(9));
  butterFly1_15_f2_mux1h_60_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, ('0'
      & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_7), INNER_LOOP3_r_11_4_sva_6_0,
      ('1' & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_8), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_2_f2_butterFly1_2_f2_mux_2_rmff <= MUX_v_32_2_2((reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd
      & reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd_1), modulo_add_15_qr_lpi_3_dfm_1, fsm_output(9));
  butterFly1_2_f2_butterFly1_2_f2_mux_3_rmff <= MUX_v_32_2_2(modulo_add_15_qr_lpi_3_dfm_1,
      (reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd_1),
      fsm_output(9));
  butterFly1_15_f2_mux1h_59_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, ('0'
      & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_8), INNER_LOOP3_r_11_4_sva_6_0,
      ('1' & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_3_f1_butterFly1_3_f1_mux_2_rmff <= MUX_v_32_2_2((reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd
      & reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd_1), modulo_add_1_qr_lpi_3_dfm_1, fsm_output(9));
  butterFly1_3_f1_butterFly1_3_f1_mux_3_rmff <= MUX_v_32_2_2(modulo_add_1_qr_lpi_3_dfm_1,
      (reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd_1),
      fsm_output(9));
  butterFly1_15_f2_mux1h_58_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, ('0'
      & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1), INNER_LOOP3_r_11_4_sva_6_0,
      ('1' & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_2), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_3_f2_butterFly1_3_f2_mux_2_rmff <= MUX_v_32_2_2((reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd
      & reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd_1), modulo_add_23_qr_lpi_3_dfm_1, fsm_output(9));
  butterFly1_3_f2_butterFly1_3_f2_mux_3_rmff <= MUX_v_32_2_2(modulo_add_23_qr_lpi_3_dfm_1,
      (reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd_1),
      fsm_output(9));
  butterFly1_15_f2_mux1h_57_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, ('0'
      & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_2), INNER_LOOP3_r_11_4_sva_6_0,
      ('1' & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_3), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_4_f1_butterFly1_4_f1_mux_2_rmff <= MUX_v_32_2_2((reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd
      & reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd_1), modulo_add_24_qr_lpi_3_dfm_1, fsm_output(9));
  butterFly1_4_f1_butterFly1_4_f1_mux_3_rmff <= MUX_v_32_2_2(modulo_add_24_qr_lpi_3_dfm_1,
      (reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd_1),
      fsm_output(9));
  butterFly1_15_f2_mux1h_56_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, ('0'
      & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_3), INNER_LOOP3_r_11_4_sva_6_0,
      ('1' & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_4), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_4_f2_butterFly1_4_f2_mux_2_rmff <= MUX_v_32_2_2((reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd
      & reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd_1), modulo_add_25_qr_lpi_3_dfm_1, fsm_output(9));
  butterFly1_4_f2_butterFly1_4_f2_mux_3_rmff <= MUX_v_32_2_2(modulo_add_25_qr_lpi_3_dfm_1,
      (reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd_1),
      fsm_output(9));
  butterFly1_15_f2_mux1h_55_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, ('0'
      & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_4), INNER_LOOP3_r_11_4_sva_6_0,
      ('1' & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_5), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_5_f1_butterFly1_5_f1_mux_2_rmff <= MUX_v_32_2_2((reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd
      & reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd_1), modulo_add_26_qr_lpi_3_dfm_1, fsm_output(9));
  butterFly1_5_f1_butterFly1_5_f1_mux_3_rmff <= MUX_v_32_2_2(modulo_add_26_qr_lpi_3_dfm_1,
      (reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd_1),
      fsm_output(9));
  butterFly1_15_f2_mux1h_54_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, ('0'
      & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_5), INNER_LOOP3_r_11_4_sva_6_0,
      ('1' & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_6), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_5_f2_butterFly1_5_f2_mux_2_rmff <= MUX_v_32_2_2((reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd
      & reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd_1), modulo_add_27_qr_lpi_3_dfm_1, fsm_output(9));
  butterFly1_5_f2_butterFly1_5_f2_mux_3_rmff <= MUX_v_32_2_2(modulo_add_27_qr_lpi_3_dfm_1,
      (reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd_1),
      fsm_output(9));
  butterFly1_15_f2_mux1h_53_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, ('0'
      & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_6), INNER_LOOP3_r_11_4_sva_6_0,
      ('1' & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_7), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_6_f1_butterFly1_6_f1_mux_2_rmff <= MUX_v_32_2_2((reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd
      & reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd_1), modulo_add_28_qr_lpi_3_dfm_1, fsm_output(9));
  butterFly1_6_f1_butterFly1_6_f1_mux_3_rmff <= MUX_v_32_2_2(modulo_add_28_qr_lpi_3_dfm_1,
      (reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd_1),
      fsm_output(9));
  butterFly1_15_f2_mux1h_52_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, ('0'
      & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_7), INNER_LOOP3_r_11_4_sva_6_0,
      ('1' & INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_9), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_6_f2_butterFly1_6_f2_mux_2_rmff <= MUX_v_32_2_2((reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd
      & reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd_1), modulo_add_29_qr_lpi_3_dfm_1, fsm_output(9));
  butterFly1_6_f2_butterFly1_6_f2_mux_3_rmff <= MUX_v_32_2_2(modulo_add_29_qr_lpi_3_dfm_1,
      (reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd_1),
      fsm_output(9));
  butterFly1_15_f2_mux1h_51_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, ('0'
      & INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_9), INNER_LOOP3_r_11_4_sva_6_0,
      ('1' & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_1), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_7_f1_butterFly1_7_f1_mux_2_rmff <= MUX_v_32_2_2((reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd
      & reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd_1), modulo_add_30_qr_lpi_3_dfm_1, fsm_output(9));
  butterFly1_7_f1_butterFly1_7_f1_mux_3_rmff <= MUX_v_32_2_2(modulo_add_30_qr_lpi_3_dfm_1,
      (reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd_1),
      fsm_output(9));
  butterFly1_15_f2_mux1h_50_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, ('0'
      & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_1), INNER_LOOP3_r_11_4_sva_6_0,
      ('1' & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_2), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_7_f2_butterFly1_7_f2_mux_2_rmff <= MUX_v_32_2_2((reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd
      & reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd_1), modulo_add_31_qr_lpi_3_dfm_1, fsm_output(9));
  butterFly1_7_f2_butterFly1_7_f2_mux_3_rmff <= MUX_v_32_2_2(modulo_add_31_qr_lpi_3_dfm_1,
      (reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd & reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd_1),
      fsm_output(9));
  INNER_LOOP1_tw_and_nl <= INNER_LOOP2_r_11_4_sva_6_0 AND INNER_LOOP1_r_11_4_sva_6_0;
  INNER_LOOP2_tw_and_nl <= operator_33_true_1_lshift_psp_9_4_sva AND (INNER_LOOP2_r_11_4_sva_6_0(5
      DOWNTO 0));
  INNER_LOOP1_tw_h_mux1h_4_rmff <= MUX1HOT_v_7_4_2(INNER_LOOP1_tw_and_nl, ((INNER_LOOP2_r_11_4_sva_6_0(6))
      & INNER_LOOP2_tw_and_nl), INNER_LOOP3_r_11_4_sva_6_0, INNER_LOOP4_r_11_4_sva_6_0,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  butterFly1_butterFly1_or_1_rmff <= or_tmp_21 OR or_tmp_25;
  butterFly1_butterFly1_mux_3_rmff <= MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_129_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_161_itm_9_cse, or_tmp_25);
  butterFly1_1_butterFly1_1_mux_3_rmff <= MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_192_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_224_itm_9_cse, or_tmp_25);
  butterFly1_2_butterFly1_2_mux_3_rmff <= MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_255_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_287_itm_9_cse, or_tmp_25);
  butterFly1_3_butterFly1_3_mux_3_rmff <= MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_318_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_350_itm_9_cse, or_tmp_25);
  butterFly1_4_butterFly1_4_mux_3_rmff <= MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_381_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse, or_tmp_25);
  butterFly1_7_butterFly1_7_mux_3_rmff <= MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_570_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_602_itm_9_cse, or_tmp_25);
  butterFly1_8_butterFly1_8_mux_3_rmff <= MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_633_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_114_itm_9_cse, or_tmp_25);
  butterFly1_butterFly1_or_rmff <= or_tmp_203 OR or_tmp_207;
  butterFly1_butterFly1_mux_4_rmff <= MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_129_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_161_itm_9_cse, or_tmp_207);
  butterFly1_1_butterFly1_1_mux_4_rmff <= MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_192_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_224_itm_9_cse, or_tmp_207);
  butterFly1_2_butterFly1_2_mux_4_rmff <= MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_255_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_287_itm_9_cse, or_tmp_207);
  butterFly1_3_butterFly1_3_mux_4_rmff <= MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_318_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_350_itm_9_cse, or_tmp_207);
  butterFly1_4_butterFly1_4_mux_4_rmff <= MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_381_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse, or_tmp_207);
  butterFly1_7_butterFly1_7_mux_4_rmff <= MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_570_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_602_itm_9_cse, or_tmp_207);
  butterFly1_8_butterFly1_8_mux_4_rmff <= MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_633_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_114_itm_9_cse, or_tmp_207);
  butterFly1_f1_butterFly1_f1_butterFly1_f1_butterFly1_f1_nor_rmff <= NOT(nor_7_cse
      OR (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10) OR INNER_LOOP1_stage_0_9);
  butterFly1_f1_butterFly1_f1_butterFly1_f1_butterFly1_8_f1_nor_rmff <= NOT(nor_7_cse
      OR (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10) OR (NOT INNER_LOOP1_stage_0_9));
  yt_rsc_0_0_i_adra_d <= butterFly1_nor_7_rmff & butterFly1_butterFly1_or_1_rmff
      & butterFly1_butterFly1_mux_3_rmff & '0' & butterFly1_butterFly1_and_17_rmff
      & butterFly1_mux1h_15_rmff;
  butterFly1_butterFly1_mux_2_nl <= MUX_v_32_2_2(yt_rsc_0_0_i_da_d_mx0w0_63_32, yt_rsc_0_0_i_da_d_mx0w2_63_32,
      or_tmp_25);
  butterFly1_butterFly1_mux_6_nl <= MUX_v_32_2_2(modulo_add_31_qr_lpi_3_dfm_1, modulo_add_10_qr_lpi_3_dfm_1,
      butterFly1_or_5_cse);
  yt_rsc_0_0_i_da_d <= butterFly1_butterFly1_mux_2_nl & butterFly1_butterFly1_mux_6_nl;
  butterFly1_butterFly1_nor_2_nl <= NOT(yt_rsc_0_0_i_wea_d_mx0c2 OR yt_rsc_0_0_i_wea_d_mx0c0);
  butterFly1_mux_15_nl <= MUX_s_1_2_2((NOT or_dcpl_200), (NOT or_dcpl_199), or_tmp_25);
  butterFly1_butterFly1_nor_3_nl <= NOT((NOT(butterFly1_mux_15_nl OR yt_rsc_0_0_i_wea_d_mx0c2))
      OR yt_rsc_0_0_i_wea_d_mx0c0);
  yt_rsc_0_0_i_wea_d_pff <= STD_LOGIC_VECTOR'( butterFly1_butterFly1_nor_2_nl & butterFly1_butterFly1_nor_3_nl);
  yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_1_i_adra_d <= butterFly1_nor_7_rmff & butterFly1_butterFly1_or_1_rmff
      & butterFly1_1_butterFly1_1_mux_3_rmff & '0' & butterFly1_butterFly1_and_17_rmff
      & butterFly1_1_mux1h_11_rmff;
  butterFly1_1_butterFly1_1_mux_2_nl <= MUX_v_32_2_2(yt_rsc_0_1_i_da_d_mx0w0_63_32,
      yt_rsc_0_1_i_da_d_mx0w2_63_32, or_tmp_25);
  butterFly1_1_butterFly1_1_mux_6_nl <= MUX_v_32_2_2(modulo_add_1_qr_lpi_3_dfm_1,
      modulo_add_11_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  yt_rsc_0_1_i_da_d <= butterFly1_1_butterFly1_1_mux_2_nl & butterFly1_1_butterFly1_1_mux_6_nl;
  yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_2_i_adra_d <= butterFly1_nor_7_rmff & butterFly1_butterFly1_or_1_rmff
      & butterFly1_2_butterFly1_2_mux_3_rmff & '0' & butterFly1_butterFly1_and_17_rmff
      & butterFly1_2_mux1h_11_rmff;
  butterFly1_2_butterFly1_2_mux_2_nl <= MUX_v_32_2_2(yt_rsc_0_2_i_da_d_mx0w0_63_32,
      yt_rsc_0_2_i_da_d_mx0w2_63_32, or_tmp_25);
  butterFly1_2_butterFly1_2_mux_6_nl <= MUX_v_32_2_2(modulo_add_23_qr_lpi_3_dfm_1,
      modulo_add_12_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  yt_rsc_0_2_i_da_d <= butterFly1_2_butterFly1_2_mux_2_nl & butterFly1_2_butterFly1_2_mux_6_nl;
  yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_3_i_adra_d <= butterFly1_nor_7_rmff & butterFly1_butterFly1_or_1_rmff
      & butterFly1_3_butterFly1_3_mux_3_rmff & '0' & butterFly1_butterFly1_and_17_rmff
      & butterFly1_3_mux1h_11_rmff;
  butterFly1_3_butterFly1_3_mux_2_nl <= MUX_v_32_2_2(yt_rsc_0_3_i_da_d_mx0w0_63_32,
      yt_rsc_0_3_i_da_d_mx0w2_63_32, or_tmp_25);
  butterFly1_3_butterFly1_3_mux_6_nl <= MUX_v_32_2_2(modulo_add_24_qr_lpi_3_dfm_1,
      modulo_add_13_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  yt_rsc_0_3_i_da_d <= butterFly1_3_butterFly1_3_mux_2_nl & butterFly1_3_butterFly1_3_mux_6_nl;
  yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_4_i_adra_d <= butterFly1_nor_7_rmff & butterFly1_butterFly1_or_1_rmff
      & butterFly1_4_butterFly1_4_mux_3_rmff & '0' & butterFly1_butterFly1_and_17_rmff
      & butterFly1_4_mux1h_11_rmff;
  butterFly1_4_butterFly1_4_mux_2_nl <= MUX_v_32_2_2(yt_rsc_0_4_i_da_d_mx0w0_63_32,
      yt_rsc_0_4_i_da_d_mx0w2_63_32, or_tmp_25);
  butterFly1_4_butterFly1_4_mux_6_nl <= MUX_v_32_2_2(modulo_add_25_qr_lpi_3_dfm_1,
      modulo_add_14_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  yt_rsc_0_4_i_da_d <= butterFly1_4_butterFly1_4_mux_2_nl & butterFly1_4_butterFly1_4_mux_6_nl;
  yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  butterFly1_5_butterFly1_5_mux_3_nl <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_9, or_tmp_25);
  butterFly1_5_mux1h_11_nl <= MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_1_cse
      & (fsm_output(4)) & butterFly1_or_5_cse & (fsm_output(9))));
  yt_rsc_0_5_i_adra_d <= butterFly1_nor_7_rmff & butterFly1_butterFly1_or_1_rmff
      & butterFly1_5_butterFly1_5_mux_3_nl & '0' & butterFly1_butterFly1_and_17_rmff
      & butterFly1_5_mux1h_11_nl;
  butterFly1_5_butterFly1_5_mux_2_nl <= MUX_v_32_2_2(modulo_sub_5_qelse_mux_cse,
      yt_rsc_0_5_i_da_d_mx0w2_63_32, or_tmp_25);
  butterFly1_5_butterFly1_5_mux_6_nl <= MUX_v_32_2_2(modulo_add_26_qr_lpi_3_dfm_1,
      modulo_add_15_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  yt_rsc_0_5_i_da_d <= butterFly1_5_butterFly1_5_mux_2_nl & butterFly1_5_butterFly1_5_mux_6_nl;
  yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  butterFly1_6_butterFly1_6_mux_3_nl <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_9, or_tmp_25);
  butterFly1_6_mux1h_11_nl <= MUX1HOT_v_6_4_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_9,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_1_cse
      & (fsm_output(4)) & butterFly1_or_5_cse & (fsm_output(9))));
  yt_rsc_0_6_i_adra_d <= butterFly1_nor_7_rmff & butterFly1_butterFly1_or_1_rmff
      & butterFly1_6_butterFly1_6_mux_3_nl & '0' & butterFly1_butterFly1_and_17_rmff
      & butterFly1_6_mux1h_11_nl;
  butterFly1_6_butterFly1_6_mux_2_nl <= MUX_v_32_2_2(yt_rsc_0_6_i_da_d_mx0w0_63_32,
      yt_rsc_0_6_i_da_d_mx0w2_63_32, or_tmp_25);
  butterFly1_6_butterFly1_6_mux_6_nl <= MUX_v_32_2_2(modulo_add_27_qr_lpi_3_dfm_1,
      modulo_add_1_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  yt_rsc_0_6_i_da_d <= butterFly1_6_butterFly1_6_mux_2_nl & butterFly1_6_butterFly1_6_mux_6_nl;
  yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  butterFly1_7_mux1h_11_nl <= MUX1HOT_v_6_4_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_9,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_1_cse
      & (fsm_output(4)) & butterFly1_or_5_cse & (fsm_output(9))));
  yt_rsc_0_7_i_adra_d <= butterFly1_nor_7_rmff & butterFly1_butterFly1_or_1_rmff
      & butterFly1_7_butterFly1_7_mux_3_rmff & '0' & butterFly1_butterFly1_and_17_rmff
      & butterFly1_7_mux1h_11_nl;
  butterFly1_7_butterFly1_7_mux_2_nl <= MUX_v_32_2_2(yt_rsc_0_7_i_da_d_mx0w0_63_32,
      modulo_sub_5_qelse_mux_cse, or_tmp_25);
  butterFly1_7_butterFly1_7_mux_6_nl <= MUX_v_32_2_2(modulo_add_28_qr_lpi_3_dfm_1,
      modulo_add_23_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  yt_rsc_0_7_i_da_d <= butterFly1_7_butterFly1_7_mux_2_nl & butterFly1_7_butterFly1_7_mux_6_nl;
  yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_8_i_adra_d <= butterFly1_nor_7_rmff & butterFly1_butterFly1_or_1_rmff
      & butterFly1_8_butterFly1_8_mux_3_rmff & '0' & butterFly1_butterFly1_and_17_rmff
      & butterFly1_8_mux1h_11_rmff;
  butterFly1_8_butterFly1_8_mux_2_nl <= MUX_v_32_2_2(yt_rsc_0_8_i_da_d_mx0w0_63_32,
      yt_rsc_0_8_i_da_d_mx0w2_63_32, or_tmp_25);
  butterFly1_8_butterFly1_8_mux_6_nl <= MUX_v_32_2_2(modulo_add_29_qr_lpi_3_dfm_1,
      modulo_add_24_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  yt_rsc_0_8_i_da_d <= butterFly1_8_butterFly1_8_mux_2_nl & butterFly1_8_butterFly1_8_mux_6_nl;
  yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_9_i_adra_d <= butterFly1_nor_7_rmff & butterFly1_butterFly1_or_1_rmff
      & butterFly1_butterFly1_mux_3_rmff & '0' & butterFly1_butterFly1_and_17_rmff
      & butterFly1_mux1h_15_rmff;
  butterFly1_9_butterFly1_9_mux_2_nl <= MUX_v_32_2_2(yt_rsc_0_9_i_da_d_mx0w0_63_32,
      yt_rsc_0_9_i_da_d_mx0w2_63_32, or_tmp_25);
  butterFly1_9_butterFly1_9_mux_6_nl <= MUX_v_32_2_2(modulo_add_30_qr_lpi_3_dfm_1,
      modulo_add_25_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  yt_rsc_0_9_i_da_d <= butterFly1_9_butterFly1_9_mux_2_nl & butterFly1_9_butterFly1_9_mux_6_nl;
  yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_10_i_adra_d <= butterFly1_nor_7_rmff & butterFly1_butterFly1_or_1_rmff
      & butterFly1_1_butterFly1_1_mux_3_rmff & '0' & butterFly1_butterFly1_and_17_rmff
      & butterFly1_1_mux1h_11_rmff;
  butterFly1_10_butterFly1_10_mux_2_nl <= MUX_v_32_2_2(yt_rsc_0_10_i_da_d_mx0w0_63_32,
      yt_rsc_0_10_i_da_d_mx0w2_63_32, or_tmp_25);
  butterFly1_10_butterFly1_10_mux_6_nl <= MUX_v_32_2_2(modulo_add_10_qr_lpi_3_dfm_1,
      modulo_add_26_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  yt_rsc_0_10_i_da_d <= butterFly1_10_butterFly1_10_mux_2_nl & butterFly1_10_butterFly1_10_mux_6_nl;
  yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_11_i_adra_d <= butterFly1_nor_7_rmff & butterFly1_butterFly1_or_1_rmff
      & butterFly1_2_butterFly1_2_mux_3_rmff & '0' & butterFly1_butterFly1_and_17_rmff
      & butterFly1_2_mux1h_11_rmff;
  butterFly1_11_butterFly1_11_mux_2_nl <= MUX_v_32_2_2(yt_rsc_0_11_i_da_d_mx0w0_63_32,
      yt_rsc_0_11_i_da_d_mx0w2_63_32, or_tmp_25);
  butterFly1_11_butterFly1_11_mux_6_nl <= MUX_v_32_2_2(modulo_add_11_qr_lpi_3_dfm_1,
      modulo_add_27_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  yt_rsc_0_11_i_da_d <= butterFly1_11_butterFly1_11_mux_2_nl & butterFly1_11_butterFly1_11_mux_6_nl;
  yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_12_i_adra_d <= butterFly1_nor_7_rmff & butterFly1_butterFly1_or_1_rmff
      & butterFly1_3_butterFly1_3_mux_3_rmff & '0' & butterFly1_butterFly1_and_17_rmff
      & butterFly1_3_mux1h_11_rmff;
  butterFly1_12_butterFly1_12_mux_2_nl <= MUX_v_32_2_2(yt_rsc_0_12_i_da_d_mx0w0_63_32,
      yt_rsc_0_12_i_da_d_mx0w2_63_32, or_tmp_25);
  butterFly1_12_butterFly1_12_mux_6_nl <= MUX_v_32_2_2(modulo_add_12_qr_lpi_3_dfm_1,
      modulo_add_28_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  yt_rsc_0_12_i_da_d <= butterFly1_12_butterFly1_12_mux_2_nl & butterFly1_12_butterFly1_12_mux_6_nl;
  yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_13_i_adra_d <= butterFly1_nor_7_rmff & butterFly1_butterFly1_or_1_rmff
      & butterFly1_4_butterFly1_4_mux_3_rmff & '0' & butterFly1_butterFly1_and_17_rmff
      & butterFly1_4_mux1h_11_rmff;
  butterFly1_13_butterFly1_13_mux_2_nl <= MUX_v_32_2_2(yt_rsc_0_13_i_da_d_mx0w0_63_32,
      yt_rsc_0_13_i_da_d_mx0w2_63_32, or_tmp_25);
  butterFly1_13_butterFly1_13_mux_6_nl <= MUX_v_32_2_2(modulo_add_13_qr_lpi_3_dfm_1,
      modulo_add_29_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  yt_rsc_0_13_i_da_d <= butterFly1_13_butterFly1_13_mux_2_nl & butterFly1_13_butterFly1_13_mux_6_nl;
  yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  butterFly1_14_mux1h_11_nl <= MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_1_cse
      & (fsm_output(4)) & butterFly1_or_5_cse & (fsm_output(9))));
  yt_rsc_0_14_i_adra_d <= butterFly1_nor_7_rmff & butterFly1_butterFly1_or_1_rmff
      & butterFly1_7_butterFly1_7_mux_3_rmff & '0' & butterFly1_butterFly1_and_17_rmff
      & butterFly1_14_mux1h_11_nl;
  butterFly1_14_butterFly1_14_mux_2_nl <= MUX_v_32_2_2(yt_rsc_0_14_i_da_d_mx0w0_63_32,
      yt_rsc_0_14_i_da_d_mx0w2_63_32, or_tmp_25);
  butterFly1_14_butterFly1_14_mux_6_nl <= MUX_v_32_2_2(modulo_add_14_qr_lpi_3_dfm_1,
      modulo_add_30_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  yt_rsc_0_14_i_da_d <= butterFly1_14_butterFly1_14_mux_2_nl & butterFly1_14_butterFly1_14_mux_6_nl;
  yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_15_i_adra_d <= butterFly1_nor_7_rmff & butterFly1_butterFly1_or_1_rmff
      & butterFly1_8_butterFly1_8_mux_3_rmff & '0' & butterFly1_butterFly1_and_17_rmff
      & butterFly1_8_mux1h_11_rmff;
  butterFly1_15_butterFly1_15_mux_2_nl <= MUX_v_32_2_2(yt_rsc_0_15_i_da_d_mx0w0_63_32,
      yt_rsc_0_15_i_da_d_mx0w2_63_32, or_tmp_25);
  butterFly1_15_butterFly1_15_mux_6_nl <= MUX_v_32_2_2(modulo_add_15_qr_lpi_3_dfm_1,
      modulo_add_31_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  yt_rsc_0_15_i_da_d <= butterFly1_15_butterFly1_15_mux_2_nl & butterFly1_15_butterFly1_15_mux_6_nl;
  yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_16_i_adra_d <= butterFly1_nor_4_rmff & butterFly1_butterFly1_or_rmff &
      butterFly1_butterFly1_mux_4_rmff & '0' & butterFly1_butterFly1_and_15_rmff
      & butterFly1_mux1h_13_rmff;
  butterFly1_butterFly1_mux_nl <= MUX_v_32_2_2(yt_rsc_0_0_i_da_d_mx0w0_63_32, yt_rsc_0_0_i_da_d_mx0w2_63_32,
      or_tmp_207);
  butterFly1_butterFly1_mux_5_nl <= MUX_v_32_2_2(modulo_add_31_qr_lpi_3_dfm_1, modulo_add_10_qr_lpi_3_dfm_1,
      butterFly1_or_4_cse);
  yt_rsc_0_16_i_da_d <= butterFly1_butterFly1_mux_nl & butterFly1_butterFly1_mux_5_nl;
  butterFly1_butterFly1_nor_nl <= NOT(yt_rsc_0_16_i_wea_d_mx0c2 OR yt_rsc_0_16_i_wea_d_mx0c0);
  butterFly1_mux_nl <= MUX_s_1_2_2((NOT or_dcpl_208), (NOT or_dcpl_207), or_tmp_207);
  butterFly1_butterFly1_nor_1_nl <= NOT((NOT(butterFly1_mux_nl OR yt_rsc_0_16_i_wea_d_mx0c2))
      OR yt_rsc_0_16_i_wea_d_mx0c0);
  yt_rsc_0_16_i_wea_d_pff <= STD_LOGIC_VECTOR'( butterFly1_butterFly1_nor_nl & butterFly1_butterFly1_nor_1_nl);
  yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_17_i_adra_d <= butterFly1_nor_4_rmff & butterFly1_butterFly1_or_rmff &
      butterFly1_1_butterFly1_1_mux_4_rmff & '0' & butterFly1_butterFly1_and_15_rmff
      & butterFly1_1_mux1h_9_rmff;
  butterFly1_1_butterFly1_1_mux_nl <= MUX_v_32_2_2(yt_rsc_0_1_i_da_d_mx0w0_63_32,
      yt_rsc_0_1_i_da_d_mx0w2_63_32, or_tmp_207);
  butterFly1_1_butterFly1_1_mux_5_nl <= MUX_v_32_2_2(modulo_add_1_qr_lpi_3_dfm_1,
      modulo_add_11_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  yt_rsc_0_17_i_da_d <= butterFly1_1_butterFly1_1_mux_nl & butterFly1_1_butterFly1_1_mux_5_nl;
  yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_18_i_adra_d <= butterFly1_nor_4_rmff & butterFly1_butterFly1_or_rmff &
      butterFly1_2_butterFly1_2_mux_4_rmff & '0' & butterFly1_butterFly1_and_15_rmff
      & butterFly1_2_mux1h_9_rmff;
  butterFly1_2_butterFly1_2_mux_nl <= MUX_v_32_2_2(yt_rsc_0_2_i_da_d_mx0w0_63_32,
      yt_rsc_0_2_i_da_d_mx0w2_63_32, or_tmp_207);
  butterFly1_2_butterFly1_2_mux_5_nl <= MUX_v_32_2_2(modulo_add_23_qr_lpi_3_dfm_1,
      modulo_add_12_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  yt_rsc_0_18_i_da_d <= butterFly1_2_butterFly1_2_mux_nl & butterFly1_2_butterFly1_2_mux_5_nl;
  yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_19_i_adra_d <= butterFly1_nor_4_rmff & butterFly1_butterFly1_or_rmff &
      butterFly1_3_butterFly1_3_mux_4_rmff & '0' & butterFly1_butterFly1_and_15_rmff
      & butterFly1_3_mux1h_9_rmff;
  butterFly1_3_butterFly1_3_mux_nl <= MUX_v_32_2_2(yt_rsc_0_3_i_da_d_mx0w0_63_32,
      yt_rsc_0_3_i_da_d_mx0w2_63_32, or_tmp_207);
  butterFly1_3_butterFly1_3_mux_5_nl <= MUX_v_32_2_2(modulo_add_24_qr_lpi_3_dfm_1,
      modulo_add_13_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  yt_rsc_0_19_i_da_d <= butterFly1_3_butterFly1_3_mux_nl & butterFly1_3_butterFly1_3_mux_5_nl;
  yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_20_i_adra_d <= butterFly1_nor_4_rmff & butterFly1_butterFly1_or_rmff &
      butterFly1_4_butterFly1_4_mux_4_rmff & '0' & butterFly1_butterFly1_and_15_rmff
      & butterFly1_4_mux1h_9_rmff;
  butterFly1_4_butterFly1_4_mux_nl <= MUX_v_32_2_2(yt_rsc_0_4_i_da_d_mx0w0_63_32,
      yt_rsc_0_4_i_da_d_mx0w2_63_32, or_tmp_207);
  butterFly1_4_butterFly1_4_mux_5_nl <= MUX_v_32_2_2(modulo_add_25_qr_lpi_3_dfm_1,
      modulo_add_14_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  yt_rsc_0_20_i_da_d <= butterFly1_4_butterFly1_4_mux_nl & butterFly1_4_butterFly1_4_mux_5_nl;
  yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  butterFly1_5_butterFly1_5_mux_4_nl <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_9, or_tmp_207);
  butterFly1_5_mux1h_9_nl <= MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_cse
      & (fsm_output(4)) & butterFly1_or_4_cse & (fsm_output(9))));
  yt_rsc_0_21_i_adra_d <= butterFly1_nor_4_rmff & butterFly1_butterFly1_or_rmff &
      butterFly1_5_butterFly1_5_mux_4_nl & '0' & butterFly1_butterFly1_and_15_rmff
      & butterFly1_5_mux1h_9_nl;
  butterFly1_5_butterFly1_5_mux_nl <= MUX_v_32_2_2(modulo_sub_5_qelse_mux_cse, yt_rsc_0_5_i_da_d_mx0w2_63_32,
      or_tmp_207);
  butterFly1_5_butterFly1_5_mux_5_nl <= MUX_v_32_2_2(modulo_add_26_qr_lpi_3_dfm_1,
      modulo_add_15_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  yt_rsc_0_21_i_da_d <= butterFly1_5_butterFly1_5_mux_nl & butterFly1_5_butterFly1_5_mux_5_nl;
  yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  butterFly1_6_butterFly1_6_mux_4_nl <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_9, or_tmp_207);
  butterFly1_6_mux1h_9_nl <= MUX1HOT_v_6_4_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_9,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_cse
      & (fsm_output(4)) & butterFly1_or_4_cse & (fsm_output(9))));
  yt_rsc_0_22_i_adra_d <= butterFly1_nor_4_rmff & butterFly1_butterFly1_or_rmff &
      butterFly1_6_butterFly1_6_mux_4_nl & '0' & butterFly1_butterFly1_and_15_rmff
      & butterFly1_6_mux1h_9_nl;
  butterFly1_6_butterFly1_6_mux_nl <= MUX_v_32_2_2(yt_rsc_0_6_i_da_d_mx0w0_63_32,
      yt_rsc_0_6_i_da_d_mx0w2_63_32, or_tmp_207);
  butterFly1_6_butterFly1_6_mux_5_nl <= MUX_v_32_2_2(modulo_add_27_qr_lpi_3_dfm_1,
      modulo_add_1_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  yt_rsc_0_22_i_da_d <= butterFly1_6_butterFly1_6_mux_nl & butterFly1_6_butterFly1_6_mux_5_nl;
  yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  butterFly1_7_mux1h_9_nl <= MUX1HOT_v_6_4_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_9,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_cse
      & (fsm_output(4)) & butterFly1_or_4_cse & (fsm_output(9))));
  yt_rsc_0_23_i_adra_d <= butterFly1_nor_4_rmff & butterFly1_butterFly1_or_rmff &
      butterFly1_7_butterFly1_7_mux_4_rmff & '0' & butterFly1_butterFly1_and_15_rmff
      & butterFly1_7_mux1h_9_nl;
  butterFly1_7_butterFly1_7_mux_nl <= MUX_v_32_2_2(yt_rsc_0_7_i_da_d_mx0w0_63_32,
      modulo_sub_5_qelse_mux_cse, or_tmp_207);
  butterFly1_7_butterFly1_7_mux_5_nl <= MUX_v_32_2_2(modulo_add_28_qr_lpi_3_dfm_1,
      modulo_add_23_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  yt_rsc_0_23_i_da_d <= butterFly1_7_butterFly1_7_mux_nl & butterFly1_7_butterFly1_7_mux_5_nl;
  yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_24_i_adra_d <= butterFly1_nor_4_rmff & butterFly1_butterFly1_or_rmff &
      butterFly1_8_butterFly1_8_mux_4_rmff & '0' & butterFly1_butterFly1_and_15_rmff
      & butterFly1_8_mux1h_9_rmff;
  butterFly1_8_butterFly1_8_mux_nl <= MUX_v_32_2_2(yt_rsc_0_8_i_da_d_mx0w0_63_32,
      yt_rsc_0_8_i_da_d_mx0w2_63_32, or_tmp_207);
  butterFly1_8_butterFly1_8_mux_5_nl <= MUX_v_32_2_2(modulo_add_29_qr_lpi_3_dfm_1,
      modulo_add_24_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  yt_rsc_0_24_i_da_d <= butterFly1_8_butterFly1_8_mux_nl & butterFly1_8_butterFly1_8_mux_5_nl;
  yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_25_i_adra_d <= butterFly1_nor_4_rmff & butterFly1_butterFly1_or_rmff &
      butterFly1_butterFly1_mux_4_rmff & '0' & butterFly1_butterFly1_and_15_rmff
      & butterFly1_mux1h_13_rmff;
  butterFly1_9_butterFly1_9_mux_nl <= MUX_v_32_2_2(yt_rsc_0_9_i_da_d_mx0w0_63_32,
      yt_rsc_0_9_i_da_d_mx0w2_63_32, or_tmp_207);
  butterFly1_9_butterFly1_9_mux_5_nl <= MUX_v_32_2_2(modulo_add_30_qr_lpi_3_dfm_1,
      modulo_add_25_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  yt_rsc_0_25_i_da_d <= butterFly1_9_butterFly1_9_mux_nl & butterFly1_9_butterFly1_9_mux_5_nl;
  yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_26_i_adra_d <= butterFly1_nor_4_rmff & butterFly1_butterFly1_or_rmff &
      butterFly1_1_butterFly1_1_mux_4_rmff & '0' & butterFly1_butterFly1_and_15_rmff
      & butterFly1_1_mux1h_9_rmff;
  butterFly1_10_butterFly1_10_mux_nl <= MUX_v_32_2_2(yt_rsc_0_10_i_da_d_mx0w0_63_32,
      yt_rsc_0_10_i_da_d_mx0w2_63_32, or_tmp_207);
  butterFly1_10_butterFly1_10_mux_5_nl <= MUX_v_32_2_2(modulo_add_10_qr_lpi_3_dfm_1,
      modulo_add_26_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  yt_rsc_0_26_i_da_d <= butterFly1_10_butterFly1_10_mux_nl & butterFly1_10_butterFly1_10_mux_5_nl;
  yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_27_i_adra_d <= butterFly1_nor_4_rmff & butterFly1_butterFly1_or_rmff &
      butterFly1_2_butterFly1_2_mux_4_rmff & '0' & butterFly1_butterFly1_and_15_rmff
      & butterFly1_2_mux1h_9_rmff;
  butterFly1_11_butterFly1_11_mux_nl <= MUX_v_32_2_2(yt_rsc_0_11_i_da_d_mx0w0_63_32,
      yt_rsc_0_11_i_da_d_mx0w2_63_32, or_tmp_207);
  butterFly1_11_butterFly1_11_mux_5_nl <= MUX_v_32_2_2(modulo_add_11_qr_lpi_3_dfm_1,
      modulo_add_27_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  yt_rsc_0_27_i_da_d <= butterFly1_11_butterFly1_11_mux_nl & butterFly1_11_butterFly1_11_mux_5_nl;
  yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_28_i_adra_d <= butterFly1_nor_4_rmff & butterFly1_butterFly1_or_rmff &
      butterFly1_3_butterFly1_3_mux_4_rmff & '0' & butterFly1_butterFly1_and_15_rmff
      & butterFly1_3_mux1h_9_rmff;
  butterFly1_12_butterFly1_12_mux_nl <= MUX_v_32_2_2(yt_rsc_0_12_i_da_d_mx0w0_63_32,
      yt_rsc_0_12_i_da_d_mx0w2_63_32, or_tmp_207);
  butterFly1_12_butterFly1_12_mux_5_nl <= MUX_v_32_2_2(modulo_add_12_qr_lpi_3_dfm_1,
      modulo_add_28_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  yt_rsc_0_28_i_da_d <= butterFly1_12_butterFly1_12_mux_nl & butterFly1_12_butterFly1_12_mux_5_nl;
  yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_29_i_adra_d <= butterFly1_nor_4_rmff & butterFly1_butterFly1_or_rmff &
      butterFly1_4_butterFly1_4_mux_4_rmff & '0' & butterFly1_butterFly1_and_15_rmff
      & butterFly1_4_mux1h_9_rmff;
  butterFly1_13_butterFly1_13_mux_nl <= MUX_v_32_2_2(yt_rsc_0_13_i_da_d_mx0w0_63_32,
      yt_rsc_0_13_i_da_d_mx0w2_63_32, or_tmp_207);
  butterFly1_13_butterFly1_13_mux_5_nl <= MUX_v_32_2_2(modulo_add_13_qr_lpi_3_dfm_1,
      modulo_add_29_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  yt_rsc_0_29_i_da_d <= butterFly1_13_butterFly1_13_mux_nl & butterFly1_13_butterFly1_13_mux_5_nl;
  yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  butterFly1_14_mux1h_9_nl <= MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0(5 DOWNTO 0)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0(5 DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_or_cse
      & (fsm_output(4)) & butterFly1_or_4_cse & (fsm_output(9))));
  yt_rsc_0_30_i_adra_d <= butterFly1_nor_4_rmff & butterFly1_butterFly1_or_rmff &
      butterFly1_7_butterFly1_7_mux_4_rmff & '0' & butterFly1_butterFly1_and_15_rmff
      & butterFly1_14_mux1h_9_nl;
  butterFly1_14_butterFly1_14_mux_nl <= MUX_v_32_2_2(yt_rsc_0_14_i_da_d_mx0w0_63_32,
      yt_rsc_0_14_i_da_d_mx0w2_63_32, or_tmp_207);
  butterFly1_14_butterFly1_14_mux_5_nl <= MUX_v_32_2_2(modulo_add_14_qr_lpi_3_dfm_1,
      modulo_add_30_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  yt_rsc_0_30_i_da_d <= butterFly1_14_butterFly1_14_mux_nl & butterFly1_14_butterFly1_14_mux_5_nl;
  yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  yt_rsc_0_31_i_adra_d <= butterFly1_nor_4_rmff & butterFly1_butterFly1_or_rmff &
      butterFly1_8_butterFly1_8_mux_4_rmff & '0' & butterFly1_butterFly1_and_15_rmff
      & butterFly1_8_mux1h_9_rmff;
  butterFly1_15_butterFly1_15_mux_nl <= MUX_v_32_2_2(yt_rsc_0_15_i_da_d_mx0w0_63_32,
      yt_rsc_0_15_i_da_d_mx0w2_63_32, or_tmp_207);
  butterFly1_15_butterFly1_15_mux_5_nl <= MUX_v_32_2_2(modulo_add_15_qr_lpi_3_dfm_1,
      modulo_add_31_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  yt_rsc_0_31_i_da_d <= butterFly1_15_butterFly1_15_mux_nl & butterFly1_15_butterFly1_15_mux_5_nl;
  yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_202_rmff);
  xt_rsc_0_0_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_3
      & '0' & butterFly1_15_f2_mux1h_65_rmff;
  xt_rsc_0_0_i_da_d <= butterFly1_f1_butterFly1_f1_mux_2_rmff & butterFly1_f1_butterFly1_f1_mux_3_rmff;
  xt_rsc_0_0_i_wea_d_pff <= STD_LOGIC_VECTOR'( butterFly1_f1_butterFly1_f1_butterFly1_f1_butterFly1_f1_nor_rmff
      & butterFly1_f1_butterFly1_f1_butterFly1_f1_butterFly1_f1_nor_rmff);
  xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_1_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_4
      & '0' & butterFly1_15_f2_mux1h_64_rmff;
  xt_rsc_0_1_i_da_d <= butterFly1_f2_butterFly1_f2_mux_2_rmff & butterFly1_f2_butterFly1_f2_mux_3_rmff;
  xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_2_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_5
      & '0' & butterFly1_15_f2_mux1h_63_rmff;
  xt_rsc_0_2_i_da_d <= butterFly1_1_f1_butterFly1_1_f1_mux_2_rmff & butterFly1_1_f1_butterFly1_1_f1_mux_3_rmff;
  xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_3_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_6
      & '0' & butterFly1_15_f2_mux1h_62_rmff;
  xt_rsc_0_3_i_da_d <= butterFly1_1_f2_butterFly1_1_f2_mux_2_rmff & butterFly1_1_f2_butterFly1_1_f2_mux_3_rmff;
  xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_4_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_7
      & '0' & butterFly1_15_f2_mux1h_61_rmff;
  xt_rsc_0_4_i_da_d <= butterFly1_2_f1_butterFly1_2_f1_mux_2_rmff & butterFly1_2_f1_butterFly1_2_f1_mux_3_rmff;
  xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_5_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_8
      & '0' & butterFly1_15_f2_mux1h_60_rmff;
  xt_rsc_0_5_i_da_d <= butterFly1_2_f2_butterFly1_2_f2_mux_2_rmff & butterFly1_2_f2_butterFly1_2_f2_mux_3_rmff;
  xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_6_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_9
      & '0' & butterFly1_15_f2_mux1h_59_rmff;
  xt_rsc_0_6_i_da_d <= butterFly1_3_f1_butterFly1_3_f1_mux_2_rmff & butterFly1_3_f1_butterFly1_3_f1_mux_3_rmff;
  xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_7_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_1
      & '0' & butterFly1_15_f2_mux1h_58_rmff;
  xt_rsc_0_7_i_da_d <= butterFly1_3_f2_butterFly1_3_f2_mux_2_rmff & butterFly1_3_f2_butterFly1_3_f2_mux_3_rmff;
  xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_8_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_2
      & '0' & butterFly1_15_f2_mux1h_57_rmff;
  xt_rsc_0_8_i_da_d <= butterFly1_4_f1_butterFly1_4_f1_mux_2_rmff & butterFly1_4_f1_butterFly1_4_f1_mux_3_rmff;
  xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_9_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_3
      & '0' & butterFly1_15_f2_mux1h_56_rmff;
  xt_rsc_0_9_i_da_d <= butterFly1_4_f2_butterFly1_4_f2_mux_2_rmff & butterFly1_4_f2_butterFly1_4_f2_mux_3_rmff;
  xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_10_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_4
      & '0' & butterFly1_15_f2_mux1h_55_rmff;
  xt_rsc_0_10_i_da_d <= butterFly1_5_f1_butterFly1_5_f1_mux_2_rmff & butterFly1_5_f1_butterFly1_5_f1_mux_3_rmff;
  xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_11_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_5
      & '0' & butterFly1_15_f2_mux1h_54_rmff;
  xt_rsc_0_11_i_da_d <= butterFly1_5_f2_butterFly1_5_f2_mux_2_rmff & butterFly1_5_f2_butterFly1_5_f2_mux_3_rmff;
  xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_12_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_6
      & '0' & butterFly1_15_f2_mux1h_53_rmff;
  xt_rsc_0_12_i_da_d <= butterFly1_6_f1_butterFly1_6_f1_mux_2_rmff & butterFly1_6_f1_butterFly1_6_f1_mux_3_rmff;
  xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_13_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_9
      & '0' & butterFly1_15_f2_mux1h_52_rmff;
  xt_rsc_0_13_i_da_d <= butterFly1_6_f2_butterFly1_6_f2_mux_2_rmff & butterFly1_6_f2_butterFly1_6_f2_mux_3_rmff;
  xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_14_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1
      & '0' & butterFly1_15_f2_mux1h_51_rmff;
  xt_rsc_0_14_i_da_d <= butterFly1_7_f1_butterFly1_7_f1_mux_2_rmff & butterFly1_7_f1_butterFly1_7_f1_mux_3_rmff;
  xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_15_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_2
      & '0' & butterFly1_15_f2_mux1h_50_rmff;
  xt_rsc_0_15_i_da_d <= butterFly1_7_f2_butterFly1_7_f2_mux_2_rmff & butterFly1_7_f2_butterFly1_7_f2_mux_3_rmff;
  xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_16_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_3
      & '0' & butterFly1_15_f2_mux1h_65_rmff;
  xt_rsc_0_16_i_da_d <= butterFly1_f1_butterFly1_f1_mux_2_rmff & butterFly1_f1_butterFly1_f1_mux_3_rmff;
  xt_rsc_0_16_i_wea_d_pff <= STD_LOGIC_VECTOR'( butterFly1_f1_butterFly1_f1_butterFly1_f1_butterFly1_8_f1_nor_rmff
      & butterFly1_f1_butterFly1_f1_butterFly1_f1_butterFly1_8_f1_nor_rmff);
  xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_17_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_4
      & '0' & butterFly1_15_f2_mux1h_64_rmff;
  xt_rsc_0_17_i_da_d <= butterFly1_f2_butterFly1_f2_mux_2_rmff & butterFly1_f2_butterFly1_f2_mux_3_rmff;
  xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_18_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_5
      & '0' & butterFly1_15_f2_mux1h_63_rmff;
  xt_rsc_0_18_i_da_d <= butterFly1_1_f1_butterFly1_1_f1_mux_2_rmff & butterFly1_1_f1_butterFly1_1_f1_mux_3_rmff;
  xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_19_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_6
      & '0' & butterFly1_15_f2_mux1h_62_rmff;
  xt_rsc_0_19_i_da_d <= butterFly1_1_f2_butterFly1_1_f2_mux_2_rmff & butterFly1_1_f2_butterFly1_1_f2_mux_3_rmff;
  xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_20_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_7
      & '0' & butterFly1_15_f2_mux1h_61_rmff;
  xt_rsc_0_20_i_da_d <= butterFly1_2_f1_butterFly1_2_f1_mux_2_rmff & butterFly1_2_f1_butterFly1_2_f1_mux_3_rmff;
  xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_21_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_8
      & '0' & butterFly1_15_f2_mux1h_60_rmff;
  xt_rsc_0_21_i_da_d <= butterFly1_2_f2_butterFly1_2_f2_mux_2_rmff & butterFly1_2_f2_butterFly1_2_f2_mux_3_rmff;
  xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_22_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_9
      & '0' & butterFly1_15_f2_mux1h_59_rmff;
  xt_rsc_0_22_i_da_d <= butterFly1_3_f1_butterFly1_3_f1_mux_2_rmff & butterFly1_3_f1_butterFly1_3_f1_mux_3_rmff;
  xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_23_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_1
      & '0' & butterFly1_15_f2_mux1h_58_rmff;
  xt_rsc_0_23_i_da_d <= butterFly1_3_f2_butterFly1_3_f2_mux_2_rmff & butterFly1_3_f2_butterFly1_3_f2_mux_3_rmff;
  xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_24_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_2
      & '0' & butterFly1_15_f2_mux1h_57_rmff;
  xt_rsc_0_24_i_da_d <= butterFly1_4_f1_butterFly1_4_f1_mux_2_rmff & butterFly1_4_f1_butterFly1_4_f1_mux_3_rmff;
  xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_25_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_3
      & '0' & butterFly1_15_f2_mux1h_56_rmff;
  xt_rsc_0_25_i_da_d <= butterFly1_4_f2_butterFly1_4_f2_mux_2_rmff & butterFly1_4_f2_butterFly1_4_f2_mux_3_rmff;
  xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_26_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_4
      & '0' & butterFly1_15_f2_mux1h_55_rmff;
  xt_rsc_0_26_i_da_d <= butterFly1_5_f1_butterFly1_5_f1_mux_2_rmff & butterFly1_5_f1_butterFly1_5_f1_mux_3_rmff;
  xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_27_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_5
      & '0' & butterFly1_15_f2_mux1h_54_rmff;
  xt_rsc_0_27_i_da_d <= butterFly1_5_f2_butterFly1_5_f2_mux_2_rmff & butterFly1_5_f2_butterFly1_5_f2_mux_3_rmff;
  xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_28_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_6
      & '0' & butterFly1_15_f2_mux1h_53_rmff;
  xt_rsc_0_28_i_da_d <= butterFly1_6_f1_butterFly1_6_f1_mux_2_rmff & butterFly1_6_f1_butterFly1_6_f1_mux_3_rmff;
  xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_29_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_9
      & '0' & butterFly1_15_f2_mux1h_52_rmff;
  xt_rsc_0_29_i_da_d <= butterFly1_6_f2_butterFly1_6_f2_mux_2_rmff & butterFly1_6_f2_butterFly1_6_f2_mux_3_rmff;
  xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_30_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1
      & '0' & butterFly1_15_f2_mux1h_51_rmff;
  xt_rsc_0_30_i_da_d <= butterFly1_7_f1_butterFly1_7_f1_mux_2_rmff & butterFly1_7_f1_butterFly1_7_f1_mux_3_rmff;
  xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  xt_rsc_0_31_i_adra_d <= nor_7_cse & (NOT (fsm_output(9))) & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_2
      & '0' & butterFly1_15_f2_mux1h_50_rmff;
  xt_rsc_0_31_i_da_d <= butterFly1_7_f2_butterFly1_7_f2_mux_2_rmff & butterFly1_7_f2_butterFly1_7_f2_mux_3_rmff;
  xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' & and_921_rmff);
  twiddle_rsc_0_0_i_adra_d <= '0' & INNER_LOOP1_tw_h_mux1h_4_rmff;
  twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      and_1435_rmff);
  twiddle_rsc_0_1_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_896_rmff);
  twiddle_rsc_0_2_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_900_rmff);
  twiddle_rsc_0_3_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_904_rmff);
  twiddle_rsc_0_4_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_908_rmff);
  twiddle_rsc_0_5_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_912_rmff);
  twiddle_rsc_0_6_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_916_rmff);
  twiddle_rsc_0_7_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_920_rmff);
  twiddle_rsc_0_8_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      and_1506_rmff);
  twiddle_rsc_0_9_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_896_rmff);
  twiddle_rsc_0_10_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_900_rmff);
  twiddle_rsc_0_11_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_904_rmff);
  twiddle_rsc_0_12_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_908_rmff);
  twiddle_rsc_0_13_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_912_rmff);
  twiddle_rsc_0_14_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_916_rmff);
  twiddle_rsc_0_15_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0' &
      or_920_rmff);
  twiddle_h_rsc_0_0_i_adra_d <= '0' & INNER_LOOP1_tw_h_mux1h_4_rmff;
  twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & and_1435_rmff);
  twiddle_h_rsc_0_1_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_896_rmff);
  twiddle_h_rsc_0_2_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_900_rmff);
  twiddle_h_rsc_0_3_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_904_rmff);
  twiddle_h_rsc_0_4_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_908_rmff);
  twiddle_h_rsc_0_5_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_912_rmff);
  twiddle_h_rsc_0_6_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_916_rmff);
  twiddle_h_rsc_0_7_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_920_rmff);
  twiddle_h_rsc_0_8_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & and_1506_rmff);
  twiddle_h_rsc_0_9_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_896_rmff);
  twiddle_h_rsc_0_10_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_900_rmff);
  twiddle_h_rsc_0_11_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_904_rmff);
  twiddle_h_rsc_0_12_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_908_rmff);
  twiddle_h_rsc_0_13_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_912_rmff);
  twiddle_h_rsc_0_14_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_916_rmff);
  twiddle_h_rsc_0_15_i_adra_d <= '0' & butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( '0'
      & or_920_rmff);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( ((fsm_output(10)) OR (fsm_output(0))) = '1' ) THEN
        p_sva <= p_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        c_1_sva <= '0';
      ELSIF ( ((fsm_output(5)) OR (fsm_output(0)) OR (fsm_output(9))) = '1' ) THEN
        c_1_sva <= c_mux_nl AND (NOT (fsm_output(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_yt_rsc_0_0_cgo_cse <= '0';
        reg_yt_rsc_0_16_cgo_cse <= '0';
        reg_xt_rsc_triosy_0_31_obj_ld_cse <= '0';
        reg_ensig_cgo_cse <= '0';
        reg_ensig_cgo_17_cse <= '0';
        butterFly2_11_tw_h_slc_operator_33_true_2_lshift_psp_2_0_1_0_itm <= STD_LOGIC_VECTOR'(
            "00");
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10 <= '0';
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9 <= '0';
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8 <= '0';
        INNER_LOOP1_stage_0 <= '0';
        INNER_LOOP1_r_11_4_sva_6_0 <= STD_LOGIC_VECTOR'( "0000000");
        INNER_LOOP1_stage_0_2 <= '0';
        INNER_LOOP1_stage_0_3 <= '0';
        INNER_LOOP1_stage_0_4 <= '0';
        INNER_LOOP1_stage_0_5 <= '0';
        INNER_LOOP1_stage_0_6 <= '0';
        INNER_LOOP1_stage_0_7 <= '0';
        INNER_LOOP1_stage_0_8 <= '0';
        INNER_LOOP1_stage_0_9 <= '0';
        INNER_LOOP1_stage_0_10 <= '0';
        INNER_LOOP1_stage_0_11 <= '0';
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 <= '0';
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 <= '0';
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 <= '0';
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 <= '0';
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 <= '0';
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 <= '0';
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 <= '0';
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm <= '0';
        INNER_LOOP3_r_11_4_sva_6_0 <= STD_LOGIC_VECTOR'( "0000000");
        INNER_LOOP4_r_11_4_sva_6_0 <= STD_LOGIC_VECTOR'( "0000000");
      ELSE
        reg_yt_rsc_0_0_cgo_cse <= or_261_rmff;
        reg_yt_rsc_0_16_cgo_cse <= or_443_rmff;
        reg_xt_rsc_triosy_0_31_obj_ld_cse <= and_dcpl_51 AND (fsm_output(9));
        reg_ensig_cgo_cse <= or_997_rmff;
        reg_ensig_cgo_17_cse <= or_1156_rmff;
        butterFly2_11_tw_h_slc_operator_33_true_2_lshift_psp_2_0_1_0_itm <= MUX_v_2_2_2(STAGE_LOOP_mux1h_nl,
            STD_LOGIC_VECTOR'("11"), nor_4_nl);
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10 <= INNER_LOOP1_r_mux_44_nl
            AND (NOT or_tmp_1138);
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9 <= MUX_s_1_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8,
            INNER_LOOP1_stage_0_9, fsm_output(7));
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8 <= INNER_LOOP1_r_mux_45_nl
            AND (NOT and_192_cse);
        INNER_LOOP1_stage_0 <= (INNER_LOOP1_stage_0 AND (NOT (z_out_2(7)))) OR or_tmp_1138;
        INNER_LOOP1_r_11_4_sva_6_0 <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"), (z_out_2(6
            DOWNTO 0)), (fsm_output(2)));
        INNER_LOOP1_stage_0_2 <= INNER_LOOP1_mux_nl AND (NOT or_tmp_1138);
        INNER_LOOP1_stage_0_3 <= INNER_LOOP1_stage_0_2 AND or_dcpl_214;
        INNER_LOOP1_stage_0_4 <= INNER_LOOP1_stage_0_3 AND or_dcpl_214;
        INNER_LOOP1_stage_0_5 <= INNER_LOOP1_stage_0_4 AND or_dcpl_214;
        INNER_LOOP1_stage_0_6 <= INNER_LOOP1_stage_0_5 AND or_dcpl_214;
        INNER_LOOP1_stage_0_7 <= INNER_LOOP1_stage_0_6 AND or_dcpl_214;
        INNER_LOOP1_stage_0_8 <= INNER_LOOP1_stage_0_7 AND or_dcpl_214;
        INNER_LOOP1_stage_0_9 <= INNER_LOOP1_stage_0_8 AND or_dcpl_214;
        INNER_LOOP1_stage_0_10 <= INNER_LOOP1_r_mux1h_46_nl AND (NOT((fsm_output(10))
            OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(0)) OR (fsm_output(1))));
        INNER_LOOP1_stage_0_11 <= INNER_LOOP1_mux_11_nl AND ((fsm_output(6)) OR (fsm_output(4))
            OR (fsm_output(2)) OR (NOT and_dcpl_90));
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6
            AND (NOT or_tmp_1138);
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5
            AND (NOT or_tmp_1138);
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4
            AND (NOT or_tmp_1138);
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3
            AND (NOT or_tmp_1138);
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2
            AND (NOT or_tmp_1138);
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1
            AND (NOT or_tmp_1138);
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm
            AND (NOT or_tmp_1138);
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm <= MUX_s_1_2_2(INNER_LOOP1_r_INNER_LOOP1_r_and_nl,
            INNER_LOOP1_stage_0, or_dcpl_218);
        INNER_LOOP3_r_11_4_sva_6_0 <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"), (z_out_2(6
            DOWNTO 0)), (fsm_output(7)));
        INNER_LOOP4_r_11_4_sva_6_0 <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"), (z_out_2(6
            DOWNTO 0)), (fsm_output(9)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      modulo_add_1_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_81, (acc_2_nl(32 DOWNTO
          1)), z_out_78, z_out_76, STD_LOGIC_VECTOR'( modulo_add_1_qelse_and_nl &
          modulo_add_1_qelse_or_1_nl & modulo_add_1_qelse_and_4_nl & modulo_add_1_qelse_and_5_nl));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_9 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_8,
          (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) & (fsm_output(9))));
      modulo_add_10_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_72, (acc_6_nl(32 DOWNTO
          1)), z_out_67, z_out_68, z_out_82, STD_LOGIC_VECTOR'( modulo_add_10_qelse_and_nl
          & modulo_add_10_qelse_or_nl & modulo_add_10_qelse_and_5_nl & modulo_add_10_qelse_and_6_nl
          & modulo_add_10_qelse_and_7_nl));
      modulo_add_11_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_71, (acc_10_nl(32 DOWNTO
          1)), z_out_77, z_out_67, z_out_81, STD_LOGIC_VECTOR'( modulo_add_11_qelse_and_nl
          & modulo_add_11_qelse_or_nl & modulo_add_11_qelse_and_5_nl & modulo_add_11_qelse_and_6_nl
          & modulo_add_11_qelse_and_7_nl));
      modulo_add_12_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_70, (acc_14_nl(32 DOWNTO
          1)), z_out_82, z_out_80, STD_LOGIC_VECTOR'( modulo_add_12_qelse_and_nl
          & modulo_add_12_qelse_or_1_nl & modulo_add_12_qelse_and_4_nl & modulo_add_12_qelse_and_5_nl));
      modulo_add_13_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_69, (acc_18_nl(32 DOWNTO
          1)), z_out_81, z_out_79, STD_LOGIC_VECTOR'( modulo_add_13_qelse_and_nl
          & modulo_add_13_qelse_or_1_nl & modulo_add_13_qelse_and_4_nl & modulo_add_13_qelse_and_5_nl));
      modulo_add_14_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_68, (acc_22_nl(32 DOWNTO
          1)), z_out_80, z_out_78, STD_LOGIC_VECTOR'( modulo_add_14_qelse_and_nl
          & modulo_add_14_qelse_or_1_nl & modulo_add_14_qelse_and_4_nl & modulo_add_14_qelse_and_5_nl));
      modulo_add_15_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_67, (acc_26_nl(32 DOWNTO
          1)), z_out_82, z_out_79, z_out_77, STD_LOGIC_VECTOR'( modulo_add_15_qelse_and_nl
          & modulo_add_15_qelse_or_nl & modulo_add_15_qelse_and_5_nl & modulo_add_15_qelse_and_6_nl
          & modulo_add_15_qelse_and_7_nl));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_8 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_7,
          (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) & (fsm_output(9))));
      mult_15_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_15_z_asn_itm_2, mult_31_z_asn_itm_2,
          mult_14_z_asn_itm_2, mult_27_z_asn_itm_2, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_14_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_14_z_asn_itm_2, mult_30_z_asn_itm_2,
          mult_26_z_asn_itm_2, mult_15_z_asn_itm_2, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_13_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_13_z_asn_itm_2, mult_29_z_asn_itm_2,
          mult_28_z_asn_itm_2, STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) &
          (fsm_output(9))));
      mult_12_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_12_z_asn_itm_2, mult_28_z_asn_itm_2,
          mult_29_z_asn_itm_2, STD_LOGIC_VECTOR'( or_tmp_1189 & (fsm_output(4)) &
          (fsm_output(7))));
      mult_11_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_11_z_asn_itm_2, mult_27_z_asn_itm_2,
          mult_15_z_asn_itm_2, mult_26_z_asn_itm_2, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_10_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_10_z_asn_itm_2, mult_26_z_asn_itm_2,
          mult_25_z_asn_itm_2, mult_1_z_asn_itm_2, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_8 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_7,
          (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_7 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_6,
          (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) & (fsm_output(9))));
      mult_15_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_2_z, mult_z_mul_cmp_22_z,
          mult_z_mul_cmp_20_z, STD_LOGIC_VECTOR'( (fsm_output(2)) & or_dcpl_217 &
          (fsm_output(9))));
      mult_14_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_4_z, mult_z_mul_cmp_24_z,
          mult_z_mul_cmp_28_z, STD_LOGIC_VECTOR'( or_tmp_1189 & (fsm_output(4)) &
          (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_7 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_6,
          (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) & (fsm_output(9))));
      mult_13_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_6_z, mult_z_mul_cmp_26_z,
          mult_z_mul_cmp_24_z, mult_z_mul_cmp_12_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_6 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_5,
          (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) & (fsm_output(9))));
      mult_12_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_8_z, mult_z_mul_cmp_28_z,
          mult_z_mul_cmp_12_z, STD_LOGIC_VECTOR'( (fsm_output(2)) & or_dcpl_194 &
          (fsm_output(7))));
      mult_11_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_10_z, mult_z_mul_cmp_30_z,
          mult_z_mul_cmp_8_z, mult_z_mul_cmp_16_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_10_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_12_z, mult_z_mul_cmp_z,
          mult_z_mul_cmp_2_z, STD_LOGIC_VECTOR'( (fsm_output(2)) & or_dcpl_194 &
          (fsm_output(7))));
      mult_1_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_30_z, mult_z_mul_cmp_20_z,
          mult_z_mul_cmp_16_z, mult_z_mul_cmp_26_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_6 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_5,
          (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_5 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_4,
          (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_5 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_4,
          (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_4 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_3,
          (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_4 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_3,
          (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_3 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_2,
          (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_2 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_1,
          (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_3 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_2,
          (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6
          DOWNTO 1)), STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_1 <= MUX1HOT_v_6_3_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_602_itm_9_cse,
          (INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2))
          & or_dcpl_194 & (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_2 <= MUX1HOT_v_6_4_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1,
          (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), (INNER_LOOP3_r_11_4_sva_6_0(6
          DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6 DOWNTO 1)), STD_LOGIC_VECTOR'(
          (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_1 <= MUX1HOT_v_6_4_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), (INNER_LOOP3_r_11_4_sva_6_0(6
          DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6 DOWNTO 1)), STD_LOGIC_VECTOR'(
          (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_2 <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_1,
          (INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 1)), fsm_output(7));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_1 <= MUX1HOT_v_6_3_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_350_itm_9_cse,
          (INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2))
          & or_dcpl_194 & (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_2 <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_1,
          (INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 1)), fsm_output(7));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_1 <= MUX1HOT_v_6_3_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_287_itm_9_cse,
          (INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2))
          & or_dcpl_194 & (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_2 <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_1,
          (INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 1)), fsm_output(7));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_1 <= MUX1HOT_v_6_3_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_224_itm_9_cse,
          (INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2))
          & or_dcpl_194 & (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_2 <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_1,
          (INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 1)), fsm_output(7));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_1 <= MUX1HOT_v_6_3_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_161_itm_9_cse,
          (INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2))
          & or_dcpl_194 & (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_2 <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_1,
          (INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 1)), fsm_output(7));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_1 <= MUX1HOT_v_6_3_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_114_itm_9_cse,
          (INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2))
          & or_dcpl_194 & (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_2 <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_1,
          (INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 1)), fsm_output(7));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_2 <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_1,
          (INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 1)), fsm_output(7));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_1 <= MUX1HOT_v_6_3_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_9, (INNER_LOOP3_r_11_4_sva_6_0(6
          DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2)) & or_dcpl_194 & (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_2 <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_1,
          (INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 1)), fsm_output(7));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_1 <= MUX1HOT_v_6_3_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse,
          (INNER_LOOP3_r_11_4_sva_6_0(6 DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2))
          & or_dcpl_194 & (fsm_output(7))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1 <= MUX_v_6_2_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_570_itm_8_cse,
          or_dcpl_218);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_1 <= MUX_v_6_2_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_381_itm_8_cse,
          or_dcpl_218);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_1 <= MUX_v_6_2_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_318_itm_8_cse,
          or_dcpl_218);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_1 <= MUX_v_6_2_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_255_itm_8_cse,
          or_dcpl_218);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_1 <= MUX_v_6_2_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_192_itm_8_cse,
          or_dcpl_218);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_1 <= MUX_v_6_2_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_129_itm_8_cse,
          or_dcpl_218);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_1 <= MUX_v_6_2_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_633_itm_8_cse,
          or_dcpl_218);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_1 <= MUX1HOT_v_6_4_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), (INNER_LOOP2_r_11_4_sva_6_0(6 DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_8,
          (INNER_LOOP4_r_11_4_sva_6_0(6 DOWNTO 1)), STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_1 <= MUX_v_6_2_2((INNER_LOOP1_r_11_4_sva_6_0(6
          DOWNTO 1)), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_8, or_dcpl_218);
      mult_16_z_asn_itm_3 <= MUX_v_32_2_2(mult_31_z_asn_itm_2, mult_10_z_asn_itm_2,
          or_dcpl_217);
      mult_17_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_1_z_asn_itm_2, mult_11_z_asn_itm_2,
          mult_31_z_asn_itm_2, mult_10_z_asn_itm_2, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_18_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_23_z_asn_itm_2, mult_12_z_asn_itm_2,
          mult_24_z_asn_itm_2, STD_LOGIC_VECTOR'( or_tmp_1189 & (fsm_output(4)) &
          (fsm_output(7))));
      mult_19_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_24_z_asn_itm_2, mult_13_z_asn_itm_2,
          mult_23_z_asn_itm_2, STD_LOGIC_VECTOR'( or_tmp_1189 & (fsm_output(4)) &
          (fsm_output(7))));
      mult_20_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_25_z_asn_itm_2, mult_14_z_asn_itm_2,
          mult_28_z_asn_itm_2, mult_13_z_asn_itm_2, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_21_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_26_z_asn_itm_2, mult_15_z_asn_itm_2,
          mult_11_z_asn_itm_2, mult_30_z_asn_itm_2, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_22_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_27_z_asn_itm_2, mult_1_z_asn_itm_2,
          mult_14_z_asn_itm_2, STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) &
          (fsm_output(9))));
      mult_23_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_28_z_asn_itm_2, mult_23_z_asn_itm_2,
          mult_1_z_asn_itm_2, mult_25_z_asn_itm_2, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_24_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_29_z_asn_itm_2, mult_24_z_asn_itm_2,
          mult_12_z_asn_itm_2, STD_LOGIC_VECTOR'( or_tmp_1189 & (fsm_output(4)) &
          (fsm_output(7))));
      mult_25_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_30_z_asn_itm_2, mult_25_z_asn_itm_2,
          mult_11_z_asn_itm_2, STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) &
          (fsm_output(9))));
      modulo_add_23_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_80, (acc_29_nl(32 DOWNTO
          1)), z_out_77, z_out_75, STD_LOGIC_VECTOR'( modulo_add_23_qelse_and_nl
          & modulo_add_23_qelse_or_1_nl & modulo_add_23_qelse_and_4_nl & modulo_add_23_qelse_and_5_nl));
      modulo_add_24_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_79, (acc_32_nl(32 DOWNTO
          1)), z_out_76, z_out_74, STD_LOGIC_VECTOR'( modulo_add_24_qelse_and_nl
          & modulo_add_24_qelse_or_1_nl & modulo_add_24_qelse_and_4_nl & modulo_add_24_qelse_and_5_nl));
      modulo_add_25_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_78, (acc_34_nl(32 DOWNTO
          1)), z_out_75, z_out_73, STD_LOGIC_VECTOR'( modulo_add_25_qelse_and_nl
          & modulo_add_25_qelse_or_1_nl & modulo_add_25_qelse_and_4_nl & modulo_add_25_qelse_and_5_nl));
      modulo_add_26_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_77, (acc_37_nl(32 DOWNTO
          1)), z_out_76, z_out_74, z_out_72, STD_LOGIC_VECTOR'( modulo_add_26_qelse_and_nl
          & modulo_add_26_qelse_or_nl & modulo_add_26_qelse_and_5_nl & modulo_add_26_qelse_and_6_nl
          & modulo_add_26_qelse_and_7_nl));
      modulo_add_27_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_76, (acc_39_nl(32 DOWNTO
          1)), z_out_75, z_out_73, z_out_71, STD_LOGIC_VECTOR'( modulo_add_27_qelse_and_nl
          & modulo_add_27_qelse_or_nl & modulo_add_27_qelse_and_5_nl & modulo_add_27_qelse_and_6_nl
          & modulo_add_27_qelse_and_7_nl));
      modulo_add_28_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_75, (acc_42_nl(32 DOWNTO
          1)), z_out_74, z_out_72, z_out_70, STD_LOGIC_VECTOR'( modulo_add_28_qelse_and_nl
          & modulo_add_28_qelse_or_nl & modulo_add_28_qelse_and_5_nl & modulo_add_28_qelse_and_6_nl
          & modulo_add_28_qelse_and_7_nl));
      modulo_add_29_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_74, (acc_44_nl(32 DOWNTO
          1)), z_out_73, z_out_71, z_out_69, STD_LOGIC_VECTOR'( modulo_add_29_qelse_and_nl
          & modulo_add_29_qelse_or_nl & modulo_add_29_qelse_and_5_nl & modulo_add_29_qelse_and_6_nl
          & modulo_add_29_qelse_and_7_nl));
      modulo_add_30_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_73, (acc_47_nl(32 DOWNTO
          1)), z_out_72, z_out_70, z_out_68, STD_LOGIC_VECTOR'( modulo_add_30_qelse_and_nl
          & modulo_add_30_qelse_or_nl & modulo_add_30_qelse_and_5_nl & modulo_add_30_qelse_and_6_nl
          & modulo_add_30_qelse_and_7_nl));
      modulo_add_31_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_82, (acc_49_nl(32 DOWNTO
          1)), z_out_71, z_out_69, z_out_67, STD_LOGIC_VECTOR'( modulo_add_31_qelse_and_nl
          & modulo_add_31_qelse_or_nl & modulo_add_31_qelse_and_5_nl & modulo_add_31_qelse_and_6_nl
          & modulo_add_31_qelse_and_7_nl));
      mult_23_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_28_z, mult_z_mul_cmp_18_z,
          mult_z_mul_cmp_6_z, mult_z_mul_cmp_10_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_24_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_26_z, mult_z_mul_cmp_16_z,
          mult_z_mul_cmp_10_z, mult_z_mul_cmp_2_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_25_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_24_z, mult_z_mul_cmp_14_z,
          mult_z_mul_cmp_18_z, mult_z_mul_cmp_8_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_26_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_22_z, mult_z_mul_cmp_12_z,
          mult_z_mul_cmp_26_z, mult_z_mul_cmp_18_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_27_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_20_z, mult_z_mul_cmp_10_z,
          mult_z_mul_cmp_30_z, mult_z_mul_cmp_24_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_28_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_18_z, mult_z_mul_cmp_8_z,
          mult_z_mul_cmp_20_z, mult_z_mul_cmp_30_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_29_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_16_z, mult_z_mul_cmp_6_z,
          mult_z_mul_cmp_14_z, mult_z_mul_cmp_22_z, STD_LOGIC_VECTOR'( (fsm_output(2))
          & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
      mult_30_z_asn_itm_1 <= MUX_v_32_2_2(mult_z_mul_cmp_14_z, mult_z_mul_cmp_4_z,
          or_dcpl_217);
      mult_31_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_z, mult_z_mul_cmp_2_z,
          mult_z_mul_cmp_6_z, STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(4)) &
          (fsm_output(9))));
      tmp_10_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_0_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_10_i_qa_d(31
          DOWNTO 0)), (xt_rsc_0_4_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_0_i_qa_d(31 DOWNTO
          0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
          & (fsm_output(9))));
      tmp_102_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_2_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_12_i_qa_d(31
          DOWNTO 0)), (xt_rsc_0_6_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_2_i_qa_d(31 DOWNTO
          0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
          & (fsm_output(9))));
      tmp_104_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_4_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_14_i_qa_d(31
          DOWNTO 0)), (xt_rsc_0_8_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_4_i_qa_d(31 DOWNTO
          0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
          & (fsm_output(9))));
      tmp_106_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_6_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_16_i_qa_d(31
          DOWNTO 0)), (xt_rsc_0_10_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_6_i_qa_d(31 DOWNTO
          0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
          & (fsm_output(9))));
      tmp_108_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_8_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_18_i_qa_d(31
          DOWNTO 0)), (xt_rsc_0_12_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_8_i_qa_d(31 DOWNTO
          0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
          & (fsm_output(9))));
      tmp_110_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_10_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_2_i_qa_d(31
          DOWNTO 0)), (xt_rsc_0_14_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_10_i_qa_d(31 DOWNTO
          0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
          & (fsm_output(9))));
      tmp_112_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_12_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_20_i_qa_d(31
          DOWNTO 0)), (xt_rsc_0_16_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_12_i_qa_d(31 DOWNTO
          0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
          & (fsm_output(9))));
      tmp_114_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_14_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_22_i_qa_d(31
          DOWNTO 0)), (xt_rsc_0_18_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_14_i_qa_d(31 DOWNTO
          0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
          & (fsm_output(9))));
      tmp_116_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_16_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_24_i_qa_d(31
          DOWNTO 0)), (xt_rsc_0_20_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_16_i_qa_d(31 DOWNTO
          0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
          & (fsm_output(9))));
      tmp_118_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_18_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_26_i_qa_d(31
          DOWNTO 0)), (xt_rsc_0_22_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_18_i_qa_d(31 DOWNTO
          0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
          & (fsm_output(9))));
      tmp_120_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_20_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_28_i_qa_d(31
          DOWNTO 0)), (xt_rsc_0_24_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_20_i_qa_d(31 DOWNTO
          0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
          & (fsm_output(9))));
      tmp_122_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_22_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_30_i_qa_d(31
          DOWNTO 0)), (xt_rsc_0_26_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_22_i_qa_d(31 DOWNTO
          0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
          & (fsm_output(9))));
      tmp_124_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_24_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_4_i_qa_d(31
          DOWNTO 0)), (xt_rsc_0_28_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_24_i_qa_d(31 DOWNTO
          0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
          & (fsm_output(9))));
      tmp_126_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_26_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_6_i_qa_d(31
          DOWNTO 0)), (xt_rsc_0_30_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_26_i_qa_d(31 DOWNTO
          0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
          & (fsm_output(9))));
      tmp_60_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_28_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_8_i_qa_d(31
          DOWNTO 0)), (xt_rsc_0_0_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_28_i_qa_d(31 DOWNTO
          0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
          & (fsm_output(9))));
      tmp_62_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_30_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_0_i_qa_d(31
          DOWNTO 0)), (xt_rsc_0_2_i_qa_d(31 DOWNTO 0)), (yt_rsc_0_30_i_qa_d(31 DOWNTO
          0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
          & (fsm_output(9))));
      reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd <= (z_out_49(31)) AND (NOT(modulo_sub_16_qelse_and_ssc
          OR modulo_sub_16_qelse_and_ssc_1));
      reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_66(30 DOWNTO
          0)), (z_out_49(30 DOWNTO 0)), (z_out_51(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_16_qelse_and_ssc & modulo_sub_16_qelse_or_nl & modulo_sub_16_qelse_and_ssc_1));
      reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd <= (z_out_47(31)) AND (NOT(modulo_sub_17_qelse_and_ssc
          OR modulo_sub_17_qelse_and_ssc_1));
      reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_56(30 DOWNTO
          0)), (z_out_47(30 DOWNTO 0)), (z_out_52(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_17_qelse_and_ssc & modulo_sub_17_qelse_or_nl & modulo_sub_17_qelse_and_ssc_1));
      reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd <= (z_out_46(31)) AND (NOT(modulo_sub_18_qelse_and_ssc
          OR modulo_sub_18_qelse_and_ssc_1));
      reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_63(30 DOWNTO
          0)), (z_out_46(30 DOWNTO 0)), (z_out_53(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_18_qelse_and_ssc & modulo_sub_18_qelse_or_nl & modulo_sub_18_qelse_and_ssc_1));
      reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd <= (z_out_44(31)) AND (NOT(modulo_sub_19_qelse_and_ssc
          OR modulo_sub_19_qelse_and_ssc_1));
      reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_64(30 DOWNTO
          0)), (z_out_44(30 DOWNTO 0)), (z_out_54(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_19_qelse_and_ssc & modulo_sub_19_qelse_or_nl & modulo_sub_19_qelse_and_ssc_1));
      reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd <= (z_out_42(31)) AND (NOT(modulo_sub_20_qelse_and_ssc
          OR modulo_sub_20_qelse_and_ssc_1));
      reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_65(30 DOWNTO
          0)), (z_out_42(30 DOWNTO 0)), (z_out_55(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_20_qelse_and_ssc & modulo_sub_20_qelse_or_nl & modulo_sub_20_qelse_and_ssc_1));
      reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd <= (z_out_41(31)) AND (NOT(modulo_sub_21_qelse_and_ssc
          OR modulo_sub_21_qelse_and_ssc_1));
      reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_51(30 DOWNTO
          0)), (z_out_41(30 DOWNTO 0)), (z_out_56(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_21_qelse_and_ssc & modulo_sub_21_qelse_or_nl & modulo_sub_21_qelse_and_ssc_1));
      reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd <= (z_out_39(31)) AND (NOT(modulo_sub_22_qelse_and_ssc
          OR modulo_sub_22_qelse_and_ssc_1));
      reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_52(30 DOWNTO
          0)), (z_out_39(30 DOWNTO 0)), (z_out_57(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_22_qelse_and_ssc & modulo_sub_22_qelse_or_nl & modulo_sub_22_qelse_and_ssc_1));
      reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd <= (z_out_37(31)) AND (NOT(modulo_sub_23_qelse_and_ssc
          OR modulo_sub_23_qelse_and_ssc_1));
      reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_53(30 DOWNTO
          0)), (z_out_37(30 DOWNTO 0)), (z_out_58(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_23_qelse_and_ssc & modulo_sub_23_qelse_or_nl & modulo_sub_23_qelse_and_ssc_1));
      reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd <= (z_out_36(31)) AND (NOT(modulo_sub_24_qelse_and_ssc
          OR modulo_sub_24_qelse_and_ssc_1));
      reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_54(30 DOWNTO
          0)), (z_out_36(30 DOWNTO 0)), (z_out_59(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_24_qelse_and_ssc & modulo_sub_24_qelse_or_nl & modulo_sub_24_qelse_and_ssc_1));
      reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd <= (z_out_34(31)) AND (NOT(modulo_sub_25_qelse_and_ssc
          OR modulo_sub_25_qelse_and_ssc_1));
      reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_55(30 DOWNTO
          0)), (z_out_34(30 DOWNTO 0)), (z_out_60(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_25_qelse_and_ssc & modulo_sub_25_qelse_or_nl & modulo_sub_25_qelse_and_ssc_1));
      reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd <= (z_out_32(31)) AND (NOT(modulo_sub_26_qelse_and_ssc
          OR modulo_sub_26_qelse_and_ssc_1));
      reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_57(30 DOWNTO
          0)), (z_out_32(30 DOWNTO 0)), (z_out_61(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_26_qelse_and_ssc & modulo_sub_26_qelse_or_nl & modulo_sub_26_qelse_and_ssc_1));
      reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd <= (z_out_31(31)) AND (NOT(modulo_sub_27_qelse_and_ssc
          OR modulo_sub_27_qelse_and_ssc_1));
      reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_58(30 DOWNTO
          0)), (z_out_31(30 DOWNTO 0)), (z_out_62(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_27_qelse_and_ssc & modulo_sub_27_qelse_or_nl & modulo_sub_27_qelse_and_ssc_1));
      reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd <= (z_out_29(31)) AND (NOT(modulo_sub_28_qelse_and_ssc
          OR modulo_sub_28_qelse_and_ssc_1));
      reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_59(30 DOWNTO
          0)), (z_out_29(30 DOWNTO 0)), (z_out_63(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_28_qelse_and_ssc & modulo_sub_28_qelse_or_nl & modulo_sub_28_qelse_and_ssc_1));
      reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd <= (z_out_26(31)) AND (NOT(modulo_sub_29_qelse_and_ssc
          OR modulo_sub_29_qelse_and_ssc_1));
      reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_60(30 DOWNTO
          0)), (z_out_26(30 DOWNTO 0)), (z_out_64(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_29_qelse_and_ssc & modulo_sub_29_qelse_or_nl & modulo_sub_29_qelse_and_ssc_1));
      reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd <= (z_out_24(31)) AND (NOT(modulo_sub_30_qelse_and_ssc
          OR modulo_sub_30_qelse_and_ssc_1));
      reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_61(30 DOWNTO
          0)), (z_out_24(30 DOWNTO 0)), (z_out_65(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_30_qelse_and_ssc & modulo_sub_30_qelse_or_nl & modulo_sub_30_qelse_and_ssc_1));
      reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd <= (z_out_21(31)) AND (NOT(modulo_sub_31_qelse_and_ssc
          OR modulo_sub_31_qelse_and_ssc_1));
      reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_62(30 DOWNTO
          0)), (z_out_21(30 DOWNTO 0)), (z_out_66(30 DOWNTO 0)), STD_LOGIC_VECTOR'(
          modulo_sub_31_qelse_and_ssc & modulo_sub_31_qelse_or_nl & modulo_sub_31_qelse_and_ssc_1));
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_3 <= reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_1 <= MUX_v_6_2_2((INNER_LOOP2_r_11_4_sva_6_0(6
          DOWNTO 1)), (INNER_LOOP4_r_11_4_sva_6_0(6 DOWNTO 1)), fsm_output(9));
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_12_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5) = '1'
          ) THEN
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_114_itm_9_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_12_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4) = '1'
          ) THEN
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_161_itm_9_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_12_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3) = '1'
          ) THEN
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_224_itm_9_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_12_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2) = '1'
          ) THEN
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_287_itm_9_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_12_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1) = '1'
          ) THEN
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_350_itm_9_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_12_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm) = '1' )
          THEN
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_12_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_9 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_12_cse = '1' ) THEN
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_602_itm_9_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_13 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4) = '1'
          ) THEN
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_129_itm_8_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_13 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3) = '1'
          ) THEN
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_192_itm_8_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_13 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2) = '1'
          ) THEN
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_255_itm_8_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_13 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1) = '1'
          ) THEN
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_318_itm_8_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_13 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm) = '1'
          ) THEN
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_381_itm_8_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_13 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_13 = '1' ) THEN
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_570_itm_8_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_7;
        tmp_10_sva_7 <= tmp_10_sva_6;
        tmp_102_sva_7 <= tmp_102_sva_6;
        tmp_104_sva_7 <= tmp_104_sva_6;
        tmp_106_sva_7 <= tmp_106_sva_6;
        tmp_108_sva_7 <= tmp_108_sva_6;
        tmp_110_sva_7 <= tmp_110_sva_6;
        tmp_112_sva_7 <= tmp_112_sva_6;
        tmp_114_sva_7 <= tmp_114_sva_6;
        tmp_116_sva_7 <= tmp_116_sva_6;
        tmp_118_sva_7 <= tmp_118_sva_6;
        tmp_120_sva_7 <= tmp_120_sva_6;
        tmp_122_sva_7 <= tmp_122_sva_6;
        tmp_124_sva_7 <= tmp_124_sva_6;
        tmp_126_sva_7 <= tmp_126_sva_6;
        tmp_60_sva_7 <= tmp_60_sva_6;
        tmp_62_sva_7 <= tmp_62_sva_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_13 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5) = '1'
          ) THEN
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_633_itm_8_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP1_stage_0_8 = '1' ) THEN
        mult_15_res_lpi_3_dfm_1 <= mult_15_res_lpi_3_dfm_1_mx0;
        mult_14_res_lpi_3_dfm_1 <= mult_14_res_lpi_3_dfm_1_mx0;
        mult_13_res_lpi_3_dfm_1 <= mult_13_res_lpi_3_dfm_1_mx0;
        mult_12_res_lpi_3_dfm_1 <= mult_12_res_lpi_3_dfm_1_mx0;
        mult_11_res_lpi_3_dfm_1 <= mult_11_res_lpi_3_dfm_1_mx0;
        mult_10_res_lpi_3_dfm_1 <= mult_10_res_lpi_3_dfm_1_mx0;
        mult_9_res_lpi_3_dfm_1 <= mult_9_res_lpi_3_dfm_1_mx0;
        mult_8_res_lpi_3_dfm_1 <= mult_8_res_lpi_3_dfm_1_mx0;
        mult_7_res_lpi_3_dfm_1 <= mult_7_res_lpi_3_dfm_1_mx0;
        mult_6_res_lpi_3_dfm_1 <= mult_6_res_lpi_3_dfm_1_mx0;
        mult_5_res_lpi_3_dfm_1 <= mult_5_res_lpi_3_dfm_1_mx0;
        mult_4_res_lpi_3_dfm_1 <= mult_4_res_lpi_3_dfm_1_mx0;
        mult_3_res_lpi_3_dfm_1 <= mult_3_res_lpi_3_dfm_1_mx0;
        mult_2_res_lpi_3_dfm_1 <= mult_2_res_lpi_3_dfm_1_mx0;
        mult_1_res_lpi_3_dfm_1 <= mult_1_res_lpi_3_dfm_1_mx0;
        mult_res_lpi_3_dfm_1 <= mult_res_lpi_3_dfm_1_mx0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_20_false_acc_cse_sva <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( (NOT(or_dcpl_233 OR or_dcpl_210)) = '1' ) THEN
        operator_20_false_acc_cse_sva <= MUX_v_3_2_2(z_out_1, (z_out(2 DOWNTO 0)),
            fsm_output(6));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_22 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_44_cse = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_45 = '1' ) THEN
        mult_15_z_asn_itm_2 <= mult_15_z_asn_itm_1;
        mult_14_z_asn_itm_2 <= mult_14_z_asn_itm_1;
        mult_13_z_asn_itm_2 <= mult_13_z_asn_itm_1;
        mult_12_z_asn_itm_2 <= mult_12_z_asn_itm_1;
        mult_11_z_asn_itm_2 <= mult_11_z_asn_itm_1;
        mult_10_z_asn_itm_2 <= mult_10_z_asn_itm_1;
        mult_1_z_asn_itm_2 <= mult_1_z_asn_itm_1;
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_5;
        mult_23_z_asn_itm_2 <= mult_23_z_asn_itm_1;
        mult_24_z_asn_itm_2 <= mult_24_z_asn_itm_1;
        mult_25_z_asn_itm_2 <= mult_25_z_asn_itm_1;
        mult_26_z_asn_itm_2 <= mult_26_z_asn_itm_1;
        mult_27_z_asn_itm_2 <= mult_27_z_asn_itm_1;
        mult_28_z_asn_itm_2 <= mult_28_z_asn_itm_1;
        mult_29_z_asn_itm_2 <= mult_29_z_asn_itm_1;
        mult_30_z_asn_itm_2 <= mult_30_z_asn_itm_1;
        mult_31_z_asn_itm_2 <= mult_31_z_asn_itm_1;
        tmp_10_sva_5 <= tmp_10_sva_4;
        tmp_102_sva_5 <= tmp_102_sva_4;
        tmp_104_sva_5 <= tmp_104_sva_4;
        tmp_106_sva_5 <= tmp_106_sva_4;
        tmp_108_sva_5 <= tmp_108_sva_4;
        tmp_110_sva_5 <= tmp_110_sva_4;
        tmp_112_sva_5 <= tmp_112_sva_4;
        tmp_114_sva_5 <= tmp_114_sva_4;
        tmp_116_sva_5 <= tmp_116_sva_4;
        tmp_118_sva_5 <= tmp_118_sva_4;
        tmp_120_sva_5 <= tmp_120_sva_4;
        tmp_122_sva_5 <= tmp_122_sva_4;
        tmp_124_sva_5 <= tmp_124_sva_4;
        tmp_126_sva_5 <= tmp_126_sva_4;
        tmp_60_sva_5 <= tmp_60_sva_4;
        tmp_62_sva_5 <= tmp_62_sva_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_22 = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_6;
        tmp_10_sva_6 <= tmp_10_sva_5;
        tmp_102_sva_6 <= tmp_102_sva_5;
        tmp_104_sva_6 <= tmp_104_sva_5;
        tmp_106_sva_6 <= tmp_106_sva_5;
        tmp_108_sva_6 <= tmp_108_sva_5;
        tmp_110_sva_6 <= tmp_110_sva_5;
        tmp_112_sva_6 <= tmp_112_sva_5;
        tmp_114_sva_6 <= tmp_114_sva_5;
        tmp_116_sva_6 <= tmp_116_sva_5;
        tmp_118_sva_6 <= tmp_118_sva_5;
        tmp_120_sva_6 <= tmp_120_sva_5;
        tmp_122_sva_6 <= tmp_122_sva_5;
        tmp_124_sva_6 <= tmp_124_sva_5;
        tmp_126_sva_6 <= tmp_126_sva_5;
        tmp_60_sva_6 <= tmp_60_sva_5;
        tmp_62_sva_6 <= tmp_62_sva_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_44_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm) = '1' )
          THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_22 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_44_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_22 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_44_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_22 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_44_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_22 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_44_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_44_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_22 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_44_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_22 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_45 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_64_cse = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_64_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_45 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_64_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm) = '1' )
          THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_45 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_64_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_45 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_64_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_45 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_64_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_64_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_45 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_64_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_45 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_65 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_84_cse = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_65 = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_4;
        tmp_10_sva_4 <= tmp_10_sva_3;
        tmp_102_sva_4 <= tmp_102_sva_3;
        tmp_104_sva_4 <= tmp_104_sva_3;
        tmp_106_sva_4 <= tmp_106_sva_3;
        tmp_108_sva_4 <= tmp_108_sva_3;
        tmp_110_sva_4 <= tmp_110_sva_3;
        tmp_112_sva_4 <= tmp_112_sva_3;
        tmp_114_sva_4 <= tmp_114_sva_3;
        tmp_116_sva_4 <= tmp_116_sva_3;
        tmp_118_sva_4 <= tmp_118_sva_3;
        tmp_120_sva_4 <= tmp_120_sva_3;
        tmp_122_sva_4 <= tmp_122_sva_3;
        tmp_124_sva_4 <= tmp_124_sva_3;
        tmp_126_sva_4 <= tmp_126_sva_3;
        tmp_60_sva_4 <= tmp_60_sva_3;
        tmp_62_sva_4 <= tmp_62_sva_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_84_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_65 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_84_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_65 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_84_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm) = '1' )
          THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_65 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_84_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_65 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_84_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_84_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_65 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_84_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_65 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_101 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_103_cse = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_101 = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_3;
        tmp_10_sva_3 <= tmp_10_sva_2;
        tmp_102_sva_3 <= tmp_102_sva_2;
        tmp_104_sva_3 <= tmp_104_sva_2;
        tmp_106_sva_3 <= tmp_106_sva_2;
        tmp_108_sva_3 <= tmp_108_sva_2;
        tmp_110_sva_3 <= tmp_110_sva_2;
        tmp_112_sva_3 <= tmp_112_sva_2;
        tmp_114_sva_3 <= tmp_114_sva_2;
        tmp_116_sva_3 <= tmp_116_sva_2;
        tmp_118_sva_3 <= tmp_118_sva_2;
        tmp_120_sva_3 <= tmp_120_sva_2;
        tmp_122_sva_3 <= tmp_122_sva_2;
        tmp_124_sva_3 <= tmp_124_sva_2;
        tmp_126_sva_3 <= tmp_126_sva_2;
        tmp_60_sva_3 <= tmp_60_sva_2;
        tmp_62_sva_3 <= tmp_62_sva_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_103_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_101 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_103_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_101 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_103_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_101 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_103_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_101 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_103_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_103_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_101 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_103_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_101 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_121 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_123_cse = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_121 = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_2;
        tmp_10_sva_2 <= tmp_10_sva_1;
        tmp_102_sva_2 <= tmp_102_sva_1;
        tmp_104_sva_2 <= tmp_104_sva_1;
        tmp_106_sva_2 <= tmp_106_sva_1;
        tmp_108_sva_2 <= tmp_108_sva_1;
        tmp_110_sva_2 <= tmp_110_sva_1;
        tmp_112_sva_2 <= tmp_112_sva_1;
        tmp_114_sva_2 <= tmp_114_sva_1;
        tmp_116_sva_2 <= tmp_116_sva_1;
        tmp_118_sva_2 <= tmp_118_sva_1;
        tmp_120_sva_2 <= tmp_120_sva_1;
        tmp_122_sva_2 <= tmp_122_sva_1;
        tmp_124_sva_2 <= tmp_124_sva_1;
        tmp_126_sva_2 <= tmp_126_sva_1;
        tmp_60_sva_2 <= tmp_60_sva_1;
        tmp_62_sva_2 <= tmp_62_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_123_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_121 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_123_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_121 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_123_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_121 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_123_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_121 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_123_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_123_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_121 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_123_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_dcpl_121 OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_142_cse = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_143_cse = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_142_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_143_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_142_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_143_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_142_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_143_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_142_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_143_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_142_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_143_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_142_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_143_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_142_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (or_143_cse OR INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2) = '1'
          ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP2_r_11_4_sva_6_0 <= STD_LOGIC_VECTOR'( "0000000");
      ELSIF ( (fsm_output(2)) = '0' ) THEN
        INNER_LOOP2_r_11_4_sva_6_0 <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"), STAGE_LOOP_base_STAGE_LOOP_base_mux_nl,
            INNER_LOOP2_r_or_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_9 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_8;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_9 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 = '1' ) THEN
        reg_mult_31_res_lpi_3_dfm_1_cse <= mult_15_res_lpi_3_dfm_1_mx0;
        reg_mult_30_res_lpi_3_dfm_1_cse <= mult_14_res_lpi_3_dfm_1_mx0;
        reg_mult_29_res_lpi_3_dfm_1_cse <= mult_13_res_lpi_3_dfm_1_mx0;
        reg_mult_28_res_lpi_3_dfm_1_cse <= mult_12_res_lpi_3_dfm_1_mx0;
        reg_mult_27_res_lpi_3_dfm_1_cse <= mult_11_res_lpi_3_dfm_1_mx0;
        reg_mult_26_res_lpi_3_dfm_1_cse <= mult_10_res_lpi_3_dfm_1_mx0;
        reg_mult_25_res_lpi_3_dfm_1_cse <= mult_9_res_lpi_3_dfm_1_mx0;
        reg_mult_24_res_lpi_3_dfm_1_cse <= mult_8_res_lpi_3_dfm_1_mx0;
        reg_mult_23_res_lpi_3_dfm_1_cse <= mult_7_res_lpi_3_dfm_1_mx0;
        reg_mult_22_res_lpi_3_dfm_1_cse <= mult_6_res_lpi_3_dfm_1_mx0;
        reg_mult_21_res_lpi_3_dfm_1_cse <= mult_5_res_lpi_3_dfm_1_mx0;
        reg_mult_20_res_lpi_3_dfm_1_cse <= mult_4_res_lpi_3_dfm_1_mx0;
        reg_mult_19_res_lpi_3_dfm_1_cse <= mult_3_res_lpi_3_dfm_1_mx0;
        reg_mult_18_res_lpi_3_dfm_1_cse <= mult_2_res_lpi_3_dfm_1_mx0;
        reg_mult_17_res_lpi_3_dfm_1_cse <= mult_1_res_lpi_3_dfm_1_mx0;
        reg_mult_16_res_lpi_3_dfm_1_cse <= mult_res_lpi_3_dfm_1_mx0;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_8 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_7;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_8 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (fsm_output(4)) = '0' ) THEN
        operator_33_true_1_lshift_psp_9_4_sva <= z_out(9 DOWNTO 4);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_7 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_6;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_7 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_6 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_5;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_6 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_5 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_4;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_5 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_4 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_3;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_4 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_3 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_2 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        butterFly2_15_tw_equal_tmp_1 <= '0';
        butterFly2_15_tw_equal_tmp_3_1 <= '0';
        butterFly2_15_tw_equal_tmp_5_1 <= '0';
        butterFly2_15_tw_equal_tmp_6_1 <= '0';
        butterFly2_15_tw_equal_tmp_7_1 <= '0';
      ELSIF ( INNER_LOOP1_stage_0 = '1' ) THEN
        butterFly2_15_tw_equal_tmp_1 <= NOT(CONV_SL_1_1(operator_20_false_acc_cse_sva/=STD_LOGIC_VECTOR'("000")));
        butterFly2_15_tw_equal_tmp_3_1 <= CONV_SL_1_1(operator_20_false_acc_cse_sva=STD_LOGIC_VECTOR'("011"));
        butterFly2_15_tw_equal_tmp_5_1 <= CONV_SL_1_1(operator_20_false_acc_cse_sva=STD_LOGIC_VECTOR'("101"));
        butterFly2_15_tw_equal_tmp_6_1 <= CONV_SL_1_1(operator_20_false_acc_cse_sva=STD_LOGIC_VECTOR'("110"));
        butterFly2_15_tw_equal_tmp_7_1 <= CONV_SL_1_1(operator_20_false_acc_cse_sva=STD_LOGIC_VECTOR'("111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_33_true_3_lshift_psp_1_0_sva <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (fsm_output(9)) = '0' ) THEN
        operator_33_true_3_lshift_psp_1_0_sva <= operator_33_true_3_lshift_psp_1_0_sva_mx0w3;
      END IF;
    END IF;
  END PROCESS;
  butterFly2_21_tw_butterFly2_21_tw_or_nl <= c_1_sva OR INNER_LOOP4_nor_tmp;
  c_mux_nl <= MUX_s_1_2_2((operator_20_false_acc_cse_sva(0)), butterFly2_21_tw_butterFly2_21_tw_or_nl,
      fsm_output(9));
  STAGE_LOOP_and_nl <= (NOT (fsm_output(7))) AND or_tmp_1134;
  STAGE_LOOP_mux1h_nl <= MUX1HOT_v_2_5_2((operator_20_false_acc_cse_sva(2 DOWNTO
      1)), (z_out(1 DOWNTO 0)), (operator_20_false_acc_cse_sva(1 DOWNTO 0)), operator_33_true_3_lshift_psp_1_0_sva_mx0w3,
      operator_33_true_3_lshift_psp_1_0_sva, STD_LOGIC_VECTOR'( (fsm_output(5)) &
      STAGE_LOOP_and_nl & (fsm_output(7)) & (fsm_output(8)) & (fsm_output(9))));
  nor_4_nl <= NOT((fsm_output(8)) OR (fsm_output(5)) OR (fsm_output(6)) OR (NOT and_dcpl_90));
  INNER_LOOP1_r_mux_44_nl <= MUX_s_1_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7, or_dcpl_218);
  modulo_add_1_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(z_out_81, z_out_78, z_out_76, STD_LOGIC_VECTOR'(
      modulo_add_1_qelse_or_m1c & (fsm_output(7)) & (fsm_output(9))));
  acc_2_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_1_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_1_qelse_and_nl <= (NOT z_out_83_32) AND modulo_add_1_qelse_or_m1c;
  modulo_add_1_qelse_or_1_nl <= (z_out_83_32 AND modulo_add_1_qelse_or_m1c) OR (z_out_83_32
      AND (fsm_output(7))) OR (z_out_85_32 AND (fsm_output(9)));
  modulo_add_1_qelse_and_4_nl <= (NOT z_out_83_32) AND (fsm_output(7));
  modulo_add_1_qelse_and_5_nl <= (NOT z_out_85_32) AND (fsm_output(9));
  modulo_add_10_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_72, z_out_67, z_out_68,
      z_out_82, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  acc_6_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_10_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_10_qelse_and_nl <= (NOT z_out_84_32) AND (fsm_output(2));
  modulo_add_10_qelse_or_nl <= (z_out_84_32 AND (fsm_output(2))) OR (z_out_84_32
      AND (fsm_output(4))) OR (z_out_84_32 AND (fsm_output(7))) OR (z_out_86_32 AND
      (fsm_output(9)));
  modulo_add_10_qelse_and_5_nl <= (NOT z_out_84_32) AND (fsm_output(4));
  modulo_add_10_qelse_and_6_nl <= (NOT z_out_84_32) AND (fsm_output(7));
  modulo_add_10_qelse_and_7_nl <= (NOT z_out_86_32) AND (fsm_output(9));
  modulo_add_11_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_71, z_out_77, z_out_67,
      z_out_81, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_11_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_11_qelse_and_nl <= (NOT z_out_86_32) AND (fsm_output(2));
  modulo_add_11_qelse_or_nl <= (z_out_86_32 AND (fsm_output(2))) OR (z_out_86_32
      AND (fsm_output(4))) OR (z_out_87_32 AND (fsm_output(7))) OR (z_out_87_32 AND
      (fsm_output(9)));
  modulo_add_11_qelse_and_5_nl <= (NOT z_out_86_32) AND (fsm_output(4));
  modulo_add_11_qelse_and_6_nl <= (NOT z_out_87_32) AND (fsm_output(7));
  modulo_add_11_qelse_and_7_nl <= (NOT z_out_87_32) AND (fsm_output(9));
  modulo_add_12_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(z_out_70, z_out_82, z_out_80,
      STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & (fsm_output(7)) & (fsm_output(9))));
  acc_14_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_12_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_12_qelse_and_nl <= (NOT z_out_87_32) AND modulo_add_1_qelse_or_m1c;
  modulo_add_12_qelse_or_1_nl <= (z_out_87_32 AND modulo_add_1_qelse_or_m1c) OR (z_out_88_32
      AND (fsm_output(7))) OR (z_out_90_32 AND (fsm_output(9)));
  modulo_add_12_qelse_and_4_nl <= (NOT z_out_88_32) AND (fsm_output(7));
  modulo_add_12_qelse_and_5_nl <= (NOT z_out_90_32) AND (fsm_output(9));
  modulo_add_13_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(z_out_69, z_out_81, z_out_79,
      STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & (fsm_output(7)) & (fsm_output(9))));
  acc_18_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_13_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_13_qelse_and_nl <= (NOT z_out_90_32) AND modulo_add_1_qelse_or_m1c;
  modulo_add_13_qelse_or_1_nl <= (z_out_90_32 AND modulo_add_1_qelse_or_m1c) OR (z_out_90_32
      AND (fsm_output(7))) OR (z_out_91_32 AND (fsm_output(9)));
  modulo_add_13_qelse_and_4_nl <= (NOT z_out_90_32) AND (fsm_output(7));
  modulo_add_13_qelse_and_5_nl <= (NOT z_out_91_32) AND (fsm_output(9));
  modulo_add_14_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(z_out_68, z_out_80, z_out_78,
      STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & (fsm_output(7)) & (fsm_output(9))));
  acc_22_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_14_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_14_qelse_and_nl <= (NOT z_out_92_32) AND modulo_add_1_qelse_or_m1c;
  modulo_add_14_qelse_or_1_nl <= (z_out_92_32 AND modulo_add_1_qelse_or_m1c) OR (z_out_93_32
      AND (fsm_output(7))) OR (z_out_94_32 AND (fsm_output(9)));
  modulo_add_14_qelse_and_4_nl <= (NOT z_out_93_32) AND (fsm_output(7));
  modulo_add_14_qelse_and_5_nl <= (NOT z_out_94_32) AND (fsm_output(9));
  modulo_add_15_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_67, z_out_82, z_out_79,
      z_out_77, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7))
      & (fsm_output(9))));
  acc_26_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_15_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_15_qelse_and_nl <= (NOT z_out_93_32) AND (fsm_output(2));
  modulo_add_15_qelse_or_nl <= (z_out_93_32 AND (fsm_output(2))) OR (z_out_93_32
      AND (fsm_output(4))) OR (z_out_94_32 AND (fsm_output(7))) OR (z_out_97_32 AND
      (fsm_output(9)));
  modulo_add_15_qelse_and_5_nl <= (NOT z_out_93_32) AND (fsm_output(4));
  modulo_add_15_qelse_and_6_nl <= (NOT z_out_94_32) AND (fsm_output(7));
  modulo_add_15_qelse_and_7_nl <= (NOT z_out_97_32) AND (fsm_output(9));
  INNER_LOOP1_r_mux_45_nl <= MUX_s_1_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10, fsm_output(7));
  INNER_LOOP1_mux_nl <= MUX_s_1_2_2(INNER_LOOP1_stage_0, INNER_LOOP1_stage_0_11,
      or_dcpl_218);
  INNER_LOOP1_r_INNER_LOOP1_r_and_1_nl <= (z_out_2(0)) AND (fsm_output(4));
  INNER_LOOP1_r_INNER_LOOP1_r_and_3_nl <= (z_out_2(0)) AND (fsm_output(9));
  or_1465_nl <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("00"));
  INNER_LOOP1_r_mux1h_46_nl <= MUX1HOT_s_1_4_2(INNER_LOOP1_stage_0_9, INNER_LOOP1_r_INNER_LOOP1_r_and_1_nl,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9, INNER_LOOP1_r_INNER_LOOP1_r_and_3_nl,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & or_dcpl_233 & (fsm_output(7)) & or_1465_nl));
  INNER_LOOP1_r_INNER_LOOP1_r_and_2_nl <= (z_out_2(0)) AND (fsm_output(7));
  INNER_LOOP1_mux_11_nl <= MUX_s_1_2_2(INNER_LOOP1_stage_0_10, INNER_LOOP1_r_INNER_LOOP1_r_and_2_nl,
      or_tmp_1134);
  INNER_LOOP1_r_INNER_LOOP1_r_and_nl <= (z_out_2(0)) AND (fsm_output(2));
  modulo_add_2_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(z_out_80, z_out_77, z_out_75, STD_LOGIC_VECTOR'(
      modulo_add_1_qelse_or_m1c & (fsm_output(7)) & (fsm_output(9))));
  acc_29_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_2_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_23_qelse_and_nl <= (NOT z_out_96_32) AND modulo_add_1_qelse_or_m1c;
  modulo_add_23_qelse_or_1_nl <= (z_out_96_32 AND modulo_add_1_qelse_or_m1c) OR (z_out_96_32
      AND (fsm_output(7))) OR (z_out_98_32 AND (fsm_output(9)));
  modulo_add_23_qelse_and_4_nl <= (NOT z_out_96_32) AND (fsm_output(7));
  modulo_add_23_qelse_and_5_nl <= (NOT z_out_98_32) AND (fsm_output(9));
  modulo_add_3_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(z_out_79, z_out_76, z_out_74, STD_LOGIC_VECTOR'(
      modulo_add_1_qelse_or_m1c & (fsm_output(7)) & (fsm_output(9))));
  acc_32_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_3_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_24_qelse_and_nl <= (NOT z_out_98_32) AND modulo_add_1_qelse_or_m1c;
  modulo_add_24_qelse_or_1_nl <= (z_out_98_32 AND modulo_add_1_qelse_or_m1c) OR (z_out_97_32
      AND (fsm_output(7))) OR (z_out_96_32 AND (fsm_output(9)));
  modulo_add_24_qelse_and_4_nl <= (NOT z_out_97_32) AND (fsm_output(7));
  modulo_add_24_qelse_and_5_nl <= (NOT z_out_96_32) AND (fsm_output(9));
  modulo_add_4_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(z_out_78, z_out_75, z_out_73, STD_LOGIC_VECTOR'(
      modulo_add_1_qelse_or_m1c & (fsm_output(7)) & (fsm_output(9))));
  acc_34_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_4_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_25_qelse_and_nl <= (NOT z_out_97_32) AND modulo_add_1_qelse_or_m1c;
  modulo_add_25_qelse_or_1_nl <= (z_out_97_32 AND modulo_add_1_qelse_or_m1c) OR (z_out_95_32
      AND (fsm_output(7))) OR (z_out_92_32 AND (fsm_output(9)));
  modulo_add_25_qelse_and_4_nl <= (NOT z_out_95_32) AND (fsm_output(7));
  modulo_add_25_qelse_and_5_nl <= (NOT z_out_92_32) AND (fsm_output(9));
  modulo_add_5_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_77, z_out_76, z_out_74, z_out_72,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_37_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_5_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_26_qelse_and_nl <= (NOT z_out_91_32) AND (fsm_output(2));
  modulo_add_26_qelse_or_nl <= (z_out_91_32 AND (fsm_output(2))) OR (z_out_91_32
      AND (fsm_output(4))) OR (z_out_91_32 AND (fsm_output(7))) OR (z_out_88_32 AND
      (fsm_output(9)));
  modulo_add_26_qelse_and_5_nl <= (NOT z_out_91_32) AND (fsm_output(4));
  modulo_add_26_qelse_and_6_nl <= (NOT z_out_91_32) AND (fsm_output(7));
  modulo_add_26_qelse_and_7_nl <= (NOT z_out_88_32) AND (fsm_output(9));
  modulo_add_6_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_76, z_out_75, z_out_73, z_out_71,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_39_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_6_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_27_qelse_and_nl <= (NOT z_out_89_32) AND (fsm_output(2));
  modulo_add_27_qelse_or_nl <= (z_out_89_32 AND (fsm_output(2))) OR (z_out_89_32
      AND (fsm_output(4))) OR (z_out_85_32 AND (fsm_output(7))) OR (z_out_84_32 AND
      (fsm_output(9)));
  modulo_add_27_qelse_and_5_nl <= (NOT z_out_89_32) AND (fsm_output(4));
  modulo_add_27_qelse_and_6_nl <= (NOT z_out_85_32) AND (fsm_output(7));
  modulo_add_27_qelse_and_7_nl <= (NOT z_out_84_32) AND (fsm_output(9));
  modulo_add_7_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_75, z_out_74, z_out_72, z_out_70,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_42_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_7_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_28_qelse_and_nl <= (NOT z_out_85_32) AND (fsm_output(2));
  modulo_add_28_qelse_or_nl <= (z_out_85_32 AND (fsm_output(2))) OR (z_out_85_32
      AND (fsm_output(4))) OR (z_out_89_32 AND (fsm_output(7))) OR (z_out_93_32 AND
      (fsm_output(9)));
  modulo_add_28_qelse_and_5_nl <= (NOT z_out_85_32) AND (fsm_output(4));
  modulo_add_28_qelse_and_6_nl <= (NOT z_out_89_32) AND (fsm_output(7));
  modulo_add_28_qelse_and_7_nl <= (NOT z_out_93_32) AND (fsm_output(9));
  modulo_add_8_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_74, z_out_73, z_out_71, z_out_69,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_44_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_8_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_29_qelse_and_nl <= (NOT z_out_95_32) AND (fsm_output(2));
  modulo_add_29_qelse_or_nl <= (z_out_95_32 AND (fsm_output(2))) OR (z_out_95_32
      AND (fsm_output(4))) OR (z_out_98_32 AND (fsm_output(7))) OR (z_out_95_32 AND
      (fsm_output(9)));
  modulo_add_29_qelse_and_5_nl <= (NOT z_out_95_32) AND (fsm_output(4));
  modulo_add_29_qelse_and_6_nl <= (NOT z_out_98_32) AND (fsm_output(7));
  modulo_add_29_qelse_and_7_nl <= (NOT z_out_95_32) AND (fsm_output(9));
  modulo_add_9_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_73, z_out_72, z_out_70, z_out_68,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_47_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_9_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_30_qelse_and_nl <= (NOT z_out_94_32) AND (fsm_output(2));
  modulo_add_30_qelse_or_nl <= (z_out_94_32 AND (fsm_output(2))) OR (z_out_94_32
      AND (fsm_output(4))) OR (z_out_92_32 AND (fsm_output(7))) OR (z_out_89_32 AND
      (fsm_output(9)));
  modulo_add_30_qelse_and_5_nl <= (NOT z_out_94_32) AND (fsm_output(4));
  modulo_add_30_qelse_and_6_nl <= (NOT z_out_92_32) AND (fsm_output(7));
  modulo_add_30_qelse_and_7_nl <= (NOT z_out_89_32) AND (fsm_output(9));
  modulo_add_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(z_out_82, z_out_71, z_out_69, z_out_67,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_49_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  modulo_add_31_qelse_and_nl <= (NOT z_out_88_32) AND (fsm_output(2));
  modulo_add_31_qelse_or_nl <= (z_out_88_32 AND (fsm_output(2))) OR (z_out_88_32
      AND (fsm_output(4))) OR (z_out_86_32 AND (fsm_output(7))) OR (z_out_83_32 AND
      (fsm_output(9)));
  modulo_add_31_qelse_and_5_nl <= (NOT z_out_88_32) AND (fsm_output(4));
  modulo_add_31_qelse_and_6_nl <= (NOT z_out_86_32) AND (fsm_output(7));
  modulo_add_31_qelse_and_7_nl <= (NOT z_out_83_32) AND (fsm_output(9));
  modulo_sub_16_qelse_or_nl <= ((z_out_66(31)) AND (NOT (fsm_output(9)))) OR ((z_out_51(31))
      AND (fsm_output(9)));
  modulo_sub_17_qelse_or_nl <= ((z_out_56(31)) AND (NOT (fsm_output(9)))) OR ((z_out_52(31))
      AND (fsm_output(9)));
  modulo_sub_18_qelse_or_nl <= ((z_out_63(31)) AND (NOT (fsm_output(9)))) OR ((z_out_53(31))
      AND (fsm_output(9)));
  modulo_sub_19_qelse_or_nl <= ((z_out_64(31)) AND (NOT (fsm_output(9)))) OR ((z_out_54(31))
      AND (fsm_output(9)));
  modulo_sub_20_qelse_or_nl <= ((z_out_65(31)) AND (NOT (fsm_output(9)))) OR ((z_out_55(31))
      AND (fsm_output(9)));
  modulo_sub_21_qelse_or_nl <= ((z_out_51(31)) AND (NOT (fsm_output(9)))) OR ((z_out_56(31))
      AND (fsm_output(9)));
  modulo_sub_22_qelse_or_nl <= ((z_out_52(31)) AND (NOT (fsm_output(9)))) OR ((z_out_57(31))
      AND (fsm_output(9)));
  modulo_sub_23_qelse_or_nl <= ((z_out_53(31)) AND (NOT (fsm_output(9)))) OR ((z_out_58(31))
      AND (fsm_output(9)));
  modulo_sub_24_qelse_or_nl <= ((z_out_54(31)) AND (NOT (fsm_output(9)))) OR ((z_out_59(31))
      AND (fsm_output(9)));
  modulo_sub_25_qelse_or_nl <= ((z_out_55(31)) AND (NOT (fsm_output(9)))) OR ((z_out_60(31))
      AND (fsm_output(9)));
  modulo_sub_26_qelse_or_nl <= ((z_out_57(31)) AND (NOT (fsm_output(9)))) OR ((z_out_61(31))
      AND (fsm_output(9)));
  modulo_sub_27_qelse_or_nl <= ((z_out_58(31)) AND (NOT (fsm_output(9)))) OR ((z_out_62(31))
      AND (fsm_output(9)));
  modulo_sub_28_qelse_or_nl <= ((z_out_59(31)) AND (NOT (fsm_output(9)))) OR ((z_out_63(31))
      AND (fsm_output(9)));
  modulo_sub_29_qelse_or_nl <= ((z_out_60(31)) AND (NOT (fsm_output(9)))) OR ((z_out_64(31))
      AND (fsm_output(9)));
  modulo_sub_30_qelse_or_nl <= ((z_out_61(31)) AND (NOT (fsm_output(9)))) OR ((z_out_65(31))
      AND (fsm_output(9)));
  modulo_sub_31_qelse_or_nl <= ((z_out_62(31)) AND (NOT (fsm_output(9)))) OR ((z_out_66(31))
      AND (fsm_output(9)));
  STAGE_LOOP_base_STAGE_LOOP_base_mux_nl <= MUX_v_7_2_2((z_out(10 DOWNTO 4)), (z_out_2(6
      DOWNTO 0)), fsm_output(4));
  INNER_LOOP2_r_or_nl <= (fsm_output(4)) OR (fsm_output(1)) OR (fsm_output(2));
  operator_20_false_mux_2_nl <= MUX_v_3_2_2((butterFly2_11_tw_h_slc_operator_33_true_2_lshift_psp_2_0_1_0_itm
      & c_1_sva), operator_20_false_acc_cse_sva, fsm_output(5));
  z_out_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(operator_20_false_mux_2_nl)
      + UNSIGNED'( '1' & (NOT (fsm_output(5))) & '1'), 3));
  operator_20_false_mux1h_2_nl <= MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0, INNER_LOOP2_r_11_4_sva_6_0,
      INNER_LOOP3_r_11_4_sva_6_0, INNER_LOOP4_r_11_4_sva_6_0, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(operator_20_false_mux1h_2_nl),
      8) + UNSIGNED'( "00000001"), 8));
  modulo_sub_6_qif_mux_2_nl <= MUX_v_31_2_2((z_out_57(30 DOWNTO 0)), (z_out_55(30
      DOWNTO 0)), fsm_output(7));
  z_out_4 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_6_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_37_qif_mux_2_nl <= MUX_v_31_2_2((z_out_54(30 DOWNTO 0)), (z_out_58(30
      DOWNTO 0)), fsm_output(2));
  z_out_5 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_37_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_36_qif_mux_2_nl <= MUX_v_31_2_2((z_out_53(30 DOWNTO 0)), (z_out_59(30
      DOWNTO 0)), fsm_output(2));
  z_out_8 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_36_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_4_qif_mux_2_nl <= MUX_v_31_2_2((z_out_55(30 DOWNTO 0)), (z_out_57(30
      DOWNTO 0)), fsm_output(7));
  z_out_9 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_4_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_35_qif_mux_2_nl <= MUX_v_31_2_2((z_out_52(30 DOWNTO 0)), (z_out_60(30
      DOWNTO 0)), fsm_output(2));
  z_out_10 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_35_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_3_qif_mux_2_nl <= MUX_v_31_2_2((z_out_54(30 DOWNTO 0)), (z_out_58(30
      DOWNTO 0)), fsm_output(7));
  z_out_12 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_3_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_34_qif_mux_2_nl <= MUX_v_31_2_2((z_out_51(30 DOWNTO 0)), (z_out_61(30
      DOWNTO 0)), fsm_output(2));
  z_out_13 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_34_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_2_qif_mux_2_nl <= MUX_v_31_2_2((z_out_53(30 DOWNTO 0)), (z_out_59(30
      DOWNTO 0)), fsm_output(7));
  z_out_14 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_2_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_33_qif_mux_2_nl <= MUX_v_31_2_2((z_out_66(30 DOWNTO 0)), (z_out_62(30
      DOWNTO 0)), fsm_output(2));
  z_out_16 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_33_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_1_qif_mux_2_nl <= MUX_v_31_2_2((z_out_52(30 DOWNTO 0)), (z_out_60(30
      DOWNTO 0)), fsm_output(7));
  z_out_17 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_1_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_32_qif_mux_2_nl <= MUX_v_31_2_2((z_out_65(30 DOWNTO 0)), (z_out_63(30
      DOWNTO 0)), fsm_output(2));
  z_out_18 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_32_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_qif_mux_2_nl <= MUX_v_31_2_2((z_out_51(30 DOWNTO 0)), (z_out_61(30 DOWNTO
      0)), fsm_output(7));
  z_out_20 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_31_qif_mux_2_nl <= MUX_v_31_2_2((z_out_62(30 DOWNTO 0)), (z_out_66(30
      DOWNTO 0)), fsm_output(9));
  z_out_21 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_31_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_13_qif_mux_2_nl <= MUX_v_31_2_2((z_out_64(30 DOWNTO 0)), (z_out_63(30
      DOWNTO 0)), fsm_output(7));
  z_out_22 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_13_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_30_qif_mux_2_nl <= MUX_v_31_2_2((z_out_61(30 DOWNTO 0)), (z_out_65(30
      DOWNTO 0)), fsm_output(9));
  z_out_24 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_30_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_45_qif_mux_2_nl <= MUX_v_31_2_2((z_out_62(30 DOWNTO 0)), (z_out_65(30
      DOWNTO 0)), fsm_output(2));
  z_out_25 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_45_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_29_qif_mux_2_nl <= MUX_v_31_2_2((z_out_60(30 DOWNTO 0)), (z_out_64(30
      DOWNTO 0)), fsm_output(9));
  z_out_26 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_29_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_15_qif_mux_2_nl <= MUX_v_31_2_2((z_out_66(30 DOWNTO 0)), (z_out_64(30
      DOWNTO 0)), fsm_output(7));
  z_out_28 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_15_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_28_qif_mux_2_nl <= MUX_v_31_2_2((z_out_59(30 DOWNTO 0)), (z_out_63(30
      DOWNTO 0)), fsm_output(9));
  z_out_29 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_28_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_27_qif_mux_2_nl <= MUX_v_31_2_2((z_out_58(30 DOWNTO 0)), (z_out_62(30
      DOWNTO 0)), fsm_output(9));
  z_out_31 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_27_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_26_qif_mux_2_nl <= MUX_v_31_2_2((z_out_57(30 DOWNTO 0)), (z_out_61(30
      DOWNTO 0)), fsm_output(9));
  z_out_32 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_26_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_25_qif_mux_2_nl <= MUX_v_31_2_2((z_out_55(30 DOWNTO 0)), (z_out_60(30
      DOWNTO 0)), fsm_output(9));
  z_out_34 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_25_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_24_qif_mux_2_nl <= MUX_v_31_2_2((z_out_54(30 DOWNTO 0)), (z_out_59(30
      DOWNTO 0)), fsm_output(9));
  z_out_36 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_24_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_23_qif_mux_2_nl <= MUX_v_31_2_2((z_out_53(30 DOWNTO 0)), (z_out_58(30
      DOWNTO 0)), fsm_output(9));
  z_out_37 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_23_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_22_qif_mux_2_nl <= MUX_v_31_2_2((z_out_52(30 DOWNTO 0)), (z_out_57(30
      DOWNTO 0)), fsm_output(9));
  z_out_39 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_22_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_21_qif_mux_2_nl <= MUX_v_31_2_2((z_out_51(30 DOWNTO 0)), (z_out_56(30
      DOWNTO 0)), fsm_output(9));
  z_out_41 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_21_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_20_qif_mux_2_nl <= MUX_v_31_2_2((z_out_65(30 DOWNTO 0)), (z_out_55(30
      DOWNTO 0)), fsm_output(9));
  z_out_42 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_20_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_19_qif_mux_2_nl <= MUX_v_31_2_2((z_out_64(30 DOWNTO 0)), (z_out_54(30
      DOWNTO 0)), fsm_output(9));
  z_out_44 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_19_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_18_qif_mux_2_nl <= MUX_v_31_2_2((z_out_63(30 DOWNTO 0)), (z_out_53(30
      DOWNTO 0)), fsm_output(9));
  z_out_46 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_18_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_17_qif_mux_2_nl <= MUX_v_31_2_2((z_out_56(30 DOWNTO 0)), (z_out_52(30
      DOWNTO 0)), fsm_output(9));
  z_out_47 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_17_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_16_qif_mux_2_nl <= MUX_v_31_2_2((z_out_66(30 DOWNTO 0)), (z_out_51(30
      DOWNTO 0)), fsm_output(9));
  z_out_49 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_16_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  butterFly1_mux1h_17_nl <= MUX1HOT_v_32_4_2((NOT mult_res_lpi_3_dfm_1), (NOT reg_mult_21_res_lpi_3_dfm_1_cse),
      (NOT reg_mult_24_res_lpi_3_dfm_1_cse), (NOT reg_mult_17_res_lpi_3_dfm_1_cse),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  acc_50_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_10_sva_7 & '1') + UNSIGNED(butterFly1_mux1h_17_nl
      & '1'), 33));
  z_out_51 <= acc_50_nl(32 DOWNTO 1);
  butterFly1_1_mux1h_13_nl <= MUX1HOT_v_32_4_2((NOT mult_1_res_lpi_3_dfm_1), (NOT
      reg_mult_22_res_lpi_3_dfm_1_cse), (NOT reg_mult_29_res_lpi_3_dfm_1_cse), (NOT
      reg_mult_25_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  acc_51_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_102_sva_7 & '1') + UNSIGNED(butterFly1_1_mux1h_13_nl
      & '1'), 33));
  z_out_52 <= acc_51_nl(32 DOWNTO 1);
  butterFly1_2_mux1h_13_nl <= MUX1HOT_v_32_4_2((NOT mult_2_res_lpi_3_dfm_1), (NOT
      reg_mult_23_res_lpi_3_dfm_1_cse), (NOT reg_mult_31_res_lpi_3_dfm_1_cse), (NOT
      reg_mult_28_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  acc_52_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_104_sva_7 & '1') + UNSIGNED(butterFly1_2_mux1h_13_nl
      & '1'), 33));
  z_out_53 <= acc_52_nl(32 DOWNTO 1);
  butterFly1_3_mux1h_13_nl <= MUX1HOT_v_32_4_2((NOT mult_3_res_lpi_3_dfm_1), (NOT
      reg_mult_24_res_lpi_3_dfm_1_cse), (NOT reg_mult_27_res_lpi_3_dfm_1_cse), (NOT
      reg_mult_20_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  acc_53_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_106_sva_7 & '1') + UNSIGNED(butterFly1_3_mux1h_13_nl
      & '1'), 33));
  z_out_54 <= acc_53_nl(32 DOWNTO 1);
  butterFly1_4_mux1h_13_nl <= MUX1HOT_v_32_4_2((NOT mult_4_res_lpi_3_dfm_1), (NOT
      reg_mult_25_res_lpi_3_dfm_1_cse), (NOT reg_mult_23_res_lpi_3_dfm_1_cse), (NOT
      reg_mult_22_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  acc_54_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_108_sva_7 & '1') + UNSIGNED(butterFly1_4_mux1h_13_nl
      & '1'), 33));
  z_out_55 <= acc_54_nl(32 DOWNTO 1);
  butterFly1_5_mux1h_13_nl <= MUX1HOT_v_32_4_2((NOT mult_5_res_lpi_3_dfm_1), (NOT
      reg_mult_17_res_lpi_3_dfm_1_cse), (NOT reg_mult_19_res_lpi_3_dfm_1_cse), (NOT
      reg_mult_30_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  acc_55_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_110_sva_7 & '1') + UNSIGNED(butterFly1_5_mux1h_13_nl
      & '1'), 33));
  z_out_56 <= acc_55_nl(32 DOWNTO 1);
  butterFly1_6_mux1h_13_nl <= MUX1HOT_v_32_3_2((NOT mult_6_res_lpi_3_dfm_1), (NOT
      reg_mult_26_res_lpi_3_dfm_1_cse), (NOT reg_mult_18_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & or_dcpl_194 & (fsm_output(7))));
  acc_56_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_112_sva_7 & '1') + UNSIGNED(butterFly1_6_mux1h_13_nl
      & '1'), 33));
  z_out_57 <= acc_56_nl(32 DOWNTO 1);
  butterFly1_7_mux1h_13_nl <= MUX1HOT_v_32_4_2((NOT mult_7_res_lpi_3_dfm_1), (NOT
      reg_mult_27_res_lpi_3_dfm_1_cse), (NOT reg_mult_26_res_lpi_3_dfm_1_cse), (NOT
      reg_mult_18_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  acc_57_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_114_sva_7 & '1') + UNSIGNED(butterFly1_7_mux1h_13_nl
      & '1'), 33));
  z_out_58 <= acc_57_nl(32 DOWNTO 1);
  butterFly1_8_mux1h_13_nl <= MUX1HOT_v_32_4_2((NOT mult_8_res_lpi_3_dfm_1), (NOT
      reg_mult_28_res_lpi_3_dfm_1_cse), (NOT reg_mult_30_res_lpi_3_dfm_1_cse), (NOT
      reg_mult_19_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  acc_58_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_116_sva_7 & '1') + UNSIGNED(butterFly1_8_mux1h_13_nl
      & '1'), 33));
  z_out_59 <= acc_58_nl(32 DOWNTO 1);
  butterFly1_9_mux1h_13_nl <= MUX1HOT_v_32_4_2((NOT mult_9_res_lpi_3_dfm_1), (NOT
      reg_mult_29_res_lpi_3_dfm_1_cse), (NOT reg_mult_22_res_lpi_3_dfm_1_cse), (NOT
      reg_mult_23_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  acc_59_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_118_sva_7 & '1') + UNSIGNED(butterFly1_9_mux1h_13_nl
      & '1'), 33));
  z_out_60 <= acc_59_nl(32 DOWNTO 1);
  butterFly1_10_mux1h_13_nl <= MUX1HOT_v_32_4_2((NOT mult_10_res_lpi_3_dfm_1), (NOT
      reg_mult_30_res_lpi_3_dfm_1_cse), (NOT reg_mult_20_res_lpi_3_dfm_1_cse), (NOT
      reg_mult_27_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  acc_60_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_120_sva_7 & '1') + UNSIGNED(butterFly1_10_mux1h_13_nl
      & '1'), 33));
  z_out_61 <= acc_60_nl(32 DOWNTO 1);
  butterFly1_11_mux1h_13_nl <= MUX1HOT_v_32_3_2((NOT mult_11_res_lpi_3_dfm_1), (NOT
      reg_mult_31_res_lpi_3_dfm_1_cse), (NOT reg_mult_28_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & or_dcpl_194 & (fsm_output(7))));
  acc_61_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_122_sva_7 & '1') + UNSIGNED(butterFly1_11_mux1h_13_nl
      & '1'), 33));
  z_out_62 <= acc_61_nl(32 DOWNTO 1);
  butterFly1_12_mux1h_13_nl <= MUX1HOT_v_32_4_2((NOT mult_12_res_lpi_3_dfm_1), (NOT
      reg_mult_18_res_lpi_3_dfm_1_cse), (NOT reg_mult_25_res_lpi_3_dfm_1_cse), (NOT
      reg_mult_29_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  acc_62_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_124_sva_7 & '1') + UNSIGNED(butterFly1_12_mux1h_13_nl
      & '1'), 33));
  z_out_63 <= acc_62_nl(32 DOWNTO 1);
  butterFly1_13_mux1h_13_nl <= MUX1HOT_v_32_4_2((NOT mult_13_res_lpi_3_dfm_1), (NOT
      reg_mult_19_res_lpi_3_dfm_1_cse), (NOT reg_mult_17_res_lpi_3_dfm_1_cse), (NOT
      reg_mult_24_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  acc_63_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_126_sva_7 & '1') + UNSIGNED(butterFly1_13_mux1h_13_nl
      & '1'), 33));
  z_out_64 <= acc_63_nl(32 DOWNTO 1);
  butterFly1_14_mux1h_13_nl <= MUX1HOT_v_32_4_2((NOT mult_14_res_lpi_3_dfm_1), (NOT
      reg_mult_20_res_lpi_3_dfm_1_cse), (NOT reg_mult_16_res_lpi_3_dfm_1_cse), (NOT
      reg_mult_21_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  acc_64_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_60_sva_7 & '1') + UNSIGNED(butterFly1_14_mux1h_13_nl
      & '1'), 33));
  z_out_65 <= acc_64_nl(32 DOWNTO 1);
  butterFly1_15_mux1h_13_nl <= MUX1HOT_v_32_3_2((NOT mult_15_res_lpi_3_dfm_1), (NOT
      reg_mult_16_res_lpi_3_dfm_1_cse), (NOT reg_mult_21_res_lpi_3_dfm_1_cse), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & or_dcpl_194 & (fsm_output(7))));
  acc_65_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_62_sva_7 & '1') + UNSIGNED(butterFly1_15_mux1h_13_nl
      & '1'), 33));
  z_out_66 <= acc_65_nl(32 DOWNTO 1);
  butterFly1_15_mux1h_14_nl <= MUX1HOT_v_32_3_2(mult_15_res_lpi_3_dfm_1, reg_mult_16_res_lpi_3_dfm_1_cse,
      reg_mult_21_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'( (fsm_output(2)) & or_dcpl_194
      & (fsm_output(7))));
  z_out_67 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_62_sva_7) + UNSIGNED(butterFly1_15_mux1h_14_nl),
      32));
  butterFly1_14_mux1h_14_nl <= MUX1HOT_v_32_4_2(mult_14_res_lpi_3_dfm_1, reg_mult_20_res_lpi_3_dfm_1_cse,
      reg_mult_16_res_lpi_3_dfm_1_cse, reg_mult_21_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_68 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_60_sva_7) + UNSIGNED(butterFly1_14_mux1h_14_nl),
      32));
  butterFly1_13_mux1h_14_nl <= MUX1HOT_v_32_4_2(mult_13_res_lpi_3_dfm_1, reg_mult_19_res_lpi_3_dfm_1_cse,
      reg_mult_17_res_lpi_3_dfm_1_cse, reg_mult_24_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_69 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_126_sva_7) + UNSIGNED(butterFly1_13_mux1h_14_nl),
      32));
  butterFly1_12_mux1h_14_nl <= MUX1HOT_v_32_4_2(mult_12_res_lpi_3_dfm_1, reg_mult_18_res_lpi_3_dfm_1_cse,
      reg_mult_25_res_lpi_3_dfm_1_cse, reg_mult_29_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_70 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_124_sva_7) + UNSIGNED(butterFly1_12_mux1h_14_nl),
      32));
  butterFly1_11_mux1h_14_nl <= MUX1HOT_v_32_3_2(mult_11_res_lpi_3_dfm_1, reg_mult_31_res_lpi_3_dfm_1_cse,
      reg_mult_28_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'( (fsm_output(2)) & or_dcpl_194
      & (fsm_output(7))));
  z_out_71 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_122_sva_7) + UNSIGNED(butterFly1_11_mux1h_14_nl),
      32));
  butterFly1_10_mux1h_14_nl <= MUX1HOT_v_32_4_2(mult_10_res_lpi_3_dfm_1, reg_mult_30_res_lpi_3_dfm_1_cse,
      reg_mult_20_res_lpi_3_dfm_1_cse, reg_mult_27_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_72 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_120_sva_7) + UNSIGNED(butterFly1_10_mux1h_14_nl),
      32));
  butterFly1_9_mux1h_14_nl <= MUX1HOT_v_32_4_2(mult_9_res_lpi_3_dfm_1, reg_mult_29_res_lpi_3_dfm_1_cse,
      reg_mult_22_res_lpi_3_dfm_1_cse, reg_mult_23_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_73 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_118_sva_7) + UNSIGNED(butterFly1_9_mux1h_14_nl),
      32));
  butterFly1_8_mux1h_14_nl <= MUX1HOT_v_32_4_2(mult_8_res_lpi_3_dfm_1, reg_mult_28_res_lpi_3_dfm_1_cse,
      reg_mult_30_res_lpi_3_dfm_1_cse, reg_mult_19_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_74 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_116_sva_7) + UNSIGNED(butterFly1_8_mux1h_14_nl),
      32));
  butterFly1_7_mux1h_14_nl <= MUX1HOT_v_32_4_2(mult_7_res_lpi_3_dfm_1, reg_mult_27_res_lpi_3_dfm_1_cse,
      reg_mult_26_res_lpi_3_dfm_1_cse, reg_mult_18_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_75 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_114_sva_7) + UNSIGNED(butterFly1_7_mux1h_14_nl),
      32));
  butterFly1_6_mux1h_14_nl <= MUX1HOT_v_32_3_2(mult_6_res_lpi_3_dfm_1, reg_mult_26_res_lpi_3_dfm_1_cse,
      reg_mult_18_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'( (fsm_output(2)) & or_dcpl_194
      & (fsm_output(7))));
  z_out_76 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_112_sva_7) + UNSIGNED(butterFly1_6_mux1h_14_nl),
      32));
  butterFly1_5_mux1h_14_nl <= MUX1HOT_v_32_4_2(mult_5_res_lpi_3_dfm_1, reg_mult_17_res_lpi_3_dfm_1_cse,
      reg_mult_19_res_lpi_3_dfm_1_cse, reg_mult_30_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_77 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_110_sva_7) + UNSIGNED(butterFly1_5_mux1h_14_nl),
      32));
  butterFly1_4_mux1h_14_nl <= MUX1HOT_v_32_4_2(mult_4_res_lpi_3_dfm_1, reg_mult_25_res_lpi_3_dfm_1_cse,
      reg_mult_23_res_lpi_3_dfm_1_cse, reg_mult_22_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_78 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_108_sva_7) + UNSIGNED(butterFly1_4_mux1h_14_nl),
      32));
  butterFly1_3_mux1h_14_nl <= MUX1HOT_v_32_4_2(mult_3_res_lpi_3_dfm_1, reg_mult_24_res_lpi_3_dfm_1_cse,
      reg_mult_27_res_lpi_3_dfm_1_cse, reg_mult_20_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_79 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_106_sva_7) + UNSIGNED(butterFly1_3_mux1h_14_nl),
      32));
  butterFly1_2_mux1h_14_nl <= MUX1HOT_v_32_4_2(mult_2_res_lpi_3_dfm_1, reg_mult_23_res_lpi_3_dfm_1_cse,
      reg_mult_31_res_lpi_3_dfm_1_cse, reg_mult_28_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_80 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_104_sva_7) + UNSIGNED(butterFly1_2_mux1h_14_nl),
      32));
  butterFly1_1_mux1h_14_nl <= MUX1HOT_v_32_4_2(mult_1_res_lpi_3_dfm_1, reg_mult_22_res_lpi_3_dfm_1_cse,
      reg_mult_29_res_lpi_3_dfm_1_cse, reg_mult_25_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_81 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_102_sva_7) + UNSIGNED(butterFly1_1_mux1h_14_nl),
      32));
  butterFly1_mux1h_18_nl <= MUX1HOT_v_32_4_2(mult_res_lpi_3_dfm_1, reg_mult_21_res_lpi_3_dfm_1_cse,
      reg_mult_24_res_lpi_3_dfm_1_cse, reg_mult_17_res_lpi_3_dfm_1_cse, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(9))));
  z_out_82 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_10_sva_7) + UNSIGNED(butterFly1_mux1h_18_nl),
      32));
  modulo_add_1_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT z_out_81), (NOT z_out_78), (NOT
      z_out_67), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & (fsm_output(7)) &
      (fsm_output(9))));
  acc_82_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_1_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_83_32 <= acc_82_nl(33);
  modulo_add_10_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT z_out_72), (NOT z_out_67), (NOT
      z_out_68), (NOT z_out_71), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  acc_83_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_10_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_84_32 <= acc_83_nl(33);
  modulo_add_54_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT z_out_76), (NOT z_out_73), (NOT
      z_out_75), (NOT z_out_74), STD_LOGIC_VECTOR'( (fsm_output(9)) & (fsm_output(7))
      & (fsm_output(2)) & (fsm_output(4))));
  acc_84_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_54_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_85_32 <= acc_84_nl(33);
  modulo_add_48_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT z_out_82), (NOT z_out_71), (NOT
      z_out_77), (NOT z_out_69), STD_LOGIC_VECTOR'( (fsm_output(9)) & (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(7))));
  acc_85_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_48_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_86_32 <= acc_85_nl(33);
  modulo_add_33_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT z_out_67), (NOT z_out_81), (NOT
      z_out_70), STD_LOGIC_VECTOR'( (fsm_output(7)) & (fsm_output(9)) & modulo_add_1_qelse_or_m1c));
  acc_86_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_33_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_87_32 <= acc_86_nl(33);
  modulo_add_34_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT z_out_82), (NOT z_out_72), (NOT
      z_out_71), STD_LOGIC_VECTOR'( or_dcpl_210 & (fsm_output(9)) & (fsm_output(4))));
  acc_87_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_34_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_88_32 <= acc_87_nl(33);
  modulo_add_6_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT z_out_76), (NOT z_out_75), (NOT
      z_out_72), (NOT z_out_68), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4))
      & (fsm_output(7)) & (fsm_output(9))));
  acc_88_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_6_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_89_32 <= acc_88_nl(33);
  modulo_add_50_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT z_out_80), (NOT z_out_69), (NOT
      z_out_81), STD_LOGIC_VECTOR'( (fsm_output(9)) & modulo_add_1_qelse_or_m1c &
      (fsm_output(7))));
  acc_89_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_50_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_90_32 <= acc_89_nl(33);
  modulo_add_51_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT z_out_79), (NOT z_out_77), (NOT
      z_out_76), (NOT z_out_74), STD_LOGIC_VECTOR'( (fsm_output(9)) & (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(7))));
  acc_90_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_51_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_91_32 <= acc_90_nl(33);
  modulo_add_14_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT z_out_68), (NOT z_out_73), (NOT
      z_out_70), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & (fsm_output(9)) &
      (fsm_output(7))));
  acc_91_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_14_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_92_32 <= acc_91_nl(33);
  modulo_add_36_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT z_out_80), (NOT z_out_67), (NOT
      z_out_82), (NOT z_out_70), STD_LOGIC_VECTOR'( (fsm_output(7)) & (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(9))));
  acc_92_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_36_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_93_32 <= acc_92_nl(33);
  modulo_add_52_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT z_out_78), (NOT z_out_79), (NOT
      z_out_73), (NOT z_out_72), STD_LOGIC_VECTOR'( (fsm_output(9)) & (fsm_output(7))
      & (fsm_output(2)) & (fsm_output(4))));
  acc_93_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_52_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_94_32 <= acc_93_nl(33);
  modulo_add_41_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT z_out_75), (NOT z_out_74), (NOT
      z_out_73), (NOT z_out_69), STD_LOGIC_VECTOR'( (fsm_output(7)) & (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(9))));
  acc_94_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_41_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_95_32 <= acc_94_nl(33);
  modulo_add_2_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT z_out_80), (NOT z_out_77), (NOT
      z_out_74), STD_LOGIC_VECTOR'( modulo_add_1_qelse_or_m1c & (fsm_output(7)) &
      (fsm_output(9))));
  acc_95_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_2_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_96_32 <= acc_95_nl(33);
  modulo_add_53_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT z_out_77), (NOT z_out_76), (NOT
      z_out_78), STD_LOGIC_VECTOR'( (fsm_output(9)) & (fsm_output(7)) & modulo_add_1_qelse_or_m1c));
  acc_96_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_53_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_97_32 <= acc_96_nl(33);
  modulo_add_55_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT z_out_75), (NOT z_out_79), (NOT
      z_out_71), STD_LOGIC_VECTOR'( (fsm_output(9)) & modulo_add_1_qelse_or_m1c &
      (fsm_output(7))));
  acc_97_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_55_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_98_32 <= acc_97_nl(33);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY peaseNTT IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_0_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_0_wea : OUT STD_LOGIC;
    xt_rsc_0_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_0_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_0_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_0_web : OUT STD_LOGIC;
    xt_rsc_0_0_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    xt_rsc_0_1_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_1_wea : OUT STD_LOGIC;
    xt_rsc_0_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_1_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_1_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_1_web : OUT STD_LOGIC;
    xt_rsc_0_1_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    xt_rsc_0_2_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_2_wea : OUT STD_LOGIC;
    xt_rsc_0_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_2_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_2_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_2_web : OUT STD_LOGIC;
    xt_rsc_0_2_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    xt_rsc_0_3_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_3_wea : OUT STD_LOGIC;
    xt_rsc_0_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_3_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_3_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_3_web : OUT STD_LOGIC;
    xt_rsc_0_3_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    xt_rsc_0_4_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_4_wea : OUT STD_LOGIC;
    xt_rsc_0_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_4_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_4_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_4_web : OUT STD_LOGIC;
    xt_rsc_0_4_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    xt_rsc_0_5_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_5_wea : OUT STD_LOGIC;
    xt_rsc_0_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_5_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_5_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_5_web : OUT STD_LOGIC;
    xt_rsc_0_5_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    xt_rsc_0_6_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_6_wea : OUT STD_LOGIC;
    xt_rsc_0_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_6_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_6_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_6_web : OUT STD_LOGIC;
    xt_rsc_0_6_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    xt_rsc_0_7_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_7_wea : OUT STD_LOGIC;
    xt_rsc_0_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_7_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_7_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_7_web : OUT STD_LOGIC;
    xt_rsc_0_7_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    xt_rsc_0_8_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_8_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_8_wea : OUT STD_LOGIC;
    xt_rsc_0_8_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_8_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_8_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_8_web : OUT STD_LOGIC;
    xt_rsc_0_8_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    xt_rsc_0_9_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_9_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_9_wea : OUT STD_LOGIC;
    xt_rsc_0_9_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_9_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_9_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_9_web : OUT STD_LOGIC;
    xt_rsc_0_9_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    xt_rsc_0_10_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_10_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_10_wea : OUT STD_LOGIC;
    xt_rsc_0_10_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_10_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_10_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_10_web : OUT STD_LOGIC;
    xt_rsc_0_10_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    xt_rsc_0_11_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_11_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_11_wea : OUT STD_LOGIC;
    xt_rsc_0_11_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_11_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_11_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_11_web : OUT STD_LOGIC;
    xt_rsc_0_11_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    xt_rsc_0_12_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_12_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_12_wea : OUT STD_LOGIC;
    xt_rsc_0_12_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_12_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_12_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_12_web : OUT STD_LOGIC;
    xt_rsc_0_12_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    xt_rsc_0_13_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_13_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_13_wea : OUT STD_LOGIC;
    xt_rsc_0_13_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_13_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_13_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_13_web : OUT STD_LOGIC;
    xt_rsc_0_13_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    xt_rsc_0_14_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_14_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_14_wea : OUT STD_LOGIC;
    xt_rsc_0_14_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_14_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_14_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_14_web : OUT STD_LOGIC;
    xt_rsc_0_14_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    xt_rsc_0_15_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_15_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_15_wea : OUT STD_LOGIC;
    xt_rsc_0_15_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_15_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_15_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_15_web : OUT STD_LOGIC;
    xt_rsc_0_15_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    xt_rsc_0_16_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_16_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_16_wea : OUT STD_LOGIC;
    xt_rsc_0_16_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_16_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_16_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_16_web : OUT STD_LOGIC;
    xt_rsc_0_16_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_16_lz : OUT STD_LOGIC;
    xt_rsc_0_17_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_17_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_17_wea : OUT STD_LOGIC;
    xt_rsc_0_17_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_17_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_17_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_17_web : OUT STD_LOGIC;
    xt_rsc_0_17_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_17_lz : OUT STD_LOGIC;
    xt_rsc_0_18_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_18_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_18_wea : OUT STD_LOGIC;
    xt_rsc_0_18_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_18_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_18_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_18_web : OUT STD_LOGIC;
    xt_rsc_0_18_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_18_lz : OUT STD_LOGIC;
    xt_rsc_0_19_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_19_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_19_wea : OUT STD_LOGIC;
    xt_rsc_0_19_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_19_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_19_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_19_web : OUT STD_LOGIC;
    xt_rsc_0_19_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_19_lz : OUT STD_LOGIC;
    xt_rsc_0_20_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_20_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_20_wea : OUT STD_LOGIC;
    xt_rsc_0_20_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_20_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_20_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_20_web : OUT STD_LOGIC;
    xt_rsc_0_20_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_20_lz : OUT STD_LOGIC;
    xt_rsc_0_21_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_21_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_21_wea : OUT STD_LOGIC;
    xt_rsc_0_21_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_21_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_21_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_21_web : OUT STD_LOGIC;
    xt_rsc_0_21_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_21_lz : OUT STD_LOGIC;
    xt_rsc_0_22_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_22_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_22_wea : OUT STD_LOGIC;
    xt_rsc_0_22_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_22_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_22_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_22_web : OUT STD_LOGIC;
    xt_rsc_0_22_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_22_lz : OUT STD_LOGIC;
    xt_rsc_0_23_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_23_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_23_wea : OUT STD_LOGIC;
    xt_rsc_0_23_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_23_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_23_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_23_web : OUT STD_LOGIC;
    xt_rsc_0_23_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_23_lz : OUT STD_LOGIC;
    xt_rsc_0_24_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_24_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_24_wea : OUT STD_LOGIC;
    xt_rsc_0_24_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_24_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_24_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_24_web : OUT STD_LOGIC;
    xt_rsc_0_24_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_24_lz : OUT STD_LOGIC;
    xt_rsc_0_25_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_25_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_25_wea : OUT STD_LOGIC;
    xt_rsc_0_25_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_25_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_25_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_25_web : OUT STD_LOGIC;
    xt_rsc_0_25_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_25_lz : OUT STD_LOGIC;
    xt_rsc_0_26_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_26_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_26_wea : OUT STD_LOGIC;
    xt_rsc_0_26_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_26_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_26_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_26_web : OUT STD_LOGIC;
    xt_rsc_0_26_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_26_lz : OUT STD_LOGIC;
    xt_rsc_0_27_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_27_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_27_wea : OUT STD_LOGIC;
    xt_rsc_0_27_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_27_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_27_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_27_web : OUT STD_LOGIC;
    xt_rsc_0_27_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_27_lz : OUT STD_LOGIC;
    xt_rsc_0_28_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_28_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_28_wea : OUT STD_LOGIC;
    xt_rsc_0_28_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_28_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_28_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_28_web : OUT STD_LOGIC;
    xt_rsc_0_28_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_28_lz : OUT STD_LOGIC;
    xt_rsc_0_29_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_29_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_29_wea : OUT STD_LOGIC;
    xt_rsc_0_29_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_29_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_29_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_29_web : OUT STD_LOGIC;
    xt_rsc_0_29_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_29_lz : OUT STD_LOGIC;
    xt_rsc_0_30_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_30_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_30_wea : OUT STD_LOGIC;
    xt_rsc_0_30_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_30_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_30_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_30_web : OUT STD_LOGIC;
    xt_rsc_0_30_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_30_lz : OUT STD_LOGIC;
    xt_rsc_0_31_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_31_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_31_wea : OUT STD_LOGIC;
    xt_rsc_0_31_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_31_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    xt_rsc_0_31_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_31_web : OUT STD_LOGIC;
    xt_rsc_0_31_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_31_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsc_0_0_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_wea : OUT STD_LOGIC;
    twiddle_rsc_0_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_0_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_web : OUT STD_LOGIC;
    twiddle_rsc_0_0_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_rsc_0_1_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_wea : OUT STD_LOGIC;
    twiddle_rsc_0_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_1_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_web : OUT STD_LOGIC;
    twiddle_rsc_0_1_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_rsc_0_2_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_wea : OUT STD_LOGIC;
    twiddle_rsc_0_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_2_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_web : OUT STD_LOGIC;
    twiddle_rsc_0_2_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_rsc_0_3_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_wea : OUT STD_LOGIC;
    twiddle_rsc_0_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_3_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_web : OUT STD_LOGIC;
    twiddle_rsc_0_3_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_rsc_0_4_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_wea : OUT STD_LOGIC;
    twiddle_rsc_0_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_4_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_web : OUT STD_LOGIC;
    twiddle_rsc_0_4_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_rsc_0_5_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_wea : OUT STD_LOGIC;
    twiddle_rsc_0_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_5_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_web : OUT STD_LOGIC;
    twiddle_rsc_0_5_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_rsc_0_6_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_wea : OUT STD_LOGIC;
    twiddle_rsc_0_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_6_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_web : OUT STD_LOGIC;
    twiddle_rsc_0_6_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_rsc_0_7_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_wea : OUT STD_LOGIC;
    twiddle_rsc_0_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_7_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_web : OUT STD_LOGIC;
    twiddle_rsc_0_7_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_rsc_0_8_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_8_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_8_wea : OUT STD_LOGIC;
    twiddle_rsc_0_8_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_8_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_8_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_8_web : OUT STD_LOGIC;
    twiddle_rsc_0_8_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_rsc_0_9_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_9_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_9_wea : OUT STD_LOGIC;
    twiddle_rsc_0_9_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_9_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_9_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_9_web : OUT STD_LOGIC;
    twiddle_rsc_0_9_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_rsc_0_10_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_10_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_10_wea : OUT STD_LOGIC;
    twiddle_rsc_0_10_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_10_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_10_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_10_web : OUT STD_LOGIC;
    twiddle_rsc_0_10_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_rsc_0_11_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_11_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_11_wea : OUT STD_LOGIC;
    twiddle_rsc_0_11_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_11_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_11_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_11_web : OUT STD_LOGIC;
    twiddle_rsc_0_11_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_rsc_0_12_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_12_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_12_wea : OUT STD_LOGIC;
    twiddle_rsc_0_12_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_12_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_12_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_12_web : OUT STD_LOGIC;
    twiddle_rsc_0_12_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_rsc_0_13_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_13_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_13_wea : OUT STD_LOGIC;
    twiddle_rsc_0_13_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_13_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_13_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_13_web : OUT STD_LOGIC;
    twiddle_rsc_0_13_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_rsc_0_14_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_14_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_14_wea : OUT STD_LOGIC;
    twiddle_rsc_0_14_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_14_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_14_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_14_web : OUT STD_LOGIC;
    twiddle_rsc_0_14_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_rsc_0_15_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_15_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_15_wea : OUT STD_LOGIC;
    twiddle_rsc_0_15_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_15_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_15_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_15_web : OUT STD_LOGIC;
    twiddle_rsc_0_15_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_0_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_1_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_2_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_3_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_4_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_5_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_6_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_7_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_8_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_8_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_8_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_8_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_8_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_9_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_9_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_9_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_9_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_9_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_10_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_10_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_10_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_10_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_10_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_11_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_11_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_11_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_11_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_11_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_12_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_12_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_12_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_12_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_12_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_13_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_13_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_13_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_13_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_13_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_14_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_14_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_14_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_14_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_14_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_15_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_15_wea : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_15_adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_15_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_15_web : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_15_lz : OUT STD_LOGIC
  );
END peaseNTT;

ARCHITECTURE v11 OF peaseNTT IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL yt_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yt_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_16_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_clka_en_d : STD_LOGIC;
  SIGNAL yt_rsc_0_16_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_17_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_18_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_19_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_20_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_21_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_22_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_23_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_24_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_25_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_26_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_27_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_28_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_29_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_30_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_31_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_16_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_17_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_18_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_19_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_20_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_21_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_22_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_23_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_24_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_25_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_26_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_27_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_28_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_29_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_30_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_31_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL twiddle_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL yt_rsc_0_0_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_0_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_web : STD_LOGIC;
  SIGNAL yt_rsc_0_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_1_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_1_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_1_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_web : STD_LOGIC;
  SIGNAL yt_rsc_0_1_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_1_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_1_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_2_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_2_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_2_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_web : STD_LOGIC;
  SIGNAL yt_rsc_0_2_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_2_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_2_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_3_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_3_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_3_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_web : STD_LOGIC;
  SIGNAL yt_rsc_0_3_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_3_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_3_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_4_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_4_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_4_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_web : STD_LOGIC;
  SIGNAL yt_rsc_0_4_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_4_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_4_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_5_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_5_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_5_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_web : STD_LOGIC;
  SIGNAL yt_rsc_0_5_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_5_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_5_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_6_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_6_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_6_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_web : STD_LOGIC;
  SIGNAL yt_rsc_0_6_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_6_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_6_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_7_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_7_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_7_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_web : STD_LOGIC;
  SIGNAL yt_rsc_0_7_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_7_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_7_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_8_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_8_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_8_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_web : STD_LOGIC;
  SIGNAL yt_rsc_0_8_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_8_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_8_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_9_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_9_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_9_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_web : STD_LOGIC;
  SIGNAL yt_rsc_0_9_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_9_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_9_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_10_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_10_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_10_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_web : STD_LOGIC;
  SIGNAL yt_rsc_0_10_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_10_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_10_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_11_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_11_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_11_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_web : STD_LOGIC;
  SIGNAL yt_rsc_0_11_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_11_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_11_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_12_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_12_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_12_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_web : STD_LOGIC;
  SIGNAL yt_rsc_0_12_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_12_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_12_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_13_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_13_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_13_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_web : STD_LOGIC;
  SIGNAL yt_rsc_0_13_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_13_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_13_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_14_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_14_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_14_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_web : STD_LOGIC;
  SIGNAL yt_rsc_0_14_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_14_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_14_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_15_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_15_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_15_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_web : STD_LOGIC;
  SIGNAL yt_rsc_0_15_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_15_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_15_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_16_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_16_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_16_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_web : STD_LOGIC;
  SIGNAL yt_rsc_0_16_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_16_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_16_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_17_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_17_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_17_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_web : STD_LOGIC;
  SIGNAL yt_rsc_0_17_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_17_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_17_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_18_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_18_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_18_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_web : STD_LOGIC;
  SIGNAL yt_rsc_0_18_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_18_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_18_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_19_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_19_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_19_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_web : STD_LOGIC;
  SIGNAL yt_rsc_0_19_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_19_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_19_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_20_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_20_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_20_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_web : STD_LOGIC;
  SIGNAL yt_rsc_0_20_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_20_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_20_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_21_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_21_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_21_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_web : STD_LOGIC;
  SIGNAL yt_rsc_0_21_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_21_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_21_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_22_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_22_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_22_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_web : STD_LOGIC;
  SIGNAL yt_rsc_0_22_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_22_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_22_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_23_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_23_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_23_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_web : STD_LOGIC;
  SIGNAL yt_rsc_0_23_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_23_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_23_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_24_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_24_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_24_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_web : STD_LOGIC;
  SIGNAL yt_rsc_0_24_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_24_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_24_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_25_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_25_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_25_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_web : STD_LOGIC;
  SIGNAL yt_rsc_0_25_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_25_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_25_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_26_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_26_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_26_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_web : STD_LOGIC;
  SIGNAL yt_rsc_0_26_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_26_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_26_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_27_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_27_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_27_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_web : STD_LOGIC;
  SIGNAL yt_rsc_0_27_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_27_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_27_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_28_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_28_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_28_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_web : STD_LOGIC;
  SIGNAL yt_rsc_0_28_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_28_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_28_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_29_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_29_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_29_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_web : STD_LOGIC;
  SIGNAL yt_rsc_0_29_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_29_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_29_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_30_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_30_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_30_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_web : STD_LOGIC;
  SIGNAL yt_rsc_0_30_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_30_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_30_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_31_clkb_en : STD_LOGIC;
  SIGNAL yt_rsc_0_31_clka_en : STD_LOGIC;
  SIGNAL yt_rsc_0_31_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_web : STD_LOGIC;
  SIGNAL yt_rsc_0_31_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_31_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_31_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_wea_d_iff : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_wea_d_iff : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_wea_d_iff : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_wea_d_iff : STD_LOGIC_VECTOR (1 DOWNTO 0);

  SIGNAL yt_rsc_0_0_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_0_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_1_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_1_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_1_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_2_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_2_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_2_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_3_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_3_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_3_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_4_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_4_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_4_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_5_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_5_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_5_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_6_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_6_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_6_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_7_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_7_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_7_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_8_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_8_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_8_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_9_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_9_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_9_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_10_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_10_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_10_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_11_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_11_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_11_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_12_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_12_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_12_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_13_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_13_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_13_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_14_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_14_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_14_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_15_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_15_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_15_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_16_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_16_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_16_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_17_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_17_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_17_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_18_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_18_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_18_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_19_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_19_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_19_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_20_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_20_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_20_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_21_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_21_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_21_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_22_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_22_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_22_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_23_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_23_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_23_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_24_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_24_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_24_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_25_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_25_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_25_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_26_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_26_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_26_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_27_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_27_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_27_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_28_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_28_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_28_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_29_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_29_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_29_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_30_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_30_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_30_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_31_comp_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_31_comp_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_31_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_7_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_8_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_1_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_9_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_2_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_10_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_3_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_11_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_4_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_12_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_5_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_13_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_6_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_14_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_7_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_15_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_8_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_16_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_9_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_17_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_10_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_18_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_11_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_19_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_12_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_20_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_13_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_21_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_14_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_22_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_15_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_23_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_16_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_16_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_24_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_17_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_17_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_25_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_18_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_18_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_26_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_19_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_19_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_27_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_20_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_20_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_28_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_21_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_21_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_29_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_22_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_22_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_30_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_23_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_23_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_31_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_24_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_24_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_32_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_25_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_25_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_33_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_26_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_26_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_34_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_27_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_27_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_35_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_28_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_28_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_36_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_29_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_29_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_37_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_30_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_30_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_38_8_32_256_256_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_31_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yt_rsc_0_31_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_39_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_40_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_1_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_41_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_2_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_42_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_3_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_43_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_4_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_44_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_5_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_45_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_6_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_46_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_7_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_47_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_8_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_48_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_9_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_49_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_10_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_50_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_11_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_51_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_12_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_52_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_13_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_53_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_14_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_54_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_15_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_55_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_16_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_16_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_56_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_17_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_17_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_57_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_18_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_18_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_58_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_19_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_19_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_59_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_20_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_20_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_60_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_21_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_21_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_61_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_22_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_22_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_62_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_23_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_23_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_63_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_24_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_24_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_64_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_25_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_25_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_65_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_26_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_26_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_66_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_27_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_27_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_67_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_28_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_28_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_68_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_29_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_29_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_69_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_30_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_30_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_70_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_31_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xt_rsc_0_31_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_71_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_72_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_1_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_73_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_2_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_74_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_3_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_75_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_4_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_76_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_5_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_77_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_6_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_78_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_7_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_79_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_8_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_80_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_9_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_81_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_10_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_82_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_11_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_83_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_12_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_84_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_13_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_85_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_14_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_86_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_15_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1
      DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_87_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_88_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_1_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_89_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_2_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_90_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_3_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_91_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_4_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_92_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_5_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_93_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_6_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_94_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_7_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_95_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_8_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_96_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_9_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_97_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_10_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_98_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_11_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_99_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_12_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_100_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_13_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_101_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_14_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_102_8_32_256_256_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_15_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_adrb : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_adra_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);

  COMPONENT peaseNTT_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_16_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_17_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_18_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_19_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_20_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_21_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_22_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_23_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_24_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_25_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_26_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_27_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_28_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_29_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_30_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_31_lz : OUT STD_LOGIC;
      p_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      p_rsc_triosy_lz : OUT STD_LOGIC;
      r_rsc_triosy_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      yt_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_0_i_clka_en_d : OUT STD_LOGIC;
      yt_rsc_0_0_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_1_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_1_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_2_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_2_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_3_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_3_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_4_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_4_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_5_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_5_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_6_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_6_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_7_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_7_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_8_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_8_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_9_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_9_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_10_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_10_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_11_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_11_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_12_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_12_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_13_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_13_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_14_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_14_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_15_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_15_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_16_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_16_i_clka_en_d : OUT STD_LOGIC;
      yt_rsc_0_16_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_16_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_17_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_17_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_17_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_18_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_18_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_18_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_19_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_19_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_19_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_20_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_20_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_20_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_21_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_21_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_21_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_22_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_22_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_22_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_23_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_23_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_23_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_24_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_24_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_24_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_25_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_25_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_25_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_26_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_26_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_26_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_27_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_27_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_27_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_28_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_28_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_28_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_29_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_29_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_29_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_30_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_30_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_30_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yt_rsc_0_31_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      yt_rsc_0_31_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_31_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_0_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_1_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_1_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_2_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_2_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_3_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_3_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_4_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_4_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_5_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_5_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_6_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_6_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_7_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_7_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_8_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_8_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_9_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_9_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_10_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_10_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_11_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_11_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_12_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_12_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_13_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_13_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_14_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_14_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_15_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_15_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_16_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_16_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_16_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_17_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_17_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_17_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_18_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_18_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_18_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_19_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_19_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_19_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_20_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_20_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_20_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_21_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_21_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_21_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_22_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_22_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_22_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_23_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_23_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_23_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_24_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_24_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_24_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_25_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_25_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_25_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_26_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_26_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_26_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_27_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_27_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_27_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_28_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_28_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_28_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_29_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_29_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_29_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_30_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_30_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_30_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xt_rsc_0_31_i_adra_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      xt_rsc_0_31_i_da_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_31_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      twiddle_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_1_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_2_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_3_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_4_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_5_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_6_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_7_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_8_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_9_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1
          DOWNTO 0);
      twiddle_rsc_0_10_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_rsc_0_11_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_rsc_0_12_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_rsc_0_13_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_rsc_0_14_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_rsc_0_15_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_1_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_2_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_3_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_4_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_5_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_6_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_7_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_8_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_9_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_10_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_11_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_12_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_13_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_14_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      twiddle_h_rsc_0_15_i_adra_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      yt_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yt_rsc_0_16_i_wea_d_pff : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xt_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xt_rsc_0_16_i_wea_d_pff : OUT STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_inst_p_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_8_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_9_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_10_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_11_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_12_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_13_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_14_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_15_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_16_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_16_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_16_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_17_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_17_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_17_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_18_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_18_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_18_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_19_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_19_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_19_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_20_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_20_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_20_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_21_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_21_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_21_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_22_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_22_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_22_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_23_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_23_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_23_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_24_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_24_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_24_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_25_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_25_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_25_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_26_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_26_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_26_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_27_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_27_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_27_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_28_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_28_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_28_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_29_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_29_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_29_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_30_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_30_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_30_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_31_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_31_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_31_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_8_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_9_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_10_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_11_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_12_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_13_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_14_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_15_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_16_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_16_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_16_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_17_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_17_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_17_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_18_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_18_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_18_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_19_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_19_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_19_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_20_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_20_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_20_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_21_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_21_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_21_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_22_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_22_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_22_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_23_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_23_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_23_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_24_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_24_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_24_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_25_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_25_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_25_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_26_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_26_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_26_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_27_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_27_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_27_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_28_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_28_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_28_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_29_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_29_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_29_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_30_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_30_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_30_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_31_i_adra_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_31_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_31_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d :
      STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_0_i_wea_d_pff : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_16_i_wea_d_pff : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_0_i_wea_d_pff : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_16_i_wea_d_pff : STD_LOGIC_VECTOR (1 DOWNTO
      0);

BEGIN
  yt_rsc_0_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_0_comp_adra,
      adrb => yt_rsc_0_0_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_0_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_0_clkb_en,
      da => yt_rsc_0_0_comp_da,
      db => yt_rsc_0_0_comp_db,
      qa => yt_rsc_0_0_comp_qa,
      qb => yt_rsc_0_0_comp_qb,
      wea => yt_rsc_0_0_wea,
      web => yt_rsc_0_0_web
    );
  yt_rsc_0_0_comp_adra <= yt_rsc_0_0_adra;
  yt_rsc_0_0_comp_adrb <= yt_rsc_0_0_adrb;
  yt_rsc_0_0_comp_da <= yt_rsc_0_0_da;
  yt_rsc_0_0_comp_db <= yt_rsc_0_0_db;
  yt_rsc_0_0_qa <= yt_rsc_0_0_comp_qa;
  yt_rsc_0_0_qb <= yt_rsc_0_0_comp_qb;

  yt_rsc_0_1_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_1_comp_adra,
      adrb => yt_rsc_0_1_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_1_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_1_clkb_en,
      da => yt_rsc_0_1_comp_da,
      db => yt_rsc_0_1_comp_db,
      qa => yt_rsc_0_1_comp_qa,
      qb => yt_rsc_0_1_comp_qb,
      wea => yt_rsc_0_1_wea,
      web => yt_rsc_0_1_web
    );
  yt_rsc_0_1_comp_adra <= yt_rsc_0_1_adra;
  yt_rsc_0_1_comp_adrb <= yt_rsc_0_1_adrb;
  yt_rsc_0_1_comp_da <= yt_rsc_0_1_da;
  yt_rsc_0_1_comp_db <= yt_rsc_0_1_db;
  yt_rsc_0_1_qa <= yt_rsc_0_1_comp_qa;
  yt_rsc_0_1_qb <= yt_rsc_0_1_comp_qb;

  yt_rsc_0_2_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_2_comp_adra,
      adrb => yt_rsc_0_2_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_2_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_2_clkb_en,
      da => yt_rsc_0_2_comp_da,
      db => yt_rsc_0_2_comp_db,
      qa => yt_rsc_0_2_comp_qa,
      qb => yt_rsc_0_2_comp_qb,
      wea => yt_rsc_0_2_wea,
      web => yt_rsc_0_2_web
    );
  yt_rsc_0_2_comp_adra <= yt_rsc_0_2_adra;
  yt_rsc_0_2_comp_adrb <= yt_rsc_0_2_adrb;
  yt_rsc_0_2_comp_da <= yt_rsc_0_2_da;
  yt_rsc_0_2_comp_db <= yt_rsc_0_2_db;
  yt_rsc_0_2_qa <= yt_rsc_0_2_comp_qa;
  yt_rsc_0_2_qb <= yt_rsc_0_2_comp_qb;

  yt_rsc_0_3_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_3_comp_adra,
      adrb => yt_rsc_0_3_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_3_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_3_clkb_en,
      da => yt_rsc_0_3_comp_da,
      db => yt_rsc_0_3_comp_db,
      qa => yt_rsc_0_3_comp_qa,
      qb => yt_rsc_0_3_comp_qb,
      wea => yt_rsc_0_3_wea,
      web => yt_rsc_0_3_web
    );
  yt_rsc_0_3_comp_adra <= yt_rsc_0_3_adra;
  yt_rsc_0_3_comp_adrb <= yt_rsc_0_3_adrb;
  yt_rsc_0_3_comp_da <= yt_rsc_0_3_da;
  yt_rsc_0_3_comp_db <= yt_rsc_0_3_db;
  yt_rsc_0_3_qa <= yt_rsc_0_3_comp_qa;
  yt_rsc_0_3_qb <= yt_rsc_0_3_comp_qb;

  yt_rsc_0_4_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_4_comp_adra,
      adrb => yt_rsc_0_4_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_4_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_4_clkb_en,
      da => yt_rsc_0_4_comp_da,
      db => yt_rsc_0_4_comp_db,
      qa => yt_rsc_0_4_comp_qa,
      qb => yt_rsc_0_4_comp_qb,
      wea => yt_rsc_0_4_wea,
      web => yt_rsc_0_4_web
    );
  yt_rsc_0_4_comp_adra <= yt_rsc_0_4_adra;
  yt_rsc_0_4_comp_adrb <= yt_rsc_0_4_adrb;
  yt_rsc_0_4_comp_da <= yt_rsc_0_4_da;
  yt_rsc_0_4_comp_db <= yt_rsc_0_4_db;
  yt_rsc_0_4_qa <= yt_rsc_0_4_comp_qa;
  yt_rsc_0_4_qb <= yt_rsc_0_4_comp_qb;

  yt_rsc_0_5_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_5_comp_adra,
      adrb => yt_rsc_0_5_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_5_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_5_clkb_en,
      da => yt_rsc_0_5_comp_da,
      db => yt_rsc_0_5_comp_db,
      qa => yt_rsc_0_5_comp_qa,
      qb => yt_rsc_0_5_comp_qb,
      wea => yt_rsc_0_5_wea,
      web => yt_rsc_0_5_web
    );
  yt_rsc_0_5_comp_adra <= yt_rsc_0_5_adra;
  yt_rsc_0_5_comp_adrb <= yt_rsc_0_5_adrb;
  yt_rsc_0_5_comp_da <= yt_rsc_0_5_da;
  yt_rsc_0_5_comp_db <= yt_rsc_0_5_db;
  yt_rsc_0_5_qa <= yt_rsc_0_5_comp_qa;
  yt_rsc_0_5_qb <= yt_rsc_0_5_comp_qb;

  yt_rsc_0_6_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_6_comp_adra,
      adrb => yt_rsc_0_6_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_6_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_6_clkb_en,
      da => yt_rsc_0_6_comp_da,
      db => yt_rsc_0_6_comp_db,
      qa => yt_rsc_0_6_comp_qa,
      qb => yt_rsc_0_6_comp_qb,
      wea => yt_rsc_0_6_wea,
      web => yt_rsc_0_6_web
    );
  yt_rsc_0_6_comp_adra <= yt_rsc_0_6_adra;
  yt_rsc_0_6_comp_adrb <= yt_rsc_0_6_adrb;
  yt_rsc_0_6_comp_da <= yt_rsc_0_6_da;
  yt_rsc_0_6_comp_db <= yt_rsc_0_6_db;
  yt_rsc_0_6_qa <= yt_rsc_0_6_comp_qa;
  yt_rsc_0_6_qb <= yt_rsc_0_6_comp_qb;

  yt_rsc_0_7_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_7_comp_adra,
      adrb => yt_rsc_0_7_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_7_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_7_clkb_en,
      da => yt_rsc_0_7_comp_da,
      db => yt_rsc_0_7_comp_db,
      qa => yt_rsc_0_7_comp_qa,
      qb => yt_rsc_0_7_comp_qb,
      wea => yt_rsc_0_7_wea,
      web => yt_rsc_0_7_web
    );
  yt_rsc_0_7_comp_adra <= yt_rsc_0_7_adra;
  yt_rsc_0_7_comp_adrb <= yt_rsc_0_7_adrb;
  yt_rsc_0_7_comp_da <= yt_rsc_0_7_da;
  yt_rsc_0_7_comp_db <= yt_rsc_0_7_db;
  yt_rsc_0_7_qa <= yt_rsc_0_7_comp_qa;
  yt_rsc_0_7_qb <= yt_rsc_0_7_comp_qb;

  yt_rsc_0_8_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_8_comp_adra,
      adrb => yt_rsc_0_8_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_8_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_8_clkb_en,
      da => yt_rsc_0_8_comp_da,
      db => yt_rsc_0_8_comp_db,
      qa => yt_rsc_0_8_comp_qa,
      qb => yt_rsc_0_8_comp_qb,
      wea => yt_rsc_0_8_wea,
      web => yt_rsc_0_8_web
    );
  yt_rsc_0_8_comp_adra <= yt_rsc_0_8_adra;
  yt_rsc_0_8_comp_adrb <= yt_rsc_0_8_adrb;
  yt_rsc_0_8_comp_da <= yt_rsc_0_8_da;
  yt_rsc_0_8_comp_db <= yt_rsc_0_8_db;
  yt_rsc_0_8_qa <= yt_rsc_0_8_comp_qa;
  yt_rsc_0_8_qb <= yt_rsc_0_8_comp_qb;

  yt_rsc_0_9_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_9_comp_adra,
      adrb => yt_rsc_0_9_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_9_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_9_clkb_en,
      da => yt_rsc_0_9_comp_da,
      db => yt_rsc_0_9_comp_db,
      qa => yt_rsc_0_9_comp_qa,
      qb => yt_rsc_0_9_comp_qb,
      wea => yt_rsc_0_9_wea,
      web => yt_rsc_0_9_web
    );
  yt_rsc_0_9_comp_adra <= yt_rsc_0_9_adra;
  yt_rsc_0_9_comp_adrb <= yt_rsc_0_9_adrb;
  yt_rsc_0_9_comp_da <= yt_rsc_0_9_da;
  yt_rsc_0_9_comp_db <= yt_rsc_0_9_db;
  yt_rsc_0_9_qa <= yt_rsc_0_9_comp_qa;
  yt_rsc_0_9_qb <= yt_rsc_0_9_comp_qb;

  yt_rsc_0_10_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_10_comp_adra,
      adrb => yt_rsc_0_10_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_10_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_10_clkb_en,
      da => yt_rsc_0_10_comp_da,
      db => yt_rsc_0_10_comp_db,
      qa => yt_rsc_0_10_comp_qa,
      qb => yt_rsc_0_10_comp_qb,
      wea => yt_rsc_0_10_wea,
      web => yt_rsc_0_10_web
    );
  yt_rsc_0_10_comp_adra <= yt_rsc_0_10_adra;
  yt_rsc_0_10_comp_adrb <= yt_rsc_0_10_adrb;
  yt_rsc_0_10_comp_da <= yt_rsc_0_10_da;
  yt_rsc_0_10_comp_db <= yt_rsc_0_10_db;
  yt_rsc_0_10_qa <= yt_rsc_0_10_comp_qa;
  yt_rsc_0_10_qb <= yt_rsc_0_10_comp_qb;

  yt_rsc_0_11_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_11_comp_adra,
      adrb => yt_rsc_0_11_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_11_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_11_clkb_en,
      da => yt_rsc_0_11_comp_da,
      db => yt_rsc_0_11_comp_db,
      qa => yt_rsc_0_11_comp_qa,
      qb => yt_rsc_0_11_comp_qb,
      wea => yt_rsc_0_11_wea,
      web => yt_rsc_0_11_web
    );
  yt_rsc_0_11_comp_adra <= yt_rsc_0_11_adra;
  yt_rsc_0_11_comp_adrb <= yt_rsc_0_11_adrb;
  yt_rsc_0_11_comp_da <= yt_rsc_0_11_da;
  yt_rsc_0_11_comp_db <= yt_rsc_0_11_db;
  yt_rsc_0_11_qa <= yt_rsc_0_11_comp_qa;
  yt_rsc_0_11_qb <= yt_rsc_0_11_comp_qb;

  yt_rsc_0_12_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_12_comp_adra,
      adrb => yt_rsc_0_12_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_12_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_12_clkb_en,
      da => yt_rsc_0_12_comp_da,
      db => yt_rsc_0_12_comp_db,
      qa => yt_rsc_0_12_comp_qa,
      qb => yt_rsc_0_12_comp_qb,
      wea => yt_rsc_0_12_wea,
      web => yt_rsc_0_12_web
    );
  yt_rsc_0_12_comp_adra <= yt_rsc_0_12_adra;
  yt_rsc_0_12_comp_adrb <= yt_rsc_0_12_adrb;
  yt_rsc_0_12_comp_da <= yt_rsc_0_12_da;
  yt_rsc_0_12_comp_db <= yt_rsc_0_12_db;
  yt_rsc_0_12_qa <= yt_rsc_0_12_comp_qa;
  yt_rsc_0_12_qb <= yt_rsc_0_12_comp_qb;

  yt_rsc_0_13_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_13_comp_adra,
      adrb => yt_rsc_0_13_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_13_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_13_clkb_en,
      da => yt_rsc_0_13_comp_da,
      db => yt_rsc_0_13_comp_db,
      qa => yt_rsc_0_13_comp_qa,
      qb => yt_rsc_0_13_comp_qb,
      wea => yt_rsc_0_13_wea,
      web => yt_rsc_0_13_web
    );
  yt_rsc_0_13_comp_adra <= yt_rsc_0_13_adra;
  yt_rsc_0_13_comp_adrb <= yt_rsc_0_13_adrb;
  yt_rsc_0_13_comp_da <= yt_rsc_0_13_da;
  yt_rsc_0_13_comp_db <= yt_rsc_0_13_db;
  yt_rsc_0_13_qa <= yt_rsc_0_13_comp_qa;
  yt_rsc_0_13_qb <= yt_rsc_0_13_comp_qb;

  yt_rsc_0_14_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_14_comp_adra,
      adrb => yt_rsc_0_14_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_14_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_14_clkb_en,
      da => yt_rsc_0_14_comp_da,
      db => yt_rsc_0_14_comp_db,
      qa => yt_rsc_0_14_comp_qa,
      qb => yt_rsc_0_14_comp_qb,
      wea => yt_rsc_0_14_wea,
      web => yt_rsc_0_14_web
    );
  yt_rsc_0_14_comp_adra <= yt_rsc_0_14_adra;
  yt_rsc_0_14_comp_adrb <= yt_rsc_0_14_adrb;
  yt_rsc_0_14_comp_da <= yt_rsc_0_14_da;
  yt_rsc_0_14_comp_db <= yt_rsc_0_14_db;
  yt_rsc_0_14_qa <= yt_rsc_0_14_comp_qa;
  yt_rsc_0_14_qb <= yt_rsc_0_14_comp_qb;

  yt_rsc_0_15_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_15_comp_adra,
      adrb => yt_rsc_0_15_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_15_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_15_clkb_en,
      da => yt_rsc_0_15_comp_da,
      db => yt_rsc_0_15_comp_db,
      qa => yt_rsc_0_15_comp_qa,
      qb => yt_rsc_0_15_comp_qb,
      wea => yt_rsc_0_15_wea,
      web => yt_rsc_0_15_web
    );
  yt_rsc_0_15_comp_adra <= yt_rsc_0_15_adra;
  yt_rsc_0_15_comp_adrb <= yt_rsc_0_15_adrb;
  yt_rsc_0_15_comp_da <= yt_rsc_0_15_da;
  yt_rsc_0_15_comp_db <= yt_rsc_0_15_db;
  yt_rsc_0_15_qa <= yt_rsc_0_15_comp_qa;
  yt_rsc_0_15_qb <= yt_rsc_0_15_comp_qb;

  yt_rsc_0_16_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_16_comp_adra,
      adrb => yt_rsc_0_16_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_16_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_16_clkb_en,
      da => yt_rsc_0_16_comp_da,
      db => yt_rsc_0_16_comp_db,
      qa => yt_rsc_0_16_comp_qa,
      qb => yt_rsc_0_16_comp_qb,
      wea => yt_rsc_0_16_wea,
      web => yt_rsc_0_16_web
    );
  yt_rsc_0_16_comp_adra <= yt_rsc_0_16_adra;
  yt_rsc_0_16_comp_adrb <= yt_rsc_0_16_adrb;
  yt_rsc_0_16_comp_da <= yt_rsc_0_16_da;
  yt_rsc_0_16_comp_db <= yt_rsc_0_16_db;
  yt_rsc_0_16_qa <= yt_rsc_0_16_comp_qa;
  yt_rsc_0_16_qb <= yt_rsc_0_16_comp_qb;

  yt_rsc_0_17_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_17_comp_adra,
      adrb => yt_rsc_0_17_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_17_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_17_clkb_en,
      da => yt_rsc_0_17_comp_da,
      db => yt_rsc_0_17_comp_db,
      qa => yt_rsc_0_17_comp_qa,
      qb => yt_rsc_0_17_comp_qb,
      wea => yt_rsc_0_17_wea,
      web => yt_rsc_0_17_web
    );
  yt_rsc_0_17_comp_adra <= yt_rsc_0_17_adra;
  yt_rsc_0_17_comp_adrb <= yt_rsc_0_17_adrb;
  yt_rsc_0_17_comp_da <= yt_rsc_0_17_da;
  yt_rsc_0_17_comp_db <= yt_rsc_0_17_db;
  yt_rsc_0_17_qa <= yt_rsc_0_17_comp_qa;
  yt_rsc_0_17_qb <= yt_rsc_0_17_comp_qb;

  yt_rsc_0_18_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_18_comp_adra,
      adrb => yt_rsc_0_18_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_18_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_18_clkb_en,
      da => yt_rsc_0_18_comp_da,
      db => yt_rsc_0_18_comp_db,
      qa => yt_rsc_0_18_comp_qa,
      qb => yt_rsc_0_18_comp_qb,
      wea => yt_rsc_0_18_wea,
      web => yt_rsc_0_18_web
    );
  yt_rsc_0_18_comp_adra <= yt_rsc_0_18_adra;
  yt_rsc_0_18_comp_adrb <= yt_rsc_0_18_adrb;
  yt_rsc_0_18_comp_da <= yt_rsc_0_18_da;
  yt_rsc_0_18_comp_db <= yt_rsc_0_18_db;
  yt_rsc_0_18_qa <= yt_rsc_0_18_comp_qa;
  yt_rsc_0_18_qb <= yt_rsc_0_18_comp_qb;

  yt_rsc_0_19_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_19_comp_adra,
      adrb => yt_rsc_0_19_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_19_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_19_clkb_en,
      da => yt_rsc_0_19_comp_da,
      db => yt_rsc_0_19_comp_db,
      qa => yt_rsc_0_19_comp_qa,
      qb => yt_rsc_0_19_comp_qb,
      wea => yt_rsc_0_19_wea,
      web => yt_rsc_0_19_web
    );
  yt_rsc_0_19_comp_adra <= yt_rsc_0_19_adra;
  yt_rsc_0_19_comp_adrb <= yt_rsc_0_19_adrb;
  yt_rsc_0_19_comp_da <= yt_rsc_0_19_da;
  yt_rsc_0_19_comp_db <= yt_rsc_0_19_db;
  yt_rsc_0_19_qa <= yt_rsc_0_19_comp_qa;
  yt_rsc_0_19_qb <= yt_rsc_0_19_comp_qb;

  yt_rsc_0_20_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_20_comp_adra,
      adrb => yt_rsc_0_20_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_20_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_20_clkb_en,
      da => yt_rsc_0_20_comp_da,
      db => yt_rsc_0_20_comp_db,
      qa => yt_rsc_0_20_comp_qa,
      qb => yt_rsc_0_20_comp_qb,
      wea => yt_rsc_0_20_wea,
      web => yt_rsc_0_20_web
    );
  yt_rsc_0_20_comp_adra <= yt_rsc_0_20_adra;
  yt_rsc_0_20_comp_adrb <= yt_rsc_0_20_adrb;
  yt_rsc_0_20_comp_da <= yt_rsc_0_20_da;
  yt_rsc_0_20_comp_db <= yt_rsc_0_20_db;
  yt_rsc_0_20_qa <= yt_rsc_0_20_comp_qa;
  yt_rsc_0_20_qb <= yt_rsc_0_20_comp_qb;

  yt_rsc_0_21_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_21_comp_adra,
      adrb => yt_rsc_0_21_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_21_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_21_clkb_en,
      da => yt_rsc_0_21_comp_da,
      db => yt_rsc_0_21_comp_db,
      qa => yt_rsc_0_21_comp_qa,
      qb => yt_rsc_0_21_comp_qb,
      wea => yt_rsc_0_21_wea,
      web => yt_rsc_0_21_web
    );
  yt_rsc_0_21_comp_adra <= yt_rsc_0_21_adra;
  yt_rsc_0_21_comp_adrb <= yt_rsc_0_21_adrb;
  yt_rsc_0_21_comp_da <= yt_rsc_0_21_da;
  yt_rsc_0_21_comp_db <= yt_rsc_0_21_db;
  yt_rsc_0_21_qa <= yt_rsc_0_21_comp_qa;
  yt_rsc_0_21_qb <= yt_rsc_0_21_comp_qb;

  yt_rsc_0_22_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_22_comp_adra,
      adrb => yt_rsc_0_22_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_22_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_22_clkb_en,
      da => yt_rsc_0_22_comp_da,
      db => yt_rsc_0_22_comp_db,
      qa => yt_rsc_0_22_comp_qa,
      qb => yt_rsc_0_22_comp_qb,
      wea => yt_rsc_0_22_wea,
      web => yt_rsc_0_22_web
    );
  yt_rsc_0_22_comp_adra <= yt_rsc_0_22_adra;
  yt_rsc_0_22_comp_adrb <= yt_rsc_0_22_adrb;
  yt_rsc_0_22_comp_da <= yt_rsc_0_22_da;
  yt_rsc_0_22_comp_db <= yt_rsc_0_22_db;
  yt_rsc_0_22_qa <= yt_rsc_0_22_comp_qa;
  yt_rsc_0_22_qb <= yt_rsc_0_22_comp_qb;

  yt_rsc_0_23_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_23_comp_adra,
      adrb => yt_rsc_0_23_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_23_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_23_clkb_en,
      da => yt_rsc_0_23_comp_da,
      db => yt_rsc_0_23_comp_db,
      qa => yt_rsc_0_23_comp_qa,
      qb => yt_rsc_0_23_comp_qb,
      wea => yt_rsc_0_23_wea,
      web => yt_rsc_0_23_web
    );
  yt_rsc_0_23_comp_adra <= yt_rsc_0_23_adra;
  yt_rsc_0_23_comp_adrb <= yt_rsc_0_23_adrb;
  yt_rsc_0_23_comp_da <= yt_rsc_0_23_da;
  yt_rsc_0_23_comp_db <= yt_rsc_0_23_db;
  yt_rsc_0_23_qa <= yt_rsc_0_23_comp_qa;
  yt_rsc_0_23_qb <= yt_rsc_0_23_comp_qb;

  yt_rsc_0_24_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_24_comp_adra,
      adrb => yt_rsc_0_24_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_24_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_24_clkb_en,
      da => yt_rsc_0_24_comp_da,
      db => yt_rsc_0_24_comp_db,
      qa => yt_rsc_0_24_comp_qa,
      qb => yt_rsc_0_24_comp_qb,
      wea => yt_rsc_0_24_wea,
      web => yt_rsc_0_24_web
    );
  yt_rsc_0_24_comp_adra <= yt_rsc_0_24_adra;
  yt_rsc_0_24_comp_adrb <= yt_rsc_0_24_adrb;
  yt_rsc_0_24_comp_da <= yt_rsc_0_24_da;
  yt_rsc_0_24_comp_db <= yt_rsc_0_24_db;
  yt_rsc_0_24_qa <= yt_rsc_0_24_comp_qa;
  yt_rsc_0_24_qb <= yt_rsc_0_24_comp_qb;

  yt_rsc_0_25_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_25_comp_adra,
      adrb => yt_rsc_0_25_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_25_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_25_clkb_en,
      da => yt_rsc_0_25_comp_da,
      db => yt_rsc_0_25_comp_db,
      qa => yt_rsc_0_25_comp_qa,
      qb => yt_rsc_0_25_comp_qb,
      wea => yt_rsc_0_25_wea,
      web => yt_rsc_0_25_web
    );
  yt_rsc_0_25_comp_adra <= yt_rsc_0_25_adra;
  yt_rsc_0_25_comp_adrb <= yt_rsc_0_25_adrb;
  yt_rsc_0_25_comp_da <= yt_rsc_0_25_da;
  yt_rsc_0_25_comp_db <= yt_rsc_0_25_db;
  yt_rsc_0_25_qa <= yt_rsc_0_25_comp_qa;
  yt_rsc_0_25_qb <= yt_rsc_0_25_comp_qb;

  yt_rsc_0_26_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_26_comp_adra,
      adrb => yt_rsc_0_26_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_26_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_26_clkb_en,
      da => yt_rsc_0_26_comp_da,
      db => yt_rsc_0_26_comp_db,
      qa => yt_rsc_0_26_comp_qa,
      qb => yt_rsc_0_26_comp_qb,
      wea => yt_rsc_0_26_wea,
      web => yt_rsc_0_26_web
    );
  yt_rsc_0_26_comp_adra <= yt_rsc_0_26_adra;
  yt_rsc_0_26_comp_adrb <= yt_rsc_0_26_adrb;
  yt_rsc_0_26_comp_da <= yt_rsc_0_26_da;
  yt_rsc_0_26_comp_db <= yt_rsc_0_26_db;
  yt_rsc_0_26_qa <= yt_rsc_0_26_comp_qa;
  yt_rsc_0_26_qb <= yt_rsc_0_26_comp_qb;

  yt_rsc_0_27_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_27_comp_adra,
      adrb => yt_rsc_0_27_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_27_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_27_clkb_en,
      da => yt_rsc_0_27_comp_da,
      db => yt_rsc_0_27_comp_db,
      qa => yt_rsc_0_27_comp_qa,
      qb => yt_rsc_0_27_comp_qb,
      wea => yt_rsc_0_27_wea,
      web => yt_rsc_0_27_web
    );
  yt_rsc_0_27_comp_adra <= yt_rsc_0_27_adra;
  yt_rsc_0_27_comp_adrb <= yt_rsc_0_27_adrb;
  yt_rsc_0_27_comp_da <= yt_rsc_0_27_da;
  yt_rsc_0_27_comp_db <= yt_rsc_0_27_db;
  yt_rsc_0_27_qa <= yt_rsc_0_27_comp_qa;
  yt_rsc_0_27_qb <= yt_rsc_0_27_comp_qb;

  yt_rsc_0_28_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_28_comp_adra,
      adrb => yt_rsc_0_28_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_28_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_28_clkb_en,
      da => yt_rsc_0_28_comp_da,
      db => yt_rsc_0_28_comp_db,
      qa => yt_rsc_0_28_comp_qa,
      qb => yt_rsc_0_28_comp_qb,
      wea => yt_rsc_0_28_wea,
      web => yt_rsc_0_28_web
    );
  yt_rsc_0_28_comp_adra <= yt_rsc_0_28_adra;
  yt_rsc_0_28_comp_adrb <= yt_rsc_0_28_adrb;
  yt_rsc_0_28_comp_da <= yt_rsc_0_28_da;
  yt_rsc_0_28_comp_db <= yt_rsc_0_28_db;
  yt_rsc_0_28_qa <= yt_rsc_0_28_comp_qa;
  yt_rsc_0_28_qb <= yt_rsc_0_28_comp_qb;

  yt_rsc_0_29_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_29_comp_adra,
      adrb => yt_rsc_0_29_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_29_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_29_clkb_en,
      da => yt_rsc_0_29_comp_da,
      db => yt_rsc_0_29_comp_db,
      qa => yt_rsc_0_29_comp_qa,
      qb => yt_rsc_0_29_comp_qb,
      wea => yt_rsc_0_29_wea,
      web => yt_rsc_0_29_web
    );
  yt_rsc_0_29_comp_adra <= yt_rsc_0_29_adra;
  yt_rsc_0_29_comp_adrb <= yt_rsc_0_29_adrb;
  yt_rsc_0_29_comp_da <= yt_rsc_0_29_da;
  yt_rsc_0_29_comp_db <= yt_rsc_0_29_db;
  yt_rsc_0_29_qa <= yt_rsc_0_29_comp_qa;
  yt_rsc_0_29_qb <= yt_rsc_0_29_comp_qb;

  yt_rsc_0_30_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_30_comp_adra,
      adrb => yt_rsc_0_30_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_30_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_30_clkb_en,
      da => yt_rsc_0_30_comp_da,
      db => yt_rsc_0_30_comp_db,
      qa => yt_rsc_0_30_comp_qa,
      qb => yt_rsc_0_30_comp_qb,
      wea => yt_rsc_0_30_wea,
      web => yt_rsc_0_30_web
    );
  yt_rsc_0_30_comp_adra <= yt_rsc_0_30_adra;
  yt_rsc_0_30_comp_adrb <= yt_rsc_0_30_adrb;
  yt_rsc_0_30_comp_da <= yt_rsc_0_30_da;
  yt_rsc_0_30_comp_db <= yt_rsc_0_30_db;
  yt_rsc_0_30_qa <= yt_rsc_0_30_comp_qa;
  yt_rsc_0_30_qb <= yt_rsc_0_30_comp_qb;

  yt_rsc_0_31_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 8,
      data_width => 32,
      depth => 256,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_31_comp_adra,
      adrb => yt_rsc_0_31_comp_adrb,
      clka => clk,
      clka_en => yt_rsc_0_31_clkb_en,
      clkb => clk,
      clkb_en => yt_rsc_0_31_clkb_en,
      da => yt_rsc_0_31_comp_da,
      db => yt_rsc_0_31_comp_db,
      qa => yt_rsc_0_31_comp_qa,
      qb => yt_rsc_0_31_comp_qb,
      wea => yt_rsc_0_31_wea,
      web => yt_rsc_0_31_web
    );
  yt_rsc_0_31_comp_adra <= yt_rsc_0_31_adra;
  yt_rsc_0_31_comp_adrb <= yt_rsc_0_31_adrb;
  yt_rsc_0_31_comp_da <= yt_rsc_0_31_da;
  yt_rsc_0_31_comp_db <= yt_rsc_0_31_db;
  yt_rsc_0_31_qa <= yt_rsc_0_31_comp_qa;
  yt_rsc_0_31_qb <= yt_rsc_0_31_comp_qb;

  yt_rsc_0_0_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_7_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_0_clkb_en,
      clka_en => yt_rsc_0_0_clka_en,
      qb => yt_rsc_0_0_i_qb,
      web => yt_rsc_0_0_web,
      db => yt_rsc_0_0_i_db,
      adrb => yt_rsc_0_0_i_adrb,
      qa => yt_rsc_0_0_i_qa,
      wea => yt_rsc_0_0_wea,
      da => yt_rsc_0_0_i_da,
      adra => yt_rsc_0_0_i_adra,
      adra_d => yt_rsc_0_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_0_i_clka_en_d,
      clkb_en_d => yt_rsc_0_0_i_clka_en_d,
      da_d => yt_rsc_0_0_i_da_d_1,
      qa_d => yt_rsc_0_0_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_0_i_qb <= yt_rsc_0_0_qb;
  yt_rsc_0_0_db <= yt_rsc_0_0_i_db;
  yt_rsc_0_0_adrb <= yt_rsc_0_0_i_adrb;
  yt_rsc_0_0_i_qa <= yt_rsc_0_0_qa;
  yt_rsc_0_0_da <= yt_rsc_0_0_i_da;
  yt_rsc_0_0_adra <= yt_rsc_0_0_i_adra;
  yt_rsc_0_0_i_adra_d_1 <= yt_rsc_0_0_i_adra_d;
  yt_rsc_0_0_i_da_d_1 <= yt_rsc_0_0_i_da_d;
  yt_rsc_0_0_i_qa_d <= yt_rsc_0_0_i_qa_d_1;
  yt_rsc_0_0_i_wea_d <= yt_rsc_0_0_i_wea_d_iff;
  yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_0_i_wea_d_iff;

  yt_rsc_0_1_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_8_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_1_clkb_en,
      clka_en => yt_rsc_0_1_clka_en,
      qb => yt_rsc_0_1_i_qb,
      web => yt_rsc_0_1_web,
      db => yt_rsc_0_1_i_db,
      adrb => yt_rsc_0_1_i_adrb,
      qa => yt_rsc_0_1_i_qa,
      wea => yt_rsc_0_1_wea,
      da => yt_rsc_0_1_i_da,
      adra => yt_rsc_0_1_i_adra,
      adra_d => yt_rsc_0_1_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_0_i_clka_en_d,
      clkb_en_d => yt_rsc_0_0_i_clka_en_d,
      da_d => yt_rsc_0_1_i_da_d_1,
      qa_d => yt_rsc_0_1_i_qa_d_1,
      wea_d => yt_rsc_0_1_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_1_i_qb <= yt_rsc_0_1_qb;
  yt_rsc_0_1_db <= yt_rsc_0_1_i_db;
  yt_rsc_0_1_adrb <= yt_rsc_0_1_i_adrb;
  yt_rsc_0_1_i_qa <= yt_rsc_0_1_qa;
  yt_rsc_0_1_da <= yt_rsc_0_1_i_da;
  yt_rsc_0_1_adra <= yt_rsc_0_1_i_adra;
  yt_rsc_0_1_i_adra_d_1 <= yt_rsc_0_1_i_adra_d;
  yt_rsc_0_1_i_da_d_1 <= yt_rsc_0_1_i_da_d;
  yt_rsc_0_1_i_qa_d <= yt_rsc_0_1_i_qa_d_1;
  yt_rsc_0_1_i_wea_d <= yt_rsc_0_0_i_wea_d_iff;
  yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_0_i_wea_d_iff;

  yt_rsc_0_2_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_9_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_2_clkb_en,
      clka_en => yt_rsc_0_2_clka_en,
      qb => yt_rsc_0_2_i_qb,
      web => yt_rsc_0_2_web,
      db => yt_rsc_0_2_i_db,
      adrb => yt_rsc_0_2_i_adrb,
      qa => yt_rsc_0_2_i_qa,
      wea => yt_rsc_0_2_wea,
      da => yt_rsc_0_2_i_da,
      adra => yt_rsc_0_2_i_adra,
      adra_d => yt_rsc_0_2_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_0_i_clka_en_d,
      clkb_en_d => yt_rsc_0_0_i_clka_en_d,
      da_d => yt_rsc_0_2_i_da_d_1,
      qa_d => yt_rsc_0_2_i_qa_d_1,
      wea_d => yt_rsc_0_2_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_2_i_qb <= yt_rsc_0_2_qb;
  yt_rsc_0_2_db <= yt_rsc_0_2_i_db;
  yt_rsc_0_2_adrb <= yt_rsc_0_2_i_adrb;
  yt_rsc_0_2_i_qa <= yt_rsc_0_2_qa;
  yt_rsc_0_2_da <= yt_rsc_0_2_i_da;
  yt_rsc_0_2_adra <= yt_rsc_0_2_i_adra;
  yt_rsc_0_2_i_adra_d_1 <= yt_rsc_0_2_i_adra_d;
  yt_rsc_0_2_i_da_d_1 <= yt_rsc_0_2_i_da_d;
  yt_rsc_0_2_i_qa_d <= yt_rsc_0_2_i_qa_d_1;
  yt_rsc_0_2_i_wea_d <= yt_rsc_0_0_i_wea_d_iff;
  yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_0_i_wea_d_iff;

  yt_rsc_0_3_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_10_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_3_clkb_en,
      clka_en => yt_rsc_0_3_clka_en,
      qb => yt_rsc_0_3_i_qb,
      web => yt_rsc_0_3_web,
      db => yt_rsc_0_3_i_db,
      adrb => yt_rsc_0_3_i_adrb,
      qa => yt_rsc_0_3_i_qa,
      wea => yt_rsc_0_3_wea,
      da => yt_rsc_0_3_i_da,
      adra => yt_rsc_0_3_i_adra,
      adra_d => yt_rsc_0_3_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_0_i_clka_en_d,
      clkb_en_d => yt_rsc_0_0_i_clka_en_d,
      da_d => yt_rsc_0_3_i_da_d_1,
      qa_d => yt_rsc_0_3_i_qa_d_1,
      wea_d => yt_rsc_0_3_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_3_i_qb <= yt_rsc_0_3_qb;
  yt_rsc_0_3_db <= yt_rsc_0_3_i_db;
  yt_rsc_0_3_adrb <= yt_rsc_0_3_i_adrb;
  yt_rsc_0_3_i_qa <= yt_rsc_0_3_qa;
  yt_rsc_0_3_da <= yt_rsc_0_3_i_da;
  yt_rsc_0_3_adra <= yt_rsc_0_3_i_adra;
  yt_rsc_0_3_i_adra_d_1 <= yt_rsc_0_3_i_adra_d;
  yt_rsc_0_3_i_da_d_1 <= yt_rsc_0_3_i_da_d;
  yt_rsc_0_3_i_qa_d <= yt_rsc_0_3_i_qa_d_1;
  yt_rsc_0_3_i_wea_d <= yt_rsc_0_0_i_wea_d_iff;
  yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_0_i_wea_d_iff;

  yt_rsc_0_4_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_11_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_4_clkb_en,
      clka_en => yt_rsc_0_4_clka_en,
      qb => yt_rsc_0_4_i_qb,
      web => yt_rsc_0_4_web,
      db => yt_rsc_0_4_i_db,
      adrb => yt_rsc_0_4_i_adrb,
      qa => yt_rsc_0_4_i_qa,
      wea => yt_rsc_0_4_wea,
      da => yt_rsc_0_4_i_da,
      adra => yt_rsc_0_4_i_adra,
      adra_d => yt_rsc_0_4_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_0_i_clka_en_d,
      clkb_en_d => yt_rsc_0_0_i_clka_en_d,
      da_d => yt_rsc_0_4_i_da_d_1,
      qa_d => yt_rsc_0_4_i_qa_d_1,
      wea_d => yt_rsc_0_4_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_4_i_qb <= yt_rsc_0_4_qb;
  yt_rsc_0_4_db <= yt_rsc_0_4_i_db;
  yt_rsc_0_4_adrb <= yt_rsc_0_4_i_adrb;
  yt_rsc_0_4_i_qa <= yt_rsc_0_4_qa;
  yt_rsc_0_4_da <= yt_rsc_0_4_i_da;
  yt_rsc_0_4_adra <= yt_rsc_0_4_i_adra;
  yt_rsc_0_4_i_adra_d_1 <= yt_rsc_0_4_i_adra_d;
  yt_rsc_0_4_i_da_d_1 <= yt_rsc_0_4_i_da_d;
  yt_rsc_0_4_i_qa_d <= yt_rsc_0_4_i_qa_d_1;
  yt_rsc_0_4_i_wea_d <= yt_rsc_0_0_i_wea_d_iff;
  yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_0_i_wea_d_iff;

  yt_rsc_0_5_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_12_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_5_clkb_en,
      clka_en => yt_rsc_0_5_clka_en,
      qb => yt_rsc_0_5_i_qb,
      web => yt_rsc_0_5_web,
      db => yt_rsc_0_5_i_db,
      adrb => yt_rsc_0_5_i_adrb,
      qa => yt_rsc_0_5_i_qa,
      wea => yt_rsc_0_5_wea,
      da => yt_rsc_0_5_i_da,
      adra => yt_rsc_0_5_i_adra,
      adra_d => yt_rsc_0_5_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_0_i_clka_en_d,
      clkb_en_d => yt_rsc_0_0_i_clka_en_d,
      da_d => yt_rsc_0_5_i_da_d_1,
      qa_d => yt_rsc_0_5_i_qa_d_1,
      wea_d => yt_rsc_0_5_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_5_i_qb <= yt_rsc_0_5_qb;
  yt_rsc_0_5_db <= yt_rsc_0_5_i_db;
  yt_rsc_0_5_adrb <= yt_rsc_0_5_i_adrb;
  yt_rsc_0_5_i_qa <= yt_rsc_0_5_qa;
  yt_rsc_0_5_da <= yt_rsc_0_5_i_da;
  yt_rsc_0_5_adra <= yt_rsc_0_5_i_adra;
  yt_rsc_0_5_i_adra_d_1 <= yt_rsc_0_5_i_adra_d;
  yt_rsc_0_5_i_da_d_1 <= yt_rsc_0_5_i_da_d;
  yt_rsc_0_5_i_qa_d <= yt_rsc_0_5_i_qa_d_1;
  yt_rsc_0_5_i_wea_d <= yt_rsc_0_0_i_wea_d_iff;
  yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_0_i_wea_d_iff;

  yt_rsc_0_6_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_13_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_6_clkb_en,
      clka_en => yt_rsc_0_6_clka_en,
      qb => yt_rsc_0_6_i_qb,
      web => yt_rsc_0_6_web,
      db => yt_rsc_0_6_i_db,
      adrb => yt_rsc_0_6_i_adrb,
      qa => yt_rsc_0_6_i_qa,
      wea => yt_rsc_0_6_wea,
      da => yt_rsc_0_6_i_da,
      adra => yt_rsc_0_6_i_adra,
      adra_d => yt_rsc_0_6_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_0_i_clka_en_d,
      clkb_en_d => yt_rsc_0_0_i_clka_en_d,
      da_d => yt_rsc_0_6_i_da_d_1,
      qa_d => yt_rsc_0_6_i_qa_d_1,
      wea_d => yt_rsc_0_6_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_6_i_qb <= yt_rsc_0_6_qb;
  yt_rsc_0_6_db <= yt_rsc_0_6_i_db;
  yt_rsc_0_6_adrb <= yt_rsc_0_6_i_adrb;
  yt_rsc_0_6_i_qa <= yt_rsc_0_6_qa;
  yt_rsc_0_6_da <= yt_rsc_0_6_i_da;
  yt_rsc_0_6_adra <= yt_rsc_0_6_i_adra;
  yt_rsc_0_6_i_adra_d_1 <= yt_rsc_0_6_i_adra_d;
  yt_rsc_0_6_i_da_d_1 <= yt_rsc_0_6_i_da_d;
  yt_rsc_0_6_i_qa_d <= yt_rsc_0_6_i_qa_d_1;
  yt_rsc_0_6_i_wea_d <= yt_rsc_0_0_i_wea_d_iff;
  yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_0_i_wea_d_iff;

  yt_rsc_0_7_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_14_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_7_clkb_en,
      clka_en => yt_rsc_0_7_clka_en,
      qb => yt_rsc_0_7_i_qb,
      web => yt_rsc_0_7_web,
      db => yt_rsc_0_7_i_db,
      adrb => yt_rsc_0_7_i_adrb,
      qa => yt_rsc_0_7_i_qa,
      wea => yt_rsc_0_7_wea,
      da => yt_rsc_0_7_i_da,
      adra => yt_rsc_0_7_i_adra,
      adra_d => yt_rsc_0_7_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_0_i_clka_en_d,
      clkb_en_d => yt_rsc_0_0_i_clka_en_d,
      da_d => yt_rsc_0_7_i_da_d_1,
      qa_d => yt_rsc_0_7_i_qa_d_1,
      wea_d => yt_rsc_0_7_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_7_i_qb <= yt_rsc_0_7_qb;
  yt_rsc_0_7_db <= yt_rsc_0_7_i_db;
  yt_rsc_0_7_adrb <= yt_rsc_0_7_i_adrb;
  yt_rsc_0_7_i_qa <= yt_rsc_0_7_qa;
  yt_rsc_0_7_da <= yt_rsc_0_7_i_da;
  yt_rsc_0_7_adra <= yt_rsc_0_7_i_adra;
  yt_rsc_0_7_i_adra_d_1 <= yt_rsc_0_7_i_adra_d;
  yt_rsc_0_7_i_da_d_1 <= yt_rsc_0_7_i_da_d;
  yt_rsc_0_7_i_qa_d <= yt_rsc_0_7_i_qa_d_1;
  yt_rsc_0_7_i_wea_d <= yt_rsc_0_0_i_wea_d_iff;
  yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_0_i_wea_d_iff;

  yt_rsc_0_8_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_15_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_8_clkb_en,
      clka_en => yt_rsc_0_8_clka_en,
      qb => yt_rsc_0_8_i_qb,
      web => yt_rsc_0_8_web,
      db => yt_rsc_0_8_i_db,
      adrb => yt_rsc_0_8_i_adrb,
      qa => yt_rsc_0_8_i_qa,
      wea => yt_rsc_0_8_wea,
      da => yt_rsc_0_8_i_da,
      adra => yt_rsc_0_8_i_adra,
      adra_d => yt_rsc_0_8_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_0_i_clka_en_d,
      clkb_en_d => yt_rsc_0_0_i_clka_en_d,
      da_d => yt_rsc_0_8_i_da_d_1,
      qa_d => yt_rsc_0_8_i_qa_d_1,
      wea_d => yt_rsc_0_8_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_8_i_qb <= yt_rsc_0_8_qb;
  yt_rsc_0_8_db <= yt_rsc_0_8_i_db;
  yt_rsc_0_8_adrb <= yt_rsc_0_8_i_adrb;
  yt_rsc_0_8_i_qa <= yt_rsc_0_8_qa;
  yt_rsc_0_8_da <= yt_rsc_0_8_i_da;
  yt_rsc_0_8_adra <= yt_rsc_0_8_i_adra;
  yt_rsc_0_8_i_adra_d_1 <= yt_rsc_0_8_i_adra_d;
  yt_rsc_0_8_i_da_d_1 <= yt_rsc_0_8_i_da_d;
  yt_rsc_0_8_i_qa_d <= yt_rsc_0_8_i_qa_d_1;
  yt_rsc_0_8_i_wea_d <= yt_rsc_0_0_i_wea_d_iff;
  yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_0_i_wea_d_iff;

  yt_rsc_0_9_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_16_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_9_clkb_en,
      clka_en => yt_rsc_0_9_clka_en,
      qb => yt_rsc_0_9_i_qb,
      web => yt_rsc_0_9_web,
      db => yt_rsc_0_9_i_db,
      adrb => yt_rsc_0_9_i_adrb,
      qa => yt_rsc_0_9_i_qa,
      wea => yt_rsc_0_9_wea,
      da => yt_rsc_0_9_i_da,
      adra => yt_rsc_0_9_i_adra,
      adra_d => yt_rsc_0_9_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_0_i_clka_en_d,
      clkb_en_d => yt_rsc_0_0_i_clka_en_d,
      da_d => yt_rsc_0_9_i_da_d_1,
      qa_d => yt_rsc_0_9_i_qa_d_1,
      wea_d => yt_rsc_0_9_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_9_i_qb <= yt_rsc_0_9_qb;
  yt_rsc_0_9_db <= yt_rsc_0_9_i_db;
  yt_rsc_0_9_adrb <= yt_rsc_0_9_i_adrb;
  yt_rsc_0_9_i_qa <= yt_rsc_0_9_qa;
  yt_rsc_0_9_da <= yt_rsc_0_9_i_da;
  yt_rsc_0_9_adra <= yt_rsc_0_9_i_adra;
  yt_rsc_0_9_i_adra_d_1 <= yt_rsc_0_9_i_adra_d;
  yt_rsc_0_9_i_da_d_1 <= yt_rsc_0_9_i_da_d;
  yt_rsc_0_9_i_qa_d <= yt_rsc_0_9_i_qa_d_1;
  yt_rsc_0_9_i_wea_d <= yt_rsc_0_0_i_wea_d_iff;
  yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_0_i_wea_d_iff;

  yt_rsc_0_10_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_17_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_10_clkb_en,
      clka_en => yt_rsc_0_10_clka_en,
      qb => yt_rsc_0_10_i_qb,
      web => yt_rsc_0_10_web,
      db => yt_rsc_0_10_i_db,
      adrb => yt_rsc_0_10_i_adrb,
      qa => yt_rsc_0_10_i_qa,
      wea => yt_rsc_0_10_wea,
      da => yt_rsc_0_10_i_da,
      adra => yt_rsc_0_10_i_adra,
      adra_d => yt_rsc_0_10_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_0_i_clka_en_d,
      clkb_en_d => yt_rsc_0_0_i_clka_en_d,
      da_d => yt_rsc_0_10_i_da_d_1,
      qa_d => yt_rsc_0_10_i_qa_d_1,
      wea_d => yt_rsc_0_10_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_10_i_qb <= yt_rsc_0_10_qb;
  yt_rsc_0_10_db <= yt_rsc_0_10_i_db;
  yt_rsc_0_10_adrb <= yt_rsc_0_10_i_adrb;
  yt_rsc_0_10_i_qa <= yt_rsc_0_10_qa;
  yt_rsc_0_10_da <= yt_rsc_0_10_i_da;
  yt_rsc_0_10_adra <= yt_rsc_0_10_i_adra;
  yt_rsc_0_10_i_adra_d_1 <= yt_rsc_0_10_i_adra_d;
  yt_rsc_0_10_i_da_d_1 <= yt_rsc_0_10_i_da_d;
  yt_rsc_0_10_i_qa_d <= yt_rsc_0_10_i_qa_d_1;
  yt_rsc_0_10_i_wea_d <= yt_rsc_0_0_i_wea_d_iff;
  yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_0_i_wea_d_iff;

  yt_rsc_0_11_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_18_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_11_clkb_en,
      clka_en => yt_rsc_0_11_clka_en,
      qb => yt_rsc_0_11_i_qb,
      web => yt_rsc_0_11_web,
      db => yt_rsc_0_11_i_db,
      adrb => yt_rsc_0_11_i_adrb,
      qa => yt_rsc_0_11_i_qa,
      wea => yt_rsc_0_11_wea,
      da => yt_rsc_0_11_i_da,
      adra => yt_rsc_0_11_i_adra,
      adra_d => yt_rsc_0_11_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_0_i_clka_en_d,
      clkb_en_d => yt_rsc_0_0_i_clka_en_d,
      da_d => yt_rsc_0_11_i_da_d_1,
      qa_d => yt_rsc_0_11_i_qa_d_1,
      wea_d => yt_rsc_0_11_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_11_i_qb <= yt_rsc_0_11_qb;
  yt_rsc_0_11_db <= yt_rsc_0_11_i_db;
  yt_rsc_0_11_adrb <= yt_rsc_0_11_i_adrb;
  yt_rsc_0_11_i_qa <= yt_rsc_0_11_qa;
  yt_rsc_0_11_da <= yt_rsc_0_11_i_da;
  yt_rsc_0_11_adra <= yt_rsc_0_11_i_adra;
  yt_rsc_0_11_i_adra_d_1 <= yt_rsc_0_11_i_adra_d;
  yt_rsc_0_11_i_da_d_1 <= yt_rsc_0_11_i_da_d;
  yt_rsc_0_11_i_qa_d <= yt_rsc_0_11_i_qa_d_1;
  yt_rsc_0_11_i_wea_d <= yt_rsc_0_0_i_wea_d_iff;
  yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_0_i_wea_d_iff;

  yt_rsc_0_12_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_19_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_12_clkb_en,
      clka_en => yt_rsc_0_12_clka_en,
      qb => yt_rsc_0_12_i_qb,
      web => yt_rsc_0_12_web,
      db => yt_rsc_0_12_i_db,
      adrb => yt_rsc_0_12_i_adrb,
      qa => yt_rsc_0_12_i_qa,
      wea => yt_rsc_0_12_wea,
      da => yt_rsc_0_12_i_da,
      adra => yt_rsc_0_12_i_adra,
      adra_d => yt_rsc_0_12_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_0_i_clka_en_d,
      clkb_en_d => yt_rsc_0_0_i_clka_en_d,
      da_d => yt_rsc_0_12_i_da_d_1,
      qa_d => yt_rsc_0_12_i_qa_d_1,
      wea_d => yt_rsc_0_12_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_12_i_qb <= yt_rsc_0_12_qb;
  yt_rsc_0_12_db <= yt_rsc_0_12_i_db;
  yt_rsc_0_12_adrb <= yt_rsc_0_12_i_adrb;
  yt_rsc_0_12_i_qa <= yt_rsc_0_12_qa;
  yt_rsc_0_12_da <= yt_rsc_0_12_i_da;
  yt_rsc_0_12_adra <= yt_rsc_0_12_i_adra;
  yt_rsc_0_12_i_adra_d_1 <= yt_rsc_0_12_i_adra_d;
  yt_rsc_0_12_i_da_d_1 <= yt_rsc_0_12_i_da_d;
  yt_rsc_0_12_i_qa_d <= yt_rsc_0_12_i_qa_d_1;
  yt_rsc_0_12_i_wea_d <= yt_rsc_0_0_i_wea_d_iff;
  yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_0_i_wea_d_iff;

  yt_rsc_0_13_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_20_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_13_clkb_en,
      clka_en => yt_rsc_0_13_clka_en,
      qb => yt_rsc_0_13_i_qb,
      web => yt_rsc_0_13_web,
      db => yt_rsc_0_13_i_db,
      adrb => yt_rsc_0_13_i_adrb,
      qa => yt_rsc_0_13_i_qa,
      wea => yt_rsc_0_13_wea,
      da => yt_rsc_0_13_i_da,
      adra => yt_rsc_0_13_i_adra,
      adra_d => yt_rsc_0_13_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_0_i_clka_en_d,
      clkb_en_d => yt_rsc_0_0_i_clka_en_d,
      da_d => yt_rsc_0_13_i_da_d_1,
      qa_d => yt_rsc_0_13_i_qa_d_1,
      wea_d => yt_rsc_0_13_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_13_i_qb <= yt_rsc_0_13_qb;
  yt_rsc_0_13_db <= yt_rsc_0_13_i_db;
  yt_rsc_0_13_adrb <= yt_rsc_0_13_i_adrb;
  yt_rsc_0_13_i_qa <= yt_rsc_0_13_qa;
  yt_rsc_0_13_da <= yt_rsc_0_13_i_da;
  yt_rsc_0_13_adra <= yt_rsc_0_13_i_adra;
  yt_rsc_0_13_i_adra_d_1 <= yt_rsc_0_13_i_adra_d;
  yt_rsc_0_13_i_da_d_1 <= yt_rsc_0_13_i_da_d;
  yt_rsc_0_13_i_qa_d <= yt_rsc_0_13_i_qa_d_1;
  yt_rsc_0_13_i_wea_d <= yt_rsc_0_0_i_wea_d_iff;
  yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_0_i_wea_d_iff;

  yt_rsc_0_14_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_21_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_14_clkb_en,
      clka_en => yt_rsc_0_14_clka_en,
      qb => yt_rsc_0_14_i_qb,
      web => yt_rsc_0_14_web,
      db => yt_rsc_0_14_i_db,
      adrb => yt_rsc_0_14_i_adrb,
      qa => yt_rsc_0_14_i_qa,
      wea => yt_rsc_0_14_wea,
      da => yt_rsc_0_14_i_da,
      adra => yt_rsc_0_14_i_adra,
      adra_d => yt_rsc_0_14_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_0_i_clka_en_d,
      clkb_en_d => yt_rsc_0_0_i_clka_en_d,
      da_d => yt_rsc_0_14_i_da_d_1,
      qa_d => yt_rsc_0_14_i_qa_d_1,
      wea_d => yt_rsc_0_14_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_14_i_qb <= yt_rsc_0_14_qb;
  yt_rsc_0_14_db <= yt_rsc_0_14_i_db;
  yt_rsc_0_14_adrb <= yt_rsc_0_14_i_adrb;
  yt_rsc_0_14_i_qa <= yt_rsc_0_14_qa;
  yt_rsc_0_14_da <= yt_rsc_0_14_i_da;
  yt_rsc_0_14_adra <= yt_rsc_0_14_i_adra;
  yt_rsc_0_14_i_adra_d_1 <= yt_rsc_0_14_i_adra_d;
  yt_rsc_0_14_i_da_d_1 <= yt_rsc_0_14_i_da_d;
  yt_rsc_0_14_i_qa_d <= yt_rsc_0_14_i_qa_d_1;
  yt_rsc_0_14_i_wea_d <= yt_rsc_0_0_i_wea_d_iff;
  yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_0_i_wea_d_iff;

  yt_rsc_0_15_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_22_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_15_clkb_en,
      clka_en => yt_rsc_0_15_clka_en,
      qb => yt_rsc_0_15_i_qb,
      web => yt_rsc_0_15_web,
      db => yt_rsc_0_15_i_db,
      adrb => yt_rsc_0_15_i_adrb,
      qa => yt_rsc_0_15_i_qa,
      wea => yt_rsc_0_15_wea,
      da => yt_rsc_0_15_i_da,
      adra => yt_rsc_0_15_i_adra,
      adra_d => yt_rsc_0_15_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_0_i_clka_en_d,
      clkb_en_d => yt_rsc_0_0_i_clka_en_d,
      da_d => yt_rsc_0_15_i_da_d_1,
      qa_d => yt_rsc_0_15_i_qa_d_1,
      wea_d => yt_rsc_0_15_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_15_i_qb <= yt_rsc_0_15_qb;
  yt_rsc_0_15_db <= yt_rsc_0_15_i_db;
  yt_rsc_0_15_adrb <= yt_rsc_0_15_i_adrb;
  yt_rsc_0_15_i_qa <= yt_rsc_0_15_qa;
  yt_rsc_0_15_da <= yt_rsc_0_15_i_da;
  yt_rsc_0_15_adra <= yt_rsc_0_15_i_adra;
  yt_rsc_0_15_i_adra_d_1 <= yt_rsc_0_15_i_adra_d;
  yt_rsc_0_15_i_da_d_1 <= yt_rsc_0_15_i_da_d;
  yt_rsc_0_15_i_qa_d <= yt_rsc_0_15_i_qa_d_1;
  yt_rsc_0_15_i_wea_d <= yt_rsc_0_0_i_wea_d_iff;
  yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_0_i_wea_d_iff;

  yt_rsc_0_16_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_23_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_16_clkb_en,
      clka_en => yt_rsc_0_16_clka_en,
      qb => yt_rsc_0_16_i_qb,
      web => yt_rsc_0_16_web,
      db => yt_rsc_0_16_i_db,
      adrb => yt_rsc_0_16_i_adrb,
      qa => yt_rsc_0_16_i_qa,
      wea => yt_rsc_0_16_wea,
      da => yt_rsc_0_16_i_da,
      adra => yt_rsc_0_16_i_adra,
      adra_d => yt_rsc_0_16_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_16_i_clka_en_d,
      clkb_en_d => yt_rsc_0_16_i_clka_en_d,
      da_d => yt_rsc_0_16_i_da_d_1,
      qa_d => yt_rsc_0_16_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_16_i_qb <= yt_rsc_0_16_qb;
  yt_rsc_0_16_db <= yt_rsc_0_16_i_db;
  yt_rsc_0_16_adrb <= yt_rsc_0_16_i_adrb;
  yt_rsc_0_16_i_qa <= yt_rsc_0_16_qa;
  yt_rsc_0_16_da <= yt_rsc_0_16_i_da;
  yt_rsc_0_16_adra <= yt_rsc_0_16_i_adra;
  yt_rsc_0_16_i_adra_d_1 <= yt_rsc_0_16_i_adra_d;
  yt_rsc_0_16_i_da_d_1 <= yt_rsc_0_16_i_da_d;
  yt_rsc_0_16_i_qa_d <= yt_rsc_0_16_i_qa_d_1;
  yt_rsc_0_16_i_wea_d <= yt_rsc_0_16_i_wea_d_iff;
  yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_16_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_16_i_wea_d_iff;

  yt_rsc_0_17_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_24_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_17_clkb_en,
      clka_en => yt_rsc_0_17_clka_en,
      qb => yt_rsc_0_17_i_qb,
      web => yt_rsc_0_17_web,
      db => yt_rsc_0_17_i_db,
      adrb => yt_rsc_0_17_i_adrb,
      qa => yt_rsc_0_17_i_qa,
      wea => yt_rsc_0_17_wea,
      da => yt_rsc_0_17_i_da,
      adra => yt_rsc_0_17_i_adra,
      adra_d => yt_rsc_0_17_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_16_i_clka_en_d,
      clkb_en_d => yt_rsc_0_16_i_clka_en_d,
      da_d => yt_rsc_0_17_i_da_d_1,
      qa_d => yt_rsc_0_17_i_qa_d_1,
      wea_d => yt_rsc_0_17_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_17_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_17_i_qb <= yt_rsc_0_17_qb;
  yt_rsc_0_17_db <= yt_rsc_0_17_i_db;
  yt_rsc_0_17_adrb <= yt_rsc_0_17_i_adrb;
  yt_rsc_0_17_i_qa <= yt_rsc_0_17_qa;
  yt_rsc_0_17_da <= yt_rsc_0_17_i_da;
  yt_rsc_0_17_adra <= yt_rsc_0_17_i_adra;
  yt_rsc_0_17_i_adra_d_1 <= yt_rsc_0_17_i_adra_d;
  yt_rsc_0_17_i_da_d_1 <= yt_rsc_0_17_i_da_d;
  yt_rsc_0_17_i_qa_d <= yt_rsc_0_17_i_qa_d_1;
  yt_rsc_0_17_i_wea_d <= yt_rsc_0_16_i_wea_d_iff;
  yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_17_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_16_i_wea_d_iff;

  yt_rsc_0_18_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_25_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_18_clkb_en,
      clka_en => yt_rsc_0_18_clka_en,
      qb => yt_rsc_0_18_i_qb,
      web => yt_rsc_0_18_web,
      db => yt_rsc_0_18_i_db,
      adrb => yt_rsc_0_18_i_adrb,
      qa => yt_rsc_0_18_i_qa,
      wea => yt_rsc_0_18_wea,
      da => yt_rsc_0_18_i_da,
      adra => yt_rsc_0_18_i_adra,
      adra_d => yt_rsc_0_18_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_16_i_clka_en_d,
      clkb_en_d => yt_rsc_0_16_i_clka_en_d,
      da_d => yt_rsc_0_18_i_da_d_1,
      qa_d => yt_rsc_0_18_i_qa_d_1,
      wea_d => yt_rsc_0_18_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_18_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_18_i_qb <= yt_rsc_0_18_qb;
  yt_rsc_0_18_db <= yt_rsc_0_18_i_db;
  yt_rsc_0_18_adrb <= yt_rsc_0_18_i_adrb;
  yt_rsc_0_18_i_qa <= yt_rsc_0_18_qa;
  yt_rsc_0_18_da <= yt_rsc_0_18_i_da;
  yt_rsc_0_18_adra <= yt_rsc_0_18_i_adra;
  yt_rsc_0_18_i_adra_d_1 <= yt_rsc_0_18_i_adra_d;
  yt_rsc_0_18_i_da_d_1 <= yt_rsc_0_18_i_da_d;
  yt_rsc_0_18_i_qa_d <= yt_rsc_0_18_i_qa_d_1;
  yt_rsc_0_18_i_wea_d <= yt_rsc_0_16_i_wea_d_iff;
  yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_18_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_16_i_wea_d_iff;

  yt_rsc_0_19_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_26_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_19_clkb_en,
      clka_en => yt_rsc_0_19_clka_en,
      qb => yt_rsc_0_19_i_qb,
      web => yt_rsc_0_19_web,
      db => yt_rsc_0_19_i_db,
      adrb => yt_rsc_0_19_i_adrb,
      qa => yt_rsc_0_19_i_qa,
      wea => yt_rsc_0_19_wea,
      da => yt_rsc_0_19_i_da,
      adra => yt_rsc_0_19_i_adra,
      adra_d => yt_rsc_0_19_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_16_i_clka_en_d,
      clkb_en_d => yt_rsc_0_16_i_clka_en_d,
      da_d => yt_rsc_0_19_i_da_d_1,
      qa_d => yt_rsc_0_19_i_qa_d_1,
      wea_d => yt_rsc_0_19_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_19_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_19_i_qb <= yt_rsc_0_19_qb;
  yt_rsc_0_19_db <= yt_rsc_0_19_i_db;
  yt_rsc_0_19_adrb <= yt_rsc_0_19_i_adrb;
  yt_rsc_0_19_i_qa <= yt_rsc_0_19_qa;
  yt_rsc_0_19_da <= yt_rsc_0_19_i_da;
  yt_rsc_0_19_adra <= yt_rsc_0_19_i_adra;
  yt_rsc_0_19_i_adra_d_1 <= yt_rsc_0_19_i_adra_d;
  yt_rsc_0_19_i_da_d_1 <= yt_rsc_0_19_i_da_d;
  yt_rsc_0_19_i_qa_d <= yt_rsc_0_19_i_qa_d_1;
  yt_rsc_0_19_i_wea_d <= yt_rsc_0_16_i_wea_d_iff;
  yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_19_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_16_i_wea_d_iff;

  yt_rsc_0_20_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_27_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_20_clkb_en,
      clka_en => yt_rsc_0_20_clka_en,
      qb => yt_rsc_0_20_i_qb,
      web => yt_rsc_0_20_web,
      db => yt_rsc_0_20_i_db,
      adrb => yt_rsc_0_20_i_adrb,
      qa => yt_rsc_0_20_i_qa,
      wea => yt_rsc_0_20_wea,
      da => yt_rsc_0_20_i_da,
      adra => yt_rsc_0_20_i_adra,
      adra_d => yt_rsc_0_20_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_16_i_clka_en_d,
      clkb_en_d => yt_rsc_0_16_i_clka_en_d,
      da_d => yt_rsc_0_20_i_da_d_1,
      qa_d => yt_rsc_0_20_i_qa_d_1,
      wea_d => yt_rsc_0_20_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_20_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_20_i_qb <= yt_rsc_0_20_qb;
  yt_rsc_0_20_db <= yt_rsc_0_20_i_db;
  yt_rsc_0_20_adrb <= yt_rsc_0_20_i_adrb;
  yt_rsc_0_20_i_qa <= yt_rsc_0_20_qa;
  yt_rsc_0_20_da <= yt_rsc_0_20_i_da;
  yt_rsc_0_20_adra <= yt_rsc_0_20_i_adra;
  yt_rsc_0_20_i_adra_d_1 <= yt_rsc_0_20_i_adra_d;
  yt_rsc_0_20_i_da_d_1 <= yt_rsc_0_20_i_da_d;
  yt_rsc_0_20_i_qa_d <= yt_rsc_0_20_i_qa_d_1;
  yt_rsc_0_20_i_wea_d <= yt_rsc_0_16_i_wea_d_iff;
  yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_20_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_16_i_wea_d_iff;

  yt_rsc_0_21_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_28_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_21_clkb_en,
      clka_en => yt_rsc_0_21_clka_en,
      qb => yt_rsc_0_21_i_qb,
      web => yt_rsc_0_21_web,
      db => yt_rsc_0_21_i_db,
      adrb => yt_rsc_0_21_i_adrb,
      qa => yt_rsc_0_21_i_qa,
      wea => yt_rsc_0_21_wea,
      da => yt_rsc_0_21_i_da,
      adra => yt_rsc_0_21_i_adra,
      adra_d => yt_rsc_0_21_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_16_i_clka_en_d,
      clkb_en_d => yt_rsc_0_16_i_clka_en_d,
      da_d => yt_rsc_0_21_i_da_d_1,
      qa_d => yt_rsc_0_21_i_qa_d_1,
      wea_d => yt_rsc_0_21_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_21_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_21_i_qb <= yt_rsc_0_21_qb;
  yt_rsc_0_21_db <= yt_rsc_0_21_i_db;
  yt_rsc_0_21_adrb <= yt_rsc_0_21_i_adrb;
  yt_rsc_0_21_i_qa <= yt_rsc_0_21_qa;
  yt_rsc_0_21_da <= yt_rsc_0_21_i_da;
  yt_rsc_0_21_adra <= yt_rsc_0_21_i_adra;
  yt_rsc_0_21_i_adra_d_1 <= yt_rsc_0_21_i_adra_d;
  yt_rsc_0_21_i_da_d_1 <= yt_rsc_0_21_i_da_d;
  yt_rsc_0_21_i_qa_d <= yt_rsc_0_21_i_qa_d_1;
  yt_rsc_0_21_i_wea_d <= yt_rsc_0_16_i_wea_d_iff;
  yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_21_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_16_i_wea_d_iff;

  yt_rsc_0_22_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_29_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_22_clkb_en,
      clka_en => yt_rsc_0_22_clka_en,
      qb => yt_rsc_0_22_i_qb,
      web => yt_rsc_0_22_web,
      db => yt_rsc_0_22_i_db,
      adrb => yt_rsc_0_22_i_adrb,
      qa => yt_rsc_0_22_i_qa,
      wea => yt_rsc_0_22_wea,
      da => yt_rsc_0_22_i_da,
      adra => yt_rsc_0_22_i_adra,
      adra_d => yt_rsc_0_22_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_16_i_clka_en_d,
      clkb_en_d => yt_rsc_0_16_i_clka_en_d,
      da_d => yt_rsc_0_22_i_da_d_1,
      qa_d => yt_rsc_0_22_i_qa_d_1,
      wea_d => yt_rsc_0_22_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_22_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_22_i_qb <= yt_rsc_0_22_qb;
  yt_rsc_0_22_db <= yt_rsc_0_22_i_db;
  yt_rsc_0_22_adrb <= yt_rsc_0_22_i_adrb;
  yt_rsc_0_22_i_qa <= yt_rsc_0_22_qa;
  yt_rsc_0_22_da <= yt_rsc_0_22_i_da;
  yt_rsc_0_22_adra <= yt_rsc_0_22_i_adra;
  yt_rsc_0_22_i_adra_d_1 <= yt_rsc_0_22_i_adra_d;
  yt_rsc_0_22_i_da_d_1 <= yt_rsc_0_22_i_da_d;
  yt_rsc_0_22_i_qa_d <= yt_rsc_0_22_i_qa_d_1;
  yt_rsc_0_22_i_wea_d <= yt_rsc_0_16_i_wea_d_iff;
  yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_22_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_16_i_wea_d_iff;

  yt_rsc_0_23_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_30_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_23_clkb_en,
      clka_en => yt_rsc_0_23_clka_en,
      qb => yt_rsc_0_23_i_qb,
      web => yt_rsc_0_23_web,
      db => yt_rsc_0_23_i_db,
      adrb => yt_rsc_0_23_i_adrb,
      qa => yt_rsc_0_23_i_qa,
      wea => yt_rsc_0_23_wea,
      da => yt_rsc_0_23_i_da,
      adra => yt_rsc_0_23_i_adra,
      adra_d => yt_rsc_0_23_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_16_i_clka_en_d,
      clkb_en_d => yt_rsc_0_16_i_clka_en_d,
      da_d => yt_rsc_0_23_i_da_d_1,
      qa_d => yt_rsc_0_23_i_qa_d_1,
      wea_d => yt_rsc_0_23_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_23_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_23_i_qb <= yt_rsc_0_23_qb;
  yt_rsc_0_23_db <= yt_rsc_0_23_i_db;
  yt_rsc_0_23_adrb <= yt_rsc_0_23_i_adrb;
  yt_rsc_0_23_i_qa <= yt_rsc_0_23_qa;
  yt_rsc_0_23_da <= yt_rsc_0_23_i_da;
  yt_rsc_0_23_adra <= yt_rsc_0_23_i_adra;
  yt_rsc_0_23_i_adra_d_1 <= yt_rsc_0_23_i_adra_d;
  yt_rsc_0_23_i_da_d_1 <= yt_rsc_0_23_i_da_d;
  yt_rsc_0_23_i_qa_d <= yt_rsc_0_23_i_qa_d_1;
  yt_rsc_0_23_i_wea_d <= yt_rsc_0_16_i_wea_d_iff;
  yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_23_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_16_i_wea_d_iff;

  yt_rsc_0_24_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_31_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_24_clkb_en,
      clka_en => yt_rsc_0_24_clka_en,
      qb => yt_rsc_0_24_i_qb,
      web => yt_rsc_0_24_web,
      db => yt_rsc_0_24_i_db,
      adrb => yt_rsc_0_24_i_adrb,
      qa => yt_rsc_0_24_i_qa,
      wea => yt_rsc_0_24_wea,
      da => yt_rsc_0_24_i_da,
      adra => yt_rsc_0_24_i_adra,
      adra_d => yt_rsc_0_24_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_16_i_clka_en_d,
      clkb_en_d => yt_rsc_0_16_i_clka_en_d,
      da_d => yt_rsc_0_24_i_da_d_1,
      qa_d => yt_rsc_0_24_i_qa_d_1,
      wea_d => yt_rsc_0_24_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_24_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_24_i_qb <= yt_rsc_0_24_qb;
  yt_rsc_0_24_db <= yt_rsc_0_24_i_db;
  yt_rsc_0_24_adrb <= yt_rsc_0_24_i_adrb;
  yt_rsc_0_24_i_qa <= yt_rsc_0_24_qa;
  yt_rsc_0_24_da <= yt_rsc_0_24_i_da;
  yt_rsc_0_24_adra <= yt_rsc_0_24_i_adra;
  yt_rsc_0_24_i_adra_d_1 <= yt_rsc_0_24_i_adra_d;
  yt_rsc_0_24_i_da_d_1 <= yt_rsc_0_24_i_da_d;
  yt_rsc_0_24_i_qa_d <= yt_rsc_0_24_i_qa_d_1;
  yt_rsc_0_24_i_wea_d <= yt_rsc_0_16_i_wea_d_iff;
  yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_24_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_16_i_wea_d_iff;

  yt_rsc_0_25_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_32_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_25_clkb_en,
      clka_en => yt_rsc_0_25_clka_en,
      qb => yt_rsc_0_25_i_qb,
      web => yt_rsc_0_25_web,
      db => yt_rsc_0_25_i_db,
      adrb => yt_rsc_0_25_i_adrb,
      qa => yt_rsc_0_25_i_qa,
      wea => yt_rsc_0_25_wea,
      da => yt_rsc_0_25_i_da,
      adra => yt_rsc_0_25_i_adra,
      adra_d => yt_rsc_0_25_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_16_i_clka_en_d,
      clkb_en_d => yt_rsc_0_16_i_clka_en_d,
      da_d => yt_rsc_0_25_i_da_d_1,
      qa_d => yt_rsc_0_25_i_qa_d_1,
      wea_d => yt_rsc_0_25_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_25_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_25_i_qb <= yt_rsc_0_25_qb;
  yt_rsc_0_25_db <= yt_rsc_0_25_i_db;
  yt_rsc_0_25_adrb <= yt_rsc_0_25_i_adrb;
  yt_rsc_0_25_i_qa <= yt_rsc_0_25_qa;
  yt_rsc_0_25_da <= yt_rsc_0_25_i_da;
  yt_rsc_0_25_adra <= yt_rsc_0_25_i_adra;
  yt_rsc_0_25_i_adra_d_1 <= yt_rsc_0_25_i_adra_d;
  yt_rsc_0_25_i_da_d_1 <= yt_rsc_0_25_i_da_d;
  yt_rsc_0_25_i_qa_d <= yt_rsc_0_25_i_qa_d_1;
  yt_rsc_0_25_i_wea_d <= yt_rsc_0_16_i_wea_d_iff;
  yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_25_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_16_i_wea_d_iff;

  yt_rsc_0_26_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_33_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_26_clkb_en,
      clka_en => yt_rsc_0_26_clka_en,
      qb => yt_rsc_0_26_i_qb,
      web => yt_rsc_0_26_web,
      db => yt_rsc_0_26_i_db,
      adrb => yt_rsc_0_26_i_adrb,
      qa => yt_rsc_0_26_i_qa,
      wea => yt_rsc_0_26_wea,
      da => yt_rsc_0_26_i_da,
      adra => yt_rsc_0_26_i_adra,
      adra_d => yt_rsc_0_26_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_16_i_clka_en_d,
      clkb_en_d => yt_rsc_0_16_i_clka_en_d,
      da_d => yt_rsc_0_26_i_da_d_1,
      qa_d => yt_rsc_0_26_i_qa_d_1,
      wea_d => yt_rsc_0_26_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_26_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_26_i_qb <= yt_rsc_0_26_qb;
  yt_rsc_0_26_db <= yt_rsc_0_26_i_db;
  yt_rsc_0_26_adrb <= yt_rsc_0_26_i_adrb;
  yt_rsc_0_26_i_qa <= yt_rsc_0_26_qa;
  yt_rsc_0_26_da <= yt_rsc_0_26_i_da;
  yt_rsc_0_26_adra <= yt_rsc_0_26_i_adra;
  yt_rsc_0_26_i_adra_d_1 <= yt_rsc_0_26_i_adra_d;
  yt_rsc_0_26_i_da_d_1 <= yt_rsc_0_26_i_da_d;
  yt_rsc_0_26_i_qa_d <= yt_rsc_0_26_i_qa_d_1;
  yt_rsc_0_26_i_wea_d <= yt_rsc_0_16_i_wea_d_iff;
  yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_26_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_16_i_wea_d_iff;

  yt_rsc_0_27_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_34_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_27_clkb_en,
      clka_en => yt_rsc_0_27_clka_en,
      qb => yt_rsc_0_27_i_qb,
      web => yt_rsc_0_27_web,
      db => yt_rsc_0_27_i_db,
      adrb => yt_rsc_0_27_i_adrb,
      qa => yt_rsc_0_27_i_qa,
      wea => yt_rsc_0_27_wea,
      da => yt_rsc_0_27_i_da,
      adra => yt_rsc_0_27_i_adra,
      adra_d => yt_rsc_0_27_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_16_i_clka_en_d,
      clkb_en_d => yt_rsc_0_16_i_clka_en_d,
      da_d => yt_rsc_0_27_i_da_d_1,
      qa_d => yt_rsc_0_27_i_qa_d_1,
      wea_d => yt_rsc_0_27_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_27_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_27_i_qb <= yt_rsc_0_27_qb;
  yt_rsc_0_27_db <= yt_rsc_0_27_i_db;
  yt_rsc_0_27_adrb <= yt_rsc_0_27_i_adrb;
  yt_rsc_0_27_i_qa <= yt_rsc_0_27_qa;
  yt_rsc_0_27_da <= yt_rsc_0_27_i_da;
  yt_rsc_0_27_adra <= yt_rsc_0_27_i_adra;
  yt_rsc_0_27_i_adra_d_1 <= yt_rsc_0_27_i_adra_d;
  yt_rsc_0_27_i_da_d_1 <= yt_rsc_0_27_i_da_d;
  yt_rsc_0_27_i_qa_d <= yt_rsc_0_27_i_qa_d_1;
  yt_rsc_0_27_i_wea_d <= yt_rsc_0_16_i_wea_d_iff;
  yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_27_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_16_i_wea_d_iff;

  yt_rsc_0_28_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_35_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_28_clkb_en,
      clka_en => yt_rsc_0_28_clka_en,
      qb => yt_rsc_0_28_i_qb,
      web => yt_rsc_0_28_web,
      db => yt_rsc_0_28_i_db,
      adrb => yt_rsc_0_28_i_adrb,
      qa => yt_rsc_0_28_i_qa,
      wea => yt_rsc_0_28_wea,
      da => yt_rsc_0_28_i_da,
      adra => yt_rsc_0_28_i_adra,
      adra_d => yt_rsc_0_28_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_16_i_clka_en_d,
      clkb_en_d => yt_rsc_0_16_i_clka_en_d,
      da_d => yt_rsc_0_28_i_da_d_1,
      qa_d => yt_rsc_0_28_i_qa_d_1,
      wea_d => yt_rsc_0_28_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_28_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_28_i_qb <= yt_rsc_0_28_qb;
  yt_rsc_0_28_db <= yt_rsc_0_28_i_db;
  yt_rsc_0_28_adrb <= yt_rsc_0_28_i_adrb;
  yt_rsc_0_28_i_qa <= yt_rsc_0_28_qa;
  yt_rsc_0_28_da <= yt_rsc_0_28_i_da;
  yt_rsc_0_28_adra <= yt_rsc_0_28_i_adra;
  yt_rsc_0_28_i_adra_d_1 <= yt_rsc_0_28_i_adra_d;
  yt_rsc_0_28_i_da_d_1 <= yt_rsc_0_28_i_da_d;
  yt_rsc_0_28_i_qa_d <= yt_rsc_0_28_i_qa_d_1;
  yt_rsc_0_28_i_wea_d <= yt_rsc_0_16_i_wea_d_iff;
  yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_28_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_16_i_wea_d_iff;

  yt_rsc_0_29_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_36_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_29_clkb_en,
      clka_en => yt_rsc_0_29_clka_en,
      qb => yt_rsc_0_29_i_qb,
      web => yt_rsc_0_29_web,
      db => yt_rsc_0_29_i_db,
      adrb => yt_rsc_0_29_i_adrb,
      qa => yt_rsc_0_29_i_qa,
      wea => yt_rsc_0_29_wea,
      da => yt_rsc_0_29_i_da,
      adra => yt_rsc_0_29_i_adra,
      adra_d => yt_rsc_0_29_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_16_i_clka_en_d,
      clkb_en_d => yt_rsc_0_16_i_clka_en_d,
      da_d => yt_rsc_0_29_i_da_d_1,
      qa_d => yt_rsc_0_29_i_qa_d_1,
      wea_d => yt_rsc_0_29_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_29_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_29_i_qb <= yt_rsc_0_29_qb;
  yt_rsc_0_29_db <= yt_rsc_0_29_i_db;
  yt_rsc_0_29_adrb <= yt_rsc_0_29_i_adrb;
  yt_rsc_0_29_i_qa <= yt_rsc_0_29_qa;
  yt_rsc_0_29_da <= yt_rsc_0_29_i_da;
  yt_rsc_0_29_adra <= yt_rsc_0_29_i_adra;
  yt_rsc_0_29_i_adra_d_1 <= yt_rsc_0_29_i_adra_d;
  yt_rsc_0_29_i_da_d_1 <= yt_rsc_0_29_i_da_d;
  yt_rsc_0_29_i_qa_d <= yt_rsc_0_29_i_qa_d_1;
  yt_rsc_0_29_i_wea_d <= yt_rsc_0_16_i_wea_d_iff;
  yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_29_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_16_i_wea_d_iff;

  yt_rsc_0_30_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_37_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_30_clkb_en,
      clka_en => yt_rsc_0_30_clka_en,
      qb => yt_rsc_0_30_i_qb,
      web => yt_rsc_0_30_web,
      db => yt_rsc_0_30_i_db,
      adrb => yt_rsc_0_30_i_adrb,
      qa => yt_rsc_0_30_i_qa,
      wea => yt_rsc_0_30_wea,
      da => yt_rsc_0_30_i_da,
      adra => yt_rsc_0_30_i_adra,
      adra_d => yt_rsc_0_30_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_16_i_clka_en_d,
      clkb_en_d => yt_rsc_0_16_i_clka_en_d,
      da_d => yt_rsc_0_30_i_da_d_1,
      qa_d => yt_rsc_0_30_i_qa_d_1,
      wea_d => yt_rsc_0_30_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_30_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_30_i_qb <= yt_rsc_0_30_qb;
  yt_rsc_0_30_db <= yt_rsc_0_30_i_db;
  yt_rsc_0_30_adrb <= yt_rsc_0_30_i_adrb;
  yt_rsc_0_30_i_qa <= yt_rsc_0_30_qa;
  yt_rsc_0_30_da <= yt_rsc_0_30_i_da;
  yt_rsc_0_30_adra <= yt_rsc_0_30_i_adra;
  yt_rsc_0_30_i_adra_d_1 <= yt_rsc_0_30_i_adra_d;
  yt_rsc_0_30_i_da_d_1 <= yt_rsc_0_30_i_da_d;
  yt_rsc_0_30_i_qa_d <= yt_rsc_0_30_i_qa_d_1;
  yt_rsc_0_30_i_wea_d <= yt_rsc_0_16_i_wea_d_iff;
  yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_30_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_16_i_wea_d_iff;

  yt_rsc_0_31_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_38_8_32_256_256_32_1_gen
    PORT MAP(
      clkb_en => yt_rsc_0_31_clkb_en,
      clka_en => yt_rsc_0_31_clka_en,
      qb => yt_rsc_0_31_i_qb,
      web => yt_rsc_0_31_web,
      db => yt_rsc_0_31_i_db,
      adrb => yt_rsc_0_31_i_adrb,
      qa => yt_rsc_0_31_i_qa,
      wea => yt_rsc_0_31_wea,
      da => yt_rsc_0_31_i_da,
      adra => yt_rsc_0_31_i_adra,
      adra_d => yt_rsc_0_31_i_adra_d_1,
      clka => clk,
      clka_en_d => yt_rsc_0_16_i_clka_en_d,
      clkb_en_d => yt_rsc_0_16_i_clka_en_d,
      da_d => yt_rsc_0_31_i_da_d_1,
      qa_d => yt_rsc_0_31_i_qa_d_1,
      wea_d => yt_rsc_0_31_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_31_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  yt_rsc_0_31_i_qb <= yt_rsc_0_31_qb;
  yt_rsc_0_31_db <= yt_rsc_0_31_i_db;
  yt_rsc_0_31_adrb <= yt_rsc_0_31_i_adrb;
  yt_rsc_0_31_i_qa <= yt_rsc_0_31_qa;
  yt_rsc_0_31_da <= yt_rsc_0_31_i_da;
  yt_rsc_0_31_adra <= yt_rsc_0_31_i_adra;
  yt_rsc_0_31_i_adra_d_1 <= yt_rsc_0_31_i_adra_d;
  yt_rsc_0_31_i_da_d_1 <= yt_rsc_0_31_i_da_d;
  yt_rsc_0_31_i_qa_d <= yt_rsc_0_31_i_qa_d_1;
  yt_rsc_0_31_i_wea_d <= yt_rsc_0_16_i_wea_d_iff;
  yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_31_i_rwA_rw_ram_ir_internal_WMASK_B_d <= yt_rsc_0_16_i_wea_d_iff;

  xt_rsc_0_0_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_39_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_0_i_qb,
      web => xt_rsc_0_0_web,
      db => xt_rsc_0_0_i_db,
      adrb => xt_rsc_0_0_i_adrb,
      qa => xt_rsc_0_0_i_qa,
      wea => xt_rsc_0_0_wea,
      da => xt_rsc_0_0_i_da,
      adra => xt_rsc_0_0_i_adra,
      adra_d => xt_rsc_0_0_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_0_i_da_d_1,
      qa_d => xt_rsc_0_0_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_0_i_qb <= xt_rsc_0_0_qb;
  xt_rsc_0_0_db <= xt_rsc_0_0_i_db;
  xt_rsc_0_0_adrb <= xt_rsc_0_0_i_adrb;
  xt_rsc_0_0_i_qa <= xt_rsc_0_0_qa;
  xt_rsc_0_0_da <= xt_rsc_0_0_i_da;
  xt_rsc_0_0_adra <= xt_rsc_0_0_i_adra;
  xt_rsc_0_0_i_adra_d_1 <= xt_rsc_0_0_i_adra_d;
  xt_rsc_0_0_i_da_d_1 <= xt_rsc_0_0_i_da_d;
  xt_rsc_0_0_i_qa_d <= xt_rsc_0_0_i_qa_d_1;
  xt_rsc_0_0_i_wea_d <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_0_i_wea_d_iff;

  xt_rsc_0_1_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_40_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_1_i_qb,
      web => xt_rsc_0_1_web,
      db => xt_rsc_0_1_i_db,
      adrb => xt_rsc_0_1_i_adrb,
      qa => xt_rsc_0_1_i_qa,
      wea => xt_rsc_0_1_wea,
      da => xt_rsc_0_1_i_da,
      adra => xt_rsc_0_1_i_adra,
      adra_d => xt_rsc_0_1_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_1_i_da_d_1,
      qa_d => xt_rsc_0_1_i_qa_d_1,
      wea_d => xt_rsc_0_1_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_1_i_qb <= xt_rsc_0_1_qb;
  xt_rsc_0_1_db <= xt_rsc_0_1_i_db;
  xt_rsc_0_1_adrb <= xt_rsc_0_1_i_adrb;
  xt_rsc_0_1_i_qa <= xt_rsc_0_1_qa;
  xt_rsc_0_1_da <= xt_rsc_0_1_i_da;
  xt_rsc_0_1_adra <= xt_rsc_0_1_i_adra;
  xt_rsc_0_1_i_adra_d_1 <= xt_rsc_0_1_i_adra_d;
  xt_rsc_0_1_i_da_d_1 <= xt_rsc_0_1_i_da_d;
  xt_rsc_0_1_i_qa_d <= xt_rsc_0_1_i_qa_d_1;
  xt_rsc_0_1_i_wea_d <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_0_i_wea_d_iff;

  xt_rsc_0_2_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_41_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_2_i_qb,
      web => xt_rsc_0_2_web,
      db => xt_rsc_0_2_i_db,
      adrb => xt_rsc_0_2_i_adrb,
      qa => xt_rsc_0_2_i_qa,
      wea => xt_rsc_0_2_wea,
      da => xt_rsc_0_2_i_da,
      adra => xt_rsc_0_2_i_adra,
      adra_d => xt_rsc_0_2_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_2_i_da_d_1,
      qa_d => xt_rsc_0_2_i_qa_d_1,
      wea_d => xt_rsc_0_2_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_2_i_qb <= xt_rsc_0_2_qb;
  xt_rsc_0_2_db <= xt_rsc_0_2_i_db;
  xt_rsc_0_2_adrb <= xt_rsc_0_2_i_adrb;
  xt_rsc_0_2_i_qa <= xt_rsc_0_2_qa;
  xt_rsc_0_2_da <= xt_rsc_0_2_i_da;
  xt_rsc_0_2_adra <= xt_rsc_0_2_i_adra;
  xt_rsc_0_2_i_adra_d_1 <= xt_rsc_0_2_i_adra_d;
  xt_rsc_0_2_i_da_d_1 <= xt_rsc_0_2_i_da_d;
  xt_rsc_0_2_i_qa_d <= xt_rsc_0_2_i_qa_d_1;
  xt_rsc_0_2_i_wea_d <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_0_i_wea_d_iff;

  xt_rsc_0_3_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_42_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_3_i_qb,
      web => xt_rsc_0_3_web,
      db => xt_rsc_0_3_i_db,
      adrb => xt_rsc_0_3_i_adrb,
      qa => xt_rsc_0_3_i_qa,
      wea => xt_rsc_0_3_wea,
      da => xt_rsc_0_3_i_da,
      adra => xt_rsc_0_3_i_adra,
      adra_d => xt_rsc_0_3_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_3_i_da_d_1,
      qa_d => xt_rsc_0_3_i_qa_d_1,
      wea_d => xt_rsc_0_3_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_3_i_qb <= xt_rsc_0_3_qb;
  xt_rsc_0_3_db <= xt_rsc_0_3_i_db;
  xt_rsc_0_3_adrb <= xt_rsc_0_3_i_adrb;
  xt_rsc_0_3_i_qa <= xt_rsc_0_3_qa;
  xt_rsc_0_3_da <= xt_rsc_0_3_i_da;
  xt_rsc_0_3_adra <= xt_rsc_0_3_i_adra;
  xt_rsc_0_3_i_adra_d_1 <= xt_rsc_0_3_i_adra_d;
  xt_rsc_0_3_i_da_d_1 <= xt_rsc_0_3_i_da_d;
  xt_rsc_0_3_i_qa_d <= xt_rsc_0_3_i_qa_d_1;
  xt_rsc_0_3_i_wea_d <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_0_i_wea_d_iff;

  xt_rsc_0_4_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_43_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_4_i_qb,
      web => xt_rsc_0_4_web,
      db => xt_rsc_0_4_i_db,
      adrb => xt_rsc_0_4_i_adrb,
      qa => xt_rsc_0_4_i_qa,
      wea => xt_rsc_0_4_wea,
      da => xt_rsc_0_4_i_da,
      adra => xt_rsc_0_4_i_adra,
      adra_d => xt_rsc_0_4_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_4_i_da_d_1,
      qa_d => xt_rsc_0_4_i_qa_d_1,
      wea_d => xt_rsc_0_4_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_4_i_qb <= xt_rsc_0_4_qb;
  xt_rsc_0_4_db <= xt_rsc_0_4_i_db;
  xt_rsc_0_4_adrb <= xt_rsc_0_4_i_adrb;
  xt_rsc_0_4_i_qa <= xt_rsc_0_4_qa;
  xt_rsc_0_4_da <= xt_rsc_0_4_i_da;
  xt_rsc_0_4_adra <= xt_rsc_0_4_i_adra;
  xt_rsc_0_4_i_adra_d_1 <= xt_rsc_0_4_i_adra_d;
  xt_rsc_0_4_i_da_d_1 <= xt_rsc_0_4_i_da_d;
  xt_rsc_0_4_i_qa_d <= xt_rsc_0_4_i_qa_d_1;
  xt_rsc_0_4_i_wea_d <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_0_i_wea_d_iff;

  xt_rsc_0_5_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_44_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_5_i_qb,
      web => xt_rsc_0_5_web,
      db => xt_rsc_0_5_i_db,
      adrb => xt_rsc_0_5_i_adrb,
      qa => xt_rsc_0_5_i_qa,
      wea => xt_rsc_0_5_wea,
      da => xt_rsc_0_5_i_da,
      adra => xt_rsc_0_5_i_adra,
      adra_d => xt_rsc_0_5_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_5_i_da_d_1,
      qa_d => xt_rsc_0_5_i_qa_d_1,
      wea_d => xt_rsc_0_5_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_5_i_qb <= xt_rsc_0_5_qb;
  xt_rsc_0_5_db <= xt_rsc_0_5_i_db;
  xt_rsc_0_5_adrb <= xt_rsc_0_5_i_adrb;
  xt_rsc_0_5_i_qa <= xt_rsc_0_5_qa;
  xt_rsc_0_5_da <= xt_rsc_0_5_i_da;
  xt_rsc_0_5_adra <= xt_rsc_0_5_i_adra;
  xt_rsc_0_5_i_adra_d_1 <= xt_rsc_0_5_i_adra_d;
  xt_rsc_0_5_i_da_d_1 <= xt_rsc_0_5_i_da_d;
  xt_rsc_0_5_i_qa_d <= xt_rsc_0_5_i_qa_d_1;
  xt_rsc_0_5_i_wea_d <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_0_i_wea_d_iff;

  xt_rsc_0_6_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_45_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_6_i_qb,
      web => xt_rsc_0_6_web,
      db => xt_rsc_0_6_i_db,
      adrb => xt_rsc_0_6_i_adrb,
      qa => xt_rsc_0_6_i_qa,
      wea => xt_rsc_0_6_wea,
      da => xt_rsc_0_6_i_da,
      adra => xt_rsc_0_6_i_adra,
      adra_d => xt_rsc_0_6_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_6_i_da_d_1,
      qa_d => xt_rsc_0_6_i_qa_d_1,
      wea_d => xt_rsc_0_6_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_6_i_qb <= xt_rsc_0_6_qb;
  xt_rsc_0_6_db <= xt_rsc_0_6_i_db;
  xt_rsc_0_6_adrb <= xt_rsc_0_6_i_adrb;
  xt_rsc_0_6_i_qa <= xt_rsc_0_6_qa;
  xt_rsc_0_6_da <= xt_rsc_0_6_i_da;
  xt_rsc_0_6_adra <= xt_rsc_0_6_i_adra;
  xt_rsc_0_6_i_adra_d_1 <= xt_rsc_0_6_i_adra_d;
  xt_rsc_0_6_i_da_d_1 <= xt_rsc_0_6_i_da_d;
  xt_rsc_0_6_i_qa_d <= xt_rsc_0_6_i_qa_d_1;
  xt_rsc_0_6_i_wea_d <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_0_i_wea_d_iff;

  xt_rsc_0_7_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_46_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_7_i_qb,
      web => xt_rsc_0_7_web,
      db => xt_rsc_0_7_i_db,
      adrb => xt_rsc_0_7_i_adrb,
      qa => xt_rsc_0_7_i_qa,
      wea => xt_rsc_0_7_wea,
      da => xt_rsc_0_7_i_da,
      adra => xt_rsc_0_7_i_adra,
      adra_d => xt_rsc_0_7_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_7_i_da_d_1,
      qa_d => xt_rsc_0_7_i_qa_d_1,
      wea_d => xt_rsc_0_7_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_7_i_qb <= xt_rsc_0_7_qb;
  xt_rsc_0_7_db <= xt_rsc_0_7_i_db;
  xt_rsc_0_7_adrb <= xt_rsc_0_7_i_adrb;
  xt_rsc_0_7_i_qa <= xt_rsc_0_7_qa;
  xt_rsc_0_7_da <= xt_rsc_0_7_i_da;
  xt_rsc_0_7_adra <= xt_rsc_0_7_i_adra;
  xt_rsc_0_7_i_adra_d_1 <= xt_rsc_0_7_i_adra_d;
  xt_rsc_0_7_i_da_d_1 <= xt_rsc_0_7_i_da_d;
  xt_rsc_0_7_i_qa_d <= xt_rsc_0_7_i_qa_d_1;
  xt_rsc_0_7_i_wea_d <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_0_i_wea_d_iff;

  xt_rsc_0_8_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_47_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_8_i_qb,
      web => xt_rsc_0_8_web,
      db => xt_rsc_0_8_i_db,
      adrb => xt_rsc_0_8_i_adrb,
      qa => xt_rsc_0_8_i_qa,
      wea => xt_rsc_0_8_wea,
      da => xt_rsc_0_8_i_da,
      adra => xt_rsc_0_8_i_adra,
      adra_d => xt_rsc_0_8_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_8_i_da_d_1,
      qa_d => xt_rsc_0_8_i_qa_d_1,
      wea_d => xt_rsc_0_8_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_8_i_qb <= xt_rsc_0_8_qb;
  xt_rsc_0_8_db <= xt_rsc_0_8_i_db;
  xt_rsc_0_8_adrb <= xt_rsc_0_8_i_adrb;
  xt_rsc_0_8_i_qa <= xt_rsc_0_8_qa;
  xt_rsc_0_8_da <= xt_rsc_0_8_i_da;
  xt_rsc_0_8_adra <= xt_rsc_0_8_i_adra;
  xt_rsc_0_8_i_adra_d_1 <= xt_rsc_0_8_i_adra_d;
  xt_rsc_0_8_i_da_d_1 <= xt_rsc_0_8_i_da_d;
  xt_rsc_0_8_i_qa_d <= xt_rsc_0_8_i_qa_d_1;
  xt_rsc_0_8_i_wea_d <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_0_i_wea_d_iff;

  xt_rsc_0_9_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_48_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_9_i_qb,
      web => xt_rsc_0_9_web,
      db => xt_rsc_0_9_i_db,
      adrb => xt_rsc_0_9_i_adrb,
      qa => xt_rsc_0_9_i_qa,
      wea => xt_rsc_0_9_wea,
      da => xt_rsc_0_9_i_da,
      adra => xt_rsc_0_9_i_adra,
      adra_d => xt_rsc_0_9_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_9_i_da_d_1,
      qa_d => xt_rsc_0_9_i_qa_d_1,
      wea_d => xt_rsc_0_9_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_9_i_qb <= xt_rsc_0_9_qb;
  xt_rsc_0_9_db <= xt_rsc_0_9_i_db;
  xt_rsc_0_9_adrb <= xt_rsc_0_9_i_adrb;
  xt_rsc_0_9_i_qa <= xt_rsc_0_9_qa;
  xt_rsc_0_9_da <= xt_rsc_0_9_i_da;
  xt_rsc_0_9_adra <= xt_rsc_0_9_i_adra;
  xt_rsc_0_9_i_adra_d_1 <= xt_rsc_0_9_i_adra_d;
  xt_rsc_0_9_i_da_d_1 <= xt_rsc_0_9_i_da_d;
  xt_rsc_0_9_i_qa_d <= xt_rsc_0_9_i_qa_d_1;
  xt_rsc_0_9_i_wea_d <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_0_i_wea_d_iff;

  xt_rsc_0_10_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_49_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_10_i_qb,
      web => xt_rsc_0_10_web,
      db => xt_rsc_0_10_i_db,
      adrb => xt_rsc_0_10_i_adrb,
      qa => xt_rsc_0_10_i_qa,
      wea => xt_rsc_0_10_wea,
      da => xt_rsc_0_10_i_da,
      adra => xt_rsc_0_10_i_adra,
      adra_d => xt_rsc_0_10_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_10_i_da_d_1,
      qa_d => xt_rsc_0_10_i_qa_d_1,
      wea_d => xt_rsc_0_10_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_10_i_qb <= xt_rsc_0_10_qb;
  xt_rsc_0_10_db <= xt_rsc_0_10_i_db;
  xt_rsc_0_10_adrb <= xt_rsc_0_10_i_adrb;
  xt_rsc_0_10_i_qa <= xt_rsc_0_10_qa;
  xt_rsc_0_10_da <= xt_rsc_0_10_i_da;
  xt_rsc_0_10_adra <= xt_rsc_0_10_i_adra;
  xt_rsc_0_10_i_adra_d_1 <= xt_rsc_0_10_i_adra_d;
  xt_rsc_0_10_i_da_d_1 <= xt_rsc_0_10_i_da_d;
  xt_rsc_0_10_i_qa_d <= xt_rsc_0_10_i_qa_d_1;
  xt_rsc_0_10_i_wea_d <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_0_i_wea_d_iff;

  xt_rsc_0_11_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_50_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_11_i_qb,
      web => xt_rsc_0_11_web,
      db => xt_rsc_0_11_i_db,
      adrb => xt_rsc_0_11_i_adrb,
      qa => xt_rsc_0_11_i_qa,
      wea => xt_rsc_0_11_wea,
      da => xt_rsc_0_11_i_da,
      adra => xt_rsc_0_11_i_adra,
      adra_d => xt_rsc_0_11_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_11_i_da_d_1,
      qa_d => xt_rsc_0_11_i_qa_d_1,
      wea_d => xt_rsc_0_11_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_11_i_qb <= xt_rsc_0_11_qb;
  xt_rsc_0_11_db <= xt_rsc_0_11_i_db;
  xt_rsc_0_11_adrb <= xt_rsc_0_11_i_adrb;
  xt_rsc_0_11_i_qa <= xt_rsc_0_11_qa;
  xt_rsc_0_11_da <= xt_rsc_0_11_i_da;
  xt_rsc_0_11_adra <= xt_rsc_0_11_i_adra;
  xt_rsc_0_11_i_adra_d_1 <= xt_rsc_0_11_i_adra_d;
  xt_rsc_0_11_i_da_d_1 <= xt_rsc_0_11_i_da_d;
  xt_rsc_0_11_i_qa_d <= xt_rsc_0_11_i_qa_d_1;
  xt_rsc_0_11_i_wea_d <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_0_i_wea_d_iff;

  xt_rsc_0_12_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_51_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_12_i_qb,
      web => xt_rsc_0_12_web,
      db => xt_rsc_0_12_i_db,
      adrb => xt_rsc_0_12_i_adrb,
      qa => xt_rsc_0_12_i_qa,
      wea => xt_rsc_0_12_wea,
      da => xt_rsc_0_12_i_da,
      adra => xt_rsc_0_12_i_adra,
      adra_d => xt_rsc_0_12_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_12_i_da_d_1,
      qa_d => xt_rsc_0_12_i_qa_d_1,
      wea_d => xt_rsc_0_12_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_12_i_qb <= xt_rsc_0_12_qb;
  xt_rsc_0_12_db <= xt_rsc_0_12_i_db;
  xt_rsc_0_12_adrb <= xt_rsc_0_12_i_adrb;
  xt_rsc_0_12_i_qa <= xt_rsc_0_12_qa;
  xt_rsc_0_12_da <= xt_rsc_0_12_i_da;
  xt_rsc_0_12_adra <= xt_rsc_0_12_i_adra;
  xt_rsc_0_12_i_adra_d_1 <= xt_rsc_0_12_i_adra_d;
  xt_rsc_0_12_i_da_d_1 <= xt_rsc_0_12_i_da_d;
  xt_rsc_0_12_i_qa_d <= xt_rsc_0_12_i_qa_d_1;
  xt_rsc_0_12_i_wea_d <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_0_i_wea_d_iff;

  xt_rsc_0_13_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_52_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_13_i_qb,
      web => xt_rsc_0_13_web,
      db => xt_rsc_0_13_i_db,
      adrb => xt_rsc_0_13_i_adrb,
      qa => xt_rsc_0_13_i_qa,
      wea => xt_rsc_0_13_wea,
      da => xt_rsc_0_13_i_da,
      adra => xt_rsc_0_13_i_adra,
      adra_d => xt_rsc_0_13_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_13_i_da_d_1,
      qa_d => xt_rsc_0_13_i_qa_d_1,
      wea_d => xt_rsc_0_13_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_13_i_qb <= xt_rsc_0_13_qb;
  xt_rsc_0_13_db <= xt_rsc_0_13_i_db;
  xt_rsc_0_13_adrb <= xt_rsc_0_13_i_adrb;
  xt_rsc_0_13_i_qa <= xt_rsc_0_13_qa;
  xt_rsc_0_13_da <= xt_rsc_0_13_i_da;
  xt_rsc_0_13_adra <= xt_rsc_0_13_i_adra;
  xt_rsc_0_13_i_adra_d_1 <= xt_rsc_0_13_i_adra_d;
  xt_rsc_0_13_i_da_d_1 <= xt_rsc_0_13_i_da_d;
  xt_rsc_0_13_i_qa_d <= xt_rsc_0_13_i_qa_d_1;
  xt_rsc_0_13_i_wea_d <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_0_i_wea_d_iff;

  xt_rsc_0_14_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_53_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_14_i_qb,
      web => xt_rsc_0_14_web,
      db => xt_rsc_0_14_i_db,
      adrb => xt_rsc_0_14_i_adrb,
      qa => xt_rsc_0_14_i_qa,
      wea => xt_rsc_0_14_wea,
      da => xt_rsc_0_14_i_da,
      adra => xt_rsc_0_14_i_adra,
      adra_d => xt_rsc_0_14_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_14_i_da_d_1,
      qa_d => xt_rsc_0_14_i_qa_d_1,
      wea_d => xt_rsc_0_14_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_14_i_qb <= xt_rsc_0_14_qb;
  xt_rsc_0_14_db <= xt_rsc_0_14_i_db;
  xt_rsc_0_14_adrb <= xt_rsc_0_14_i_adrb;
  xt_rsc_0_14_i_qa <= xt_rsc_0_14_qa;
  xt_rsc_0_14_da <= xt_rsc_0_14_i_da;
  xt_rsc_0_14_adra <= xt_rsc_0_14_i_adra;
  xt_rsc_0_14_i_adra_d_1 <= xt_rsc_0_14_i_adra_d;
  xt_rsc_0_14_i_da_d_1 <= xt_rsc_0_14_i_da_d;
  xt_rsc_0_14_i_qa_d <= xt_rsc_0_14_i_qa_d_1;
  xt_rsc_0_14_i_wea_d <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_0_i_wea_d_iff;

  xt_rsc_0_15_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_54_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_15_i_qb,
      web => xt_rsc_0_15_web,
      db => xt_rsc_0_15_i_db,
      adrb => xt_rsc_0_15_i_adrb,
      qa => xt_rsc_0_15_i_qa,
      wea => xt_rsc_0_15_wea,
      da => xt_rsc_0_15_i_da,
      adra => xt_rsc_0_15_i_adra,
      adra_d => xt_rsc_0_15_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_15_i_da_d_1,
      qa_d => xt_rsc_0_15_i_qa_d_1,
      wea_d => xt_rsc_0_15_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_15_i_qb <= xt_rsc_0_15_qb;
  xt_rsc_0_15_db <= xt_rsc_0_15_i_db;
  xt_rsc_0_15_adrb <= xt_rsc_0_15_i_adrb;
  xt_rsc_0_15_i_qa <= xt_rsc_0_15_qa;
  xt_rsc_0_15_da <= xt_rsc_0_15_i_da;
  xt_rsc_0_15_adra <= xt_rsc_0_15_i_adra;
  xt_rsc_0_15_i_adra_d_1 <= xt_rsc_0_15_i_adra_d;
  xt_rsc_0_15_i_da_d_1 <= xt_rsc_0_15_i_da_d;
  xt_rsc_0_15_i_qa_d <= xt_rsc_0_15_i_qa_d_1;
  xt_rsc_0_15_i_wea_d <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_0_i_wea_d_iff;

  xt_rsc_0_16_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_55_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_16_i_qb,
      web => xt_rsc_0_16_web,
      db => xt_rsc_0_16_i_db,
      adrb => xt_rsc_0_16_i_adrb,
      qa => xt_rsc_0_16_i_qa,
      wea => xt_rsc_0_16_wea,
      da => xt_rsc_0_16_i_da,
      adra => xt_rsc_0_16_i_adra,
      adra_d => xt_rsc_0_16_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_16_i_da_d_1,
      qa_d => xt_rsc_0_16_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_16_i_qb <= xt_rsc_0_16_qb;
  xt_rsc_0_16_db <= xt_rsc_0_16_i_db;
  xt_rsc_0_16_adrb <= xt_rsc_0_16_i_adrb;
  xt_rsc_0_16_i_qa <= xt_rsc_0_16_qa;
  xt_rsc_0_16_da <= xt_rsc_0_16_i_da;
  xt_rsc_0_16_adra <= xt_rsc_0_16_i_adra;
  xt_rsc_0_16_i_adra_d_1 <= xt_rsc_0_16_i_adra_d;
  xt_rsc_0_16_i_da_d_1 <= xt_rsc_0_16_i_da_d;
  xt_rsc_0_16_i_qa_d <= xt_rsc_0_16_i_qa_d_1;
  xt_rsc_0_16_i_wea_d <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_16_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_16_i_wea_d_iff;

  xt_rsc_0_17_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_56_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_17_i_qb,
      web => xt_rsc_0_17_web,
      db => xt_rsc_0_17_i_db,
      adrb => xt_rsc_0_17_i_adrb,
      qa => xt_rsc_0_17_i_qa,
      wea => xt_rsc_0_17_wea,
      da => xt_rsc_0_17_i_da,
      adra => xt_rsc_0_17_i_adra,
      adra_d => xt_rsc_0_17_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_17_i_da_d_1,
      qa_d => xt_rsc_0_17_i_qa_d_1,
      wea_d => xt_rsc_0_17_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_17_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_17_i_qb <= xt_rsc_0_17_qb;
  xt_rsc_0_17_db <= xt_rsc_0_17_i_db;
  xt_rsc_0_17_adrb <= xt_rsc_0_17_i_adrb;
  xt_rsc_0_17_i_qa <= xt_rsc_0_17_qa;
  xt_rsc_0_17_da <= xt_rsc_0_17_i_da;
  xt_rsc_0_17_adra <= xt_rsc_0_17_i_adra;
  xt_rsc_0_17_i_adra_d_1 <= xt_rsc_0_17_i_adra_d;
  xt_rsc_0_17_i_da_d_1 <= xt_rsc_0_17_i_da_d;
  xt_rsc_0_17_i_qa_d <= xt_rsc_0_17_i_qa_d_1;
  xt_rsc_0_17_i_wea_d <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_17_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_16_i_wea_d_iff;

  xt_rsc_0_18_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_57_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_18_i_qb,
      web => xt_rsc_0_18_web,
      db => xt_rsc_0_18_i_db,
      adrb => xt_rsc_0_18_i_adrb,
      qa => xt_rsc_0_18_i_qa,
      wea => xt_rsc_0_18_wea,
      da => xt_rsc_0_18_i_da,
      adra => xt_rsc_0_18_i_adra,
      adra_d => xt_rsc_0_18_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_18_i_da_d_1,
      qa_d => xt_rsc_0_18_i_qa_d_1,
      wea_d => xt_rsc_0_18_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_18_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_18_i_qb <= xt_rsc_0_18_qb;
  xt_rsc_0_18_db <= xt_rsc_0_18_i_db;
  xt_rsc_0_18_adrb <= xt_rsc_0_18_i_adrb;
  xt_rsc_0_18_i_qa <= xt_rsc_0_18_qa;
  xt_rsc_0_18_da <= xt_rsc_0_18_i_da;
  xt_rsc_0_18_adra <= xt_rsc_0_18_i_adra;
  xt_rsc_0_18_i_adra_d_1 <= xt_rsc_0_18_i_adra_d;
  xt_rsc_0_18_i_da_d_1 <= xt_rsc_0_18_i_da_d;
  xt_rsc_0_18_i_qa_d <= xt_rsc_0_18_i_qa_d_1;
  xt_rsc_0_18_i_wea_d <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_18_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_16_i_wea_d_iff;

  xt_rsc_0_19_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_58_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_19_i_qb,
      web => xt_rsc_0_19_web,
      db => xt_rsc_0_19_i_db,
      adrb => xt_rsc_0_19_i_adrb,
      qa => xt_rsc_0_19_i_qa,
      wea => xt_rsc_0_19_wea,
      da => xt_rsc_0_19_i_da,
      adra => xt_rsc_0_19_i_adra,
      adra_d => xt_rsc_0_19_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_19_i_da_d_1,
      qa_d => xt_rsc_0_19_i_qa_d_1,
      wea_d => xt_rsc_0_19_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_19_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_19_i_qb <= xt_rsc_0_19_qb;
  xt_rsc_0_19_db <= xt_rsc_0_19_i_db;
  xt_rsc_0_19_adrb <= xt_rsc_0_19_i_adrb;
  xt_rsc_0_19_i_qa <= xt_rsc_0_19_qa;
  xt_rsc_0_19_da <= xt_rsc_0_19_i_da;
  xt_rsc_0_19_adra <= xt_rsc_0_19_i_adra;
  xt_rsc_0_19_i_adra_d_1 <= xt_rsc_0_19_i_adra_d;
  xt_rsc_0_19_i_da_d_1 <= xt_rsc_0_19_i_da_d;
  xt_rsc_0_19_i_qa_d <= xt_rsc_0_19_i_qa_d_1;
  xt_rsc_0_19_i_wea_d <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_19_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_16_i_wea_d_iff;

  xt_rsc_0_20_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_59_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_20_i_qb,
      web => xt_rsc_0_20_web,
      db => xt_rsc_0_20_i_db,
      adrb => xt_rsc_0_20_i_adrb,
      qa => xt_rsc_0_20_i_qa,
      wea => xt_rsc_0_20_wea,
      da => xt_rsc_0_20_i_da,
      adra => xt_rsc_0_20_i_adra,
      adra_d => xt_rsc_0_20_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_20_i_da_d_1,
      qa_d => xt_rsc_0_20_i_qa_d_1,
      wea_d => xt_rsc_0_20_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_20_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_20_i_qb <= xt_rsc_0_20_qb;
  xt_rsc_0_20_db <= xt_rsc_0_20_i_db;
  xt_rsc_0_20_adrb <= xt_rsc_0_20_i_adrb;
  xt_rsc_0_20_i_qa <= xt_rsc_0_20_qa;
  xt_rsc_0_20_da <= xt_rsc_0_20_i_da;
  xt_rsc_0_20_adra <= xt_rsc_0_20_i_adra;
  xt_rsc_0_20_i_adra_d_1 <= xt_rsc_0_20_i_adra_d;
  xt_rsc_0_20_i_da_d_1 <= xt_rsc_0_20_i_da_d;
  xt_rsc_0_20_i_qa_d <= xt_rsc_0_20_i_qa_d_1;
  xt_rsc_0_20_i_wea_d <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_20_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_16_i_wea_d_iff;

  xt_rsc_0_21_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_60_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_21_i_qb,
      web => xt_rsc_0_21_web,
      db => xt_rsc_0_21_i_db,
      adrb => xt_rsc_0_21_i_adrb,
      qa => xt_rsc_0_21_i_qa,
      wea => xt_rsc_0_21_wea,
      da => xt_rsc_0_21_i_da,
      adra => xt_rsc_0_21_i_adra,
      adra_d => xt_rsc_0_21_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_21_i_da_d_1,
      qa_d => xt_rsc_0_21_i_qa_d_1,
      wea_d => xt_rsc_0_21_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_21_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_21_i_qb <= xt_rsc_0_21_qb;
  xt_rsc_0_21_db <= xt_rsc_0_21_i_db;
  xt_rsc_0_21_adrb <= xt_rsc_0_21_i_adrb;
  xt_rsc_0_21_i_qa <= xt_rsc_0_21_qa;
  xt_rsc_0_21_da <= xt_rsc_0_21_i_da;
  xt_rsc_0_21_adra <= xt_rsc_0_21_i_adra;
  xt_rsc_0_21_i_adra_d_1 <= xt_rsc_0_21_i_adra_d;
  xt_rsc_0_21_i_da_d_1 <= xt_rsc_0_21_i_da_d;
  xt_rsc_0_21_i_qa_d <= xt_rsc_0_21_i_qa_d_1;
  xt_rsc_0_21_i_wea_d <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_21_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_16_i_wea_d_iff;

  xt_rsc_0_22_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_61_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_22_i_qb,
      web => xt_rsc_0_22_web,
      db => xt_rsc_0_22_i_db,
      adrb => xt_rsc_0_22_i_adrb,
      qa => xt_rsc_0_22_i_qa,
      wea => xt_rsc_0_22_wea,
      da => xt_rsc_0_22_i_da,
      adra => xt_rsc_0_22_i_adra,
      adra_d => xt_rsc_0_22_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_22_i_da_d_1,
      qa_d => xt_rsc_0_22_i_qa_d_1,
      wea_d => xt_rsc_0_22_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_22_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_22_i_qb <= xt_rsc_0_22_qb;
  xt_rsc_0_22_db <= xt_rsc_0_22_i_db;
  xt_rsc_0_22_adrb <= xt_rsc_0_22_i_adrb;
  xt_rsc_0_22_i_qa <= xt_rsc_0_22_qa;
  xt_rsc_0_22_da <= xt_rsc_0_22_i_da;
  xt_rsc_0_22_adra <= xt_rsc_0_22_i_adra;
  xt_rsc_0_22_i_adra_d_1 <= xt_rsc_0_22_i_adra_d;
  xt_rsc_0_22_i_da_d_1 <= xt_rsc_0_22_i_da_d;
  xt_rsc_0_22_i_qa_d <= xt_rsc_0_22_i_qa_d_1;
  xt_rsc_0_22_i_wea_d <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_22_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_16_i_wea_d_iff;

  xt_rsc_0_23_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_62_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_23_i_qb,
      web => xt_rsc_0_23_web,
      db => xt_rsc_0_23_i_db,
      adrb => xt_rsc_0_23_i_adrb,
      qa => xt_rsc_0_23_i_qa,
      wea => xt_rsc_0_23_wea,
      da => xt_rsc_0_23_i_da,
      adra => xt_rsc_0_23_i_adra,
      adra_d => xt_rsc_0_23_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_23_i_da_d_1,
      qa_d => xt_rsc_0_23_i_qa_d_1,
      wea_d => xt_rsc_0_23_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_23_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_23_i_qb <= xt_rsc_0_23_qb;
  xt_rsc_0_23_db <= xt_rsc_0_23_i_db;
  xt_rsc_0_23_adrb <= xt_rsc_0_23_i_adrb;
  xt_rsc_0_23_i_qa <= xt_rsc_0_23_qa;
  xt_rsc_0_23_da <= xt_rsc_0_23_i_da;
  xt_rsc_0_23_adra <= xt_rsc_0_23_i_adra;
  xt_rsc_0_23_i_adra_d_1 <= xt_rsc_0_23_i_adra_d;
  xt_rsc_0_23_i_da_d_1 <= xt_rsc_0_23_i_da_d;
  xt_rsc_0_23_i_qa_d <= xt_rsc_0_23_i_qa_d_1;
  xt_rsc_0_23_i_wea_d <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_23_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_16_i_wea_d_iff;

  xt_rsc_0_24_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_63_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_24_i_qb,
      web => xt_rsc_0_24_web,
      db => xt_rsc_0_24_i_db,
      adrb => xt_rsc_0_24_i_adrb,
      qa => xt_rsc_0_24_i_qa,
      wea => xt_rsc_0_24_wea,
      da => xt_rsc_0_24_i_da,
      adra => xt_rsc_0_24_i_adra,
      adra_d => xt_rsc_0_24_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_24_i_da_d_1,
      qa_d => xt_rsc_0_24_i_qa_d_1,
      wea_d => xt_rsc_0_24_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_24_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_24_i_qb <= xt_rsc_0_24_qb;
  xt_rsc_0_24_db <= xt_rsc_0_24_i_db;
  xt_rsc_0_24_adrb <= xt_rsc_0_24_i_adrb;
  xt_rsc_0_24_i_qa <= xt_rsc_0_24_qa;
  xt_rsc_0_24_da <= xt_rsc_0_24_i_da;
  xt_rsc_0_24_adra <= xt_rsc_0_24_i_adra;
  xt_rsc_0_24_i_adra_d_1 <= xt_rsc_0_24_i_adra_d;
  xt_rsc_0_24_i_da_d_1 <= xt_rsc_0_24_i_da_d;
  xt_rsc_0_24_i_qa_d <= xt_rsc_0_24_i_qa_d_1;
  xt_rsc_0_24_i_wea_d <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_24_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_16_i_wea_d_iff;

  xt_rsc_0_25_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_64_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_25_i_qb,
      web => xt_rsc_0_25_web,
      db => xt_rsc_0_25_i_db,
      adrb => xt_rsc_0_25_i_adrb,
      qa => xt_rsc_0_25_i_qa,
      wea => xt_rsc_0_25_wea,
      da => xt_rsc_0_25_i_da,
      adra => xt_rsc_0_25_i_adra,
      adra_d => xt_rsc_0_25_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_25_i_da_d_1,
      qa_d => xt_rsc_0_25_i_qa_d_1,
      wea_d => xt_rsc_0_25_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_25_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_25_i_qb <= xt_rsc_0_25_qb;
  xt_rsc_0_25_db <= xt_rsc_0_25_i_db;
  xt_rsc_0_25_adrb <= xt_rsc_0_25_i_adrb;
  xt_rsc_0_25_i_qa <= xt_rsc_0_25_qa;
  xt_rsc_0_25_da <= xt_rsc_0_25_i_da;
  xt_rsc_0_25_adra <= xt_rsc_0_25_i_adra;
  xt_rsc_0_25_i_adra_d_1 <= xt_rsc_0_25_i_adra_d;
  xt_rsc_0_25_i_da_d_1 <= xt_rsc_0_25_i_da_d;
  xt_rsc_0_25_i_qa_d <= xt_rsc_0_25_i_qa_d_1;
  xt_rsc_0_25_i_wea_d <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_25_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_16_i_wea_d_iff;

  xt_rsc_0_26_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_65_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_26_i_qb,
      web => xt_rsc_0_26_web,
      db => xt_rsc_0_26_i_db,
      adrb => xt_rsc_0_26_i_adrb,
      qa => xt_rsc_0_26_i_qa,
      wea => xt_rsc_0_26_wea,
      da => xt_rsc_0_26_i_da,
      adra => xt_rsc_0_26_i_adra,
      adra_d => xt_rsc_0_26_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_26_i_da_d_1,
      qa_d => xt_rsc_0_26_i_qa_d_1,
      wea_d => xt_rsc_0_26_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_26_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_26_i_qb <= xt_rsc_0_26_qb;
  xt_rsc_0_26_db <= xt_rsc_0_26_i_db;
  xt_rsc_0_26_adrb <= xt_rsc_0_26_i_adrb;
  xt_rsc_0_26_i_qa <= xt_rsc_0_26_qa;
  xt_rsc_0_26_da <= xt_rsc_0_26_i_da;
  xt_rsc_0_26_adra <= xt_rsc_0_26_i_adra;
  xt_rsc_0_26_i_adra_d_1 <= xt_rsc_0_26_i_adra_d;
  xt_rsc_0_26_i_da_d_1 <= xt_rsc_0_26_i_da_d;
  xt_rsc_0_26_i_qa_d <= xt_rsc_0_26_i_qa_d_1;
  xt_rsc_0_26_i_wea_d <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_26_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_16_i_wea_d_iff;

  xt_rsc_0_27_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_66_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_27_i_qb,
      web => xt_rsc_0_27_web,
      db => xt_rsc_0_27_i_db,
      adrb => xt_rsc_0_27_i_adrb,
      qa => xt_rsc_0_27_i_qa,
      wea => xt_rsc_0_27_wea,
      da => xt_rsc_0_27_i_da,
      adra => xt_rsc_0_27_i_adra,
      adra_d => xt_rsc_0_27_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_27_i_da_d_1,
      qa_d => xt_rsc_0_27_i_qa_d_1,
      wea_d => xt_rsc_0_27_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_27_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_27_i_qb <= xt_rsc_0_27_qb;
  xt_rsc_0_27_db <= xt_rsc_0_27_i_db;
  xt_rsc_0_27_adrb <= xt_rsc_0_27_i_adrb;
  xt_rsc_0_27_i_qa <= xt_rsc_0_27_qa;
  xt_rsc_0_27_da <= xt_rsc_0_27_i_da;
  xt_rsc_0_27_adra <= xt_rsc_0_27_i_adra;
  xt_rsc_0_27_i_adra_d_1 <= xt_rsc_0_27_i_adra_d;
  xt_rsc_0_27_i_da_d_1 <= xt_rsc_0_27_i_da_d;
  xt_rsc_0_27_i_qa_d <= xt_rsc_0_27_i_qa_d_1;
  xt_rsc_0_27_i_wea_d <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_27_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_16_i_wea_d_iff;

  xt_rsc_0_28_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_67_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_28_i_qb,
      web => xt_rsc_0_28_web,
      db => xt_rsc_0_28_i_db,
      adrb => xt_rsc_0_28_i_adrb,
      qa => xt_rsc_0_28_i_qa,
      wea => xt_rsc_0_28_wea,
      da => xt_rsc_0_28_i_da,
      adra => xt_rsc_0_28_i_adra,
      adra_d => xt_rsc_0_28_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_28_i_da_d_1,
      qa_d => xt_rsc_0_28_i_qa_d_1,
      wea_d => xt_rsc_0_28_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_28_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_28_i_qb <= xt_rsc_0_28_qb;
  xt_rsc_0_28_db <= xt_rsc_0_28_i_db;
  xt_rsc_0_28_adrb <= xt_rsc_0_28_i_adrb;
  xt_rsc_0_28_i_qa <= xt_rsc_0_28_qa;
  xt_rsc_0_28_da <= xt_rsc_0_28_i_da;
  xt_rsc_0_28_adra <= xt_rsc_0_28_i_adra;
  xt_rsc_0_28_i_adra_d_1 <= xt_rsc_0_28_i_adra_d;
  xt_rsc_0_28_i_da_d_1 <= xt_rsc_0_28_i_da_d;
  xt_rsc_0_28_i_qa_d <= xt_rsc_0_28_i_qa_d_1;
  xt_rsc_0_28_i_wea_d <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_28_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_16_i_wea_d_iff;

  xt_rsc_0_29_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_68_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_29_i_qb,
      web => xt_rsc_0_29_web,
      db => xt_rsc_0_29_i_db,
      adrb => xt_rsc_0_29_i_adrb,
      qa => xt_rsc_0_29_i_qa,
      wea => xt_rsc_0_29_wea,
      da => xt_rsc_0_29_i_da,
      adra => xt_rsc_0_29_i_adra,
      adra_d => xt_rsc_0_29_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_29_i_da_d_1,
      qa_d => xt_rsc_0_29_i_qa_d_1,
      wea_d => xt_rsc_0_29_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_29_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_29_i_qb <= xt_rsc_0_29_qb;
  xt_rsc_0_29_db <= xt_rsc_0_29_i_db;
  xt_rsc_0_29_adrb <= xt_rsc_0_29_i_adrb;
  xt_rsc_0_29_i_qa <= xt_rsc_0_29_qa;
  xt_rsc_0_29_da <= xt_rsc_0_29_i_da;
  xt_rsc_0_29_adra <= xt_rsc_0_29_i_adra;
  xt_rsc_0_29_i_adra_d_1 <= xt_rsc_0_29_i_adra_d;
  xt_rsc_0_29_i_da_d_1 <= xt_rsc_0_29_i_da_d;
  xt_rsc_0_29_i_qa_d <= xt_rsc_0_29_i_qa_d_1;
  xt_rsc_0_29_i_wea_d <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_29_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_16_i_wea_d_iff;

  xt_rsc_0_30_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_69_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_30_i_qb,
      web => xt_rsc_0_30_web,
      db => xt_rsc_0_30_i_db,
      adrb => xt_rsc_0_30_i_adrb,
      qa => xt_rsc_0_30_i_qa,
      wea => xt_rsc_0_30_wea,
      da => xt_rsc_0_30_i_da,
      adra => xt_rsc_0_30_i_adra,
      adra_d => xt_rsc_0_30_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_30_i_da_d_1,
      qa_d => xt_rsc_0_30_i_qa_d_1,
      wea_d => xt_rsc_0_30_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_30_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_30_i_qb <= xt_rsc_0_30_qb;
  xt_rsc_0_30_db <= xt_rsc_0_30_i_db;
  xt_rsc_0_30_adrb <= xt_rsc_0_30_i_adrb;
  xt_rsc_0_30_i_qa <= xt_rsc_0_30_qa;
  xt_rsc_0_30_da <= xt_rsc_0_30_i_da;
  xt_rsc_0_30_adra <= xt_rsc_0_30_i_adra;
  xt_rsc_0_30_i_adra_d_1 <= xt_rsc_0_30_i_adra_d;
  xt_rsc_0_30_i_da_d_1 <= xt_rsc_0_30_i_da_d;
  xt_rsc_0_30_i_qa_d <= xt_rsc_0_30_i_qa_d_1;
  xt_rsc_0_30_i_wea_d <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_30_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_16_i_wea_d_iff;

  xt_rsc_0_31_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_70_8_32_256_256_32_1_gen
    PORT MAP(
      qb => xt_rsc_0_31_i_qb,
      web => xt_rsc_0_31_web,
      db => xt_rsc_0_31_i_db,
      adrb => xt_rsc_0_31_i_adrb,
      qa => xt_rsc_0_31_i_qa,
      wea => xt_rsc_0_31_wea,
      da => xt_rsc_0_31_i_da,
      adra => xt_rsc_0_31_i_adra,
      adra_d => xt_rsc_0_31_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => xt_rsc_0_31_i_da_d_1,
      qa_d => xt_rsc_0_31_i_qa_d_1,
      wea_d => xt_rsc_0_31_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_31_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  xt_rsc_0_31_i_qb <= xt_rsc_0_31_qb;
  xt_rsc_0_31_db <= xt_rsc_0_31_i_db;
  xt_rsc_0_31_adrb <= xt_rsc_0_31_i_adrb;
  xt_rsc_0_31_i_qa <= xt_rsc_0_31_qa;
  xt_rsc_0_31_da <= xt_rsc_0_31_i_da;
  xt_rsc_0_31_adra <= xt_rsc_0_31_i_adra;
  xt_rsc_0_31_i_adra_d_1 <= xt_rsc_0_31_i_adra_d;
  xt_rsc_0_31_i_da_d_1 <= xt_rsc_0_31_i_da_d;
  xt_rsc_0_31_i_qa_d <= xt_rsc_0_31_i_qa_d_1;
  xt_rsc_0_31_i_wea_d <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_31_i_rwA_rw_ram_ir_internal_WMASK_B_d <= xt_rsc_0_16_i_wea_d_iff;

  twiddle_rsc_0_0_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_71_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_0_i_qb,
      web => twiddle_rsc_0_0_web,
      db => twiddle_rsc_0_0_i_db,
      adrb => twiddle_rsc_0_0_i_adrb,
      qa => twiddle_rsc_0_0_i_qa,
      wea => twiddle_rsc_0_0_wea,
      da => twiddle_rsc_0_0_i_da,
      adra => twiddle_rsc_0_0_i_adra,
      adra_d => twiddle_rsc_0_0_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_0_i_da_d,
      qa_d => twiddle_rsc_0_0_i_qa_d_1,
      wea_d => twiddle_rsc_0_0_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_0_i_qb <= twiddle_rsc_0_0_qb;
  twiddle_rsc_0_0_db <= twiddle_rsc_0_0_i_db;
  twiddle_rsc_0_0_adrb <= twiddle_rsc_0_0_i_adrb;
  twiddle_rsc_0_0_i_qa <= twiddle_rsc_0_0_qa;
  twiddle_rsc_0_0_da <= twiddle_rsc_0_0_i_da;
  twiddle_rsc_0_0_adra <= twiddle_rsc_0_0_i_adra;
  twiddle_rsc_0_0_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_0_i_adra_d;
  twiddle_rsc_0_0_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_0_i_qa_d <= twiddle_rsc_0_0_i_qa_d_1;
  twiddle_rsc_0_0_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_1_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_72_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_1_i_qb,
      web => twiddle_rsc_0_1_web,
      db => twiddle_rsc_0_1_i_db,
      adrb => twiddle_rsc_0_1_i_adrb,
      qa => twiddle_rsc_0_1_i_qa,
      wea => twiddle_rsc_0_1_wea,
      da => twiddle_rsc_0_1_i_da,
      adra => twiddle_rsc_0_1_i_adra,
      adra_d => twiddle_rsc_0_1_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_1_i_da_d,
      qa_d => twiddle_rsc_0_1_i_qa_d_1,
      wea_d => twiddle_rsc_0_1_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_1_i_qb <= twiddle_rsc_0_1_qb;
  twiddle_rsc_0_1_db <= twiddle_rsc_0_1_i_db;
  twiddle_rsc_0_1_adrb <= twiddle_rsc_0_1_i_adrb;
  twiddle_rsc_0_1_i_qa <= twiddle_rsc_0_1_qa;
  twiddle_rsc_0_1_da <= twiddle_rsc_0_1_i_da;
  twiddle_rsc_0_1_adra <= twiddle_rsc_0_1_i_adra;
  twiddle_rsc_0_1_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_1_i_adra_d;
  twiddle_rsc_0_1_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_1_i_qa_d <= twiddle_rsc_0_1_i_qa_d_1;
  twiddle_rsc_0_1_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_2_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_73_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_2_i_qb,
      web => twiddle_rsc_0_2_web,
      db => twiddle_rsc_0_2_i_db,
      adrb => twiddle_rsc_0_2_i_adrb,
      qa => twiddle_rsc_0_2_i_qa,
      wea => twiddle_rsc_0_2_wea,
      da => twiddle_rsc_0_2_i_da,
      adra => twiddle_rsc_0_2_i_adra,
      adra_d => twiddle_rsc_0_2_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_2_i_da_d,
      qa_d => twiddle_rsc_0_2_i_qa_d_1,
      wea_d => twiddle_rsc_0_2_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_2_i_qb <= twiddle_rsc_0_2_qb;
  twiddle_rsc_0_2_db <= twiddle_rsc_0_2_i_db;
  twiddle_rsc_0_2_adrb <= twiddle_rsc_0_2_i_adrb;
  twiddle_rsc_0_2_i_qa <= twiddle_rsc_0_2_qa;
  twiddle_rsc_0_2_da <= twiddle_rsc_0_2_i_da;
  twiddle_rsc_0_2_adra <= twiddle_rsc_0_2_i_adra;
  twiddle_rsc_0_2_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_2_i_adra_d;
  twiddle_rsc_0_2_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_2_i_qa_d <= twiddle_rsc_0_2_i_qa_d_1;
  twiddle_rsc_0_2_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_3_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_74_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_3_i_qb,
      web => twiddle_rsc_0_3_web,
      db => twiddle_rsc_0_3_i_db,
      adrb => twiddle_rsc_0_3_i_adrb,
      qa => twiddle_rsc_0_3_i_qa,
      wea => twiddle_rsc_0_3_wea,
      da => twiddle_rsc_0_3_i_da,
      adra => twiddle_rsc_0_3_i_adra,
      adra_d => twiddle_rsc_0_3_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_3_i_da_d,
      qa_d => twiddle_rsc_0_3_i_qa_d_1,
      wea_d => twiddle_rsc_0_3_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_3_i_qb <= twiddle_rsc_0_3_qb;
  twiddle_rsc_0_3_db <= twiddle_rsc_0_3_i_db;
  twiddle_rsc_0_3_adrb <= twiddle_rsc_0_3_i_adrb;
  twiddle_rsc_0_3_i_qa <= twiddle_rsc_0_3_qa;
  twiddle_rsc_0_3_da <= twiddle_rsc_0_3_i_da;
  twiddle_rsc_0_3_adra <= twiddle_rsc_0_3_i_adra;
  twiddle_rsc_0_3_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_3_i_adra_d;
  twiddle_rsc_0_3_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_3_i_qa_d <= twiddle_rsc_0_3_i_qa_d_1;
  twiddle_rsc_0_3_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_4_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_75_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_4_i_qb,
      web => twiddle_rsc_0_4_web,
      db => twiddle_rsc_0_4_i_db,
      adrb => twiddle_rsc_0_4_i_adrb,
      qa => twiddle_rsc_0_4_i_qa,
      wea => twiddle_rsc_0_4_wea,
      da => twiddle_rsc_0_4_i_da,
      adra => twiddle_rsc_0_4_i_adra,
      adra_d => twiddle_rsc_0_4_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_4_i_da_d,
      qa_d => twiddle_rsc_0_4_i_qa_d_1,
      wea_d => twiddle_rsc_0_4_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_4_i_qb <= twiddle_rsc_0_4_qb;
  twiddle_rsc_0_4_db <= twiddle_rsc_0_4_i_db;
  twiddle_rsc_0_4_adrb <= twiddle_rsc_0_4_i_adrb;
  twiddle_rsc_0_4_i_qa <= twiddle_rsc_0_4_qa;
  twiddle_rsc_0_4_da <= twiddle_rsc_0_4_i_da;
  twiddle_rsc_0_4_adra <= twiddle_rsc_0_4_i_adra;
  twiddle_rsc_0_4_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_4_i_adra_d;
  twiddle_rsc_0_4_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_4_i_qa_d <= twiddle_rsc_0_4_i_qa_d_1;
  twiddle_rsc_0_4_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_5_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_76_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_5_i_qb,
      web => twiddle_rsc_0_5_web,
      db => twiddle_rsc_0_5_i_db,
      adrb => twiddle_rsc_0_5_i_adrb,
      qa => twiddle_rsc_0_5_i_qa,
      wea => twiddle_rsc_0_5_wea,
      da => twiddle_rsc_0_5_i_da,
      adra => twiddle_rsc_0_5_i_adra,
      adra_d => twiddle_rsc_0_5_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_5_i_da_d,
      qa_d => twiddle_rsc_0_5_i_qa_d_1,
      wea_d => twiddle_rsc_0_5_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_5_i_qb <= twiddle_rsc_0_5_qb;
  twiddle_rsc_0_5_db <= twiddle_rsc_0_5_i_db;
  twiddle_rsc_0_5_adrb <= twiddle_rsc_0_5_i_adrb;
  twiddle_rsc_0_5_i_qa <= twiddle_rsc_0_5_qa;
  twiddle_rsc_0_5_da <= twiddle_rsc_0_5_i_da;
  twiddle_rsc_0_5_adra <= twiddle_rsc_0_5_i_adra;
  twiddle_rsc_0_5_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_5_i_adra_d;
  twiddle_rsc_0_5_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_5_i_qa_d <= twiddle_rsc_0_5_i_qa_d_1;
  twiddle_rsc_0_5_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_6_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_77_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_6_i_qb,
      web => twiddle_rsc_0_6_web,
      db => twiddle_rsc_0_6_i_db,
      adrb => twiddle_rsc_0_6_i_adrb,
      qa => twiddle_rsc_0_6_i_qa,
      wea => twiddle_rsc_0_6_wea,
      da => twiddle_rsc_0_6_i_da,
      adra => twiddle_rsc_0_6_i_adra,
      adra_d => twiddle_rsc_0_6_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_6_i_da_d,
      qa_d => twiddle_rsc_0_6_i_qa_d_1,
      wea_d => twiddle_rsc_0_6_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_6_i_qb <= twiddle_rsc_0_6_qb;
  twiddle_rsc_0_6_db <= twiddle_rsc_0_6_i_db;
  twiddle_rsc_0_6_adrb <= twiddle_rsc_0_6_i_adrb;
  twiddle_rsc_0_6_i_qa <= twiddle_rsc_0_6_qa;
  twiddle_rsc_0_6_da <= twiddle_rsc_0_6_i_da;
  twiddle_rsc_0_6_adra <= twiddle_rsc_0_6_i_adra;
  twiddle_rsc_0_6_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_6_i_adra_d;
  twiddle_rsc_0_6_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_6_i_qa_d <= twiddle_rsc_0_6_i_qa_d_1;
  twiddle_rsc_0_6_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_7_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_78_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_7_i_qb,
      web => twiddle_rsc_0_7_web,
      db => twiddle_rsc_0_7_i_db,
      adrb => twiddle_rsc_0_7_i_adrb,
      qa => twiddle_rsc_0_7_i_qa,
      wea => twiddle_rsc_0_7_wea,
      da => twiddle_rsc_0_7_i_da,
      adra => twiddle_rsc_0_7_i_adra,
      adra_d => twiddle_rsc_0_7_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_7_i_da_d,
      qa_d => twiddle_rsc_0_7_i_qa_d_1,
      wea_d => twiddle_rsc_0_7_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_7_i_qb <= twiddle_rsc_0_7_qb;
  twiddle_rsc_0_7_db <= twiddle_rsc_0_7_i_db;
  twiddle_rsc_0_7_adrb <= twiddle_rsc_0_7_i_adrb;
  twiddle_rsc_0_7_i_qa <= twiddle_rsc_0_7_qa;
  twiddle_rsc_0_7_da <= twiddle_rsc_0_7_i_da;
  twiddle_rsc_0_7_adra <= twiddle_rsc_0_7_i_adra;
  twiddle_rsc_0_7_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_7_i_adra_d;
  twiddle_rsc_0_7_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_7_i_qa_d <= twiddle_rsc_0_7_i_qa_d_1;
  twiddle_rsc_0_7_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_8_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_79_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_8_i_qb,
      web => twiddle_rsc_0_8_web,
      db => twiddle_rsc_0_8_i_db,
      adrb => twiddle_rsc_0_8_i_adrb,
      qa => twiddle_rsc_0_8_i_qa,
      wea => twiddle_rsc_0_8_wea,
      da => twiddle_rsc_0_8_i_da,
      adra => twiddle_rsc_0_8_i_adra,
      adra_d => twiddle_rsc_0_8_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_8_i_da_d,
      qa_d => twiddle_rsc_0_8_i_qa_d_1,
      wea_d => twiddle_rsc_0_8_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_8_i_qb <= twiddle_rsc_0_8_qb;
  twiddle_rsc_0_8_db <= twiddle_rsc_0_8_i_db;
  twiddle_rsc_0_8_adrb <= twiddle_rsc_0_8_i_adrb;
  twiddle_rsc_0_8_i_qa <= twiddle_rsc_0_8_qa;
  twiddle_rsc_0_8_da <= twiddle_rsc_0_8_i_da;
  twiddle_rsc_0_8_adra <= twiddle_rsc_0_8_i_adra;
  twiddle_rsc_0_8_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_8_i_adra_d;
  twiddle_rsc_0_8_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_8_i_qa_d <= twiddle_rsc_0_8_i_qa_d_1;
  twiddle_rsc_0_8_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_9_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_80_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_9_i_qb,
      web => twiddle_rsc_0_9_web,
      db => twiddle_rsc_0_9_i_db,
      adrb => twiddle_rsc_0_9_i_adrb,
      qa => twiddle_rsc_0_9_i_qa,
      wea => twiddle_rsc_0_9_wea,
      da => twiddle_rsc_0_9_i_da,
      adra => twiddle_rsc_0_9_i_adra,
      adra_d => twiddle_rsc_0_9_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_9_i_da_d,
      qa_d => twiddle_rsc_0_9_i_qa_d_1,
      wea_d => twiddle_rsc_0_9_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_9_i_qb <= twiddle_rsc_0_9_qb;
  twiddle_rsc_0_9_db <= twiddle_rsc_0_9_i_db;
  twiddle_rsc_0_9_adrb <= twiddle_rsc_0_9_i_adrb;
  twiddle_rsc_0_9_i_qa <= twiddle_rsc_0_9_qa;
  twiddle_rsc_0_9_da <= twiddle_rsc_0_9_i_da;
  twiddle_rsc_0_9_adra <= twiddle_rsc_0_9_i_adra;
  twiddle_rsc_0_9_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_9_i_adra_d;
  twiddle_rsc_0_9_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_9_i_qa_d <= twiddle_rsc_0_9_i_qa_d_1;
  twiddle_rsc_0_9_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_10_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_81_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_10_i_qb,
      web => twiddle_rsc_0_10_web,
      db => twiddle_rsc_0_10_i_db,
      adrb => twiddle_rsc_0_10_i_adrb,
      qa => twiddle_rsc_0_10_i_qa,
      wea => twiddle_rsc_0_10_wea,
      da => twiddle_rsc_0_10_i_da,
      adra => twiddle_rsc_0_10_i_adra,
      adra_d => twiddle_rsc_0_10_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_10_i_da_d,
      qa_d => twiddle_rsc_0_10_i_qa_d_1,
      wea_d => twiddle_rsc_0_10_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_10_i_qb <= twiddle_rsc_0_10_qb;
  twiddle_rsc_0_10_db <= twiddle_rsc_0_10_i_db;
  twiddle_rsc_0_10_adrb <= twiddle_rsc_0_10_i_adrb;
  twiddle_rsc_0_10_i_qa <= twiddle_rsc_0_10_qa;
  twiddle_rsc_0_10_da <= twiddle_rsc_0_10_i_da;
  twiddle_rsc_0_10_adra <= twiddle_rsc_0_10_i_adra;
  twiddle_rsc_0_10_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_10_i_adra_d;
  twiddle_rsc_0_10_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_10_i_qa_d <= twiddle_rsc_0_10_i_qa_d_1;
  twiddle_rsc_0_10_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_11_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_82_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_11_i_qb,
      web => twiddle_rsc_0_11_web,
      db => twiddle_rsc_0_11_i_db,
      adrb => twiddle_rsc_0_11_i_adrb,
      qa => twiddle_rsc_0_11_i_qa,
      wea => twiddle_rsc_0_11_wea,
      da => twiddle_rsc_0_11_i_da,
      adra => twiddle_rsc_0_11_i_adra,
      adra_d => twiddle_rsc_0_11_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_11_i_da_d,
      qa_d => twiddle_rsc_0_11_i_qa_d_1,
      wea_d => twiddle_rsc_0_11_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_11_i_qb <= twiddle_rsc_0_11_qb;
  twiddle_rsc_0_11_db <= twiddle_rsc_0_11_i_db;
  twiddle_rsc_0_11_adrb <= twiddle_rsc_0_11_i_adrb;
  twiddle_rsc_0_11_i_qa <= twiddle_rsc_0_11_qa;
  twiddle_rsc_0_11_da <= twiddle_rsc_0_11_i_da;
  twiddle_rsc_0_11_adra <= twiddle_rsc_0_11_i_adra;
  twiddle_rsc_0_11_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_11_i_adra_d;
  twiddle_rsc_0_11_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_11_i_qa_d <= twiddle_rsc_0_11_i_qa_d_1;
  twiddle_rsc_0_11_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_12_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_83_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_12_i_qb,
      web => twiddle_rsc_0_12_web,
      db => twiddle_rsc_0_12_i_db,
      adrb => twiddle_rsc_0_12_i_adrb,
      qa => twiddle_rsc_0_12_i_qa,
      wea => twiddle_rsc_0_12_wea,
      da => twiddle_rsc_0_12_i_da,
      adra => twiddle_rsc_0_12_i_adra,
      adra_d => twiddle_rsc_0_12_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_12_i_da_d,
      qa_d => twiddle_rsc_0_12_i_qa_d_1,
      wea_d => twiddle_rsc_0_12_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_12_i_qb <= twiddle_rsc_0_12_qb;
  twiddle_rsc_0_12_db <= twiddle_rsc_0_12_i_db;
  twiddle_rsc_0_12_adrb <= twiddle_rsc_0_12_i_adrb;
  twiddle_rsc_0_12_i_qa <= twiddle_rsc_0_12_qa;
  twiddle_rsc_0_12_da <= twiddle_rsc_0_12_i_da;
  twiddle_rsc_0_12_adra <= twiddle_rsc_0_12_i_adra;
  twiddle_rsc_0_12_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_12_i_adra_d;
  twiddle_rsc_0_12_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_12_i_qa_d <= twiddle_rsc_0_12_i_qa_d_1;
  twiddle_rsc_0_12_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_13_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_84_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_13_i_qb,
      web => twiddle_rsc_0_13_web,
      db => twiddle_rsc_0_13_i_db,
      adrb => twiddle_rsc_0_13_i_adrb,
      qa => twiddle_rsc_0_13_i_qa,
      wea => twiddle_rsc_0_13_wea,
      da => twiddle_rsc_0_13_i_da,
      adra => twiddle_rsc_0_13_i_adra,
      adra_d => twiddle_rsc_0_13_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_13_i_da_d,
      qa_d => twiddle_rsc_0_13_i_qa_d_1,
      wea_d => twiddle_rsc_0_13_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_13_i_qb <= twiddle_rsc_0_13_qb;
  twiddle_rsc_0_13_db <= twiddle_rsc_0_13_i_db;
  twiddle_rsc_0_13_adrb <= twiddle_rsc_0_13_i_adrb;
  twiddle_rsc_0_13_i_qa <= twiddle_rsc_0_13_qa;
  twiddle_rsc_0_13_da <= twiddle_rsc_0_13_i_da;
  twiddle_rsc_0_13_adra <= twiddle_rsc_0_13_i_adra;
  twiddle_rsc_0_13_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_13_i_adra_d;
  twiddle_rsc_0_13_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_13_i_qa_d <= twiddle_rsc_0_13_i_qa_d_1;
  twiddle_rsc_0_13_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_14_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_85_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_14_i_qb,
      web => twiddle_rsc_0_14_web,
      db => twiddle_rsc_0_14_i_db,
      adrb => twiddle_rsc_0_14_i_adrb,
      qa => twiddle_rsc_0_14_i_qa,
      wea => twiddle_rsc_0_14_wea,
      da => twiddle_rsc_0_14_i_da,
      adra => twiddle_rsc_0_14_i_adra,
      adra_d => twiddle_rsc_0_14_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_14_i_da_d,
      qa_d => twiddle_rsc_0_14_i_qa_d_1,
      wea_d => twiddle_rsc_0_14_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_14_i_qb <= twiddle_rsc_0_14_qb;
  twiddle_rsc_0_14_db <= twiddle_rsc_0_14_i_db;
  twiddle_rsc_0_14_adrb <= twiddle_rsc_0_14_i_adrb;
  twiddle_rsc_0_14_i_qa <= twiddle_rsc_0_14_qa;
  twiddle_rsc_0_14_da <= twiddle_rsc_0_14_i_da;
  twiddle_rsc_0_14_adra <= twiddle_rsc_0_14_i_adra;
  twiddle_rsc_0_14_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_14_i_adra_d;
  twiddle_rsc_0_14_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_14_i_qa_d <= twiddle_rsc_0_14_i_qa_d_1;
  twiddle_rsc_0_14_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_rsc_0_15_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_86_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_15_i_qb,
      web => twiddle_rsc_0_15_web,
      db => twiddle_rsc_0_15_i_db,
      adrb => twiddle_rsc_0_15_i_adrb,
      qa => twiddle_rsc_0_15_i_qa,
      wea => twiddle_rsc_0_15_wea,
      da => twiddle_rsc_0_15_i_da,
      adra => twiddle_rsc_0_15_i_adra,
      adra_d => twiddle_rsc_0_15_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_rsc_0_15_i_da_d,
      qa_d => twiddle_rsc_0_15_i_qa_d_1,
      wea_d => twiddle_rsc_0_15_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_rsc_0_15_i_qb <= twiddle_rsc_0_15_qb;
  twiddle_rsc_0_15_db <= twiddle_rsc_0_15_i_db;
  twiddle_rsc_0_15_adrb <= twiddle_rsc_0_15_i_adrb;
  twiddle_rsc_0_15_i_qa <= twiddle_rsc_0_15_qa;
  twiddle_rsc_0_15_da <= twiddle_rsc_0_15_i_da;
  twiddle_rsc_0_15_adra <= twiddle_rsc_0_15_i_adra;
  twiddle_rsc_0_15_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_rsc_0_15_i_adra_d;
  twiddle_rsc_0_15_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_rsc_0_15_i_qa_d <= twiddle_rsc_0_15_i_qa_d_1;
  twiddle_rsc_0_15_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_0_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_87_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_0_i_qb,
      web => twiddle_h_rsc_0_0_web,
      db => twiddle_h_rsc_0_0_i_db,
      adrb => twiddle_h_rsc_0_0_i_adrb,
      qa => twiddle_h_rsc_0_0_i_qa,
      wea => twiddle_h_rsc_0_0_wea,
      da => twiddle_h_rsc_0_0_i_da,
      adra => twiddle_h_rsc_0_0_i_adra,
      adra_d => twiddle_h_rsc_0_0_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_0_i_da_d,
      qa_d => twiddle_h_rsc_0_0_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_0_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_0_i_qb <= twiddle_h_rsc_0_0_qb;
  twiddle_h_rsc_0_0_db <= twiddle_h_rsc_0_0_i_db;
  twiddle_h_rsc_0_0_adrb <= twiddle_h_rsc_0_0_i_adrb;
  twiddle_h_rsc_0_0_i_qa <= twiddle_h_rsc_0_0_qa;
  twiddle_h_rsc_0_0_da <= twiddle_h_rsc_0_0_i_da;
  twiddle_h_rsc_0_0_adra <= twiddle_h_rsc_0_0_i_adra;
  twiddle_h_rsc_0_0_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_0_i_adra_d;
  twiddle_h_rsc_0_0_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_0_i_qa_d <= twiddle_h_rsc_0_0_i_qa_d_1;
  twiddle_h_rsc_0_0_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_1_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_88_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_1_i_qb,
      web => twiddle_h_rsc_0_1_web,
      db => twiddle_h_rsc_0_1_i_db,
      adrb => twiddle_h_rsc_0_1_i_adrb,
      qa => twiddle_h_rsc_0_1_i_qa,
      wea => twiddle_h_rsc_0_1_wea,
      da => twiddle_h_rsc_0_1_i_da,
      adra => twiddle_h_rsc_0_1_i_adra,
      adra_d => twiddle_h_rsc_0_1_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_1_i_da_d,
      qa_d => twiddle_h_rsc_0_1_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_1_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_1_i_qb <= twiddle_h_rsc_0_1_qb;
  twiddle_h_rsc_0_1_db <= twiddle_h_rsc_0_1_i_db;
  twiddle_h_rsc_0_1_adrb <= twiddle_h_rsc_0_1_i_adrb;
  twiddle_h_rsc_0_1_i_qa <= twiddle_h_rsc_0_1_qa;
  twiddle_h_rsc_0_1_da <= twiddle_h_rsc_0_1_i_da;
  twiddle_h_rsc_0_1_adra <= twiddle_h_rsc_0_1_i_adra;
  twiddle_h_rsc_0_1_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_1_i_adra_d;
  twiddle_h_rsc_0_1_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_1_i_qa_d <= twiddle_h_rsc_0_1_i_qa_d_1;
  twiddle_h_rsc_0_1_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_2_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_89_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_2_i_qb,
      web => twiddle_h_rsc_0_2_web,
      db => twiddle_h_rsc_0_2_i_db,
      adrb => twiddle_h_rsc_0_2_i_adrb,
      qa => twiddle_h_rsc_0_2_i_qa,
      wea => twiddle_h_rsc_0_2_wea,
      da => twiddle_h_rsc_0_2_i_da,
      adra => twiddle_h_rsc_0_2_i_adra,
      adra_d => twiddle_h_rsc_0_2_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_2_i_da_d,
      qa_d => twiddle_h_rsc_0_2_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_2_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_2_i_qb <= twiddle_h_rsc_0_2_qb;
  twiddle_h_rsc_0_2_db <= twiddle_h_rsc_0_2_i_db;
  twiddle_h_rsc_0_2_adrb <= twiddle_h_rsc_0_2_i_adrb;
  twiddle_h_rsc_0_2_i_qa <= twiddle_h_rsc_0_2_qa;
  twiddle_h_rsc_0_2_da <= twiddle_h_rsc_0_2_i_da;
  twiddle_h_rsc_0_2_adra <= twiddle_h_rsc_0_2_i_adra;
  twiddle_h_rsc_0_2_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_2_i_adra_d;
  twiddle_h_rsc_0_2_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_2_i_qa_d <= twiddle_h_rsc_0_2_i_qa_d_1;
  twiddle_h_rsc_0_2_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_3_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_90_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_3_i_qb,
      web => twiddle_h_rsc_0_3_web,
      db => twiddle_h_rsc_0_3_i_db,
      adrb => twiddle_h_rsc_0_3_i_adrb,
      qa => twiddle_h_rsc_0_3_i_qa,
      wea => twiddle_h_rsc_0_3_wea,
      da => twiddle_h_rsc_0_3_i_da,
      adra => twiddle_h_rsc_0_3_i_adra,
      adra_d => twiddle_h_rsc_0_3_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_3_i_da_d,
      qa_d => twiddle_h_rsc_0_3_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_3_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_3_i_qb <= twiddle_h_rsc_0_3_qb;
  twiddle_h_rsc_0_3_db <= twiddle_h_rsc_0_3_i_db;
  twiddle_h_rsc_0_3_adrb <= twiddle_h_rsc_0_3_i_adrb;
  twiddle_h_rsc_0_3_i_qa <= twiddle_h_rsc_0_3_qa;
  twiddle_h_rsc_0_3_da <= twiddle_h_rsc_0_3_i_da;
  twiddle_h_rsc_0_3_adra <= twiddle_h_rsc_0_3_i_adra;
  twiddle_h_rsc_0_3_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_3_i_adra_d;
  twiddle_h_rsc_0_3_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_3_i_qa_d <= twiddle_h_rsc_0_3_i_qa_d_1;
  twiddle_h_rsc_0_3_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_4_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_91_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_4_i_qb,
      web => twiddle_h_rsc_0_4_web,
      db => twiddle_h_rsc_0_4_i_db,
      adrb => twiddle_h_rsc_0_4_i_adrb,
      qa => twiddle_h_rsc_0_4_i_qa,
      wea => twiddle_h_rsc_0_4_wea,
      da => twiddle_h_rsc_0_4_i_da,
      adra => twiddle_h_rsc_0_4_i_adra,
      adra_d => twiddle_h_rsc_0_4_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_4_i_da_d,
      qa_d => twiddle_h_rsc_0_4_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_4_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_4_i_qb <= twiddle_h_rsc_0_4_qb;
  twiddle_h_rsc_0_4_db <= twiddle_h_rsc_0_4_i_db;
  twiddle_h_rsc_0_4_adrb <= twiddle_h_rsc_0_4_i_adrb;
  twiddle_h_rsc_0_4_i_qa <= twiddle_h_rsc_0_4_qa;
  twiddle_h_rsc_0_4_da <= twiddle_h_rsc_0_4_i_da;
  twiddle_h_rsc_0_4_adra <= twiddle_h_rsc_0_4_i_adra;
  twiddle_h_rsc_0_4_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_4_i_adra_d;
  twiddle_h_rsc_0_4_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_4_i_qa_d <= twiddle_h_rsc_0_4_i_qa_d_1;
  twiddle_h_rsc_0_4_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_5_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_92_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_5_i_qb,
      web => twiddle_h_rsc_0_5_web,
      db => twiddle_h_rsc_0_5_i_db,
      adrb => twiddle_h_rsc_0_5_i_adrb,
      qa => twiddle_h_rsc_0_5_i_qa,
      wea => twiddle_h_rsc_0_5_wea,
      da => twiddle_h_rsc_0_5_i_da,
      adra => twiddle_h_rsc_0_5_i_adra,
      adra_d => twiddle_h_rsc_0_5_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_5_i_da_d,
      qa_d => twiddle_h_rsc_0_5_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_5_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_5_i_qb <= twiddle_h_rsc_0_5_qb;
  twiddle_h_rsc_0_5_db <= twiddle_h_rsc_0_5_i_db;
  twiddle_h_rsc_0_5_adrb <= twiddle_h_rsc_0_5_i_adrb;
  twiddle_h_rsc_0_5_i_qa <= twiddle_h_rsc_0_5_qa;
  twiddle_h_rsc_0_5_da <= twiddle_h_rsc_0_5_i_da;
  twiddle_h_rsc_0_5_adra <= twiddle_h_rsc_0_5_i_adra;
  twiddle_h_rsc_0_5_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_5_i_adra_d;
  twiddle_h_rsc_0_5_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_5_i_qa_d <= twiddle_h_rsc_0_5_i_qa_d_1;
  twiddle_h_rsc_0_5_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_6_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_93_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_6_i_qb,
      web => twiddle_h_rsc_0_6_web,
      db => twiddle_h_rsc_0_6_i_db,
      adrb => twiddle_h_rsc_0_6_i_adrb,
      qa => twiddle_h_rsc_0_6_i_qa,
      wea => twiddle_h_rsc_0_6_wea,
      da => twiddle_h_rsc_0_6_i_da,
      adra => twiddle_h_rsc_0_6_i_adra,
      adra_d => twiddle_h_rsc_0_6_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_6_i_da_d,
      qa_d => twiddle_h_rsc_0_6_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_6_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_6_i_qb <= twiddle_h_rsc_0_6_qb;
  twiddle_h_rsc_0_6_db <= twiddle_h_rsc_0_6_i_db;
  twiddle_h_rsc_0_6_adrb <= twiddle_h_rsc_0_6_i_adrb;
  twiddle_h_rsc_0_6_i_qa <= twiddle_h_rsc_0_6_qa;
  twiddle_h_rsc_0_6_da <= twiddle_h_rsc_0_6_i_da;
  twiddle_h_rsc_0_6_adra <= twiddle_h_rsc_0_6_i_adra;
  twiddle_h_rsc_0_6_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_6_i_adra_d;
  twiddle_h_rsc_0_6_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_6_i_qa_d <= twiddle_h_rsc_0_6_i_qa_d_1;
  twiddle_h_rsc_0_6_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_7_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_94_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_7_i_qb,
      web => twiddle_h_rsc_0_7_web,
      db => twiddle_h_rsc_0_7_i_db,
      adrb => twiddle_h_rsc_0_7_i_adrb,
      qa => twiddle_h_rsc_0_7_i_qa,
      wea => twiddle_h_rsc_0_7_wea,
      da => twiddle_h_rsc_0_7_i_da,
      adra => twiddle_h_rsc_0_7_i_adra,
      adra_d => twiddle_h_rsc_0_7_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_7_i_da_d,
      qa_d => twiddle_h_rsc_0_7_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_7_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_7_i_qb <= twiddle_h_rsc_0_7_qb;
  twiddle_h_rsc_0_7_db <= twiddle_h_rsc_0_7_i_db;
  twiddle_h_rsc_0_7_adrb <= twiddle_h_rsc_0_7_i_adrb;
  twiddle_h_rsc_0_7_i_qa <= twiddle_h_rsc_0_7_qa;
  twiddle_h_rsc_0_7_da <= twiddle_h_rsc_0_7_i_da;
  twiddle_h_rsc_0_7_adra <= twiddle_h_rsc_0_7_i_adra;
  twiddle_h_rsc_0_7_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_7_i_adra_d;
  twiddle_h_rsc_0_7_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_7_i_qa_d <= twiddle_h_rsc_0_7_i_qa_d_1;
  twiddle_h_rsc_0_7_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_8_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_95_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_8_i_qb,
      web => twiddle_h_rsc_0_8_web,
      db => twiddle_h_rsc_0_8_i_db,
      adrb => twiddle_h_rsc_0_8_i_adrb,
      qa => twiddle_h_rsc_0_8_i_qa,
      wea => twiddle_h_rsc_0_8_wea,
      da => twiddle_h_rsc_0_8_i_da,
      adra => twiddle_h_rsc_0_8_i_adra,
      adra_d => twiddle_h_rsc_0_8_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_8_i_da_d,
      qa_d => twiddle_h_rsc_0_8_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_8_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_8_i_qb <= twiddle_h_rsc_0_8_qb;
  twiddle_h_rsc_0_8_db <= twiddle_h_rsc_0_8_i_db;
  twiddle_h_rsc_0_8_adrb <= twiddle_h_rsc_0_8_i_adrb;
  twiddle_h_rsc_0_8_i_qa <= twiddle_h_rsc_0_8_qa;
  twiddle_h_rsc_0_8_da <= twiddle_h_rsc_0_8_i_da;
  twiddle_h_rsc_0_8_adra <= twiddle_h_rsc_0_8_i_adra;
  twiddle_h_rsc_0_8_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_8_i_adra_d;
  twiddle_h_rsc_0_8_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_8_i_qa_d <= twiddle_h_rsc_0_8_i_qa_d_1;
  twiddle_h_rsc_0_8_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_9_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_96_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_9_i_qb,
      web => twiddle_h_rsc_0_9_web,
      db => twiddle_h_rsc_0_9_i_db,
      adrb => twiddle_h_rsc_0_9_i_adrb,
      qa => twiddle_h_rsc_0_9_i_qa,
      wea => twiddle_h_rsc_0_9_wea,
      da => twiddle_h_rsc_0_9_i_da,
      adra => twiddle_h_rsc_0_9_i_adra,
      adra_d => twiddle_h_rsc_0_9_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_9_i_da_d,
      qa_d => twiddle_h_rsc_0_9_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_9_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_9_i_qb <= twiddle_h_rsc_0_9_qb;
  twiddle_h_rsc_0_9_db <= twiddle_h_rsc_0_9_i_db;
  twiddle_h_rsc_0_9_adrb <= twiddle_h_rsc_0_9_i_adrb;
  twiddle_h_rsc_0_9_i_qa <= twiddle_h_rsc_0_9_qa;
  twiddle_h_rsc_0_9_da <= twiddle_h_rsc_0_9_i_da;
  twiddle_h_rsc_0_9_adra <= twiddle_h_rsc_0_9_i_adra;
  twiddle_h_rsc_0_9_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_9_i_adra_d;
  twiddle_h_rsc_0_9_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_9_i_qa_d <= twiddle_h_rsc_0_9_i_qa_d_1;
  twiddle_h_rsc_0_9_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_10_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_97_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_10_i_qb,
      web => twiddle_h_rsc_0_10_web,
      db => twiddle_h_rsc_0_10_i_db,
      adrb => twiddle_h_rsc_0_10_i_adrb,
      qa => twiddle_h_rsc_0_10_i_qa,
      wea => twiddle_h_rsc_0_10_wea,
      da => twiddle_h_rsc_0_10_i_da,
      adra => twiddle_h_rsc_0_10_i_adra,
      adra_d => twiddle_h_rsc_0_10_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_10_i_da_d,
      qa_d => twiddle_h_rsc_0_10_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_10_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_10_i_qb <= twiddle_h_rsc_0_10_qb;
  twiddle_h_rsc_0_10_db <= twiddle_h_rsc_0_10_i_db;
  twiddle_h_rsc_0_10_adrb <= twiddle_h_rsc_0_10_i_adrb;
  twiddle_h_rsc_0_10_i_qa <= twiddle_h_rsc_0_10_qa;
  twiddle_h_rsc_0_10_da <= twiddle_h_rsc_0_10_i_da;
  twiddle_h_rsc_0_10_adra <= twiddle_h_rsc_0_10_i_adra;
  twiddle_h_rsc_0_10_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_10_i_adra_d;
  twiddle_h_rsc_0_10_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_10_i_qa_d <= twiddle_h_rsc_0_10_i_qa_d_1;
  twiddle_h_rsc_0_10_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_11_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_98_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_11_i_qb,
      web => twiddle_h_rsc_0_11_web,
      db => twiddle_h_rsc_0_11_i_db,
      adrb => twiddle_h_rsc_0_11_i_adrb,
      qa => twiddle_h_rsc_0_11_i_qa,
      wea => twiddle_h_rsc_0_11_wea,
      da => twiddle_h_rsc_0_11_i_da,
      adra => twiddle_h_rsc_0_11_i_adra,
      adra_d => twiddle_h_rsc_0_11_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_11_i_da_d,
      qa_d => twiddle_h_rsc_0_11_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_11_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_11_i_qb <= twiddle_h_rsc_0_11_qb;
  twiddle_h_rsc_0_11_db <= twiddle_h_rsc_0_11_i_db;
  twiddle_h_rsc_0_11_adrb <= twiddle_h_rsc_0_11_i_adrb;
  twiddle_h_rsc_0_11_i_qa <= twiddle_h_rsc_0_11_qa;
  twiddle_h_rsc_0_11_da <= twiddle_h_rsc_0_11_i_da;
  twiddle_h_rsc_0_11_adra <= twiddle_h_rsc_0_11_i_adra;
  twiddle_h_rsc_0_11_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_11_i_adra_d;
  twiddle_h_rsc_0_11_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_11_i_qa_d <= twiddle_h_rsc_0_11_i_qa_d_1;
  twiddle_h_rsc_0_11_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_12_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_99_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_12_i_qb,
      web => twiddle_h_rsc_0_12_web,
      db => twiddle_h_rsc_0_12_i_db,
      adrb => twiddle_h_rsc_0_12_i_adrb,
      qa => twiddle_h_rsc_0_12_i_qa,
      wea => twiddle_h_rsc_0_12_wea,
      da => twiddle_h_rsc_0_12_i_da,
      adra => twiddle_h_rsc_0_12_i_adra,
      adra_d => twiddle_h_rsc_0_12_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_12_i_da_d,
      qa_d => twiddle_h_rsc_0_12_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_12_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_12_i_qb <= twiddle_h_rsc_0_12_qb;
  twiddle_h_rsc_0_12_db <= twiddle_h_rsc_0_12_i_db;
  twiddle_h_rsc_0_12_adrb <= twiddle_h_rsc_0_12_i_adrb;
  twiddle_h_rsc_0_12_i_qa <= twiddle_h_rsc_0_12_qa;
  twiddle_h_rsc_0_12_da <= twiddle_h_rsc_0_12_i_da;
  twiddle_h_rsc_0_12_adra <= twiddle_h_rsc_0_12_i_adra;
  twiddle_h_rsc_0_12_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_12_i_adra_d;
  twiddle_h_rsc_0_12_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_12_i_qa_d <= twiddle_h_rsc_0_12_i_qa_d_1;
  twiddle_h_rsc_0_12_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_13_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_100_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_13_i_qb,
      web => twiddle_h_rsc_0_13_web,
      db => twiddle_h_rsc_0_13_i_db,
      adrb => twiddle_h_rsc_0_13_i_adrb,
      qa => twiddle_h_rsc_0_13_i_qa,
      wea => twiddle_h_rsc_0_13_wea,
      da => twiddle_h_rsc_0_13_i_da,
      adra => twiddle_h_rsc_0_13_i_adra,
      adra_d => twiddle_h_rsc_0_13_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_13_i_da_d,
      qa_d => twiddle_h_rsc_0_13_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_13_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_13_i_qb <= twiddle_h_rsc_0_13_qb;
  twiddle_h_rsc_0_13_db <= twiddle_h_rsc_0_13_i_db;
  twiddle_h_rsc_0_13_adrb <= twiddle_h_rsc_0_13_i_adrb;
  twiddle_h_rsc_0_13_i_qa <= twiddle_h_rsc_0_13_qa;
  twiddle_h_rsc_0_13_da <= twiddle_h_rsc_0_13_i_da;
  twiddle_h_rsc_0_13_adra <= twiddle_h_rsc_0_13_i_adra;
  twiddle_h_rsc_0_13_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_13_i_adra_d;
  twiddle_h_rsc_0_13_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_13_i_qa_d <= twiddle_h_rsc_0_13_i_qa_d_1;
  twiddle_h_rsc_0_13_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_14_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_101_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_14_i_qb,
      web => twiddle_h_rsc_0_14_web,
      db => twiddle_h_rsc_0_14_i_db,
      adrb => twiddle_h_rsc_0_14_i_adrb,
      qa => twiddle_h_rsc_0_14_i_qa,
      wea => twiddle_h_rsc_0_14_wea,
      da => twiddle_h_rsc_0_14_i_da,
      adra => twiddle_h_rsc_0_14_i_adra,
      adra_d => twiddle_h_rsc_0_14_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_14_i_da_d,
      qa_d => twiddle_h_rsc_0_14_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_14_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_14_i_qb <= twiddle_h_rsc_0_14_qb;
  twiddle_h_rsc_0_14_db <= twiddle_h_rsc_0_14_i_db;
  twiddle_h_rsc_0_14_adrb <= twiddle_h_rsc_0_14_i_adrb;
  twiddle_h_rsc_0_14_i_qa <= twiddle_h_rsc_0_14_qa;
  twiddle_h_rsc_0_14_da <= twiddle_h_rsc_0_14_i_da;
  twiddle_h_rsc_0_14_adra <= twiddle_h_rsc_0_14_i_adra;
  twiddle_h_rsc_0_14_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_14_i_adra_d;
  twiddle_h_rsc_0_14_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_14_i_qa_d <= twiddle_h_rsc_0_14_i_qa_d_1;
  twiddle_h_rsc_0_14_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  twiddle_h_rsc_0_15_i : peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_102_8_32_256_256_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_15_i_qb,
      web => twiddle_h_rsc_0_15_web,
      db => twiddle_h_rsc_0_15_i_db,
      adrb => twiddle_h_rsc_0_15_i_adrb,
      qa => twiddle_h_rsc_0_15_i_qa,
      wea => twiddle_h_rsc_0_15_wea,
      da => twiddle_h_rsc_0_15_i_da,
      adra => twiddle_h_rsc_0_15_i_adra,
      adra_d => twiddle_h_rsc_0_15_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => twiddle_h_rsc_0_15_i_da_d,
      qa_d => twiddle_h_rsc_0_15_i_qa_d_1,
      wea_d => twiddle_h_rsc_0_15_i_wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d
    );
  twiddle_h_rsc_0_15_i_qb <= twiddle_h_rsc_0_15_qb;
  twiddle_h_rsc_0_15_db <= twiddle_h_rsc_0_15_i_db;
  twiddle_h_rsc_0_15_adrb <= twiddle_h_rsc_0_15_i_adrb;
  twiddle_h_rsc_0_15_i_qa <= twiddle_h_rsc_0_15_qa;
  twiddle_h_rsc_0_15_da <= twiddle_h_rsc_0_15_i_da;
  twiddle_h_rsc_0_15_adra <= twiddle_h_rsc_0_15_i_adra;
  twiddle_h_rsc_0_15_i_adra_d_1 <= STD_LOGIC_VECTOR'( "00000000") & twiddle_h_rsc_0_15_i_adra_d;
  twiddle_h_rsc_0_15_i_da_d <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
  twiddle_h_rsc_0_15_i_qa_d <= twiddle_h_rsc_0_15_i_qa_d_1;
  twiddle_h_rsc_0_15_i_wea_d <= STD_LOGIC_VECTOR'( "00");
  twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( "00");

  peaseNTT_core_inst : peaseNTT_core
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_triosy_0_0_lz => xt_rsc_triosy_0_0_lz,
      xt_rsc_triosy_0_1_lz => xt_rsc_triosy_0_1_lz,
      xt_rsc_triosy_0_2_lz => xt_rsc_triosy_0_2_lz,
      xt_rsc_triosy_0_3_lz => xt_rsc_triosy_0_3_lz,
      xt_rsc_triosy_0_4_lz => xt_rsc_triosy_0_4_lz,
      xt_rsc_triosy_0_5_lz => xt_rsc_triosy_0_5_lz,
      xt_rsc_triosy_0_6_lz => xt_rsc_triosy_0_6_lz,
      xt_rsc_triosy_0_7_lz => xt_rsc_triosy_0_7_lz,
      xt_rsc_triosy_0_8_lz => xt_rsc_triosy_0_8_lz,
      xt_rsc_triosy_0_9_lz => xt_rsc_triosy_0_9_lz,
      xt_rsc_triosy_0_10_lz => xt_rsc_triosy_0_10_lz,
      xt_rsc_triosy_0_11_lz => xt_rsc_triosy_0_11_lz,
      xt_rsc_triosy_0_12_lz => xt_rsc_triosy_0_12_lz,
      xt_rsc_triosy_0_13_lz => xt_rsc_triosy_0_13_lz,
      xt_rsc_triosy_0_14_lz => xt_rsc_triosy_0_14_lz,
      xt_rsc_triosy_0_15_lz => xt_rsc_triosy_0_15_lz,
      xt_rsc_triosy_0_16_lz => xt_rsc_triosy_0_16_lz,
      xt_rsc_triosy_0_17_lz => xt_rsc_triosy_0_17_lz,
      xt_rsc_triosy_0_18_lz => xt_rsc_triosy_0_18_lz,
      xt_rsc_triosy_0_19_lz => xt_rsc_triosy_0_19_lz,
      xt_rsc_triosy_0_20_lz => xt_rsc_triosy_0_20_lz,
      xt_rsc_triosy_0_21_lz => xt_rsc_triosy_0_21_lz,
      xt_rsc_triosy_0_22_lz => xt_rsc_triosy_0_22_lz,
      xt_rsc_triosy_0_23_lz => xt_rsc_triosy_0_23_lz,
      xt_rsc_triosy_0_24_lz => xt_rsc_triosy_0_24_lz,
      xt_rsc_triosy_0_25_lz => xt_rsc_triosy_0_25_lz,
      xt_rsc_triosy_0_26_lz => xt_rsc_triosy_0_26_lz,
      xt_rsc_triosy_0_27_lz => xt_rsc_triosy_0_27_lz,
      xt_rsc_triosy_0_28_lz => xt_rsc_triosy_0_28_lz,
      xt_rsc_triosy_0_29_lz => xt_rsc_triosy_0_29_lz,
      xt_rsc_triosy_0_30_lz => xt_rsc_triosy_0_30_lz,
      xt_rsc_triosy_0_31_lz => xt_rsc_triosy_0_31_lz,
      p_rsc_dat => peaseNTT_core_inst_p_rsc_dat,
      p_rsc_triosy_lz => p_rsc_triosy_lz,
      r_rsc_triosy_lz => r_rsc_triosy_lz,
      twiddle_rsc_triosy_0_0_lz => twiddle_rsc_triosy_0_0_lz,
      twiddle_rsc_triosy_0_1_lz => twiddle_rsc_triosy_0_1_lz,
      twiddle_rsc_triosy_0_2_lz => twiddle_rsc_triosy_0_2_lz,
      twiddle_rsc_triosy_0_3_lz => twiddle_rsc_triosy_0_3_lz,
      twiddle_rsc_triosy_0_4_lz => twiddle_rsc_triosy_0_4_lz,
      twiddle_rsc_triosy_0_5_lz => twiddle_rsc_triosy_0_5_lz,
      twiddle_rsc_triosy_0_6_lz => twiddle_rsc_triosy_0_6_lz,
      twiddle_rsc_triosy_0_7_lz => twiddle_rsc_triosy_0_7_lz,
      twiddle_rsc_triosy_0_8_lz => twiddle_rsc_triosy_0_8_lz,
      twiddle_rsc_triosy_0_9_lz => twiddle_rsc_triosy_0_9_lz,
      twiddle_rsc_triosy_0_10_lz => twiddle_rsc_triosy_0_10_lz,
      twiddle_rsc_triosy_0_11_lz => twiddle_rsc_triosy_0_11_lz,
      twiddle_rsc_triosy_0_12_lz => twiddle_rsc_triosy_0_12_lz,
      twiddle_rsc_triosy_0_13_lz => twiddle_rsc_triosy_0_13_lz,
      twiddle_rsc_triosy_0_14_lz => twiddle_rsc_triosy_0_14_lz,
      twiddle_rsc_triosy_0_15_lz => twiddle_rsc_triosy_0_15_lz,
      twiddle_h_rsc_triosy_0_0_lz => twiddle_h_rsc_triosy_0_0_lz,
      twiddle_h_rsc_triosy_0_1_lz => twiddle_h_rsc_triosy_0_1_lz,
      twiddle_h_rsc_triosy_0_2_lz => twiddle_h_rsc_triosy_0_2_lz,
      twiddle_h_rsc_triosy_0_3_lz => twiddle_h_rsc_triosy_0_3_lz,
      twiddle_h_rsc_triosy_0_4_lz => twiddle_h_rsc_triosy_0_4_lz,
      twiddle_h_rsc_triosy_0_5_lz => twiddle_h_rsc_triosy_0_5_lz,
      twiddle_h_rsc_triosy_0_6_lz => twiddle_h_rsc_triosy_0_6_lz,
      twiddle_h_rsc_triosy_0_7_lz => twiddle_h_rsc_triosy_0_7_lz,
      twiddle_h_rsc_triosy_0_8_lz => twiddle_h_rsc_triosy_0_8_lz,
      twiddle_h_rsc_triosy_0_9_lz => twiddle_h_rsc_triosy_0_9_lz,
      twiddle_h_rsc_triosy_0_10_lz => twiddle_h_rsc_triosy_0_10_lz,
      twiddle_h_rsc_triosy_0_11_lz => twiddle_h_rsc_triosy_0_11_lz,
      twiddle_h_rsc_triosy_0_12_lz => twiddle_h_rsc_triosy_0_12_lz,
      twiddle_h_rsc_triosy_0_13_lz => twiddle_h_rsc_triosy_0_13_lz,
      twiddle_h_rsc_triosy_0_14_lz => twiddle_h_rsc_triosy_0_14_lz,
      twiddle_h_rsc_triosy_0_15_lz => twiddle_h_rsc_triosy_0_15_lz,
      yt_rsc_0_0_i_adra_d => peaseNTT_core_inst_yt_rsc_0_0_i_adra_d,
      yt_rsc_0_0_i_clka_en_d => yt_rsc_0_0_i_clka_en_d,
      yt_rsc_0_0_i_da_d => peaseNTT_core_inst_yt_rsc_0_0_i_da_d,
      yt_rsc_0_0_i_qa_d => peaseNTT_core_inst_yt_rsc_0_0_i_qa_d,
      yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_1_i_adra_d => peaseNTT_core_inst_yt_rsc_0_1_i_adra_d,
      yt_rsc_0_1_i_da_d => peaseNTT_core_inst_yt_rsc_0_1_i_da_d,
      yt_rsc_0_1_i_qa_d => peaseNTT_core_inst_yt_rsc_0_1_i_qa_d,
      yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_2_i_adra_d => peaseNTT_core_inst_yt_rsc_0_2_i_adra_d,
      yt_rsc_0_2_i_da_d => peaseNTT_core_inst_yt_rsc_0_2_i_da_d,
      yt_rsc_0_2_i_qa_d => peaseNTT_core_inst_yt_rsc_0_2_i_qa_d,
      yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_3_i_adra_d => peaseNTT_core_inst_yt_rsc_0_3_i_adra_d,
      yt_rsc_0_3_i_da_d => peaseNTT_core_inst_yt_rsc_0_3_i_da_d,
      yt_rsc_0_3_i_qa_d => peaseNTT_core_inst_yt_rsc_0_3_i_qa_d,
      yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_4_i_adra_d => peaseNTT_core_inst_yt_rsc_0_4_i_adra_d,
      yt_rsc_0_4_i_da_d => peaseNTT_core_inst_yt_rsc_0_4_i_da_d,
      yt_rsc_0_4_i_qa_d => peaseNTT_core_inst_yt_rsc_0_4_i_qa_d,
      yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_5_i_adra_d => peaseNTT_core_inst_yt_rsc_0_5_i_adra_d,
      yt_rsc_0_5_i_da_d => peaseNTT_core_inst_yt_rsc_0_5_i_da_d,
      yt_rsc_0_5_i_qa_d => peaseNTT_core_inst_yt_rsc_0_5_i_qa_d,
      yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_6_i_adra_d => peaseNTT_core_inst_yt_rsc_0_6_i_adra_d,
      yt_rsc_0_6_i_da_d => peaseNTT_core_inst_yt_rsc_0_6_i_da_d,
      yt_rsc_0_6_i_qa_d => peaseNTT_core_inst_yt_rsc_0_6_i_qa_d,
      yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_7_i_adra_d => peaseNTT_core_inst_yt_rsc_0_7_i_adra_d,
      yt_rsc_0_7_i_da_d => peaseNTT_core_inst_yt_rsc_0_7_i_da_d,
      yt_rsc_0_7_i_qa_d => peaseNTT_core_inst_yt_rsc_0_7_i_qa_d,
      yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_8_i_adra_d => peaseNTT_core_inst_yt_rsc_0_8_i_adra_d,
      yt_rsc_0_8_i_da_d => peaseNTT_core_inst_yt_rsc_0_8_i_da_d,
      yt_rsc_0_8_i_qa_d => peaseNTT_core_inst_yt_rsc_0_8_i_qa_d,
      yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_9_i_adra_d => peaseNTT_core_inst_yt_rsc_0_9_i_adra_d,
      yt_rsc_0_9_i_da_d => peaseNTT_core_inst_yt_rsc_0_9_i_da_d,
      yt_rsc_0_9_i_qa_d => peaseNTT_core_inst_yt_rsc_0_9_i_qa_d,
      yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_10_i_adra_d => peaseNTT_core_inst_yt_rsc_0_10_i_adra_d,
      yt_rsc_0_10_i_da_d => peaseNTT_core_inst_yt_rsc_0_10_i_da_d,
      yt_rsc_0_10_i_qa_d => peaseNTT_core_inst_yt_rsc_0_10_i_qa_d,
      yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_11_i_adra_d => peaseNTT_core_inst_yt_rsc_0_11_i_adra_d,
      yt_rsc_0_11_i_da_d => peaseNTT_core_inst_yt_rsc_0_11_i_da_d,
      yt_rsc_0_11_i_qa_d => peaseNTT_core_inst_yt_rsc_0_11_i_qa_d,
      yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_12_i_adra_d => peaseNTT_core_inst_yt_rsc_0_12_i_adra_d,
      yt_rsc_0_12_i_da_d => peaseNTT_core_inst_yt_rsc_0_12_i_da_d,
      yt_rsc_0_12_i_qa_d => peaseNTT_core_inst_yt_rsc_0_12_i_qa_d,
      yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_13_i_adra_d => peaseNTT_core_inst_yt_rsc_0_13_i_adra_d,
      yt_rsc_0_13_i_da_d => peaseNTT_core_inst_yt_rsc_0_13_i_da_d,
      yt_rsc_0_13_i_qa_d => peaseNTT_core_inst_yt_rsc_0_13_i_qa_d,
      yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_14_i_adra_d => peaseNTT_core_inst_yt_rsc_0_14_i_adra_d,
      yt_rsc_0_14_i_da_d => peaseNTT_core_inst_yt_rsc_0_14_i_da_d,
      yt_rsc_0_14_i_qa_d => peaseNTT_core_inst_yt_rsc_0_14_i_qa_d,
      yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_15_i_adra_d => peaseNTT_core_inst_yt_rsc_0_15_i_adra_d,
      yt_rsc_0_15_i_da_d => peaseNTT_core_inst_yt_rsc_0_15_i_da_d,
      yt_rsc_0_15_i_qa_d => peaseNTT_core_inst_yt_rsc_0_15_i_qa_d,
      yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_16_i_adra_d => peaseNTT_core_inst_yt_rsc_0_16_i_adra_d,
      yt_rsc_0_16_i_clka_en_d => yt_rsc_0_16_i_clka_en_d,
      yt_rsc_0_16_i_da_d => peaseNTT_core_inst_yt_rsc_0_16_i_da_d,
      yt_rsc_0_16_i_qa_d => peaseNTT_core_inst_yt_rsc_0_16_i_qa_d,
      yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_17_i_adra_d => peaseNTT_core_inst_yt_rsc_0_17_i_adra_d,
      yt_rsc_0_17_i_da_d => peaseNTT_core_inst_yt_rsc_0_17_i_da_d,
      yt_rsc_0_17_i_qa_d => peaseNTT_core_inst_yt_rsc_0_17_i_qa_d,
      yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_18_i_adra_d => peaseNTT_core_inst_yt_rsc_0_18_i_adra_d,
      yt_rsc_0_18_i_da_d => peaseNTT_core_inst_yt_rsc_0_18_i_da_d,
      yt_rsc_0_18_i_qa_d => peaseNTT_core_inst_yt_rsc_0_18_i_qa_d,
      yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_19_i_adra_d => peaseNTT_core_inst_yt_rsc_0_19_i_adra_d,
      yt_rsc_0_19_i_da_d => peaseNTT_core_inst_yt_rsc_0_19_i_da_d,
      yt_rsc_0_19_i_qa_d => peaseNTT_core_inst_yt_rsc_0_19_i_qa_d,
      yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_20_i_adra_d => peaseNTT_core_inst_yt_rsc_0_20_i_adra_d,
      yt_rsc_0_20_i_da_d => peaseNTT_core_inst_yt_rsc_0_20_i_da_d,
      yt_rsc_0_20_i_qa_d => peaseNTT_core_inst_yt_rsc_0_20_i_qa_d,
      yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_21_i_adra_d => peaseNTT_core_inst_yt_rsc_0_21_i_adra_d,
      yt_rsc_0_21_i_da_d => peaseNTT_core_inst_yt_rsc_0_21_i_da_d,
      yt_rsc_0_21_i_qa_d => peaseNTT_core_inst_yt_rsc_0_21_i_qa_d,
      yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_22_i_adra_d => peaseNTT_core_inst_yt_rsc_0_22_i_adra_d,
      yt_rsc_0_22_i_da_d => peaseNTT_core_inst_yt_rsc_0_22_i_da_d,
      yt_rsc_0_22_i_qa_d => peaseNTT_core_inst_yt_rsc_0_22_i_qa_d,
      yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_23_i_adra_d => peaseNTT_core_inst_yt_rsc_0_23_i_adra_d,
      yt_rsc_0_23_i_da_d => peaseNTT_core_inst_yt_rsc_0_23_i_da_d,
      yt_rsc_0_23_i_qa_d => peaseNTT_core_inst_yt_rsc_0_23_i_qa_d,
      yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_24_i_adra_d => peaseNTT_core_inst_yt_rsc_0_24_i_adra_d,
      yt_rsc_0_24_i_da_d => peaseNTT_core_inst_yt_rsc_0_24_i_da_d,
      yt_rsc_0_24_i_qa_d => peaseNTT_core_inst_yt_rsc_0_24_i_qa_d,
      yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_25_i_adra_d => peaseNTT_core_inst_yt_rsc_0_25_i_adra_d,
      yt_rsc_0_25_i_da_d => peaseNTT_core_inst_yt_rsc_0_25_i_da_d,
      yt_rsc_0_25_i_qa_d => peaseNTT_core_inst_yt_rsc_0_25_i_qa_d,
      yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_26_i_adra_d => peaseNTT_core_inst_yt_rsc_0_26_i_adra_d,
      yt_rsc_0_26_i_da_d => peaseNTT_core_inst_yt_rsc_0_26_i_da_d,
      yt_rsc_0_26_i_qa_d => peaseNTT_core_inst_yt_rsc_0_26_i_qa_d,
      yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_27_i_adra_d => peaseNTT_core_inst_yt_rsc_0_27_i_adra_d,
      yt_rsc_0_27_i_da_d => peaseNTT_core_inst_yt_rsc_0_27_i_da_d,
      yt_rsc_0_27_i_qa_d => peaseNTT_core_inst_yt_rsc_0_27_i_qa_d,
      yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_28_i_adra_d => peaseNTT_core_inst_yt_rsc_0_28_i_adra_d,
      yt_rsc_0_28_i_da_d => peaseNTT_core_inst_yt_rsc_0_28_i_da_d,
      yt_rsc_0_28_i_qa_d => peaseNTT_core_inst_yt_rsc_0_28_i_qa_d,
      yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_29_i_adra_d => peaseNTT_core_inst_yt_rsc_0_29_i_adra_d,
      yt_rsc_0_29_i_da_d => peaseNTT_core_inst_yt_rsc_0_29_i_da_d,
      yt_rsc_0_29_i_qa_d => peaseNTT_core_inst_yt_rsc_0_29_i_qa_d,
      yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_30_i_adra_d => peaseNTT_core_inst_yt_rsc_0_30_i_adra_d,
      yt_rsc_0_30_i_da_d => peaseNTT_core_inst_yt_rsc_0_30_i_da_d,
      yt_rsc_0_30_i_qa_d => peaseNTT_core_inst_yt_rsc_0_30_i_qa_d,
      yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_31_i_adra_d => peaseNTT_core_inst_yt_rsc_0_31_i_adra_d,
      yt_rsc_0_31_i_da_d => peaseNTT_core_inst_yt_rsc_0_31_i_da_d,
      yt_rsc_0_31_i_qa_d => peaseNTT_core_inst_yt_rsc_0_31_i_qa_d,
      yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_0_i_adra_d => peaseNTT_core_inst_xt_rsc_0_0_i_adra_d,
      xt_rsc_0_0_i_da_d => peaseNTT_core_inst_xt_rsc_0_0_i_da_d,
      xt_rsc_0_0_i_qa_d => peaseNTT_core_inst_xt_rsc_0_0_i_qa_d,
      xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_1_i_adra_d => peaseNTT_core_inst_xt_rsc_0_1_i_adra_d,
      xt_rsc_0_1_i_da_d => peaseNTT_core_inst_xt_rsc_0_1_i_da_d,
      xt_rsc_0_1_i_qa_d => peaseNTT_core_inst_xt_rsc_0_1_i_qa_d,
      xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_2_i_adra_d => peaseNTT_core_inst_xt_rsc_0_2_i_adra_d,
      xt_rsc_0_2_i_da_d => peaseNTT_core_inst_xt_rsc_0_2_i_da_d,
      xt_rsc_0_2_i_qa_d => peaseNTT_core_inst_xt_rsc_0_2_i_qa_d,
      xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_3_i_adra_d => peaseNTT_core_inst_xt_rsc_0_3_i_adra_d,
      xt_rsc_0_3_i_da_d => peaseNTT_core_inst_xt_rsc_0_3_i_da_d,
      xt_rsc_0_3_i_qa_d => peaseNTT_core_inst_xt_rsc_0_3_i_qa_d,
      xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_4_i_adra_d => peaseNTT_core_inst_xt_rsc_0_4_i_adra_d,
      xt_rsc_0_4_i_da_d => peaseNTT_core_inst_xt_rsc_0_4_i_da_d,
      xt_rsc_0_4_i_qa_d => peaseNTT_core_inst_xt_rsc_0_4_i_qa_d,
      xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_5_i_adra_d => peaseNTT_core_inst_xt_rsc_0_5_i_adra_d,
      xt_rsc_0_5_i_da_d => peaseNTT_core_inst_xt_rsc_0_5_i_da_d,
      xt_rsc_0_5_i_qa_d => peaseNTT_core_inst_xt_rsc_0_5_i_qa_d,
      xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_6_i_adra_d => peaseNTT_core_inst_xt_rsc_0_6_i_adra_d,
      xt_rsc_0_6_i_da_d => peaseNTT_core_inst_xt_rsc_0_6_i_da_d,
      xt_rsc_0_6_i_qa_d => peaseNTT_core_inst_xt_rsc_0_6_i_qa_d,
      xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_7_i_adra_d => peaseNTT_core_inst_xt_rsc_0_7_i_adra_d,
      xt_rsc_0_7_i_da_d => peaseNTT_core_inst_xt_rsc_0_7_i_da_d,
      xt_rsc_0_7_i_qa_d => peaseNTT_core_inst_xt_rsc_0_7_i_qa_d,
      xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_8_i_adra_d => peaseNTT_core_inst_xt_rsc_0_8_i_adra_d,
      xt_rsc_0_8_i_da_d => peaseNTT_core_inst_xt_rsc_0_8_i_da_d,
      xt_rsc_0_8_i_qa_d => peaseNTT_core_inst_xt_rsc_0_8_i_qa_d,
      xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_9_i_adra_d => peaseNTT_core_inst_xt_rsc_0_9_i_adra_d,
      xt_rsc_0_9_i_da_d => peaseNTT_core_inst_xt_rsc_0_9_i_da_d,
      xt_rsc_0_9_i_qa_d => peaseNTT_core_inst_xt_rsc_0_9_i_qa_d,
      xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_10_i_adra_d => peaseNTT_core_inst_xt_rsc_0_10_i_adra_d,
      xt_rsc_0_10_i_da_d => peaseNTT_core_inst_xt_rsc_0_10_i_da_d,
      xt_rsc_0_10_i_qa_d => peaseNTT_core_inst_xt_rsc_0_10_i_qa_d,
      xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_11_i_adra_d => peaseNTT_core_inst_xt_rsc_0_11_i_adra_d,
      xt_rsc_0_11_i_da_d => peaseNTT_core_inst_xt_rsc_0_11_i_da_d,
      xt_rsc_0_11_i_qa_d => peaseNTT_core_inst_xt_rsc_0_11_i_qa_d,
      xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_12_i_adra_d => peaseNTT_core_inst_xt_rsc_0_12_i_adra_d,
      xt_rsc_0_12_i_da_d => peaseNTT_core_inst_xt_rsc_0_12_i_da_d,
      xt_rsc_0_12_i_qa_d => peaseNTT_core_inst_xt_rsc_0_12_i_qa_d,
      xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_13_i_adra_d => peaseNTT_core_inst_xt_rsc_0_13_i_adra_d,
      xt_rsc_0_13_i_da_d => peaseNTT_core_inst_xt_rsc_0_13_i_da_d,
      xt_rsc_0_13_i_qa_d => peaseNTT_core_inst_xt_rsc_0_13_i_qa_d,
      xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_14_i_adra_d => peaseNTT_core_inst_xt_rsc_0_14_i_adra_d,
      xt_rsc_0_14_i_da_d => peaseNTT_core_inst_xt_rsc_0_14_i_da_d,
      xt_rsc_0_14_i_qa_d => peaseNTT_core_inst_xt_rsc_0_14_i_qa_d,
      xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_15_i_adra_d => peaseNTT_core_inst_xt_rsc_0_15_i_adra_d,
      xt_rsc_0_15_i_da_d => peaseNTT_core_inst_xt_rsc_0_15_i_da_d,
      xt_rsc_0_15_i_qa_d => peaseNTT_core_inst_xt_rsc_0_15_i_qa_d,
      xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_16_i_adra_d => peaseNTT_core_inst_xt_rsc_0_16_i_adra_d,
      xt_rsc_0_16_i_da_d => peaseNTT_core_inst_xt_rsc_0_16_i_da_d,
      xt_rsc_0_16_i_qa_d => peaseNTT_core_inst_xt_rsc_0_16_i_qa_d,
      xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_17_i_adra_d => peaseNTT_core_inst_xt_rsc_0_17_i_adra_d,
      xt_rsc_0_17_i_da_d => peaseNTT_core_inst_xt_rsc_0_17_i_da_d,
      xt_rsc_0_17_i_qa_d => peaseNTT_core_inst_xt_rsc_0_17_i_qa_d,
      xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_18_i_adra_d => peaseNTT_core_inst_xt_rsc_0_18_i_adra_d,
      xt_rsc_0_18_i_da_d => peaseNTT_core_inst_xt_rsc_0_18_i_da_d,
      xt_rsc_0_18_i_qa_d => peaseNTT_core_inst_xt_rsc_0_18_i_qa_d,
      xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_19_i_adra_d => peaseNTT_core_inst_xt_rsc_0_19_i_adra_d,
      xt_rsc_0_19_i_da_d => peaseNTT_core_inst_xt_rsc_0_19_i_da_d,
      xt_rsc_0_19_i_qa_d => peaseNTT_core_inst_xt_rsc_0_19_i_qa_d,
      xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_20_i_adra_d => peaseNTT_core_inst_xt_rsc_0_20_i_adra_d,
      xt_rsc_0_20_i_da_d => peaseNTT_core_inst_xt_rsc_0_20_i_da_d,
      xt_rsc_0_20_i_qa_d => peaseNTT_core_inst_xt_rsc_0_20_i_qa_d,
      xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_21_i_adra_d => peaseNTT_core_inst_xt_rsc_0_21_i_adra_d,
      xt_rsc_0_21_i_da_d => peaseNTT_core_inst_xt_rsc_0_21_i_da_d,
      xt_rsc_0_21_i_qa_d => peaseNTT_core_inst_xt_rsc_0_21_i_qa_d,
      xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_22_i_adra_d => peaseNTT_core_inst_xt_rsc_0_22_i_adra_d,
      xt_rsc_0_22_i_da_d => peaseNTT_core_inst_xt_rsc_0_22_i_da_d,
      xt_rsc_0_22_i_qa_d => peaseNTT_core_inst_xt_rsc_0_22_i_qa_d,
      xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_23_i_adra_d => peaseNTT_core_inst_xt_rsc_0_23_i_adra_d,
      xt_rsc_0_23_i_da_d => peaseNTT_core_inst_xt_rsc_0_23_i_da_d,
      xt_rsc_0_23_i_qa_d => peaseNTT_core_inst_xt_rsc_0_23_i_qa_d,
      xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_24_i_adra_d => peaseNTT_core_inst_xt_rsc_0_24_i_adra_d,
      xt_rsc_0_24_i_da_d => peaseNTT_core_inst_xt_rsc_0_24_i_da_d,
      xt_rsc_0_24_i_qa_d => peaseNTT_core_inst_xt_rsc_0_24_i_qa_d,
      xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_25_i_adra_d => peaseNTT_core_inst_xt_rsc_0_25_i_adra_d,
      xt_rsc_0_25_i_da_d => peaseNTT_core_inst_xt_rsc_0_25_i_da_d,
      xt_rsc_0_25_i_qa_d => peaseNTT_core_inst_xt_rsc_0_25_i_qa_d,
      xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_26_i_adra_d => peaseNTT_core_inst_xt_rsc_0_26_i_adra_d,
      xt_rsc_0_26_i_da_d => peaseNTT_core_inst_xt_rsc_0_26_i_da_d,
      xt_rsc_0_26_i_qa_d => peaseNTT_core_inst_xt_rsc_0_26_i_qa_d,
      xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_27_i_adra_d => peaseNTT_core_inst_xt_rsc_0_27_i_adra_d,
      xt_rsc_0_27_i_da_d => peaseNTT_core_inst_xt_rsc_0_27_i_da_d,
      xt_rsc_0_27_i_qa_d => peaseNTT_core_inst_xt_rsc_0_27_i_qa_d,
      xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_28_i_adra_d => peaseNTT_core_inst_xt_rsc_0_28_i_adra_d,
      xt_rsc_0_28_i_da_d => peaseNTT_core_inst_xt_rsc_0_28_i_da_d,
      xt_rsc_0_28_i_qa_d => peaseNTT_core_inst_xt_rsc_0_28_i_qa_d,
      xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_29_i_adra_d => peaseNTT_core_inst_xt_rsc_0_29_i_adra_d,
      xt_rsc_0_29_i_da_d => peaseNTT_core_inst_xt_rsc_0_29_i_da_d,
      xt_rsc_0_29_i_qa_d => peaseNTT_core_inst_xt_rsc_0_29_i_qa_d,
      xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_30_i_adra_d => peaseNTT_core_inst_xt_rsc_0_30_i_adra_d,
      xt_rsc_0_30_i_da_d => peaseNTT_core_inst_xt_rsc_0_30_i_da_d,
      xt_rsc_0_30_i_qa_d => peaseNTT_core_inst_xt_rsc_0_30_i_qa_d,
      xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_31_i_adra_d => peaseNTT_core_inst_xt_rsc_0_31_i_adra_d,
      xt_rsc_0_31_i_da_d => peaseNTT_core_inst_xt_rsc_0_31_i_da_d,
      xt_rsc_0_31_i_qa_d => peaseNTT_core_inst_xt_rsc_0_31_i_qa_d,
      xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_0_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_0_i_adra_d,
      twiddle_rsc_0_0_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_0_i_qa_d,
      twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_1_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_1_i_adra_d,
      twiddle_rsc_0_1_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_1_i_qa_d,
      twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_2_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_2_i_adra_d,
      twiddle_rsc_0_2_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_2_i_qa_d,
      twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_3_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_3_i_adra_d,
      twiddle_rsc_0_3_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_3_i_qa_d,
      twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_4_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_4_i_adra_d,
      twiddle_rsc_0_4_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_4_i_qa_d,
      twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_5_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_5_i_adra_d,
      twiddle_rsc_0_5_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_5_i_qa_d,
      twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_6_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_6_i_adra_d,
      twiddle_rsc_0_6_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_6_i_qa_d,
      twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_7_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_7_i_adra_d,
      twiddle_rsc_0_7_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_7_i_qa_d,
      twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_8_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_8_i_adra_d,
      twiddle_rsc_0_8_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_8_i_qa_d,
      twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_9_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_9_i_adra_d,
      twiddle_rsc_0_9_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_9_i_qa_d,
      twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_10_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_10_i_adra_d,
      twiddle_rsc_0_10_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_10_i_qa_d,
      twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_11_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_11_i_adra_d,
      twiddle_rsc_0_11_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_11_i_qa_d,
      twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_12_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_12_i_adra_d,
      twiddle_rsc_0_12_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_12_i_qa_d,
      twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_13_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_13_i_adra_d,
      twiddle_rsc_0_13_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_13_i_qa_d,
      twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_14_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_14_i_adra_d,
      twiddle_rsc_0_14_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_14_i_qa_d,
      twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_15_i_adra_d => peaseNTT_core_inst_twiddle_rsc_0_15_i_adra_d,
      twiddle_rsc_0_15_i_qa_d => peaseNTT_core_inst_twiddle_rsc_0_15_i_qa_d,
      twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_0_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_0_i_adra_d,
      twiddle_h_rsc_0_0_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_0_i_qa_d,
      twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_1_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_1_i_adra_d,
      twiddle_h_rsc_0_1_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_1_i_qa_d,
      twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_2_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_2_i_adra_d,
      twiddle_h_rsc_0_2_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_2_i_qa_d,
      twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_3_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_3_i_adra_d,
      twiddle_h_rsc_0_3_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_3_i_qa_d,
      twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_4_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_4_i_adra_d,
      twiddle_h_rsc_0_4_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_4_i_qa_d,
      twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_5_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_5_i_adra_d,
      twiddle_h_rsc_0_5_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_5_i_qa_d,
      twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_6_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_6_i_adra_d,
      twiddle_h_rsc_0_6_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_6_i_qa_d,
      twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_7_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_7_i_adra_d,
      twiddle_h_rsc_0_7_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_7_i_qa_d,
      twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_8_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_8_i_adra_d,
      twiddle_h_rsc_0_8_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_8_i_qa_d,
      twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_9_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_9_i_adra_d,
      twiddle_h_rsc_0_9_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_9_i_qa_d,
      twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_10_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_10_i_adra_d,
      twiddle_h_rsc_0_10_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_10_i_qa_d,
      twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_11_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_11_i_adra_d,
      twiddle_h_rsc_0_11_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_11_i_qa_d,
      twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_12_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_12_i_adra_d,
      twiddle_h_rsc_0_12_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_12_i_qa_d,
      twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_13_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_13_i_adra_d,
      twiddle_h_rsc_0_13_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_13_i_qa_d,
      twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_14_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_14_i_adra_d,
      twiddle_h_rsc_0_14_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_14_i_qa_d,
      twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_15_i_adra_d => peaseNTT_core_inst_twiddle_h_rsc_0_15_i_adra_d,
      twiddle_h_rsc_0_15_i_qa_d => peaseNTT_core_inst_twiddle_h_rsc_0_15_i_qa_d,
      twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d => peaseNTT_core_inst_twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_0_i_wea_d_pff => peaseNTT_core_inst_yt_rsc_0_0_i_wea_d_pff,
      yt_rsc_0_16_i_wea_d_pff => peaseNTT_core_inst_yt_rsc_0_16_i_wea_d_pff,
      xt_rsc_0_0_i_wea_d_pff => peaseNTT_core_inst_xt_rsc_0_0_i_wea_d_pff,
      xt_rsc_0_16_i_wea_d_pff => peaseNTT_core_inst_xt_rsc_0_16_i_wea_d_pff
    );
  peaseNTT_core_inst_p_rsc_dat <= p_rsc_dat;
  yt_rsc_0_0_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_0_i_adra_d;
  yt_rsc_0_0_i_da_d <= peaseNTT_core_inst_yt_rsc_0_0_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_0_i_qa_d <= yt_rsc_0_0_i_qa_d;
  yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_1_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_1_i_adra_d;
  yt_rsc_0_1_i_da_d <= peaseNTT_core_inst_yt_rsc_0_1_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_1_i_qa_d <= yt_rsc_0_1_i_qa_d;
  yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_2_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_2_i_adra_d;
  yt_rsc_0_2_i_da_d <= peaseNTT_core_inst_yt_rsc_0_2_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_2_i_qa_d <= yt_rsc_0_2_i_qa_d;
  yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_3_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_3_i_adra_d;
  yt_rsc_0_3_i_da_d <= peaseNTT_core_inst_yt_rsc_0_3_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_3_i_qa_d <= yt_rsc_0_3_i_qa_d;
  yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_4_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_4_i_adra_d;
  yt_rsc_0_4_i_da_d <= peaseNTT_core_inst_yt_rsc_0_4_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_4_i_qa_d <= yt_rsc_0_4_i_qa_d;
  yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_5_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_5_i_adra_d;
  yt_rsc_0_5_i_da_d <= peaseNTT_core_inst_yt_rsc_0_5_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_5_i_qa_d <= yt_rsc_0_5_i_qa_d;
  yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_6_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_6_i_adra_d;
  yt_rsc_0_6_i_da_d <= peaseNTT_core_inst_yt_rsc_0_6_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_6_i_qa_d <= yt_rsc_0_6_i_qa_d;
  yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_7_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_7_i_adra_d;
  yt_rsc_0_7_i_da_d <= peaseNTT_core_inst_yt_rsc_0_7_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_7_i_qa_d <= yt_rsc_0_7_i_qa_d;
  yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_8_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_8_i_adra_d;
  yt_rsc_0_8_i_da_d <= peaseNTT_core_inst_yt_rsc_0_8_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_8_i_qa_d <= yt_rsc_0_8_i_qa_d;
  yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_9_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_9_i_adra_d;
  yt_rsc_0_9_i_da_d <= peaseNTT_core_inst_yt_rsc_0_9_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_9_i_qa_d <= yt_rsc_0_9_i_qa_d;
  yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_10_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_10_i_adra_d;
  yt_rsc_0_10_i_da_d <= peaseNTT_core_inst_yt_rsc_0_10_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_10_i_qa_d <= yt_rsc_0_10_i_qa_d;
  yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_11_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_11_i_adra_d;
  yt_rsc_0_11_i_da_d <= peaseNTT_core_inst_yt_rsc_0_11_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_11_i_qa_d <= yt_rsc_0_11_i_qa_d;
  yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_12_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_12_i_adra_d;
  yt_rsc_0_12_i_da_d <= peaseNTT_core_inst_yt_rsc_0_12_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_12_i_qa_d <= yt_rsc_0_12_i_qa_d;
  yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_13_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_13_i_adra_d;
  yt_rsc_0_13_i_da_d <= peaseNTT_core_inst_yt_rsc_0_13_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_13_i_qa_d <= yt_rsc_0_13_i_qa_d;
  yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_14_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_14_i_adra_d;
  yt_rsc_0_14_i_da_d <= peaseNTT_core_inst_yt_rsc_0_14_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_14_i_qa_d <= yt_rsc_0_14_i_qa_d;
  yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_15_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_15_i_adra_d;
  yt_rsc_0_15_i_da_d <= peaseNTT_core_inst_yt_rsc_0_15_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_15_i_qa_d <= yt_rsc_0_15_i_qa_d;
  yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_16_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_16_i_adra_d;
  yt_rsc_0_16_i_da_d <= peaseNTT_core_inst_yt_rsc_0_16_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_16_i_qa_d <= yt_rsc_0_16_i_qa_d;
  yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_17_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_17_i_adra_d;
  yt_rsc_0_17_i_da_d <= peaseNTT_core_inst_yt_rsc_0_17_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_17_i_qa_d <= yt_rsc_0_17_i_qa_d;
  yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_18_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_18_i_adra_d;
  yt_rsc_0_18_i_da_d <= peaseNTT_core_inst_yt_rsc_0_18_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_18_i_qa_d <= yt_rsc_0_18_i_qa_d;
  yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_19_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_19_i_adra_d;
  yt_rsc_0_19_i_da_d <= peaseNTT_core_inst_yt_rsc_0_19_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_19_i_qa_d <= yt_rsc_0_19_i_qa_d;
  yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_20_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_20_i_adra_d;
  yt_rsc_0_20_i_da_d <= peaseNTT_core_inst_yt_rsc_0_20_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_20_i_qa_d <= yt_rsc_0_20_i_qa_d;
  yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_21_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_21_i_adra_d;
  yt_rsc_0_21_i_da_d <= peaseNTT_core_inst_yt_rsc_0_21_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_21_i_qa_d <= yt_rsc_0_21_i_qa_d;
  yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_22_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_22_i_adra_d;
  yt_rsc_0_22_i_da_d <= peaseNTT_core_inst_yt_rsc_0_22_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_22_i_qa_d <= yt_rsc_0_22_i_qa_d;
  yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_23_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_23_i_adra_d;
  yt_rsc_0_23_i_da_d <= peaseNTT_core_inst_yt_rsc_0_23_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_23_i_qa_d <= yt_rsc_0_23_i_qa_d;
  yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_24_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_24_i_adra_d;
  yt_rsc_0_24_i_da_d <= peaseNTT_core_inst_yt_rsc_0_24_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_24_i_qa_d <= yt_rsc_0_24_i_qa_d;
  yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_25_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_25_i_adra_d;
  yt_rsc_0_25_i_da_d <= peaseNTT_core_inst_yt_rsc_0_25_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_25_i_qa_d <= yt_rsc_0_25_i_qa_d;
  yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_26_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_26_i_adra_d;
  yt_rsc_0_26_i_da_d <= peaseNTT_core_inst_yt_rsc_0_26_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_26_i_qa_d <= yt_rsc_0_26_i_qa_d;
  yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_27_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_27_i_adra_d;
  yt_rsc_0_27_i_da_d <= peaseNTT_core_inst_yt_rsc_0_27_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_27_i_qa_d <= yt_rsc_0_27_i_qa_d;
  yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_28_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_28_i_adra_d;
  yt_rsc_0_28_i_da_d <= peaseNTT_core_inst_yt_rsc_0_28_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_28_i_qa_d <= yt_rsc_0_28_i_qa_d;
  yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_29_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_29_i_adra_d;
  yt_rsc_0_29_i_da_d <= peaseNTT_core_inst_yt_rsc_0_29_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_29_i_qa_d <= yt_rsc_0_29_i_qa_d;
  yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_30_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_30_i_adra_d;
  yt_rsc_0_30_i_da_d <= peaseNTT_core_inst_yt_rsc_0_30_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_30_i_qa_d <= yt_rsc_0_30_i_qa_d;
  yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_31_i_adra_d <= peaseNTT_core_inst_yt_rsc_0_31_i_adra_d;
  yt_rsc_0_31_i_da_d <= peaseNTT_core_inst_yt_rsc_0_31_i_da_d;
  peaseNTT_core_inst_yt_rsc_0_31_i_qa_d <= yt_rsc_0_31_i_qa_d;
  yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_0_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_0_i_adra_d;
  xt_rsc_0_0_i_da_d <= peaseNTT_core_inst_xt_rsc_0_0_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_0_i_qa_d <= xt_rsc_0_0_i_qa_d;
  xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_1_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_1_i_adra_d;
  xt_rsc_0_1_i_da_d <= peaseNTT_core_inst_xt_rsc_0_1_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_1_i_qa_d <= xt_rsc_0_1_i_qa_d;
  xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_2_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_2_i_adra_d;
  xt_rsc_0_2_i_da_d <= peaseNTT_core_inst_xt_rsc_0_2_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_2_i_qa_d <= xt_rsc_0_2_i_qa_d;
  xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_3_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_3_i_adra_d;
  xt_rsc_0_3_i_da_d <= peaseNTT_core_inst_xt_rsc_0_3_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_3_i_qa_d <= xt_rsc_0_3_i_qa_d;
  xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_4_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_4_i_adra_d;
  xt_rsc_0_4_i_da_d <= peaseNTT_core_inst_xt_rsc_0_4_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_4_i_qa_d <= xt_rsc_0_4_i_qa_d;
  xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_5_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_5_i_adra_d;
  xt_rsc_0_5_i_da_d <= peaseNTT_core_inst_xt_rsc_0_5_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_5_i_qa_d <= xt_rsc_0_5_i_qa_d;
  xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_6_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_6_i_adra_d;
  xt_rsc_0_6_i_da_d <= peaseNTT_core_inst_xt_rsc_0_6_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_6_i_qa_d <= xt_rsc_0_6_i_qa_d;
  xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_7_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_7_i_adra_d;
  xt_rsc_0_7_i_da_d <= peaseNTT_core_inst_xt_rsc_0_7_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_7_i_qa_d <= xt_rsc_0_7_i_qa_d;
  xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_8_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_8_i_adra_d;
  xt_rsc_0_8_i_da_d <= peaseNTT_core_inst_xt_rsc_0_8_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_8_i_qa_d <= xt_rsc_0_8_i_qa_d;
  xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_9_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_9_i_adra_d;
  xt_rsc_0_9_i_da_d <= peaseNTT_core_inst_xt_rsc_0_9_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_9_i_qa_d <= xt_rsc_0_9_i_qa_d;
  xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_10_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_10_i_adra_d;
  xt_rsc_0_10_i_da_d <= peaseNTT_core_inst_xt_rsc_0_10_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_10_i_qa_d <= xt_rsc_0_10_i_qa_d;
  xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_11_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_11_i_adra_d;
  xt_rsc_0_11_i_da_d <= peaseNTT_core_inst_xt_rsc_0_11_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_11_i_qa_d <= xt_rsc_0_11_i_qa_d;
  xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_12_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_12_i_adra_d;
  xt_rsc_0_12_i_da_d <= peaseNTT_core_inst_xt_rsc_0_12_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_12_i_qa_d <= xt_rsc_0_12_i_qa_d;
  xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_13_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_13_i_adra_d;
  xt_rsc_0_13_i_da_d <= peaseNTT_core_inst_xt_rsc_0_13_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_13_i_qa_d <= xt_rsc_0_13_i_qa_d;
  xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_14_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_14_i_adra_d;
  xt_rsc_0_14_i_da_d <= peaseNTT_core_inst_xt_rsc_0_14_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_14_i_qa_d <= xt_rsc_0_14_i_qa_d;
  xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_15_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_15_i_adra_d;
  xt_rsc_0_15_i_da_d <= peaseNTT_core_inst_xt_rsc_0_15_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_15_i_qa_d <= xt_rsc_0_15_i_qa_d;
  xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_16_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_16_i_adra_d;
  xt_rsc_0_16_i_da_d <= peaseNTT_core_inst_xt_rsc_0_16_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_16_i_qa_d <= xt_rsc_0_16_i_qa_d;
  xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_17_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_17_i_adra_d;
  xt_rsc_0_17_i_da_d <= peaseNTT_core_inst_xt_rsc_0_17_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_17_i_qa_d <= xt_rsc_0_17_i_qa_d;
  xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_18_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_18_i_adra_d;
  xt_rsc_0_18_i_da_d <= peaseNTT_core_inst_xt_rsc_0_18_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_18_i_qa_d <= xt_rsc_0_18_i_qa_d;
  xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_19_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_19_i_adra_d;
  xt_rsc_0_19_i_da_d <= peaseNTT_core_inst_xt_rsc_0_19_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_19_i_qa_d <= xt_rsc_0_19_i_qa_d;
  xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_20_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_20_i_adra_d;
  xt_rsc_0_20_i_da_d <= peaseNTT_core_inst_xt_rsc_0_20_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_20_i_qa_d <= xt_rsc_0_20_i_qa_d;
  xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_21_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_21_i_adra_d;
  xt_rsc_0_21_i_da_d <= peaseNTT_core_inst_xt_rsc_0_21_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_21_i_qa_d <= xt_rsc_0_21_i_qa_d;
  xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_22_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_22_i_adra_d;
  xt_rsc_0_22_i_da_d <= peaseNTT_core_inst_xt_rsc_0_22_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_22_i_qa_d <= xt_rsc_0_22_i_qa_d;
  xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_23_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_23_i_adra_d;
  xt_rsc_0_23_i_da_d <= peaseNTT_core_inst_xt_rsc_0_23_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_23_i_qa_d <= xt_rsc_0_23_i_qa_d;
  xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_24_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_24_i_adra_d;
  xt_rsc_0_24_i_da_d <= peaseNTT_core_inst_xt_rsc_0_24_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_24_i_qa_d <= xt_rsc_0_24_i_qa_d;
  xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_25_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_25_i_adra_d;
  xt_rsc_0_25_i_da_d <= peaseNTT_core_inst_xt_rsc_0_25_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_25_i_qa_d <= xt_rsc_0_25_i_qa_d;
  xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_26_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_26_i_adra_d;
  xt_rsc_0_26_i_da_d <= peaseNTT_core_inst_xt_rsc_0_26_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_26_i_qa_d <= xt_rsc_0_26_i_qa_d;
  xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_27_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_27_i_adra_d;
  xt_rsc_0_27_i_da_d <= peaseNTT_core_inst_xt_rsc_0_27_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_27_i_qa_d <= xt_rsc_0_27_i_qa_d;
  xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_28_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_28_i_adra_d;
  xt_rsc_0_28_i_da_d <= peaseNTT_core_inst_xt_rsc_0_28_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_28_i_qa_d <= xt_rsc_0_28_i_qa_d;
  xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_29_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_29_i_adra_d;
  xt_rsc_0_29_i_da_d <= peaseNTT_core_inst_xt_rsc_0_29_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_29_i_qa_d <= xt_rsc_0_29_i_qa_d;
  xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_30_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_30_i_adra_d;
  xt_rsc_0_30_i_da_d <= peaseNTT_core_inst_xt_rsc_0_30_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_30_i_qa_d <= xt_rsc_0_30_i_qa_d;
  xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xt_rsc_0_31_i_adra_d <= peaseNTT_core_inst_xt_rsc_0_31_i_adra_d;
  xt_rsc_0_31_i_da_d <= peaseNTT_core_inst_xt_rsc_0_31_i_da_d;
  peaseNTT_core_inst_xt_rsc_0_31_i_qa_d <= xt_rsc_0_31_i_qa_d;
  xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_0_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_0_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_0_i_qa_d <= twiddle_rsc_0_0_i_qa_d;
  twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_1_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_1_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_1_i_qa_d <= twiddle_rsc_0_1_i_qa_d;
  twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_2_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_2_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_2_i_qa_d <= twiddle_rsc_0_2_i_qa_d;
  twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_3_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_3_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_3_i_qa_d <= twiddle_rsc_0_3_i_qa_d;
  twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_4_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_4_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_4_i_qa_d <= twiddle_rsc_0_4_i_qa_d;
  twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_5_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_5_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_5_i_qa_d <= twiddle_rsc_0_5_i_qa_d;
  twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_6_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_6_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_6_i_qa_d <= twiddle_rsc_0_6_i_qa_d;
  twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_7_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_7_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_7_i_qa_d <= twiddle_rsc_0_7_i_qa_d;
  twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_8_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_8_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_8_i_qa_d <= twiddle_rsc_0_8_i_qa_d;
  twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_9_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_9_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_9_i_qa_d <= twiddle_rsc_0_9_i_qa_d;
  twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_10_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_10_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_10_i_qa_d <= twiddle_rsc_0_10_i_qa_d;
  twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_11_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_11_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_11_i_qa_d <= twiddle_rsc_0_11_i_qa_d;
  twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_12_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_12_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_12_i_qa_d <= twiddle_rsc_0_12_i_qa_d;
  twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_13_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_13_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_13_i_qa_d <= twiddle_rsc_0_13_i_qa_d;
  twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_14_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_14_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_14_i_qa_d <= twiddle_rsc_0_14_i_qa_d;
  twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_rsc_0_15_i_adra_d <= peaseNTT_core_inst_twiddle_rsc_0_15_i_adra_d;
  peaseNTT_core_inst_twiddle_rsc_0_15_i_qa_d <= twiddle_rsc_0_15_i_qa_d;
  twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_0_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_0_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_i_qa_d <= twiddle_h_rsc_0_0_i_qa_d;
  twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_1_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_1_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_i_qa_d <= twiddle_h_rsc_0_1_i_qa_d;
  twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_2_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_2_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_i_qa_d <= twiddle_h_rsc_0_2_i_qa_d;
  twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_3_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_3_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_i_qa_d <= twiddle_h_rsc_0_3_i_qa_d;
  twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_4_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_4_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_i_qa_d <= twiddle_h_rsc_0_4_i_qa_d;
  twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_5_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_5_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_i_qa_d <= twiddle_h_rsc_0_5_i_qa_d;
  twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_6_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_6_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_i_qa_d <= twiddle_h_rsc_0_6_i_qa_d;
  twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_7_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_7_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_i_qa_d <= twiddle_h_rsc_0_7_i_qa_d;
  twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_8_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_8_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_i_qa_d <= twiddle_h_rsc_0_8_i_qa_d;
  twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_9_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_9_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_i_qa_d <= twiddle_h_rsc_0_9_i_qa_d;
  twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_10_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_10_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_i_qa_d <= twiddle_h_rsc_0_10_i_qa_d;
  twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_11_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_11_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_i_qa_d <= twiddle_h_rsc_0_11_i_qa_d;
  twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_12_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_12_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_i_qa_d <= twiddle_h_rsc_0_12_i_qa_d;
  twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_13_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_13_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_i_qa_d <= twiddle_h_rsc_0_13_i_qa_d;
  twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_14_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_14_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_i_qa_d <= twiddle_h_rsc_0_14_i_qa_d;
  twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  twiddle_h_rsc_0_15_i_adra_d <= peaseNTT_core_inst_twiddle_h_rsc_0_15_i_adra_d;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_i_qa_d <= twiddle_h_rsc_0_15_i_qa_d;
  twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= peaseNTT_core_inst_twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yt_rsc_0_0_i_wea_d_iff <= peaseNTT_core_inst_yt_rsc_0_0_i_wea_d_pff;
  yt_rsc_0_16_i_wea_d_iff <= peaseNTT_core_inst_yt_rsc_0_16_i_wea_d_pff;
  xt_rsc_0_0_i_wea_d_iff <= peaseNTT_core_inst_xt_rsc_0_0_i_wea_d_pff;
  xt_rsc_0_16_i_wea_d_iff <= peaseNTT_core_inst_xt_rsc_0_16_i_wea_d_pff;

END v11;



