
--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_sync_in_wait_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_sync_in_wait_pkg_v1 IS

COMPONENT ccs_sync_in_wait_v1 
  GENERIC (
    rscid    : INTEGER
  );
  PORT (
    rdy : OUT   std_logic;
    vld : IN    std_logic;
    irdy : IN    std_logic;
    ivld : OUT   std_logic
  );
END COMPONENT;

END ccs_sync_in_wait_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_sync_in_wait_v1 IS
  GENERIC (
    rscid    : INTEGER
  );
  PORT (
    rdy : OUT   std_logic;
    vld : IN    std_logic;
    irdy : IN    std_logic;
    ivld : OUT   std_logic
  );
END ccs_sync_in_wait_v1;

ARCHITECTURE beh OF ccs_sync_in_wait_v1 IS
BEGIN
   rdy <= irdy;
   ivld <= vld;
END beh; 

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_sync_out_wait_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_sync_out_wait_pkg_v1 IS

COMPONENT ccs_sync_out_wait_v1
  GENERIC (
    rscid    : INTEGER
  );
  PORT (
    ivld : IN    std_logic;
    irdy : OUT   std_logic;
    vld : OUT   std_logic;
    rdy : IN    std_logic
  );
END COMPONENT;

END ccs_sync_out_wait_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_sync_out_wait_v1 IS
  GENERIC (
    rscid    : INTEGER
  );
  PORT (
    ivld : IN    std_logic;
    irdy : OUT   std_logic;
    vld : OUT   std_logic;
    rdy : IN    std_logic
  );
END ccs_sync_out_wait_v1;

ARCHITECTURE beh OF ccs_sync_out_wait_v1 IS
BEGIN
   irdy <= rdy;
   vld <= ivld;
END beh; 

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_pkg_v1 IS

COMPONENT ccs_in_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    dat    : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_in_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    dat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_in_v1;

ARCHITECTURE beh OF ccs_in_v1 IS
BEGIN

  idat <= dat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_out_dreg_pkg_v2 IS

COMPONENT mgc_out_dreg_v2
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    d        : IN  std_logic_vector(width-1 DOWNTO 0);
    z        : OUT std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_out_dreg_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_out_dreg_v2 IS
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    d        : IN  std_logic_vector(width-1 DOWNTO 0);
    z        : OUT std_logic_vector(width-1 DOWNTO 0)
  );
END mgc_out_dreg_v2;

ARCHITECTURE beh OF mgc_out_dreg_v2 IS
BEGIN

  z <= d;

END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/src/funcs.vhd 

-- a package of attributes that give verification tools a hint about
-- the function being implemented
PACKAGE attributes IS
  ATTRIBUTE CALYPTO_FUNC : string;
  ATTRIBUTE CALYPTO_DATA_ORDER : string;
end attributes;

-----------------------------------------------------------------------
-- Package that declares synthesizable functions needed for RTL output
-----------------------------------------------------------------------

LIBRARY ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

PACKAGE funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

   FUNCTION maximum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION minimum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2 : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;
   
-----------------------------------------------------------------
-- logic functions
-----------------------------------------------------------------

   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION or_v (inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- mux functions
-----------------------------------------------------------------

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC_VECTOR;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- latch functions
-----------------------------------------------------------------
   FUNCTION lat_s(dinput: STD_LOGIC       ; clk: STD_LOGIC; doutput: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- tristate functions
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC       ; control: STD_LOGIC) RETURN STD_LOGIC;
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: SIGNED  ) RETURN STD_LOGIC;

   -- RETURN 2 bits (left => lt, right => eq)
   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED;
 
   FUNCTION fabs(arg1: SIGNED  ) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "**" (l, r: UNSIGNED) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "**" (l, r: SIGNED  ) RETURN SIGNED  ;

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-- *_stdar functions use shift functions from std_logic_arith
-----------------------------------------------------------------

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;

   -----------------------------------------------------------------
   -- *_stdar functions use shift functions from std_logic_arith
   -----------------------------------------------------------------
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC;
   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE;
   --FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR ;

   FUNCTION ceil_log2(size : NATURAL) return NATURAL;
   FUNCTION bits(size : NATURAL) return NATURAL;    

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   
END funcs;


--------------------------- B O D Y ----------------------------


PACKAGE BODY funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC IS
     BEGIN IF arg1 THEN RETURN '1'; ELSE RETURN '0'; END IF; END;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
--     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;

   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
     VARIABLE result: STD_LOGIC_VECTOR(0 DOWNTO 0);
   BEGIN
     result := (0 => arg1);
     RETURN result;
   END;

   FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 > arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION minimum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 < arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;

   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := input1'LENGTH;
     ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
     ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     --synopsys translate_off
     FOR i IN len-1 DOWNTO 0 LOOP
       result(i) := resolved(input1a(i) & input2a(i));
     END LOOP;
     --synopsys translate_on
     RETURN result;
   END;

   FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED) RETURN UNSIGNED IS
   BEGIN RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

   FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED) RETURN SIGNED IS
   BEGIN RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

-----------------------------------------------------------------
-- Logic Functions
-----------------------------------------------------------------

   FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;
   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(and_v(inputs, 1)); END;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(or_v(inputs, 1)); END;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(xor_v(inputs, 1)); END;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result AND inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

   FUNCTION or_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     -- this if is added as a quick fix for a bug in catapult evaluating the loop even if inputs'LENGTH==1
     -- see dts0100971279
     IF icnt2 > 1 THEN
       FOR i IN icnt2-1 DOWNTO 1 LOOP
         inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
         result := result OR inputsx(olenM1 DOWNTO 0);
       END LOOP;
     END IF;
     RETURN result;
   END;

   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result XOR inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

-----------------------------------------------------------------
-- Muxes
-----------------------------------------------------------------
   
   FUNCTION mux_sel2_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(1 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 4;
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector( size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "01" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "10" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "11" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel3_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(2 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 8;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "001" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "010" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "011" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN "100" =>
       result := inputs0(5*size-1 DOWNTO 4*size);
     WHEN "101" =>
       result := inputs0(6*size-1 DOWNTO 5*size);
     WHEN "110" =>
       result := inputs0(7*size-1 DOWNTO 6*size);
     WHEN "111" =>
       result := inputs0(8*size-1 DOWNTO 7*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel4_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(3 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 16;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "0000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "0001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "0010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "0011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "0100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "0101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "0110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "0111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "1000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "1001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "1010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "1011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "1100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "1101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "1110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "1111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel5_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(4 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 32;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0 );
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "00001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "00010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "00011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "00100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "00101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "00110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "00111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "01000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "01001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "01010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "01011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "01100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "01101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "01110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "01111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "10000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "10001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "10010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "10011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "10100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "10101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "10110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "10111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "11000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "11001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "11010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "11011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "11100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "11101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "11110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "11111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel6_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(5 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 64;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "000001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "000010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "000011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "000100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "000101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "000110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "000111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "001000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "001001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "001010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "001011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "001100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "001101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "001110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "001111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "010000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "010001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "010010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "010011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "010100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "010101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "010110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "010111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "011000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "011001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "011010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "011011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "011100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "011101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "011110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "011111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN "100000" =>
       result := inputs0( 33*size-1 DOWNTO 32*size);
     WHEN "100001" =>
       result := inputs0( 34*size-1 DOWNTO 33*size);
     WHEN "100010" =>
       result := inputs0( 35*size-1 DOWNTO 34*size);
     WHEN "100011" =>
       result := inputs0( 36*size-1 DOWNTO 35*size);
     WHEN "100100" =>
       result := inputs0( 37*size-1 DOWNTO 36*size);
     WHEN "100101" =>
       result := inputs0( 38*size-1 DOWNTO 37*size);
     WHEN "100110" =>
       result := inputs0( 39*size-1 DOWNTO 38*size);
     WHEN "100111" =>
       result := inputs0( 40*size-1 DOWNTO 39*size);
     WHEN "101000" =>
       result := inputs0( 41*size-1 DOWNTO 40*size);
     WHEN "101001" =>
       result := inputs0( 42*size-1 DOWNTO 41*size);
     WHEN "101010" =>
       result := inputs0( 43*size-1 DOWNTO 42*size);
     WHEN "101011" =>
       result := inputs0( 44*size-1 DOWNTO 43*size);
     WHEN "101100" =>
       result := inputs0( 45*size-1 DOWNTO 44*size);
     WHEN "101101" =>
       result := inputs0( 46*size-1 DOWNTO 45*size);
     WHEN "101110" =>
       result := inputs0( 47*size-1 DOWNTO 46*size);
     WHEN "101111" =>
       result := inputs0( 48*size-1 DOWNTO 47*size);
     WHEN "110000" =>
       result := inputs0( 49*size-1 DOWNTO 48*size);
     WHEN "110001" =>
       result := inputs0( 50*size-1 DOWNTO 49*size);
     WHEN "110010" =>
       result := inputs0( 51*size-1 DOWNTO 50*size);
     WHEN "110011" =>
       result := inputs0( 52*size-1 DOWNTO 51*size);
     WHEN "110100" =>
       result := inputs0( 53*size-1 DOWNTO 52*size);
     WHEN "110101" =>
       result := inputs0( 54*size-1 DOWNTO 53*size);
     WHEN "110110" =>
       result := inputs0( 55*size-1 DOWNTO 54*size);
     WHEN "110111" =>
       result := inputs0( 56*size-1 DOWNTO 55*size);
     WHEN "111000" =>
       result := inputs0( 57*size-1 DOWNTO 56*size);
     WHEN "111001" =>
       result := inputs0( 58*size-1 DOWNTO 57*size);
     WHEN "111010" =>
       result := inputs0( 59*size-1 DOWNTO 58*size);
     WHEN "111011" =>
       result := inputs0( 60*size-1 DOWNTO 59*size);
     WHEN "111100" =>
       result := inputs0( 61*size-1 DOWNTO 60*size);
     WHEN "111101" =>
       result := inputs0( 62*size-1 DOWNTO 61*size);
     WHEN "111110" =>
       result := inputs0( 63*size-1 DOWNTO 62*size);
     WHEN "111111" =>
       result := inputs0( 64*size-1 DOWNTO 63*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS  --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2 SEVERITY FAILURE;
     --synopsys translate_on
       CASE sel IS
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0( size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1  DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0(size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
       RETURN result;
   END;
--   BEGIN RETURN mux_v(inputs, TO_STDLOGICVECTOR(sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     ALIAS    sel0   : STD_LOGIC_VECTOR( sel'LENGTH-1 DOWNTO 0 ) IS sel;

     VARIABLE sellen : INTEGER RANGE 2-sel'LENGTH TO sel'LENGTH;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2**sel'LENGTH;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
     TYPE inputs_array_type is array(natural range <>) of std_logic_vector( olen - 1 DOWNTO 0);
     VARIABLE inputs_array : inputs_array_type( 2**sel'LENGTH - 1 DOWNTO 0);
   BEGIN
     sellen := sel'LENGTH;
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2**sellen SEVERITY FAILURE;
     sellen := 2-sellen;
     --synopsys translate_on
     CASE sellen IS
     WHEN 1 =>
       CASE sel0(0) IS

       WHEN '1' 
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0(  size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1 DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0( size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
     WHEN 2 =>
       result := mux_sel2_v(inputs, not sel);
     WHEN 3 =>
       result := mux_sel3_v(inputs, not sel);
     WHEN 4 =>
       result := mux_sel4_v(inputs, not sel);
     WHEN 5 =>
       result := mux_sel5_v(inputs, not sel);
     WHEN 6 =>
       result := mux_sel6_v(inputs, not sel);
     WHEN others =>
       -- synopsys translate_off
       IF(Is_X(sel0)) THEN
         result := (others => 'X');
       ELSE
       -- synopsys translate_on
         FOR i in 0 to 2**sel'LENGTH - 1 LOOP
           inputs_array(i) := inputs0( ((i + 1) * olen) - 1  DOWNTO i*olen);
         END LOOP;
         result := inputs_array(CONV_INTEGER( (UNSIGNED(NOT sel0)) ));
       -- synopsys translate_off
       END IF;
       -- synopsys translate_on
     END CASE;
     RETURN result;
   END;

 
-----------------------------------------------------------------
-- Latches
-----------------------------------------------------------------

   FUNCTION lat_s(dinput: STD_LOGIC; clk: STD_LOGIC; doutput: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN mux_s(STD_LOGIC_VECTOR'(doutput & dinput), clk); END;

   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR ; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR ) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     --synopsys translate_off
     ASSERT dinput'LENGTH = doutput'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN mux_v(doutput & dinput, clk);
   END;

-----------------------------------------------------------------
-- Tri-States
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC; control: STD_LOGIC) RETURN STD_LOGIC IS
--   BEGIN RETURN TO_STDLOGIC(tri_v(TO_STDLOGICVECTOR(dinput), control)); END;
--
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR ; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
--     VARIABLE result: STD_LOGIC_VECTOR(dinput'range);
--   BEGIN
--     CASE control IS
--     WHEN '0' | 'L' =>
--       result := (others => 'Z');
--     WHEN '1' | 'H' =>
--       FOR i IN dinput'range LOOP
--         result(i) := to_UX01(dinput(i));
--       END LOOP;
--     WHEN others =>
--       -- synopsys translate_off
--       result := (others => 'X');
--       -- synopsys translate_on
--     END CASE;
--     RETURN result;
--   END;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;

   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     VARIABLE diff: UNSIGNED(l'LENGTH DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     diff := ('0'&l) - ('0'&r);
     RETURN diff(l'LENGTH);
   END;
   FUNCTION "<"(l, r: SIGNED  ) RETURN STD_LOGIC IS
   BEGIN
     RETURN (UNSIGNED(l) < UNSIGNED(r)) xor (l(l'LEFT) xor r(r'LEFT));
   END;

   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION "<=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">"(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;
   FUNCTION ">=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;

   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN not or_s(l xor r);
   END;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   --some functions to placate spyglass
   FUNCTION mult_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a*b;
   END mult_natural;

   FUNCTION div_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a/b;
   END div_natural;

   FUNCTION mod_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a mod b;
   END mod_natural;

   FUNCTION add_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a+b;
   END add_unsigned;

   FUNCTION sub_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a-b;
   END sub_unsigned;

   FUNCTION sub_int(a,b : INTEGER) RETURN INTEGER IS
   BEGIN
     return a-b;
   END sub_int;

   FUNCTION concat_0(b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return '0' & b;
   END concat_0;

   FUNCTION concat_uns(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a&b;
   END concat_uns;

   FUNCTION concat_vect(a,b : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     return a&b;
   END concat_vect;





   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED IS
     CONSTANT ninps : NATURAL := arg'LENGTH / width;
     ALIAS    arg0  : UNSIGNED(arg'LENGTH-1 DOWNTO 0) IS arg;
     VARIABLE result: UNSIGNED(width-1 DOWNTO 0);
     VARIABLE from  : INTEGER;
     VARIABLE dto   : INTEGER;
   BEGIN
     --synopsys translate_off
     ASSERT arg'LENGTH = width * ninps SEVERITY FAILURE;
     --synopsys translate_on
     result := (OTHERS => '0');
     FOR i IN ninps-1 DOWNTO 0 LOOP
       --result := result + arg0((i+1)*width-1 DOWNTO i*width);
       from := mult_natural((i+1), width)-1; --2.1.6.3
       dto  := mult_natural(i,width); --2.1.6.3
       result := add_unsigned(result , arg0(from DOWNTO dto) );
     END LOOP;
     RETURN result;
   END faccu;

   FUNCTION  fabs (arg1: SIGNED) RETURN UNSIGNED IS
   BEGIN
     CASE arg1(arg1'LEFT) IS
     WHEN '1'
     --synopsys translate_off
          | 'H'
     --synopsys translate_on
       =>
       RETURN UNSIGNED'("0") - UNSIGNED(arg1);
     WHEN '0'
     --synopsys translate_off
          | 'L'
     --synopsys translate_on
       =>
       RETURN UNSIGNED(arg1);
     WHEN others =>
       RETURN resolve_unsigned(UNSIGNED(arg1), UNSIGNED'("0") - UNSIGNED(arg1));
     END CASE;
   END;

   PROCEDURE divmod(l, r: UNSIGNED; rdiv, rmod: OUT UNSIGNED) IS
     CONSTANT llen: INTEGER := l'LENGTH;
     CONSTANT rlen: INTEGER := r'LENGTH;
     CONSTANT llen_plus_rlen: INTEGER := llen + rlen;
     VARIABLE lbuf: UNSIGNED(llen+rlen-1 DOWNTO 0);
     VARIABLE diff: UNSIGNED(rlen DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT rdiv'LENGTH = llen AND rmod'LENGTH = rlen SEVERITY FAILURE;
     --synopsys translate_on
     lbuf := (others => '0');
     lbuf(llen-1 DOWNTO 0) := l;
     FOR i IN rdiv'range LOOP
       diff := sub_unsigned(lbuf(llen_plus_rlen-1 DOWNTO llen-1) ,(concat_0(r)));
       rdiv(i) := not diff(rlen);
       IF diff(rlen) = '0' THEN
         lbuf(llen_plus_rlen-1 DOWNTO llen-1) := diff;
       END IF;
       lbuf(llen_plus_rlen-1 DOWNTO 1) := lbuf(llen_plus_rlen-2 DOWNTO 0);
     END LOOP;
     rmod := lbuf(llen_plus_rlen-1 DOWNTO llen);
   END divmod;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rdiv;
   END "/";

   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rmod;
   END;

   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN l MOD r; END;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rdiv := UNSIGNED'("0") - rdiv;
     END IF;
     RETURN SIGNED(rdiv); -- overflow problem "1000" / "11"
   END "/";

   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
     CONSTANT rnul: UNSIGNED(r'LENGTH-1 DOWNTO 0) := (others => '0');
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     IF rmod /= rnul AND to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rmod := UNSIGNED(r) + rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "MOD";

   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "REM";

   FUNCTION mult_unsigned(l,r : UNSIGNED) return UNSIGNED is
   BEGIN
     return l*r; 
   END mult_unsigned;

   FUNCTION "**" (l, r : UNSIGNED) RETURN UNSIGNED IS
     CONSTANT llen  : NATURAL := l'LENGTH;
     VARIABLE result: UNSIGNED(llen-1 DOWNTO 0);
     VARIABLE fak   : UNSIGNED(llen-1 DOWNTO 0);
   BEGIN
     fak := l;
     result := (others => '0'); result(0) := '1';
     FOR i IN r'reverse_range LOOP
       --was:result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(result & (result*fak)), r(i)));
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR( concat_uns(result , mult_unsigned(result,fak) )), r(i)));

       fak := mult_unsigned(fak , fak);
     END LOOP;
     RETURN result;
   END "**";

   FUNCTION "**" (l, r : SIGNED) RETURN SIGNED IS
     CONSTANT rlen  : NATURAL := r'LENGTH;
     ALIAS    r0    : SIGNED(0 TO r'LENGTH-1) IS r;
     VARIABLE result: SIGNED(l'range);
   BEGIN
     CASE r(r'LEFT) IS
     WHEN '0'
   --synopsys translate_off
          | 'L'
   --synopsys translate_on
     =>
       result := SIGNED(UNSIGNED(l) ** UNSIGNED(r0(1 TO r'LENGTH-1)));
     WHEN '1'
   --synopsys translate_off
          | 'H'
   --synopsys translate_on
     =>
       result := (others => '0');
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END "**";

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-----------------------------------------------------------------

   FUNCTION add_nat(arg1 : NATURAL; arg2 : NATURAL ) RETURN NATURAL IS
   BEGIN
     return (arg1 + arg2);
   END;
   
--   FUNCTION UNSIGNED_2_BIT_VECTOR(arg1 : NATURAL; arg2 : NATURAL ) RETURN BIT_VECTOR IS
--   BEGIN
--     return (arg1 + arg2);
--   END;
   
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(SIGNED(result), arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
        =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
        =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;


   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     --SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: NATURAL range 1 TO len;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => '0');
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         --was:temp(i2+sw) := result(i2);
         temp_idx := add_nat(i2,sw);
         temp(temp_idx) := result(i2);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: sw_range;
     VARIABLE result_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => sbit);
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         -- was: temp(i2) := result(i2+sw);
         result_idx := add_nat(i2,sw);
         temp(i2) := result(result_idx);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;


   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := arg1'LENGTH;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     VARIABLE temp: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     SUBTYPE sw_range IS NATURAL range 0 TO len-1;
     VARIABLE sw: sw_range;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     result := (others=>'0');
     result := arg1;
     sw := sdir MOD len;
     FOR i IN arg2'reverse_range LOOP
       EXIT WHEN sw = 0;
       IF signd2 AND i = arg2'LEFT THEN 
         sw := sub_int(len,sw); 
       END IF;
       -- temp := result(len-sw-1 DOWNTO 0) & result(len-1 DOWNTO len-sw)
       FOR i2 IN len-1 DOWNTO 0 LOOP
         --was: temp((i2+sw) MOD len) := result(i2);
         temp_idx := add_nat(i2,sw) MOD len;
         temp(temp_idx) := result(i2);
       END LOOP;
       result := mux_v(STD_LOGIC_VECTOR(concat_vect(result,temp)), arg2(i));
       sw := mod_natural(mult_natural(sw,2), len);
     END LOOP;
     RETURN result;
   END frot;

   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, -1); END;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, -1); END;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC IS
     CONSTANT len : INTEGER := vec'LENGTH;
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
   BEGIN
     IF index >= len OR index < 0 THEN
       RETURN 'X';
     END IF;
     RETURN vec0(index);
   END;

   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     CONSTANT indexPwidthM1 : INTEGER := index+width-1; --2.1.6.3
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
     CONSTANT xxx : STD_LOGIC_VECTOR(width-1 DOWNTO 0) := (others => 'X');
   BEGIN
     IF index+width > len OR index < 0 THEN
       RETURN xxx;
     END IF;
     RETURN vec0(indexPwidthM1 DOWNTO index);
   END;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     VARIABLE vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     CONSTANT xxx : STD_LOGIC_VECTOR(len-1 DOWNTO 0) := (others => 'X');
   BEGIN
     vec0 := vec;
     IF index >= len OR index < 0 THEN
       RETURN xxx;
     END IF;
     vec0(index) := dinput;
     RETURN vec0;
   END;

   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE IS
     VARIABLE n_b : POSITIVE;
     VARIABLE p_v : NATURAL;
   BEGIN
     p_v := p;
     FOR i IN 1 TO 32 LOOP
       p_v := div_natural(p_v,2);
       n_b := i;
       EXIT WHEN (p_v = 0);
     END LOOP;
     RETURN n_b;
   END;


--   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
--
--     CONSTANT vlen: INTEGER := vec'LENGTH;
--     CONSTANT ilen: INTEGER := dinput'LENGTH;
--     CONSTANT max_shift: INTEGER := vlen-ilen;
--     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
--     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
--     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
--     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
--     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
--     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
--   BEGIN
--     inp := (others => '0');
--     mask := (others => '0');
--
--     IF index > max_shift OR index < 0 THEN
--       RETURN xxx;
--     END IF;
--
--     shift := CONV_UNSIGNED(index, shift'LENGTH);
--     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
--     mask(ilen-1 DOWNTO 0) := ones;
--     inp := fshl(inp, shift, vlen);
--     mask := fshl(mask, shift, vlen);
--     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
--     RETURN vec0;
--   END;

   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR IS

     type enable_matrix is array (0 to enable'LENGTH-1 ) of std_logic_vector(byte_width-1 downto 0);
     CONSTANT vlen: INTEGER := vec'LENGTH;
     CONSTANT ilen: INTEGER := dinput'LENGTH;
     CONSTANT max_shift: INTEGER := vlen-ilen;
     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask2: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE enables: enable_matrix;
     VARIABLE cat_enables: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0 );
     VARIABLE lsbi : INTEGER;
     VARIABLE msbi : INTEGER;

   BEGIN
     cat_enables := (others => '0');
     lsbi := 0;
     msbi := byte_width-1;
     inp := (others => '0');
     mask := (others => '0');

     IF index > max_shift OR index < 0 THEN
       RETURN xxx;
     END IF;

     --initialize enables
     for i in 0 TO (enable'LENGTH-1) loop
       enables(i)  := (others => enable(i));
       cat_enables(msbi downto lsbi) := enables(i) ;
       lsbi := msbi+1;
       msbi := msbi+byte_width;
     end loop;


     shift := CONV_UNSIGNED(index, shift'LENGTH);
     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
     mask(ilen-1 DOWNTO 0) := UNSIGNED((STD_LOGIC_VECTOR(ones) AND cat_enables));
     inp := fshl(inp, shift, vlen);
     mask := fshl(mask, shift, vlen);
     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
     RETURN vec0;
   END;


   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;
   
   FUNCTION bits(size : NATURAL) return NATURAL is
   begin
     return ceil_log2(size);
   END;

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH) xor conv_std_logic_vector(c, s'LENGTH);
     cout := ( (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH)) or (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) or (conv_std_logic_vector(b, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) );
   END PROCEDURE csa;

   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH);
     cout := (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH));
   END PROCEDURE csha;

END funcs;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_comps.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_comps IS
 
FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
FUNCTION ceil_log2(size : NATURAL) return NATURAL;
 

COMPONENT mgc_not
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_and
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nand
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_or
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xnor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux
  GENERIC (
    width  :  NATURAL;
    ctrlw  :  NATURAL;
    p2ctrlw : NATURAL := 0
  );
  PORT (
    a: in  std_logic_vector(width*(2**ctrlw) - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw            - 1 DOWNTO 0);
    z: out std_logic_vector(width            - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux1hot
  GENERIC (
    width  : NATURAL;
    ctrlw  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ctrlw - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw       - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_reg_pos
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;  -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL  -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_reg_neg
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;   -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_generic_reg
  GENERIC(
   width: natural := 8;
   ph_clk: integer range 0 to 1 := 1; -- clock polarity, 1=rising_edge
   ph_en: integer range 0 to 1 := 1;
   ph_a_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   ph_s_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   a_rst_used: integer range 0 to 1 := 1;
   s_rst_used: integer range 0 to 1 := 0;
   en_used: integer range 0 to 1 := 1
  );
  PORT(
   d: std_logic_vector(width-1 downto 0);
   clk: in std_logic;
   en: in std_logic;
   a_rst: in std_logic;
   s_rst: in std_logic;
   q: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_equal
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a : in  std_logic_vector(width-1 DOWNTO 0);
    b : in  std_logic_vector(width-1 DOWNTO 0);
    eq: out std_logic;
    ne: out std_logic
  );
END COMPONENT;

COMPONENT mgc_shift_l
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rot
  GENERIC (
    width  : NATURAL;
    width_s: NATURAL;
    signd_s: NATURAL;      -- 0:unsigned 1:signed
    sleft  : NATURAL;      -- 0:right 1:left;
    log2w  : NATURAL := 0; -- LOG2(width)
    l2wp2  : NATURAL := 0  --2**LOG2(width)
  );
  PORT (
    a : in  std_logic_vector(width  -1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width  -1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_sub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_ci
  GENERIC (
    width_a : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width_a, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width_a, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width_a,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width_a,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_addc
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add3
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_c : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_c : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(ifeqsel(width_c,0,width,width_c)-1 DOWNTO 0);
    d: in  std_logic_vector(0 DOWNTO 0);
    e: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_sub_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addc_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     c: in std_logic_vector(0 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addsub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    add: in  std_logic;
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_accu
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_abs
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_fast
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_pipe
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2  : NATURAL;
    add_d2  : NATURAL
  );
  PORT (
    a   : in  std_logic_vector(width_a-1 DOWNTO 0);
    b   : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2  : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c   : in  std_logic_vector(width_c-1 DOWNTO 0);
    d   : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2  : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst : in  std_logic_vector(width_e-1 DOWNTO 0);
    z   : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1_pipe
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2   : NATURAL;
    add_d2   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2     : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2     : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_e-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL
  );
  PORT (
    a:   in  std_logic_vector(width_a-1 DOWNTO 0);
    b:   in  std_logic_vector(width_b-1 DOWNTO 0);
    c:   in  std_logic_vector(width_c-1 DOWNTO 0);
    cst: in  std_logic_vector(width_cst-1 DOWNTO 0);
    d:   in  std_logic_vector(width_d-1 DOWNTO 0);
    z:   out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1_pipe
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_cst-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mulacc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2acc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    add_cxd : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    d         : in  std_logic_vector(width_d-1 DOWNTO 0);
    e         : in  std_logic_vector(width_e-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_div
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mod
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rem
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_csa
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     c: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_csha
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_rom
    GENERIC (
      rom_id : natural := 1;
      size : natural := 33;
      width : natural := 32
      );
    PORT (
      data_in : std_logic_vector((size*width)-1 downto 0);
      addr : std_logic_vector(ceil_log2(size)-1 downto 0);
      data_out : out std_logic_vector(width-1 downto 0)
    );
END COMPONENT;

END mgc_comps;

PACKAGE BODY mgc_comps IS
 
   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;
 
END mgc_comps;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_mul_pipe IS
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_mul_pipe;

LIBRARY IEEE;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_mul_pipe IS
  TYPE reg_array_type is array(natural range<>) of std_logic_vector(width_z-1 DOWNTO 0); 
  SIGNAL xz : std_logic_vector(width_a+width_b DOWNTO 0);

--MF Added pipelined input
    signal a_f     : STD_LOGIC_VECTOR(width_a-1 downto 0); 
    signal b_f     : STD_LOGIC_VECTOR(width_b-1 downto 0);
   type a_array is array (natural range <>) of STD_LOGIC_VECTOR(width_a-1 downto 0);
   type b_array is array (natural range <>) of STD_LOGIC_VECTOR(width_b-1 downto 0);
BEGIN
  n_inreg_gt_0: if n_inreg > 0 generate
    GENPOS_INREG: IF clock_edge = 1 GENERATE
     I0: process(clk)
        variable a_in_reg: a_array(n_inreg-1 downto 0);
        variable b_in_reg: b_array(n_inreg-1 downto 0);
      begin
        if (clk'event and clk = '1' ) then
          if (conv_integer(en) = enable_active) then
            for i in n_inreg - 2 downto 0 loop
              a_in_reg(i+1) := a_in_reg(i);
              b_in_reg(i+1) := b_in_reg(i);
            end loop;                                                                                                                             
            a_in_reg(0) := a;
            b_in_reg(0) := b;

            a_f <= a_in_reg(n_inreg-1);             
            b_f <= b_in_reg(n_inreg-1);    
                                                   
          end if;
        end if;
      end process;
    END GENERATE;
  
   GENNEG_INREG: IF clock_edge = 0 GENERATE
     I0: process(clk)
        variable a_in_reg: a_array(n_inreg-1 downto 0);
        variable b_in_reg: b_array(n_inreg-1 downto 0);
      begin
        if (clk'event and clk = '0' ) then
          if (conv_integer(en) = enable_active) then
            for i in n_inreg - 2 downto 0 loop
              a_in_reg(i+1) := a_in_reg(i);
              b_in_reg(i+1) := b_in_reg(i);
            end loop;                                                                                                                             
            a_in_reg(0) := a;
            b_in_reg(0) := b;            
                                 
            a_f <= a_in_reg(n_inreg-1);             
            b_f <= b_in_reg(n_inreg-1);
                                                        
          end if;
        end if;
      end process;
    END GENERATE;
  END GENERATE;

  n_inreg_eq_0: if n_inreg = 0 generate
    a_f <= a;
    b_f <= b;
  end generate n_inreg_eq_0;

  xz <= '0'&(unsigned(a_f) * unsigned(b_f)) WHEN signd_a = 0 AND signd_b = 0 ELSE
            (  signed(a_f) * unsigned(b_f)) WHEN signd_a = 1 AND signd_b = 0 ELSE
            (unsigned(a_f) *   signed(b_f)) WHEN signd_a = 0 AND signd_b = 1 ELSE
        '0'&(  signed(a_f) *   signed(b_f));

  GENPOS: IF clock_edge = 1 GENERATE
    PROCESS (clk)
    VARIABLE reg_array: reg_array_type(stages-2 DOWNTO 0);
    BEGIN
      IF ( clk'EVENT AND clk = '1') THEN
        IF ( conv_integer(en) = enable_active) THEN
          FOR I IN stages-2 DOWNTO 1 LOOP
            reg_array(I) := reg_array(I-1);
          END LOOP;
          reg_array(0) := xz(width_z-1 DOWNTO 0);
          z <= reg_array(stages-2);
        END IF;
      END IF;
    END PROCESS;
  END GENERATE;

  GENNEG: IF clock_edge = 0 GENERATE
    PROCESS (clk)
    VARIABLE reg_array: reg_array_type(stages-2 DOWNTO 0);
    BEGIN
      IF ( clk'EVENT AND clk = '0') THEN
        IF ( conv_integer(en) = enable_active) THEN
          FOR I IN stages-2 DOWNTO 1 LOOP
            reg_array(I) := reg_array(I-1);
          END LOOP;
          reg_array(0) := xz(width_z-1 DOWNTO 0);
          z <= reg_array(stages-2);
        END IF;
      END IF;
    END PROCESS;
  END GENERATE;
END beh;

--------> ../td_ccore_solutions/mult_b3d4a0c17af05a92530fe047f70695c970ca_0/rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Mon Sep 13 16:20:57 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    mult_core_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;
USE work.mgc_comps.ALL;


ENTITY mult_core_wait_dp IS
  PORT(
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC;
    ensig_cgo_iro : IN STD_LOGIC;
    z_mul_cmp_z : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    z_mul_cmp_1_z : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    ensig_cgo : IN STD_LOGIC;
    t_mul_cmp_en : OUT STD_LOGIC;
    z_mul_cmp_z_oreg : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    z_mul_cmp_1_z_oreg : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END mult_core_wait_dp;

ARCHITECTURE v1 OF mult_core_wait_dp IS
  -- Default Constants

BEGIN
  t_mul_cmp_en <= ccs_ccore_en AND (ensig_cgo OR ensig_cgo_iro);
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( ccs_ccore_en = '1' ) THEN
        z_mul_cmp_z_oreg <= z_mul_cmp_z;
        z_mul_cmp_1_z_oreg <= z_mul_cmp_1_z;
      END IF;
    END IF;
  END PROCESS;
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    mult_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;
USE work.mgc_comps.ALL;


ENTITY mult_core IS
  PORT(
    x_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    y_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    y_rsc_dat_1 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    p_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    return_rsc_z : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    ccs_ccore_start_rsc_dat : IN STD_LOGIC;
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_srst : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC;
    z_mul_cmp_a : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    z_mul_cmp_b : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    z_mul_cmp_z : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    z_mul_cmp_1_a : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    z_mul_cmp_1_b : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    z_mul_cmp_1_z : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END mult_core;

ARCHITECTURE v1 OF mult_core IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Output Reader Declarations
  SIGNAL z_mul_cmp_1_b_drv : STD_LOGIC_VECTOR (31 DOWNTO 0);

  -- Interconnect Declarations
  SIGNAL x_rsci_idat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL y_rsci_idat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL y_rsci_idat_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL p_rsci_idat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL return_rsci_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL ccs_ccore_start_rsci_idat : STD_LOGIC;
  SIGNAL t_mul_cmp_en : STD_LOGIC;
  SIGNAL t_mul_cmp_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL z_mul_cmp_z_oreg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_mul_cmp_1_z_oreg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL and_dcpl : STD_LOGIC;
  SIGNAL main_stage_0_2 : STD_LOGIC;
  SIGNAL VEC_LOOP_asn_itm_1 : STD_LOGIC;
  SIGNAL main_stage_0_4 : STD_LOGIC;
  SIGNAL VEC_LOOP_asn_itm_3 : STD_LOGIC;
  SIGNAL slc_32_svs_1 : STD_LOGIC;
  SIGNAL VEC_LOOP_asn_itm_2 : STD_LOGIC;
  SIGNAL main_stage_0_3 : STD_LOGIC;
  SIGNAL reg_CGHpart_irsig_cse : STD_LOGIC;
  SIGNAL reg_t_mul_cmp_a_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL and_4_cse : STD_LOGIC;
  SIGNAL and_8_cse : STD_LOGIC;
  SIGNAL t_or_rmff : STD_LOGIC;
  SIGNAL main_stage_0_5 : STD_LOGIC;
  SIGNAL main_stage_0_6 : STD_LOGIC;
  SIGNAL p_buf_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL p_buf_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL p_buf_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL p_buf_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL p_buf_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_asn_itm_4 : STD_LOGIC;
  SIGNAL VEC_LOOP_asn_itm_5 : STD_LOGIC;
  SIGNAL res_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL res_and_cse : STD_LOGIC;
  SIGNAL p_and_2_cse : STD_LOGIC;
  SIGNAL p_and_1_cse : STD_LOGIC;
  SIGNAL if_acc_1_itm_32_1 : STD_LOGIC;

  SIGNAL if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL x_rsci_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsci_idat_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL y_rsci_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL y_rsci_idat_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL y_rsci_1_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL y_rsci_1_idat : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL p_rsci_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL p_rsci_idat_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL return_rsci_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL return_rsci_z : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL ccs_ccore_start_rsci_dat : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL ccs_ccore_start_rsci_idat_1 : STD_LOGIC_VECTOR (0 DOWNTO 0);

  SIGNAL t_mul_cmp_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL t_mul_cmp_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL t_mul_cmp_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT mult_core_wait_dp
    PORT(
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC;
      ensig_cgo_iro : IN STD_LOGIC;
      z_mul_cmp_z : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      z_mul_cmp_1_z : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      ensig_cgo : IN STD_LOGIC;
      t_mul_cmp_en : OUT STD_LOGIC;
      z_mul_cmp_z_oreg : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      z_mul_cmp_1_z_oreg : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL mult_core_wait_dp_inst_z_mul_cmp_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_core_wait_dp_inst_z_mul_cmp_1_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_core_wait_dp_inst_z_mul_cmp_z_oreg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_core_wait_dp_inst_z_mul_cmp_1_z_oreg : STD_LOGIC_VECTOR (31 DOWNTO
      0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  z_mul_cmp_1_b <= z_mul_cmp_1_b_drv;

  x_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 7,
      width => 32
      )
    PORT MAP(
      dat => x_rsci_dat,
      idat => x_rsci_idat_1
    );
  x_rsci_dat <= x_rsc_dat;
  x_rsci_idat <= x_rsci_idat_1;

  y_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 8,
      width => 32
      )
    PORT MAP(
      dat => y_rsci_dat,
      idat => y_rsci_idat_2
    );
  y_rsci_dat <= y_rsc_dat;
  y_rsci_idat <= y_rsci_idat_2;

  y_rsci_1 : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 9,
      width => 32
      )
    PORT MAP(
      dat => y_rsci_1_dat,
      idat => y_rsci_1_idat
    );
  y_rsci_1_dat <= y_rsc_dat_1;
  y_rsci_idat_1 <= y_rsci_1_idat;

  p_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 10,
      width => 32
      )
    PORT MAP(
      dat => p_rsci_dat,
      idat => p_rsci_idat_1
    );
  p_rsci_dat <= p_rsc_dat;
  p_rsci_idat <= p_rsci_idat_1;

  return_rsci : work.mgc_out_dreg_pkg_v2.mgc_out_dreg_v2
    GENERIC MAP(
      rscid => 11,
      width => 32
      )
    PORT MAP(
      d => return_rsci_d_1,
      z => return_rsci_z
    );
  return_rsci_d_1 <= return_rsci_d;
  return_rsc_z <= return_rsci_z;

  ccs_ccore_start_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 19,
      width => 1
      )
    PORT MAP(
      dat => ccs_ccore_start_rsci_dat,
      idat => ccs_ccore_start_rsci_idat_1
    );
  ccs_ccore_start_rsci_dat(0) <= ccs_ccore_start_rsc_dat;
  ccs_ccore_start_rsci_idat <= ccs_ccore_start_rsci_idat_1(0);

  t_mul_cmp : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 64,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => t_mul_cmp_a,
      b => t_mul_cmp_b,
      clk => ccs_ccore_clk,
      en => t_mul_cmp_en,
      a_rst => '1',
      s_rst => ccs_ccore_srst,
      z => t_mul_cmp_z_1
    );
  t_mul_cmp_a <= x_rsci_idat;
  t_mul_cmp_b <= y_rsci_idat_1;
  t_mul_cmp_z <= t_mul_cmp_z_1;

  mult_core_wait_dp_inst : mult_core_wait_dp
    PORT MAP(
      ccs_ccore_clk => ccs_ccore_clk,
      ccs_ccore_en => ccs_ccore_en,
      ensig_cgo_iro => t_or_rmff,
      z_mul_cmp_z => mult_core_wait_dp_inst_z_mul_cmp_z,
      z_mul_cmp_1_z => mult_core_wait_dp_inst_z_mul_cmp_1_z,
      ensig_cgo => reg_CGHpart_irsig_cse,
      t_mul_cmp_en => t_mul_cmp_en,
      z_mul_cmp_z_oreg => mult_core_wait_dp_inst_z_mul_cmp_z_oreg,
      z_mul_cmp_1_z_oreg => mult_core_wait_dp_inst_z_mul_cmp_1_z_oreg
    );
  mult_core_wait_dp_inst_z_mul_cmp_z <= z_mul_cmp_z;
  mult_core_wait_dp_inst_z_mul_cmp_1_z <= z_mul_cmp_1_z;
  z_mul_cmp_z_oreg <= mult_core_wait_dp_inst_z_mul_cmp_z_oreg;
  z_mul_cmp_1_z_oreg <= mult_core_wait_dp_inst_z_mul_cmp_1_z_oreg;

  res_and_cse <= ccs_ccore_en AND and_dcpl;
  p_and_1_cse <= ccs_ccore_en AND and_8_cse;
  t_or_rmff <= and_8_cse OR and_4_cse OR ccs_ccore_start_rsci_idat;
  z_mul_cmp_a <= reg_t_mul_cmp_a_cse;
  p_and_2_cse <= ccs_ccore_en AND main_stage_0_5 AND VEC_LOOP_asn_itm_4;
  and_4_cse <= main_stage_0_2 AND VEC_LOOP_asn_itm_1;
  res_sva_3 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(z_asn_itm_3) - UNSIGNED(z_mul_cmp_1_z_oreg),
      32));
  if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & res_sva_3) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT
      p_buf_sva_5), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"), 33));
  if_acc_1_itm_32_1 <= if_acc_1_nl(32);
  and_8_cse <= main_stage_0_3 AND VEC_LOOP_asn_itm_2;
  and_dcpl <= main_stage_0_6 AND VEC_LOOP_asn_itm_5;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( ccs_ccore_en = '1' ) THEN
        return_rsci_d <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(if_acc_nl),
            32)), res_sva_1, slc_32_svs_1);
        z_mul_cmp_1_b_drv <= p_buf_sva_3;
        z_mul_cmp_1_a <= t_mul_cmp_z(63 DOWNTO 32);
        reg_t_mul_cmp_a_cse <= x_rsci_idat;
        z_mul_cmp_b <= y_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        VEC_LOOP_asn_itm_5 <= '0';
        VEC_LOOP_asn_itm_3 <= '0';
        reg_CGHpart_irsig_cse <= '0';
        VEC_LOOP_asn_itm_2 <= '0';
        VEC_LOOP_asn_itm_1 <= '0';
        main_stage_0_2 <= '0';
        main_stage_0_3 <= '0';
        main_stage_0_4 <= '0';
        main_stage_0_6 <= '0';
        VEC_LOOP_asn_itm_4 <= '0';
        main_stage_0_5 <= '0';
      ELSIF ( ccs_ccore_en = '1' ) THEN
        VEC_LOOP_asn_itm_5 <= VEC_LOOP_asn_itm_4;
        VEC_LOOP_asn_itm_3 <= VEC_LOOP_asn_itm_2;
        reg_CGHpart_irsig_cse <= t_or_rmff;
        VEC_LOOP_asn_itm_2 <= VEC_LOOP_asn_itm_1;
        VEC_LOOP_asn_itm_1 <= ccs_ccore_start_rsci_idat;
        main_stage_0_2 <= '1';
        main_stage_0_3 <= main_stage_0_2;
        main_stage_0_4 <= main_stage_0_3;
        main_stage_0_6 <= main_stage_0_5;
        VEC_LOOP_asn_itm_4 <= VEC_LOOP_asn_itm_3;
        main_stage_0_5 <= main_stage_0_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( res_and_cse = '1' ) THEN
        res_sva_1 <= res_sva_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        slc_32_svs_1 <= '0';
      ELSIF ( res_and_cse = '1' ) THEN
        slc_32_svs_1 <= if_acc_1_itm_32_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( (ccs_ccore_en AND and_dcpl AND (NOT if_acc_1_itm_32_1)) = '1' ) THEN
        p_buf_sva_6 <= p_buf_sva_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( p_and_1_cse = '1' ) THEN
        p_buf_sva_3 <= p_buf_sva_2;
        z_asn_itm_1 <= z_mul_cmp_z_oreg;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( p_and_2_cse = '1' ) THEN
        p_buf_sva_5 <= z_mul_cmp_1_b_drv;
        z_asn_itm_3 <= z_asn_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( (ccs_ccore_en AND and_4_cse) = '1' ) THEN
        p_buf_sva_2 <= p_buf_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( (ccs_ccore_en AND main_stage_0_4 AND VEC_LOOP_asn_itm_3) = '1' ) THEN
        z_asn_itm_2 <= z_asn_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( (ccs_ccore_en AND ccs_ccore_start_rsci_idat) = '1' ) THEN
        p_buf_sva_1 <= p_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(res_sva_1) - UNSIGNED(p_buf_sva_6),
      32));
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    mult
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;
USE work.mgc_comps.ALL;


ENTITY mult IS
  PORT(
    x_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    y_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    y_rsc_dat_1 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    p_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    return_rsc_z : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    ccs_ccore_start_rsc_dat : IN STD_LOGIC;
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_srst : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC
  );
END mult;

ARCHITECTURE v1 OF mult IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL z_mul_cmp_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_mul_cmp_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_mul_cmp_1_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_mul_cmp_1_b : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT mult_core
    PORT(
      x_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      y_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      y_rsc_dat_1 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      p_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      return_rsc_z : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      ccs_ccore_start_rsc_dat : IN STD_LOGIC;
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_srst : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC;
      z_mul_cmp_a : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      z_mul_cmp_b : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      z_mul_cmp_z : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      z_mul_cmp_1_a : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      z_mul_cmp_1_b : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      z_mul_cmp_1_z : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL mult_core_inst_x_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_core_inst_y_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_core_inst_y_rsc_dat_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_core_inst_p_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_core_inst_return_rsc_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_core_inst_z_mul_cmp_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_core_inst_z_mul_cmp_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_core_inst_z_mul_cmp_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_core_inst_z_mul_cmp_1_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_core_inst_z_mul_cmp_1_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_core_inst_z_mul_cmp_1_z : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  mult_core_inst : mult_core
    PORT MAP(
      x_rsc_dat => mult_core_inst_x_rsc_dat,
      y_rsc_dat => mult_core_inst_y_rsc_dat,
      y_rsc_dat_1 => mult_core_inst_y_rsc_dat_1,
      p_rsc_dat => mult_core_inst_p_rsc_dat,
      return_rsc_z => mult_core_inst_return_rsc_z,
      ccs_ccore_start_rsc_dat => ccs_ccore_start_rsc_dat,
      ccs_ccore_clk => ccs_ccore_clk,
      ccs_ccore_srst => ccs_ccore_srst,
      ccs_ccore_en => ccs_ccore_en,
      z_mul_cmp_a => mult_core_inst_z_mul_cmp_a,
      z_mul_cmp_b => mult_core_inst_z_mul_cmp_b,
      z_mul_cmp_z => mult_core_inst_z_mul_cmp_z,
      z_mul_cmp_1_a => mult_core_inst_z_mul_cmp_1_a,
      z_mul_cmp_1_b => mult_core_inst_z_mul_cmp_1_b,
      z_mul_cmp_1_z => mult_core_inst_z_mul_cmp_1_z
    );
  mult_core_inst_x_rsc_dat <= x_rsc_dat;
  mult_core_inst_y_rsc_dat <= y_rsc_dat;
  mult_core_inst_y_rsc_dat_1 <= y_rsc_dat_1;
  mult_core_inst_p_rsc_dat <= p_rsc_dat;
  return_rsc_z <= mult_core_inst_return_rsc_z;
  z_mul_cmp_a <= mult_core_inst_z_mul_cmp_a;
  z_mul_cmp_b <= mult_core_inst_z_mul_cmp_b;
  mult_core_inst_z_mul_cmp_z <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( UNSIGNED(z_mul_cmp_a)
      * UNSIGNED(z_mul_cmp_b)), 32));
  z_mul_cmp_1_a <= mult_core_inst_z_mul_cmp_1_a;
  z_mul_cmp_1_b <= mult_core_inst_z_mul_cmp_1_b;
  mult_core_inst_z_mul_cmp_1_z <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( UNSIGNED(z_mul_cmp_1_a)
      * UNSIGNED(z_mul_cmp_1_b)), 32));

END v1;




--------> ../td_ccore_solutions/modulo_sub_cc250ff62aef060f45cde5681b558542635b_0/rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Mon Sep 13 16:20:58 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    modulo_sub_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;


ENTITY modulo_sub_core IS
  PORT(
    base_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    m_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    return_rsc_z : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC
  );
END modulo_sub_core;

ARCHITECTURE v1 OF modulo_sub_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL base_rsci_idat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL m_rsci_idat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL return_rsci_d : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL qif_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL base_rsci_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL base_rsci_idat_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL m_rsci_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL m_rsci_idat_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL return_rsci_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL return_rsci_z : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  base_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 4,
      width => 32
      )
    PORT MAP(
      dat => base_rsci_dat,
      idat => base_rsci_idat_1
    );
  base_rsci_dat <= base_rsc_dat;
  base_rsci_idat <= base_rsci_idat_1;

  m_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 5,
      width => 32
      )
    PORT MAP(
      dat => m_rsci_dat,
      idat => m_rsci_idat_1
    );
  m_rsci_dat <= m_rsc_dat;
  m_rsci_idat <= m_rsci_idat_1;

  return_rsci : work.mgc_out_dreg_pkg_v2.mgc_out_dreg_v2
    GENERIC MAP(
      rscid => 6,
      width => 32
      )
    PORT MAP(
      d => return_rsci_d_1,
      z => return_rsci_z
    );
  return_rsci_d_1 <= return_rsci_d;
  return_rsc_z <= return_rsci_z;

  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( ccs_ccore_en = '1' ) THEN
        return_rsci_d <= MUX_v_32_2_2(('0' & (base_rsci_idat(30 DOWNTO 0))), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(qif_acc_nl),
            32)), base_rsci_idat(31));
      END IF;
    END IF;
  END PROCESS;
  qif_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & (base_rsci_idat(30
      DOWNTO 0))) + UNSIGNED(m_rsci_idat), 32));
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    modulo_sub
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;


ENTITY modulo_sub IS
  PORT(
    base_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    m_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    return_rsc_z : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    ccs_ccore_start_rsc_dat : IN STD_LOGIC;
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_srst : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC
  );
END modulo_sub;

ARCHITECTURE v1 OF modulo_sub IS
  -- Default Constants

  COMPONENT modulo_sub_core
    PORT(
      base_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      m_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      return_rsc_z : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL modulo_sub_core_inst_base_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_core_inst_m_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_core_inst_return_rsc_z : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  modulo_sub_core_inst : modulo_sub_core
    PORT MAP(
      base_rsc_dat => modulo_sub_core_inst_base_rsc_dat,
      m_rsc_dat => modulo_sub_core_inst_m_rsc_dat,
      return_rsc_z => modulo_sub_core_inst_return_rsc_z,
      ccs_ccore_clk => ccs_ccore_clk,
      ccs_ccore_en => ccs_ccore_en
    );
  modulo_sub_core_inst_base_rsc_dat <= base_rsc_dat;
  modulo_sub_core_inst_m_rsc_dat <= m_rsc_dat;
  return_rsc_z <= modulo_sub_core_inst_return_rsc_z;

END v1;




--------> ../td_ccore_solutions/modulo_add_12aaf73a68dd9ce714254cc9a57be62160d2_0/rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Mon Sep 13 16:21:00 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    modulo_add_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;


ENTITY modulo_add_core IS
  PORT(
    base_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    m_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    return_rsc_z : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC
  );
END modulo_add_core;

ARCHITECTURE v1 OF modulo_add_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL base_rsci_idat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL m_rsci_idat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL return_rsci_d : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL qif_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL base_rsci_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL base_rsci_idat_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL m_rsci_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL m_rsci_idat_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL return_rsci_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL return_rsci_z : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  base_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 1,
      width => 32
      )
    PORT MAP(
      dat => base_rsci_dat,
      idat => base_rsci_idat_1
    );
  base_rsci_dat <= base_rsc_dat;
  base_rsci_idat <= base_rsci_idat_1;

  m_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 2,
      width => 32
      )
    PORT MAP(
      dat => m_rsci_dat,
      idat => m_rsci_idat_1
    );
  m_rsci_dat <= m_rsc_dat;
  m_rsci_idat <= m_rsci_idat_1;

  return_rsci : work.mgc_out_dreg_pkg_v2.mgc_out_dreg_v2
    GENERIC MAP(
      rscid => 3,
      width => 32
      )
    PORT MAP(
      d => return_rsci_d_1,
      z => return_rsci_z
    );
  return_rsci_d_1 <= return_rsci_d;
  return_rsc_z <= return_rsci_z;

  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( ccs_ccore_en = '1' ) THEN
        return_rsci_d <= MUX_v_32_2_2(base_rsci_idat, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(qif_acc_nl),
            32)), acc_nl(33));
      END IF;
    END IF;
  END PROCESS;
  qif_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(base_rsci_idat) - UNSIGNED(m_rsci_idat),
      32));
  acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(m_rsci_idat),
      32), 34) - CONV_UNSIGNED(CONV_SIGNED(SIGNED(base_rsci_idat), 32), 34), 34));
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    modulo_add
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;


ENTITY modulo_add IS
  PORT(
    base_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    m_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    return_rsc_z : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    ccs_ccore_start_rsc_dat : IN STD_LOGIC;
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_srst : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC
  );
END modulo_add;

ARCHITECTURE v1 OF modulo_add IS
  -- Default Constants

  COMPONENT modulo_add_core
    PORT(
      base_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      m_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      return_rsc_z : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL modulo_add_core_inst_base_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_core_inst_m_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_core_inst_return_rsc_z : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  modulo_add_core_inst : modulo_add_core
    PORT MAP(
      base_rsc_dat => modulo_add_core_inst_base_rsc_dat,
      m_rsc_dat => modulo_add_core_inst_m_rsc_dat,
      return_rsc_z => modulo_add_core_inst_return_rsc_z,
      ccs_ccore_clk => ccs_ccore_clk,
      ccs_ccore_en => ccs_ccore_en
    );
  modulo_add_core_inst_base_rsc_dat <= base_rsc_dat;
  modulo_add_core_inst_m_rsc_dat <= m_rsc_dat;
  return_rsc_z <= modulo_add_core_inst_return_rsc_z;

END v1;




--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_comps_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_shift_comps_v5 IS

COMPONENT mgc_shift_l_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_shift_comps_v5;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_shift_l_v5 IS
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_shift_l_v5;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_shift_l_v5 IS

  FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1 > arg2) THEN
      RETURN(arg1) ;
    ELSE
      RETURN(arg2) ;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(SIGNED(result), arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE)
  RETURN UNSIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, '0', olen);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE)
  RETURN SIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen);
  END;

BEGIN
UNSGNED:  IF signd_a = 0 GENERATE
    z <= std_logic_vector(fshl_stdar(unsigned(a), unsigned(s), width_z));
  END GENERATE;
SGNED:  IF signd_a /= 0 GENERATE
    z <= std_logic_vector(fshl_stdar(  signed(a), unsigned(s), width_z));
  END GENERATE;
END beh;

--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Mon Sep 13 19:31:44 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_69_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_69_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_69_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_69_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_68_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_68_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_68_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_68_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_67_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_67_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_67_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_67_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_66_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_66_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_66_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_66_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_65_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_65_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_65_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_65_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_64_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_64_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_64_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_64_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_63_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_63_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_63_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_63_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_62_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_62_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_62_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_62_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_61_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_61_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_61_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_61_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_60_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_60_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_60_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_60_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_59_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_59_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_59_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_59_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_58_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_58_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_58_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_58_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_57_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_57_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_57_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_57_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_56_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_56_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_56_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_56_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_55_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_55_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_55_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_55_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_54_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_54_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_54_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_54_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_53_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_53_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_53_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_53_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_52_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_52_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_52_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_52_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_51_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_51_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_51_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_51_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_50_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_50_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_50_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_50_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_49_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_49_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_49_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_49_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_48_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_48_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_48_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_48_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_47_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_47_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_47_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_47_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_46_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_46_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_46_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_46_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_45_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_45_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_45_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_45_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_44_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_44_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_44_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_44_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_43_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_43_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_43_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_43_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_42_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_42_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_42_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_42_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_41_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_41_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_41_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_41_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_40_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_40_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_40_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_40_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_39_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_39_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_39_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_39_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_38_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_38_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_38_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_38_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_37_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_37_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_37_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_37_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(11 DOWNTO 6));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(5 DOWNTO 0));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_36_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_36_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_36_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_36_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(11 DOWNTO 6));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(5 DOWNTO 0));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_35_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_35_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_35_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_35_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(11 DOWNTO 6));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(5 DOWNTO 0));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_34_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_34_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_34_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_34_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(11 DOWNTO 6));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(5 DOWNTO 0));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_33_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_33_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_33_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_33_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(11 DOWNTO 6));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(5 DOWNTO 0));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_32_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_32_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_32_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_32_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(11 DOWNTO 6));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(5 DOWNTO 0));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_31_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_31_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_31_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_31_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(11 DOWNTO 6));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(5 DOWNTO 0));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_30_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_30_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_30_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_30_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(11 DOWNTO 6));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(5 DOWNTO 0));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_29_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_29_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_29_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_29_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(11 DOWNTO 6));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(5 DOWNTO 0));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_28_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_28_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_28_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_28_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(11 DOWNTO 6));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(5 DOWNTO 0));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_27_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_27_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_27_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_27_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(11 DOWNTO 6));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(5 DOWNTO 0));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_26_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_26_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_26_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_26_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(11 DOWNTO 6));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(5 DOWNTO 0));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_25_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_25_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_25_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_25_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(11 DOWNTO 6));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(5 DOWNTO 0));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_24_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_24_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_24_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_24_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(11 DOWNTO 6));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(5 DOWNTO 0));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_23_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_23_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_23_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_23_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(11 DOWNTO 6));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(5 DOWNTO 0));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_22_6_32_64_64_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_22_6_32_64_64_32_1_gen
    IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_22_6_32_64_64_32_1_gen;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_22_6_32_64_64_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(11 DOWNTO 6));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(5 DOWNTO 0));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    complete_rsci_wen_comp : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
    main_C_0_tr0 : IN STD_LOGIC;
    VEC_LOOP_C_11_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_4_tr0 : IN STD_LOGIC;
    STAGE_LOOP_C_1_tr0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_core_fsm;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for inPlaceNTT_DIF_precomp_core_core_fsm_1
  TYPE inPlaceNTT_DIF_precomp_core_core_fsm_1_ST IS (main_C_0, STAGE_LOOP_C_0, COMP_LOOP_C_0,
      COMP_LOOP_C_1, COMP_LOOP_C_2, COMP_LOOP_C_3, VEC_LOOP_C_0, VEC_LOOP_C_1, VEC_LOOP_C_2,
      VEC_LOOP_C_3, VEC_LOOP_C_4, VEC_LOOP_C_5, VEC_LOOP_C_6, VEC_LOOP_C_7, VEC_LOOP_C_8,
      VEC_LOOP_C_9, VEC_LOOP_C_10, VEC_LOOP_C_11, COMP_LOOP_C_4, STAGE_LOOP_C_1,
      main_C_1, main_C_2);

  SIGNAL state_var : inPlaceNTT_DIF_precomp_core_core_fsm_1_ST;
  SIGNAL state_var_NS : inPlaceNTT_DIF_precomp_core_core_fsm_1_ST;

BEGIN
  inPlaceNTT_DIF_precomp_core_core_fsm_1 : PROCESS (main_C_0_tr0, VEC_LOOP_C_11_tr0,
      COMP_LOOP_C_4_tr0, STAGE_LOOP_C_1_tr0, state_var)
  BEGIN
    CASE state_var IS
      WHEN STAGE_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000000000000010");
        state_var_NS <= COMP_LOOP_C_0;
      WHEN COMP_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000000000000100");
        state_var_NS <= COMP_LOOP_C_1;
      WHEN COMP_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000000000001000");
        state_var_NS <= COMP_LOOP_C_2;
      WHEN COMP_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000000000010000");
        state_var_NS <= COMP_LOOP_C_3;
      WHEN COMP_LOOP_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000000000100000");
        state_var_NS <= VEC_LOOP_C_0;
      WHEN VEC_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000000001000000");
        state_var_NS <= VEC_LOOP_C_1;
      WHEN VEC_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000000010000000");
        state_var_NS <= VEC_LOOP_C_2;
      WHEN VEC_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000000100000000");
        state_var_NS <= VEC_LOOP_C_3;
      WHEN VEC_LOOP_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000001000000000");
        state_var_NS <= VEC_LOOP_C_4;
      WHEN VEC_LOOP_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000010000000000");
        state_var_NS <= VEC_LOOP_C_5;
      WHEN VEC_LOOP_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000100000000000");
        state_var_NS <= VEC_LOOP_C_6;
      WHEN VEC_LOOP_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000001000000000000");
        state_var_NS <= VEC_LOOP_C_7;
      WHEN VEC_LOOP_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000010000000000000");
        state_var_NS <= VEC_LOOP_C_8;
      WHEN VEC_LOOP_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000100000000000000");
        state_var_NS <= VEC_LOOP_C_9;
      WHEN VEC_LOOP_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001000000000000000");
        state_var_NS <= VEC_LOOP_C_10;
      WHEN VEC_LOOP_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010000000000000000");
        state_var_NS <= VEC_LOOP_C_11;
      WHEN VEC_LOOP_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100000000000000000");
        IF ( VEC_LOOP_C_11_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_4;
        ELSE
          state_var_NS <= VEC_LOOP_C_0;
        END IF;
      WHEN COMP_LOOP_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000000000000000000");
        IF ( COMP_LOOP_C_4_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN STAGE_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000000000000000000");
        IF ( STAGE_LOOP_C_1_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSE
          state_var_NS <= STAGE_LOOP_C_0;
        END IF;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000000000000000000");
        state_var_NS <= main_C_2;
      WHEN main_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000000000000000000");
        state_var_NS <= main_C_0;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000000000000001");
        IF ( main_C_0_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSE
          state_var_NS <= STAGE_LOOP_C_0;
        END IF;
    END CASE;
  END PROCESS inPlaceNTT_DIF_precomp_core_core_fsm_1;

  inPlaceNTT_DIF_precomp_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        IF ( complete_rsci_wen_comp = '1' ) THEN
          state_var <= state_var_NS;
        END IF;
      END IF;
    END IF;
  END PROCESS inPlaceNTT_DIF_precomp_core_core_fsm_1_REG;

END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_staller
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_staller IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    core_wten : OUT STD_LOGIC;
    complete_rsci_wen_comp : IN STD_LOGIC;
    core_wten_pff : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_staller;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_staller IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL core_wten_reg : STD_LOGIC;

BEGIN
  core_wten <= core_wten_reg;
  core_wten_pff <= NOT complete_rsci_wen_comp;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        core_wten_reg <= '0';
      ELSE
        core_wten_reg <= NOT complete_rsci_wen_comp;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_0_obj_twiddle_h_rsc_triosy_0_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_0_obj_twiddle_h_rsc_triosy_0_0_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_0_obj_twiddle_h_rsc_triosy_0_0_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_0_obj_twiddle_h_rsc_triosy_0_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_0_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_0_obj_iswt0
      AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_1_obj_twiddle_h_rsc_triosy_0_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_1_obj_twiddle_h_rsc_triosy_0_1_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_1_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_1_obj_twiddle_h_rsc_triosy_0_1_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_1_obj_twiddle_h_rsc_triosy_0_1_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_1_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_1_obj_iswt0
      AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_2_obj_twiddle_h_rsc_triosy_0_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_2_obj_twiddle_h_rsc_triosy_0_2_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_2_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_2_obj_twiddle_h_rsc_triosy_0_2_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_2_obj_twiddle_h_rsc_triosy_0_2_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_2_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_2_obj_iswt0
      AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_3_obj_twiddle_h_rsc_triosy_0_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_3_obj_twiddle_h_rsc_triosy_0_3_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_3_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_3_obj_twiddle_h_rsc_triosy_0_3_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_3_obj_twiddle_h_rsc_triosy_0_3_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_3_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_3_obj_iswt0
      AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_4_obj_twiddle_h_rsc_triosy_0_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_4_obj_twiddle_h_rsc_triosy_0_4_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_4_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_4_obj_twiddle_h_rsc_triosy_0_4_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_4_obj_twiddle_h_rsc_triosy_0_4_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_4_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_4_obj_iswt0
      AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_5_obj_twiddle_h_rsc_triosy_0_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_5_obj_twiddle_h_rsc_triosy_0_5_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_5_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_5_obj_twiddle_h_rsc_triosy_0_5_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_5_obj_twiddle_h_rsc_triosy_0_5_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_5_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_5_obj_iswt0
      AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_6_obj_twiddle_h_rsc_triosy_0_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_6_obj_twiddle_h_rsc_triosy_0_6_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_6_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_6_obj_twiddle_h_rsc_triosy_0_6_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_6_obj_twiddle_h_rsc_triosy_0_6_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_6_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_6_obj_iswt0
      AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_7_obj_twiddle_h_rsc_triosy_0_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_7_obj_twiddle_h_rsc_triosy_0_7_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_7_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_7_obj_twiddle_h_rsc_triosy_0_7_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_7_obj_twiddle_h_rsc_triosy_0_7_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_7_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_7_obj_iswt0
      AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_0_obj_twiddle_h_rsc_triosy_1_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_0_obj_twiddle_h_rsc_triosy_1_0_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_0_obj_twiddle_h_rsc_triosy_1_0_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_0_obj_twiddle_h_rsc_triosy_1_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_1_0_obj_ld_core_sct <= twiddle_h_rsc_triosy_1_0_obj_iswt0
      AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_1_obj_twiddle_h_rsc_triosy_1_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_1_obj_twiddle_h_rsc_triosy_1_1_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_1_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_1_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_1_obj_twiddle_h_rsc_triosy_1_1_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_1_obj_twiddle_h_rsc_triosy_1_1_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_1_1_obj_ld_core_sct <= twiddle_h_rsc_triosy_1_1_obj_iswt0
      AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_2_obj_twiddle_h_rsc_triosy_1_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_2_obj_twiddle_h_rsc_triosy_1_2_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_2_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_2_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_2_obj_twiddle_h_rsc_triosy_1_2_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_2_obj_twiddle_h_rsc_triosy_1_2_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_1_2_obj_ld_core_sct <= twiddle_h_rsc_triosy_1_2_obj_iswt0
      AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_3_obj_twiddle_h_rsc_triosy_1_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_3_obj_twiddle_h_rsc_triosy_1_3_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_3_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_3_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_3_obj_twiddle_h_rsc_triosy_1_3_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_3_obj_twiddle_h_rsc_triosy_1_3_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_1_3_obj_ld_core_sct <= twiddle_h_rsc_triosy_1_3_obj_iswt0
      AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_4_obj_twiddle_h_rsc_triosy_1_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_4_obj_twiddle_h_rsc_triosy_1_4_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_4_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_4_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_4_obj_twiddle_h_rsc_triosy_1_4_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_4_obj_twiddle_h_rsc_triosy_1_4_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_1_4_obj_ld_core_sct <= twiddle_h_rsc_triosy_1_4_obj_iswt0
      AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_5_obj_twiddle_h_rsc_triosy_1_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_5_obj_twiddle_h_rsc_triosy_1_5_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_5_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_5_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_5_obj_twiddle_h_rsc_triosy_1_5_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_5_obj_twiddle_h_rsc_triosy_1_5_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_1_5_obj_ld_core_sct <= twiddle_h_rsc_triosy_1_5_obj_iswt0
      AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_6_obj_twiddle_h_rsc_triosy_1_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_6_obj_twiddle_h_rsc_triosy_1_6_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_6_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_6_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_6_obj_twiddle_h_rsc_triosy_1_6_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_6_obj_twiddle_h_rsc_triosy_1_6_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_1_6_obj_ld_core_sct <= twiddle_h_rsc_triosy_1_6_obj_iswt0
      AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_7_obj_twiddle_h_rsc_triosy_1_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_7_obj_twiddle_h_rsc_triosy_1_7_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_7_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_7_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_7_obj_twiddle_h_rsc_triosy_1_7_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_7_obj_twiddle_h_rsc_triosy_1_7_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_1_7_obj_ld_core_sct <= twiddle_h_rsc_triosy_1_7_obj_iswt0
      AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_0_obj_twiddle_rsc_triosy_0_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_0_obj_twiddle_rsc_triosy_0_0_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_0_obj_twiddle_rsc_triosy_0_0_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_0_obj_twiddle_rsc_triosy_0_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_0_obj_ld_core_sct <= twiddle_rsc_triosy_0_0_obj_iswt0 AND
      (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_1_obj_twiddle_rsc_triosy_0_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_1_obj_twiddle_rsc_triosy_0_1_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_1_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_1_obj_twiddle_rsc_triosy_0_1_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_1_obj_twiddle_rsc_triosy_0_1_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_1_obj_ld_core_sct <= twiddle_rsc_triosy_0_1_obj_iswt0 AND
      (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_2_obj_twiddle_rsc_triosy_0_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_2_obj_twiddle_rsc_triosy_0_2_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_2_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_2_obj_twiddle_rsc_triosy_0_2_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_2_obj_twiddle_rsc_triosy_0_2_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_2_obj_ld_core_sct <= twiddle_rsc_triosy_0_2_obj_iswt0 AND
      (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_3_obj_twiddle_rsc_triosy_0_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_3_obj_twiddle_rsc_triosy_0_3_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_3_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_3_obj_twiddle_rsc_triosy_0_3_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_3_obj_twiddle_rsc_triosy_0_3_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_3_obj_ld_core_sct <= twiddle_rsc_triosy_0_3_obj_iswt0 AND
      (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_4_obj_twiddle_rsc_triosy_0_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_4_obj_twiddle_rsc_triosy_0_4_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_4_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_4_obj_twiddle_rsc_triosy_0_4_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_4_obj_twiddle_rsc_triosy_0_4_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_4_obj_ld_core_sct <= twiddle_rsc_triosy_0_4_obj_iswt0 AND
      (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_5_obj_twiddle_rsc_triosy_0_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_5_obj_twiddle_rsc_triosy_0_5_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_5_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_5_obj_twiddle_rsc_triosy_0_5_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_5_obj_twiddle_rsc_triosy_0_5_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_5_obj_ld_core_sct <= twiddle_rsc_triosy_0_5_obj_iswt0 AND
      (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_6_obj_twiddle_rsc_triosy_0_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_6_obj_twiddle_rsc_triosy_0_6_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_6_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_6_obj_twiddle_rsc_triosy_0_6_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_6_obj_twiddle_rsc_triosy_0_6_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_6_obj_ld_core_sct <= twiddle_rsc_triosy_0_6_obj_iswt0 AND
      (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_7_obj_twiddle_rsc_triosy_0_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_7_obj_twiddle_rsc_triosy_0_7_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_7_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_7_obj_twiddle_rsc_triosy_0_7_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_7_obj_twiddle_rsc_triosy_0_7_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_7_obj_ld_core_sct <= twiddle_rsc_triosy_0_7_obj_iswt0 AND
      (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_0_obj_twiddle_rsc_triosy_1_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_0_obj_twiddle_rsc_triosy_1_0_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_1_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_0_obj_twiddle_rsc_triosy_1_0_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_0_obj_twiddle_rsc_triosy_1_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_1_0_obj_ld_core_sct <= twiddle_rsc_triosy_1_0_obj_iswt0 AND
      (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_1_obj_twiddle_rsc_triosy_1_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_1_obj_twiddle_rsc_triosy_1_1_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_1_1_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_1_1_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_1_obj_twiddle_rsc_triosy_1_1_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_1_obj_twiddle_rsc_triosy_1_1_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_1_1_obj_ld_core_sct <= twiddle_rsc_triosy_1_1_obj_iswt0 AND
      (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_2_obj_twiddle_rsc_triosy_1_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_2_obj_twiddle_rsc_triosy_1_2_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_1_2_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_1_2_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_2_obj_twiddle_rsc_triosy_1_2_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_2_obj_twiddle_rsc_triosy_1_2_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_1_2_obj_ld_core_sct <= twiddle_rsc_triosy_1_2_obj_iswt0 AND
      (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_3_obj_twiddle_rsc_triosy_1_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_3_obj_twiddle_rsc_triosy_1_3_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_1_3_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_1_3_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_3_obj_twiddle_rsc_triosy_1_3_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_3_obj_twiddle_rsc_triosy_1_3_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_1_3_obj_ld_core_sct <= twiddle_rsc_triosy_1_3_obj_iswt0 AND
      (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_4_obj_twiddle_rsc_triosy_1_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_4_obj_twiddle_rsc_triosy_1_4_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_1_4_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_1_4_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_4_obj_twiddle_rsc_triosy_1_4_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_4_obj_twiddle_rsc_triosy_1_4_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_1_4_obj_ld_core_sct <= twiddle_rsc_triosy_1_4_obj_iswt0 AND
      (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_5_obj_twiddle_rsc_triosy_1_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_5_obj_twiddle_rsc_triosy_1_5_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_1_5_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_1_5_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_5_obj_twiddle_rsc_triosy_1_5_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_5_obj_twiddle_rsc_triosy_1_5_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_1_5_obj_ld_core_sct <= twiddle_rsc_triosy_1_5_obj_iswt0 AND
      (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_6_obj_twiddle_rsc_triosy_1_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_6_obj_twiddle_rsc_triosy_1_6_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_1_6_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_1_6_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_6_obj_twiddle_rsc_triosy_1_6_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_6_obj_twiddle_rsc_triosy_1_6_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_1_6_obj_ld_core_sct <= twiddle_rsc_triosy_1_6_obj_iswt0 AND
      (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_7_obj_twiddle_rsc_triosy_1_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_7_obj_twiddle_rsc_triosy_1_7_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_1_7_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_1_7_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_7_obj_twiddle_rsc_triosy_1_7_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_7_obj_twiddle_rsc_triosy_1_7_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_1_7_obj_ld_core_sct <= twiddle_rsc_triosy_1_7_obj_iswt0 AND
      (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_r_rsc_triosy_obj_r_rsc_triosy_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_r_rsc_triosy_obj_r_rsc_triosy_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    r_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
    r_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_r_rsc_triosy_obj_r_rsc_triosy_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_r_rsc_triosy_obj_r_rsc_triosy_wait_ctrl
    IS
  -- Default Constants

BEGIN
  r_rsc_triosy_obj_ld_core_sct <= r_rsc_triosy_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_p_rsc_triosy_obj_p_rsc_triosy_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_p_rsc_triosy_obj_p_rsc_triosy_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    p_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
    p_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_p_rsc_triosy_obj_p_rsc_triosy_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_p_rsc_triosy_obj_p_rsc_triosy_wait_ctrl
    IS
  -- Default Constants

BEGIN
  p_rsc_triosy_obj_ld_core_sct <= p_rsc_triosy_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_0_obj_vec_rsc_triosy_0_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_0_obj_vec_rsc_triosy_0_0_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC;
    vec_rsc_triosy_0_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_0_obj_vec_rsc_triosy_0_0_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_0_obj_vec_rsc_triosy_0_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  vec_rsc_triosy_0_0_obj_ld_core_sct <= vec_rsc_triosy_0_0_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_1_obj_vec_rsc_triosy_0_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_1_obj_vec_rsc_triosy_0_1_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC;
    vec_rsc_triosy_0_1_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_1_obj_vec_rsc_triosy_0_1_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_1_obj_vec_rsc_triosy_0_1_wait_ctrl
    IS
  -- Default Constants

BEGIN
  vec_rsc_triosy_0_1_obj_ld_core_sct <= vec_rsc_triosy_0_1_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_2_obj_vec_rsc_triosy_0_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_2_obj_vec_rsc_triosy_0_2_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC;
    vec_rsc_triosy_0_2_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_2_obj_vec_rsc_triosy_0_2_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_2_obj_vec_rsc_triosy_0_2_wait_ctrl
    IS
  -- Default Constants

BEGIN
  vec_rsc_triosy_0_2_obj_ld_core_sct <= vec_rsc_triosy_0_2_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_3_obj_vec_rsc_triosy_0_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_3_obj_vec_rsc_triosy_0_3_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC;
    vec_rsc_triosy_0_3_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_3_obj_vec_rsc_triosy_0_3_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_3_obj_vec_rsc_triosy_0_3_wait_ctrl
    IS
  -- Default Constants

BEGIN
  vec_rsc_triosy_0_3_obj_ld_core_sct <= vec_rsc_triosy_0_3_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_4_obj_vec_rsc_triosy_0_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_4_obj_vec_rsc_triosy_0_4_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC;
    vec_rsc_triosy_0_4_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_4_obj_vec_rsc_triosy_0_4_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_4_obj_vec_rsc_triosy_0_4_wait_ctrl
    IS
  -- Default Constants

BEGIN
  vec_rsc_triosy_0_4_obj_ld_core_sct <= vec_rsc_triosy_0_4_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_5_obj_vec_rsc_triosy_0_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_5_obj_vec_rsc_triosy_0_5_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC;
    vec_rsc_triosy_0_5_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_5_obj_vec_rsc_triosy_0_5_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_5_obj_vec_rsc_triosy_0_5_wait_ctrl
    IS
  -- Default Constants

BEGIN
  vec_rsc_triosy_0_5_obj_ld_core_sct <= vec_rsc_triosy_0_5_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_6_obj_vec_rsc_triosy_0_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_6_obj_vec_rsc_triosy_0_6_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC;
    vec_rsc_triosy_0_6_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_6_obj_vec_rsc_triosy_0_6_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_6_obj_vec_rsc_triosy_0_6_wait_ctrl
    IS
  -- Default Constants

BEGIN
  vec_rsc_triosy_0_6_obj_ld_core_sct <= vec_rsc_triosy_0_6_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_7_obj_vec_rsc_triosy_0_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_7_obj_vec_rsc_triosy_0_7_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC;
    vec_rsc_triosy_0_7_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_7_obj_vec_rsc_triosy_0_7_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_7_obj_vec_rsc_triosy_0_7_wait_ctrl
    IS
  -- Default Constants

BEGIN
  vec_rsc_triosy_0_7_obj_ld_core_sct <= vec_rsc_triosy_0_7_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_0_obj_vec_rsc_triosy_1_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_0_obj_vec_rsc_triosy_1_0_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC;
    vec_rsc_triosy_1_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_0_obj_vec_rsc_triosy_1_0_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_0_obj_vec_rsc_triosy_1_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  vec_rsc_triosy_1_0_obj_ld_core_sct <= vec_rsc_triosy_1_0_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_1_obj_vec_rsc_triosy_1_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_1_obj_vec_rsc_triosy_1_1_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_1_1_obj_iswt0 : IN STD_LOGIC;
    vec_rsc_triosy_1_1_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_1_obj_vec_rsc_triosy_1_1_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_1_obj_vec_rsc_triosy_1_1_wait_ctrl
    IS
  -- Default Constants

BEGIN
  vec_rsc_triosy_1_1_obj_ld_core_sct <= vec_rsc_triosy_1_1_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_2_obj_vec_rsc_triosy_1_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_2_obj_vec_rsc_triosy_1_2_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_1_2_obj_iswt0 : IN STD_LOGIC;
    vec_rsc_triosy_1_2_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_2_obj_vec_rsc_triosy_1_2_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_2_obj_vec_rsc_triosy_1_2_wait_ctrl
    IS
  -- Default Constants

BEGIN
  vec_rsc_triosy_1_2_obj_ld_core_sct <= vec_rsc_triosy_1_2_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_3_obj_vec_rsc_triosy_1_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_3_obj_vec_rsc_triosy_1_3_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_1_3_obj_iswt0 : IN STD_LOGIC;
    vec_rsc_triosy_1_3_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_3_obj_vec_rsc_triosy_1_3_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_3_obj_vec_rsc_triosy_1_3_wait_ctrl
    IS
  -- Default Constants

BEGIN
  vec_rsc_triosy_1_3_obj_ld_core_sct <= vec_rsc_triosy_1_3_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_4_obj_vec_rsc_triosy_1_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_4_obj_vec_rsc_triosy_1_4_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_1_4_obj_iswt0 : IN STD_LOGIC;
    vec_rsc_triosy_1_4_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_4_obj_vec_rsc_triosy_1_4_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_4_obj_vec_rsc_triosy_1_4_wait_ctrl
    IS
  -- Default Constants

BEGIN
  vec_rsc_triosy_1_4_obj_ld_core_sct <= vec_rsc_triosy_1_4_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_5_obj_vec_rsc_triosy_1_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_5_obj_vec_rsc_triosy_1_5_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_1_5_obj_iswt0 : IN STD_LOGIC;
    vec_rsc_triosy_1_5_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_5_obj_vec_rsc_triosy_1_5_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_5_obj_vec_rsc_triosy_1_5_wait_ctrl
    IS
  -- Default Constants

BEGIN
  vec_rsc_triosy_1_5_obj_ld_core_sct <= vec_rsc_triosy_1_5_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_6_obj_vec_rsc_triosy_1_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_6_obj_vec_rsc_triosy_1_6_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_1_6_obj_iswt0 : IN STD_LOGIC;
    vec_rsc_triosy_1_6_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_6_obj_vec_rsc_triosy_1_6_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_6_obj_vec_rsc_triosy_1_6_wait_ctrl
    IS
  -- Default Constants

BEGIN
  vec_rsc_triosy_1_6_obj_ld_core_sct <= vec_rsc_triosy_1_6_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_7_obj_vec_rsc_triosy_1_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_7_obj_vec_rsc_triosy_1_7_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_1_7_obj_iswt0 : IN STD_LOGIC;
    vec_rsc_triosy_1_7_obj_ld_core_sct : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_7_obj_vec_rsc_triosy_1_7_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_7_obj_vec_rsc_triosy_1_7_wait_ctrl
    IS
  -- Default Constants

BEGIN
  vec_rsc_triosy_1_7_obj_ld_core_sct <= vec_rsc_triosy_1_7_obj_iswt0 AND (NOT core_wten);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_dp
    IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_1_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_7_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_7_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_1_7_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_1_7_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_7_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsc_1_7_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_1_7_i_qb_d, twiddle_h_rsc_1_7_i_qb_d_bfwt,
      twiddle_h_rsc_1_7_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_1_7_i_bcwt <= '0';
      ELSE
        twiddle_h_rsc_1_7_i_bcwt <= NOT((NOT(twiddle_h_rsc_1_7_i_bcwt OR twiddle_h_rsc_1_7_i_biwt))
            OR twiddle_h_rsc_1_7_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_1_7_i_biwt = '1' ) THEN
        twiddle_h_rsc_1_7_i_qb_d_bfwt <= twiddle_h_rsc_1_7_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_1_7_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_1_7_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_1_7_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_1_7_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_1_7_i_bdwt <= twiddle_h_rsc_1_7_i_oswt AND core_wen;
  twiddle_h_rsc_1_7_i_biwt <= (NOT core_wten) AND twiddle_h_rsc_1_7_i_oswt;
  twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_h_rsc_1_7_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_dp
    IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_1_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_6_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_6_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_1_6_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_1_6_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_6_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsc_1_6_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_1_6_i_qb_d, twiddle_h_rsc_1_6_i_qb_d_bfwt,
      twiddle_h_rsc_1_6_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_1_6_i_bcwt <= '0';
      ELSE
        twiddle_h_rsc_1_6_i_bcwt <= NOT((NOT(twiddle_h_rsc_1_6_i_bcwt OR twiddle_h_rsc_1_6_i_biwt))
            OR twiddle_h_rsc_1_6_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_1_6_i_biwt = '1' ) THEN
        twiddle_h_rsc_1_6_i_qb_d_bfwt <= twiddle_h_rsc_1_6_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_1_6_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_1_6_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_1_6_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_1_6_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_1_6_i_bdwt <= twiddle_h_rsc_1_6_i_oswt AND core_wen;
  twiddle_h_rsc_1_6_i_biwt <= (NOT core_wten) AND twiddle_h_rsc_1_6_i_oswt;
  twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_h_rsc_1_6_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_dp
    IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_1_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_5_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_5_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_1_5_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_1_5_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_5_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsc_1_5_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_1_5_i_qb_d, twiddle_h_rsc_1_5_i_qb_d_bfwt,
      twiddle_h_rsc_1_5_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_1_5_i_bcwt <= '0';
      ELSE
        twiddle_h_rsc_1_5_i_bcwt <= NOT((NOT(twiddle_h_rsc_1_5_i_bcwt OR twiddle_h_rsc_1_5_i_biwt))
            OR twiddle_h_rsc_1_5_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_1_5_i_biwt = '1' ) THEN
        twiddle_h_rsc_1_5_i_qb_d_bfwt <= twiddle_h_rsc_1_5_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_1_5_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_1_5_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_1_5_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_1_5_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_1_5_i_bdwt <= twiddle_h_rsc_1_5_i_oswt AND core_wen;
  twiddle_h_rsc_1_5_i_biwt <= (NOT core_wten) AND twiddle_h_rsc_1_5_i_oswt;
  twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_h_rsc_1_5_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_dp
    IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_1_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_4_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_4_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_1_4_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_1_4_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_4_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsc_1_4_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_1_4_i_qb_d, twiddle_h_rsc_1_4_i_qb_d_bfwt,
      twiddle_h_rsc_1_4_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_1_4_i_bcwt <= '0';
      ELSE
        twiddle_h_rsc_1_4_i_bcwt <= NOT((NOT(twiddle_h_rsc_1_4_i_bcwt OR twiddle_h_rsc_1_4_i_biwt))
            OR twiddle_h_rsc_1_4_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_1_4_i_biwt = '1' ) THEN
        twiddle_h_rsc_1_4_i_qb_d_bfwt <= twiddle_h_rsc_1_4_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_1_4_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_1_4_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_1_4_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_1_4_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_1_4_i_bdwt <= twiddle_h_rsc_1_4_i_oswt AND core_wen;
  twiddle_h_rsc_1_4_i_biwt <= (NOT core_wten) AND twiddle_h_rsc_1_4_i_oswt;
  twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_h_rsc_1_4_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_dp
    IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_1_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_3_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_3_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_1_3_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_1_3_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_3_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsc_1_3_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_1_3_i_qb_d, twiddle_h_rsc_1_3_i_qb_d_bfwt,
      twiddle_h_rsc_1_3_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_1_3_i_bcwt <= '0';
      ELSE
        twiddle_h_rsc_1_3_i_bcwt <= NOT((NOT(twiddle_h_rsc_1_3_i_bcwt OR twiddle_h_rsc_1_3_i_biwt))
            OR twiddle_h_rsc_1_3_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_1_3_i_biwt = '1' ) THEN
        twiddle_h_rsc_1_3_i_qb_d_bfwt <= twiddle_h_rsc_1_3_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_1_3_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_1_3_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_1_3_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_1_3_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_1_3_i_bdwt <= twiddle_h_rsc_1_3_i_oswt AND core_wen;
  twiddle_h_rsc_1_3_i_biwt <= (NOT core_wten) AND twiddle_h_rsc_1_3_i_oswt;
  twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_h_rsc_1_3_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_dp
    IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_1_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_2_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_2_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_1_2_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_1_2_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_2_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsc_1_2_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_1_2_i_qb_d, twiddle_h_rsc_1_2_i_qb_d_bfwt,
      twiddle_h_rsc_1_2_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_1_2_i_bcwt <= '0';
      ELSE
        twiddle_h_rsc_1_2_i_bcwt <= NOT((NOT(twiddle_h_rsc_1_2_i_bcwt OR twiddle_h_rsc_1_2_i_biwt))
            OR twiddle_h_rsc_1_2_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_1_2_i_biwt = '1' ) THEN
        twiddle_h_rsc_1_2_i_qb_d_bfwt <= twiddle_h_rsc_1_2_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_1_2_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_1_2_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_1_2_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_1_2_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_1_2_i_bdwt <= twiddle_h_rsc_1_2_i_oswt AND core_wen;
  twiddle_h_rsc_1_2_i_biwt <= (NOT core_wten) AND twiddle_h_rsc_1_2_i_oswt;
  twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_h_rsc_1_2_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_dp
    IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_1_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_1_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_1_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_1_1_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_1_1_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_1_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsc_1_1_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_1_1_i_qb_d, twiddle_h_rsc_1_1_i_qb_d_bfwt,
      twiddle_h_rsc_1_1_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_1_1_i_bcwt <= '0';
      ELSE
        twiddle_h_rsc_1_1_i_bcwt <= NOT((NOT(twiddle_h_rsc_1_1_i_bcwt OR twiddle_h_rsc_1_1_i_biwt))
            OR twiddle_h_rsc_1_1_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_1_1_i_biwt = '1' ) THEN
        twiddle_h_rsc_1_1_i_qb_d_bfwt <= twiddle_h_rsc_1_1_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_1_1_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_1_1_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_1_1_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_1_1_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_1_1_i_bdwt <= twiddle_h_rsc_1_1_i_oswt AND core_wen;
  twiddle_h_rsc_1_1_i_biwt <= (NOT core_wten) AND twiddle_h_rsc_1_1_i_oswt;
  twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_h_rsc_1_1_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_dp
    IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_1_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_0_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_0_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_1_0_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_1_0_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_0_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsc_1_0_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_1_0_i_qb_d, twiddle_h_rsc_1_0_i_qb_d_bfwt,
      twiddle_h_rsc_1_0_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_1_0_i_bcwt <= '0';
      ELSE
        twiddle_h_rsc_1_0_i_bcwt <= NOT((NOT(twiddle_h_rsc_1_0_i_bcwt OR twiddle_h_rsc_1_0_i_biwt))
            OR twiddle_h_rsc_1_0_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_1_0_i_biwt = '1' ) THEN
        twiddle_h_rsc_1_0_i_qb_d_bfwt <= twiddle_h_rsc_1_0_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_1_0_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_1_0_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_1_0_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_1_0_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_1_0_i_bdwt <= twiddle_h_rsc_1_0_i_oswt AND core_wen;
  twiddle_h_rsc_1_0_i_biwt <= (NOT core_wten) AND twiddle_h_rsc_1_0_i_oswt;
  twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_h_rsc_1_0_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_dp
    IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_7_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_7_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsc_0_7_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_7_i_qb_d, twiddle_h_rsc_0_7_i_qb_d_bfwt,
      twiddle_h_rsc_0_7_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_7_i_bcwt <= '0';
      ELSE
        twiddle_h_rsc_0_7_i_bcwt <= NOT((NOT(twiddle_h_rsc_0_7_i_bcwt OR twiddle_h_rsc_0_7_i_biwt))
            OR twiddle_h_rsc_0_7_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_7_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_7_i_qb_d_bfwt <= twiddle_h_rsc_0_7_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_0_7_i_bdwt <= twiddle_h_rsc_0_7_i_oswt AND core_wen;
  twiddle_h_rsc_0_7_i_biwt <= (NOT core_wten) AND twiddle_h_rsc_0_7_i_oswt;
  twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_h_rsc_0_7_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_dp
    IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_6_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_6_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsc_0_6_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_6_i_qb_d, twiddle_h_rsc_0_6_i_qb_d_bfwt,
      twiddle_h_rsc_0_6_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_6_i_bcwt <= '0';
      ELSE
        twiddle_h_rsc_0_6_i_bcwt <= NOT((NOT(twiddle_h_rsc_0_6_i_bcwt OR twiddle_h_rsc_0_6_i_biwt))
            OR twiddle_h_rsc_0_6_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_6_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_6_i_qb_d_bfwt <= twiddle_h_rsc_0_6_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_0_6_i_bdwt <= twiddle_h_rsc_0_6_i_oswt AND core_wen;
  twiddle_h_rsc_0_6_i_biwt <= (NOT core_wten) AND twiddle_h_rsc_0_6_i_oswt;
  twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_h_rsc_0_6_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_dp
    IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_5_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_5_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsc_0_5_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_5_i_qb_d, twiddle_h_rsc_0_5_i_qb_d_bfwt,
      twiddle_h_rsc_0_5_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_5_i_bcwt <= '0';
      ELSE
        twiddle_h_rsc_0_5_i_bcwt <= NOT((NOT(twiddle_h_rsc_0_5_i_bcwt OR twiddle_h_rsc_0_5_i_biwt))
            OR twiddle_h_rsc_0_5_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_5_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_5_i_qb_d_bfwt <= twiddle_h_rsc_0_5_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_0_5_i_bdwt <= twiddle_h_rsc_0_5_i_oswt AND core_wen;
  twiddle_h_rsc_0_5_i_biwt <= (NOT core_wten) AND twiddle_h_rsc_0_5_i_oswt;
  twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_h_rsc_0_5_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_dp
    IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_4_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_4_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsc_0_4_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_4_i_qb_d, twiddle_h_rsc_0_4_i_qb_d_bfwt,
      twiddle_h_rsc_0_4_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_4_i_bcwt <= '0';
      ELSE
        twiddle_h_rsc_0_4_i_bcwt <= NOT((NOT(twiddle_h_rsc_0_4_i_bcwt OR twiddle_h_rsc_0_4_i_biwt))
            OR twiddle_h_rsc_0_4_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_4_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_4_i_qb_d_bfwt <= twiddle_h_rsc_0_4_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_0_4_i_bdwt <= twiddle_h_rsc_0_4_i_oswt AND core_wen;
  twiddle_h_rsc_0_4_i_biwt <= (NOT core_wten) AND twiddle_h_rsc_0_4_i_oswt;
  twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_h_rsc_0_4_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_dp
    IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_3_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_3_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsc_0_3_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_3_i_qb_d, twiddle_h_rsc_0_3_i_qb_d_bfwt,
      twiddle_h_rsc_0_3_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_3_i_bcwt <= '0';
      ELSE
        twiddle_h_rsc_0_3_i_bcwt <= NOT((NOT(twiddle_h_rsc_0_3_i_bcwt OR twiddle_h_rsc_0_3_i_biwt))
            OR twiddle_h_rsc_0_3_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_3_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_3_i_qb_d_bfwt <= twiddle_h_rsc_0_3_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_0_3_i_bdwt <= twiddle_h_rsc_0_3_i_oswt AND core_wen;
  twiddle_h_rsc_0_3_i_biwt <= (NOT core_wten) AND twiddle_h_rsc_0_3_i_oswt;
  twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_h_rsc_0_3_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_dp
    IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_2_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_2_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsc_0_2_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_2_i_qb_d, twiddle_h_rsc_0_2_i_qb_d_bfwt,
      twiddle_h_rsc_0_2_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_2_i_bcwt <= '0';
      ELSE
        twiddle_h_rsc_0_2_i_bcwt <= NOT((NOT(twiddle_h_rsc_0_2_i_bcwt OR twiddle_h_rsc_0_2_i_biwt))
            OR twiddle_h_rsc_0_2_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_2_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_2_i_qb_d_bfwt <= twiddle_h_rsc_0_2_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_0_2_i_bdwt <= twiddle_h_rsc_0_2_i_oswt AND core_wen;
  twiddle_h_rsc_0_2_i_biwt <= (NOT core_wten) AND twiddle_h_rsc_0_2_i_oswt;
  twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_h_rsc_0_2_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_dp
    IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_1_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_1_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsc_0_1_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_1_i_qb_d, twiddle_h_rsc_0_1_i_qb_d_bfwt,
      twiddle_h_rsc_0_1_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_1_i_bcwt <= '0';
      ELSE
        twiddle_h_rsc_0_1_i_bcwt <= NOT((NOT(twiddle_h_rsc_0_1_i_bcwt OR twiddle_h_rsc_0_1_i_biwt))
            OR twiddle_h_rsc_0_1_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_1_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_1_i_qb_d_bfwt <= twiddle_h_rsc_0_1_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_0_1_i_bdwt <= twiddle_h_rsc_0_1_i_oswt AND core_wen;
  twiddle_h_rsc_0_1_i_biwt <= (NOT core_wten) AND twiddle_h_rsc_0_1_i_oswt;
  twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_h_rsc_0_1_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_dp
    IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_0_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_0_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsc_0_0_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_0_i_qb_d, twiddle_h_rsc_0_0_i_qb_d_bfwt,
      twiddle_h_rsc_0_0_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_0_i_bcwt <= '0';
      ELSE
        twiddle_h_rsc_0_0_i_bcwt <= NOT((NOT(twiddle_h_rsc_0_0_i_bcwt OR twiddle_h_rsc_0_0_i_biwt))
            OR twiddle_h_rsc_0_0_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_0_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_0_i_qb_d_bfwt <= twiddle_h_rsc_0_0_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_0_0_i_bdwt <= twiddle_h_rsc_0_0_i_oswt AND core_wen;
  twiddle_h_rsc_0_0_i_biwt <= (NOT core_wten) AND twiddle_h_rsc_0_0_i_oswt;
  twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_h_rsc_0_0_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_1_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_7_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_7_i_biwt : IN STD_LOGIC;
    twiddle_rsc_1_7_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_1_7_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_7_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsc_1_7_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsc_1_7_i_qb_d, twiddle_rsc_1_7_i_qb_d_bfwt,
      twiddle_rsc_1_7_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_1_7_i_bcwt <= '0';
      ELSE
        twiddle_rsc_1_7_i_bcwt <= NOT((NOT(twiddle_rsc_1_7_i_bcwt OR twiddle_rsc_1_7_i_biwt))
            OR twiddle_rsc_1_7_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_1_7_i_biwt = '1' ) THEN
        twiddle_rsc_1_7_i_qb_d_bfwt <= twiddle_rsc_1_7_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_1_7_i_oswt : IN STD_LOGIC;
    twiddle_rsc_1_7_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_1_7_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_rsc_1_7_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_1_7_i_bdwt <= twiddle_rsc_1_7_i_oswt AND core_wen;
  twiddle_rsc_1_7_i_biwt <= (NOT core_wten) AND twiddle_rsc_1_7_i_oswt;
  twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_rsc_1_7_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_1_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_6_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_6_i_biwt : IN STD_LOGIC;
    twiddle_rsc_1_6_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_1_6_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_6_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsc_1_6_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsc_1_6_i_qb_d, twiddle_rsc_1_6_i_qb_d_bfwt,
      twiddle_rsc_1_6_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_1_6_i_bcwt <= '0';
      ELSE
        twiddle_rsc_1_6_i_bcwt <= NOT((NOT(twiddle_rsc_1_6_i_bcwt OR twiddle_rsc_1_6_i_biwt))
            OR twiddle_rsc_1_6_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_1_6_i_biwt = '1' ) THEN
        twiddle_rsc_1_6_i_qb_d_bfwt <= twiddle_rsc_1_6_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_1_6_i_oswt : IN STD_LOGIC;
    twiddle_rsc_1_6_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_1_6_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_rsc_1_6_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_1_6_i_bdwt <= twiddle_rsc_1_6_i_oswt AND core_wen;
  twiddle_rsc_1_6_i_biwt <= (NOT core_wten) AND twiddle_rsc_1_6_i_oswt;
  twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_rsc_1_6_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_1_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_5_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_5_i_biwt : IN STD_LOGIC;
    twiddle_rsc_1_5_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_1_5_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_5_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsc_1_5_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsc_1_5_i_qb_d, twiddle_rsc_1_5_i_qb_d_bfwt,
      twiddle_rsc_1_5_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_1_5_i_bcwt <= '0';
      ELSE
        twiddle_rsc_1_5_i_bcwt <= NOT((NOT(twiddle_rsc_1_5_i_bcwt OR twiddle_rsc_1_5_i_biwt))
            OR twiddle_rsc_1_5_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_1_5_i_biwt = '1' ) THEN
        twiddle_rsc_1_5_i_qb_d_bfwt <= twiddle_rsc_1_5_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_1_5_i_oswt : IN STD_LOGIC;
    twiddle_rsc_1_5_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_1_5_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_rsc_1_5_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_1_5_i_bdwt <= twiddle_rsc_1_5_i_oswt AND core_wen;
  twiddle_rsc_1_5_i_biwt <= (NOT core_wten) AND twiddle_rsc_1_5_i_oswt;
  twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_rsc_1_5_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_1_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_4_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_4_i_biwt : IN STD_LOGIC;
    twiddle_rsc_1_4_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_1_4_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_4_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsc_1_4_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsc_1_4_i_qb_d, twiddle_rsc_1_4_i_qb_d_bfwt,
      twiddle_rsc_1_4_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_1_4_i_bcwt <= '0';
      ELSE
        twiddle_rsc_1_4_i_bcwt <= NOT((NOT(twiddle_rsc_1_4_i_bcwt OR twiddle_rsc_1_4_i_biwt))
            OR twiddle_rsc_1_4_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_1_4_i_biwt = '1' ) THEN
        twiddle_rsc_1_4_i_qb_d_bfwt <= twiddle_rsc_1_4_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_1_4_i_oswt : IN STD_LOGIC;
    twiddle_rsc_1_4_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_1_4_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_rsc_1_4_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_1_4_i_bdwt <= twiddle_rsc_1_4_i_oswt AND core_wen;
  twiddle_rsc_1_4_i_biwt <= (NOT core_wten) AND twiddle_rsc_1_4_i_oswt;
  twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_rsc_1_4_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_1_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_3_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_3_i_biwt : IN STD_LOGIC;
    twiddle_rsc_1_3_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_1_3_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_3_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsc_1_3_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsc_1_3_i_qb_d, twiddle_rsc_1_3_i_qb_d_bfwt,
      twiddle_rsc_1_3_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_1_3_i_bcwt <= '0';
      ELSE
        twiddle_rsc_1_3_i_bcwt <= NOT((NOT(twiddle_rsc_1_3_i_bcwt OR twiddle_rsc_1_3_i_biwt))
            OR twiddle_rsc_1_3_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_1_3_i_biwt = '1' ) THEN
        twiddle_rsc_1_3_i_qb_d_bfwt <= twiddle_rsc_1_3_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_1_3_i_oswt : IN STD_LOGIC;
    twiddle_rsc_1_3_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_1_3_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_rsc_1_3_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_1_3_i_bdwt <= twiddle_rsc_1_3_i_oswt AND core_wen;
  twiddle_rsc_1_3_i_biwt <= (NOT core_wten) AND twiddle_rsc_1_3_i_oswt;
  twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_rsc_1_3_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_1_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_2_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_2_i_biwt : IN STD_LOGIC;
    twiddle_rsc_1_2_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_1_2_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_2_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsc_1_2_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsc_1_2_i_qb_d, twiddle_rsc_1_2_i_qb_d_bfwt,
      twiddle_rsc_1_2_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_1_2_i_bcwt <= '0';
      ELSE
        twiddle_rsc_1_2_i_bcwt <= NOT((NOT(twiddle_rsc_1_2_i_bcwt OR twiddle_rsc_1_2_i_biwt))
            OR twiddle_rsc_1_2_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_1_2_i_biwt = '1' ) THEN
        twiddle_rsc_1_2_i_qb_d_bfwt <= twiddle_rsc_1_2_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_1_2_i_oswt : IN STD_LOGIC;
    twiddle_rsc_1_2_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_1_2_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_rsc_1_2_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_1_2_i_bdwt <= twiddle_rsc_1_2_i_oswt AND core_wen;
  twiddle_rsc_1_2_i_biwt <= (NOT core_wten) AND twiddle_rsc_1_2_i_oswt;
  twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_rsc_1_2_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_1_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_1_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_1_i_biwt : IN STD_LOGIC;
    twiddle_rsc_1_1_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_1_1_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_1_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsc_1_1_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsc_1_1_i_qb_d, twiddle_rsc_1_1_i_qb_d_bfwt,
      twiddle_rsc_1_1_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_1_1_i_bcwt <= '0';
      ELSE
        twiddle_rsc_1_1_i_bcwt <= NOT((NOT(twiddle_rsc_1_1_i_bcwt OR twiddle_rsc_1_1_i_biwt))
            OR twiddle_rsc_1_1_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_1_1_i_biwt = '1' ) THEN
        twiddle_rsc_1_1_i_qb_d_bfwt <= twiddle_rsc_1_1_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_1_1_i_oswt : IN STD_LOGIC;
    twiddle_rsc_1_1_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_1_1_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_rsc_1_1_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_1_1_i_bdwt <= twiddle_rsc_1_1_i_oswt AND core_wen;
  twiddle_rsc_1_1_i_biwt <= (NOT core_wten) AND twiddle_rsc_1_1_i_oswt;
  twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_rsc_1_1_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_1_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_0_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_0_i_biwt : IN STD_LOGIC;
    twiddle_rsc_1_0_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_1_0_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_0_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsc_1_0_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsc_1_0_i_qb_d, twiddle_rsc_1_0_i_qb_d_bfwt,
      twiddle_rsc_1_0_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_1_0_i_bcwt <= '0';
      ELSE
        twiddle_rsc_1_0_i_bcwt <= NOT((NOT(twiddle_rsc_1_0_i_bcwt OR twiddle_rsc_1_0_i_biwt))
            OR twiddle_rsc_1_0_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_1_0_i_biwt = '1' ) THEN
        twiddle_rsc_1_0_i_qb_d_bfwt <= twiddle_rsc_1_0_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_1_0_i_oswt : IN STD_LOGIC;
    twiddle_rsc_1_0_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_1_0_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_rsc_1_0_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_1_0_i_bdwt <= twiddle_rsc_1_0_i_oswt AND core_wen;
  twiddle_rsc_1_0_i_biwt <= (NOT core_wten) AND twiddle_rsc_1_0_i_oswt;
  twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_rsc_1_0_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_7_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_7_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_7_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsc_0_7_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_7_i_qb_d, twiddle_rsc_0_7_i_qb_d_bfwt,
      twiddle_rsc_0_7_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_7_i_bcwt <= '0';
      ELSE
        twiddle_rsc_0_7_i_bcwt <= NOT((NOT(twiddle_rsc_0_7_i_bcwt OR twiddle_rsc_0_7_i_biwt))
            OR twiddle_rsc_0_7_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_7_i_biwt = '1' ) THEN
        twiddle_rsc_0_7_i_qb_d_bfwt <= twiddle_rsc_0_7_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_0_7_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_7_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_7_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_7_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_0_7_i_bdwt <= twiddle_rsc_0_7_i_oswt AND core_wen;
  twiddle_rsc_0_7_i_biwt <= (NOT core_wten) AND twiddle_rsc_0_7_i_oswt;
  twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_rsc_0_7_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_6_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_6_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_6_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsc_0_6_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_6_i_qb_d, twiddle_rsc_0_6_i_qb_d_bfwt,
      twiddle_rsc_0_6_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_6_i_bcwt <= '0';
      ELSE
        twiddle_rsc_0_6_i_bcwt <= NOT((NOT(twiddle_rsc_0_6_i_bcwt OR twiddle_rsc_0_6_i_biwt))
            OR twiddle_rsc_0_6_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_6_i_biwt = '1' ) THEN
        twiddle_rsc_0_6_i_qb_d_bfwt <= twiddle_rsc_0_6_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_0_6_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_6_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_6_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_6_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_0_6_i_bdwt <= twiddle_rsc_0_6_i_oswt AND core_wen;
  twiddle_rsc_0_6_i_biwt <= (NOT core_wten) AND twiddle_rsc_0_6_i_oswt;
  twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_rsc_0_6_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_5_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_5_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_5_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsc_0_5_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_5_i_qb_d, twiddle_rsc_0_5_i_qb_d_bfwt,
      twiddle_rsc_0_5_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_5_i_bcwt <= '0';
      ELSE
        twiddle_rsc_0_5_i_bcwt <= NOT((NOT(twiddle_rsc_0_5_i_bcwt OR twiddle_rsc_0_5_i_biwt))
            OR twiddle_rsc_0_5_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_5_i_biwt = '1' ) THEN
        twiddle_rsc_0_5_i_qb_d_bfwt <= twiddle_rsc_0_5_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_0_5_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_5_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_5_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_5_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_0_5_i_bdwt <= twiddle_rsc_0_5_i_oswt AND core_wen;
  twiddle_rsc_0_5_i_biwt <= (NOT core_wten) AND twiddle_rsc_0_5_i_oswt;
  twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_rsc_0_5_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_4_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_4_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_4_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsc_0_4_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_4_i_qb_d, twiddle_rsc_0_4_i_qb_d_bfwt,
      twiddle_rsc_0_4_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_4_i_bcwt <= '0';
      ELSE
        twiddle_rsc_0_4_i_bcwt <= NOT((NOT(twiddle_rsc_0_4_i_bcwt OR twiddle_rsc_0_4_i_biwt))
            OR twiddle_rsc_0_4_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_4_i_biwt = '1' ) THEN
        twiddle_rsc_0_4_i_qb_d_bfwt <= twiddle_rsc_0_4_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_0_4_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_4_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_4_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_4_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_0_4_i_bdwt <= twiddle_rsc_0_4_i_oswt AND core_wen;
  twiddle_rsc_0_4_i_biwt <= (NOT core_wten) AND twiddle_rsc_0_4_i_oswt;
  twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_rsc_0_4_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_3_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_3_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_3_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsc_0_3_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_3_i_qb_d, twiddle_rsc_0_3_i_qb_d_bfwt,
      twiddle_rsc_0_3_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_3_i_bcwt <= '0';
      ELSE
        twiddle_rsc_0_3_i_bcwt <= NOT((NOT(twiddle_rsc_0_3_i_bcwt OR twiddle_rsc_0_3_i_biwt))
            OR twiddle_rsc_0_3_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_3_i_biwt = '1' ) THEN
        twiddle_rsc_0_3_i_qb_d_bfwt <= twiddle_rsc_0_3_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_0_3_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_3_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_3_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_3_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_0_3_i_bdwt <= twiddle_rsc_0_3_i_oswt AND core_wen;
  twiddle_rsc_0_3_i_biwt <= (NOT core_wten) AND twiddle_rsc_0_3_i_oswt;
  twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_rsc_0_3_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_2_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_2_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_2_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsc_0_2_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_2_i_qb_d, twiddle_rsc_0_2_i_qb_d_bfwt,
      twiddle_rsc_0_2_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_2_i_bcwt <= '0';
      ELSE
        twiddle_rsc_0_2_i_bcwt <= NOT((NOT(twiddle_rsc_0_2_i_bcwt OR twiddle_rsc_0_2_i_biwt))
            OR twiddle_rsc_0_2_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_2_i_biwt = '1' ) THEN
        twiddle_rsc_0_2_i_qb_d_bfwt <= twiddle_rsc_0_2_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_0_2_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_2_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_2_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_2_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_0_2_i_bdwt <= twiddle_rsc_0_2_i_oswt AND core_wen;
  twiddle_rsc_0_2_i_biwt <= (NOT core_wten) AND twiddle_rsc_0_2_i_oswt;
  twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_rsc_0_2_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_1_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_1_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_1_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsc_0_1_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_1_i_qb_d, twiddle_rsc_0_1_i_qb_d_bfwt,
      twiddle_rsc_0_1_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_1_i_bcwt <= '0';
      ELSE
        twiddle_rsc_0_1_i_bcwt <= NOT((NOT(twiddle_rsc_0_1_i_bcwt OR twiddle_rsc_0_1_i_biwt))
            OR twiddle_rsc_0_1_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_1_i_biwt = '1' ) THEN
        twiddle_rsc_0_1_i_qb_d_bfwt <= twiddle_rsc_0_1_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_0_1_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_1_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_1_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_1_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_0_1_i_bdwt <= twiddle_rsc_0_1_i_oswt AND core_wen;
  twiddle_rsc_0_1_i_biwt <= (NOT core_wten) AND twiddle_rsc_0_1_i_oswt;
  twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_rsc_0_1_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_0_i_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_0_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_0_i_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsc_0_0_i_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_0_i_qb_d, twiddle_rsc_0_0_i_qb_d_bfwt,
      twiddle_rsc_0_0_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_0_i_bcwt <= '0';
      ELSE
        twiddle_rsc_0_0_i_bcwt <= NOT((NOT(twiddle_rsc_0_0_i_bcwt OR twiddle_rsc_0_0_i_biwt))
            OR twiddle_rsc_0_0_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_0_i_biwt = '1' ) THEN
        twiddle_rsc_0_0_i_qb_d_bfwt <= twiddle_rsc_0_0_i_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_ctrl
    IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_0_0_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_0_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_0_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_0_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_0_0_i_bdwt <= twiddle_rsc_0_0_i_oswt AND core_wen;
  twiddle_rsc_0_0_i_biwt <= (NOT core_wten) AND twiddle_rsc_0_0_i_oswt;
  twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct <= twiddle_rsc_0_0_i_oswt_pff
      AND (NOT core_wten_pff);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_1_7_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_7_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_7_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_7_i_biwt : IN STD_LOGIC;
    vec_rsc_1_7_i_bdwt : IN STD_LOGIC;
    vec_rsc_1_7_i_biwt_1 : IN STD_LOGIC;
    vec_rsc_1_7_i_bdwt_2 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_7_i_bcwt : STD_LOGIC;
  SIGNAL vec_rsc_1_7_i_bcwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_1_7_i_qa_d_bfwt_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_qa_d_bfwt_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL VEC_LOOP_mux_62_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_63_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  VEC_LOOP_mux_62_nl <= MUX_v_32_2_2((vec_rsc_1_7_i_qa_d(63 DOWNTO 32)), vec_rsc_1_7_i_qa_d_bfwt_63_32,
      vec_rsc_1_7_i_bcwt_1);
  VEC_LOOP_mux_63_nl <= MUX_v_32_2_2((vec_rsc_1_7_i_qa_d(31 DOWNTO 0)), vec_rsc_1_7_i_qa_d_bfwt_31_0,
      vec_rsc_1_7_i_bcwt);
  vec_rsc_1_7_i_qa_d_mxwt <= VEC_LOOP_mux_62_nl & VEC_LOOP_mux_63_nl;
  vec_rsc_1_7_i_da_d <= vec_rsc_1_7_i_da_d_core(31 DOWNTO 0);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        vec_rsc_1_7_i_bcwt <= '0';
        vec_rsc_1_7_i_bcwt_1 <= '0';
      ELSE
        vec_rsc_1_7_i_bcwt <= NOT((NOT(vec_rsc_1_7_i_bcwt OR vec_rsc_1_7_i_biwt))
            OR vec_rsc_1_7_i_bdwt);
        vec_rsc_1_7_i_bcwt_1 <= NOT((NOT(vec_rsc_1_7_i_bcwt_1 OR vec_rsc_1_7_i_biwt_1))
            OR vec_rsc_1_7_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_1_7_i_biwt_1 = '1' ) THEN
        vec_rsc_1_7_i_qa_d_bfwt_63_32 <= vec_rsc_1_7_i_qa_d(63 DOWNTO 32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_1_7_i_biwt = '1' ) THEN
        vec_rsc_1_7_i_qa_d_bfwt_31_0 <= vec_rsc_1_7_i_qa_d(31 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_1_7_i_oswt : IN STD_LOGIC;
    vec_rsc_1_7_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_1_7_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_7_i_biwt : OUT STD_LOGIC;
    vec_rsc_1_7_i_bdwt : OUT STD_LOGIC;
    vec_rsc_1_7_i_biwt_1 : OUT STD_LOGIC;
    vec_rsc_1_7_i_bdwt_2 : OUT STD_LOGIC;
    vec_rsc_1_7_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_1_7_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_1_7_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_7_i_dswt_pff : STD_LOGIC;

  SIGNAL VEC_LOOP_and_173_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_177_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_175_nl : STD_LOGIC;
BEGIN
  vec_rsc_1_7_i_bdwt <= vec_rsc_1_7_i_oswt AND core_wen;
  vec_rsc_1_7_i_biwt <= (NOT core_wten) AND vec_rsc_1_7_i_oswt;
  vec_rsc_1_7_i_bdwt_2 <= vec_rsc_1_7_i_oswt_1 AND core_wen;
  vec_rsc_1_7_i_biwt_1 <= (NOT core_wten) AND vec_rsc_1_7_i_oswt_1;
  VEC_LOOP_and_173_nl <= (vec_rsc_1_7_i_wea_d_core_psct(0)) AND vec_rsc_1_7_i_dswt_pff;
  vec_rsc_1_7_i_wea_d_core_sct <= STD_LOGIC_VECTOR'( '0' & VEC_LOOP_and_173_nl);
  vec_rsc_1_7_i_dswt_pff <= (NOT core_wten_pff) AND vec_rsc_1_7_i_oswt_pff;
  VEC_LOOP_and_177_nl <= (NOT core_wten_pff) AND vec_rsc_1_7_i_oswt_1_pff;
  vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND STD_LOGIC_VECTOR'( VEC_LOOP_and_177_nl & vec_rsc_1_7_i_dswt_pff);
  VEC_LOOP_and_175_nl <= (vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0))
      AND vec_rsc_1_7_i_dswt_pff;
  vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= STD_LOGIC_VECTOR'( '0'
      & VEC_LOOP_and_175_nl);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_1_6_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_6_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_6_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_6_i_biwt : IN STD_LOGIC;
    vec_rsc_1_6_i_bdwt : IN STD_LOGIC;
    vec_rsc_1_6_i_biwt_1 : IN STD_LOGIC;
    vec_rsc_1_6_i_bdwt_2 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_6_i_bcwt : STD_LOGIC;
  SIGNAL vec_rsc_1_6_i_bcwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_1_6_i_qa_d_bfwt_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_qa_d_bfwt_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL VEC_LOOP_mux_58_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_59_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  VEC_LOOP_mux_58_nl <= MUX_v_32_2_2((vec_rsc_1_6_i_qa_d(63 DOWNTO 32)), vec_rsc_1_6_i_qa_d_bfwt_63_32,
      vec_rsc_1_6_i_bcwt_1);
  VEC_LOOP_mux_59_nl <= MUX_v_32_2_2((vec_rsc_1_6_i_qa_d(31 DOWNTO 0)), vec_rsc_1_6_i_qa_d_bfwt_31_0,
      vec_rsc_1_6_i_bcwt);
  vec_rsc_1_6_i_qa_d_mxwt <= VEC_LOOP_mux_58_nl & VEC_LOOP_mux_59_nl;
  vec_rsc_1_6_i_da_d <= vec_rsc_1_6_i_da_d_core(31 DOWNTO 0);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        vec_rsc_1_6_i_bcwt <= '0';
        vec_rsc_1_6_i_bcwt_1 <= '0';
      ELSE
        vec_rsc_1_6_i_bcwt <= NOT((NOT(vec_rsc_1_6_i_bcwt OR vec_rsc_1_6_i_biwt))
            OR vec_rsc_1_6_i_bdwt);
        vec_rsc_1_6_i_bcwt_1 <= NOT((NOT(vec_rsc_1_6_i_bcwt_1 OR vec_rsc_1_6_i_biwt_1))
            OR vec_rsc_1_6_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_1_6_i_biwt_1 = '1' ) THEN
        vec_rsc_1_6_i_qa_d_bfwt_63_32 <= vec_rsc_1_6_i_qa_d(63 DOWNTO 32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_1_6_i_biwt = '1' ) THEN
        vec_rsc_1_6_i_qa_d_bfwt_31_0 <= vec_rsc_1_6_i_qa_d(31 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_1_6_i_oswt : IN STD_LOGIC;
    vec_rsc_1_6_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_1_6_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_6_i_biwt : OUT STD_LOGIC;
    vec_rsc_1_6_i_bdwt : OUT STD_LOGIC;
    vec_rsc_1_6_i_biwt_1 : OUT STD_LOGIC;
    vec_rsc_1_6_i_bdwt_2 : OUT STD_LOGIC;
    vec_rsc_1_6_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_1_6_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_1_6_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_6_i_dswt_pff : STD_LOGIC;

  SIGNAL VEC_LOOP_and_162_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_166_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_164_nl : STD_LOGIC;
BEGIN
  vec_rsc_1_6_i_bdwt <= vec_rsc_1_6_i_oswt AND core_wen;
  vec_rsc_1_6_i_biwt <= (NOT core_wten) AND vec_rsc_1_6_i_oswt;
  vec_rsc_1_6_i_bdwt_2 <= vec_rsc_1_6_i_oswt_1 AND core_wen;
  vec_rsc_1_6_i_biwt_1 <= (NOT core_wten) AND vec_rsc_1_6_i_oswt_1;
  VEC_LOOP_and_162_nl <= (vec_rsc_1_6_i_wea_d_core_psct(0)) AND vec_rsc_1_6_i_dswt_pff;
  vec_rsc_1_6_i_wea_d_core_sct <= STD_LOGIC_VECTOR'( '0' & VEC_LOOP_and_162_nl);
  vec_rsc_1_6_i_dswt_pff <= (NOT core_wten_pff) AND vec_rsc_1_6_i_oswt_pff;
  VEC_LOOP_and_166_nl <= (NOT core_wten_pff) AND vec_rsc_1_6_i_oswt_1_pff;
  vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND STD_LOGIC_VECTOR'( VEC_LOOP_and_166_nl & vec_rsc_1_6_i_dswt_pff);
  VEC_LOOP_and_164_nl <= (vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0))
      AND vec_rsc_1_6_i_dswt_pff;
  vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= STD_LOGIC_VECTOR'( '0'
      & VEC_LOOP_and_164_nl);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_1_5_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_5_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_5_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_5_i_biwt : IN STD_LOGIC;
    vec_rsc_1_5_i_bdwt : IN STD_LOGIC;
    vec_rsc_1_5_i_biwt_1 : IN STD_LOGIC;
    vec_rsc_1_5_i_bdwt_2 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_5_i_bcwt : STD_LOGIC;
  SIGNAL vec_rsc_1_5_i_bcwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_1_5_i_qa_d_bfwt_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_qa_d_bfwt_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL VEC_LOOP_mux_54_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_55_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  VEC_LOOP_mux_54_nl <= MUX_v_32_2_2((vec_rsc_1_5_i_qa_d(63 DOWNTO 32)), vec_rsc_1_5_i_qa_d_bfwt_63_32,
      vec_rsc_1_5_i_bcwt_1);
  VEC_LOOP_mux_55_nl <= MUX_v_32_2_2((vec_rsc_1_5_i_qa_d(31 DOWNTO 0)), vec_rsc_1_5_i_qa_d_bfwt_31_0,
      vec_rsc_1_5_i_bcwt);
  vec_rsc_1_5_i_qa_d_mxwt <= VEC_LOOP_mux_54_nl & VEC_LOOP_mux_55_nl;
  vec_rsc_1_5_i_da_d <= vec_rsc_1_5_i_da_d_core(31 DOWNTO 0);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        vec_rsc_1_5_i_bcwt <= '0';
        vec_rsc_1_5_i_bcwt_1 <= '0';
      ELSE
        vec_rsc_1_5_i_bcwt <= NOT((NOT(vec_rsc_1_5_i_bcwt OR vec_rsc_1_5_i_biwt))
            OR vec_rsc_1_5_i_bdwt);
        vec_rsc_1_5_i_bcwt_1 <= NOT((NOT(vec_rsc_1_5_i_bcwt_1 OR vec_rsc_1_5_i_biwt_1))
            OR vec_rsc_1_5_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_1_5_i_biwt_1 = '1' ) THEN
        vec_rsc_1_5_i_qa_d_bfwt_63_32 <= vec_rsc_1_5_i_qa_d(63 DOWNTO 32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_1_5_i_biwt = '1' ) THEN
        vec_rsc_1_5_i_qa_d_bfwt_31_0 <= vec_rsc_1_5_i_qa_d(31 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_1_5_i_oswt : IN STD_LOGIC;
    vec_rsc_1_5_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_1_5_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_5_i_biwt : OUT STD_LOGIC;
    vec_rsc_1_5_i_bdwt : OUT STD_LOGIC;
    vec_rsc_1_5_i_biwt_1 : OUT STD_LOGIC;
    vec_rsc_1_5_i_bdwt_2 : OUT STD_LOGIC;
    vec_rsc_1_5_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_1_5_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_1_5_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_5_i_dswt_pff : STD_LOGIC;

  SIGNAL VEC_LOOP_and_151_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_155_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_153_nl : STD_LOGIC;
BEGIN
  vec_rsc_1_5_i_bdwt <= vec_rsc_1_5_i_oswt AND core_wen;
  vec_rsc_1_5_i_biwt <= (NOT core_wten) AND vec_rsc_1_5_i_oswt;
  vec_rsc_1_5_i_bdwt_2 <= vec_rsc_1_5_i_oswt_1 AND core_wen;
  vec_rsc_1_5_i_biwt_1 <= (NOT core_wten) AND vec_rsc_1_5_i_oswt_1;
  VEC_LOOP_and_151_nl <= (vec_rsc_1_5_i_wea_d_core_psct(0)) AND vec_rsc_1_5_i_dswt_pff;
  vec_rsc_1_5_i_wea_d_core_sct <= STD_LOGIC_VECTOR'( '0' & VEC_LOOP_and_151_nl);
  vec_rsc_1_5_i_dswt_pff <= (NOT core_wten_pff) AND vec_rsc_1_5_i_oswt_pff;
  VEC_LOOP_and_155_nl <= (NOT core_wten_pff) AND vec_rsc_1_5_i_oswt_1_pff;
  vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND STD_LOGIC_VECTOR'( VEC_LOOP_and_155_nl & vec_rsc_1_5_i_dswt_pff);
  VEC_LOOP_and_153_nl <= (vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0))
      AND vec_rsc_1_5_i_dswt_pff;
  vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= STD_LOGIC_VECTOR'( '0'
      & VEC_LOOP_and_153_nl);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_1_4_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_4_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_4_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_4_i_biwt : IN STD_LOGIC;
    vec_rsc_1_4_i_bdwt : IN STD_LOGIC;
    vec_rsc_1_4_i_biwt_1 : IN STD_LOGIC;
    vec_rsc_1_4_i_bdwt_2 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_4_i_bcwt : STD_LOGIC;
  SIGNAL vec_rsc_1_4_i_bcwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_1_4_i_qa_d_bfwt_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_qa_d_bfwt_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL VEC_LOOP_mux_50_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_51_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  VEC_LOOP_mux_50_nl <= MUX_v_32_2_2((vec_rsc_1_4_i_qa_d(63 DOWNTO 32)), vec_rsc_1_4_i_qa_d_bfwt_63_32,
      vec_rsc_1_4_i_bcwt_1);
  VEC_LOOP_mux_51_nl <= MUX_v_32_2_2((vec_rsc_1_4_i_qa_d(31 DOWNTO 0)), vec_rsc_1_4_i_qa_d_bfwt_31_0,
      vec_rsc_1_4_i_bcwt);
  vec_rsc_1_4_i_qa_d_mxwt <= VEC_LOOP_mux_50_nl & VEC_LOOP_mux_51_nl;
  vec_rsc_1_4_i_da_d <= vec_rsc_1_4_i_da_d_core(31 DOWNTO 0);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        vec_rsc_1_4_i_bcwt <= '0';
        vec_rsc_1_4_i_bcwt_1 <= '0';
      ELSE
        vec_rsc_1_4_i_bcwt <= NOT((NOT(vec_rsc_1_4_i_bcwt OR vec_rsc_1_4_i_biwt))
            OR vec_rsc_1_4_i_bdwt);
        vec_rsc_1_4_i_bcwt_1 <= NOT((NOT(vec_rsc_1_4_i_bcwt_1 OR vec_rsc_1_4_i_biwt_1))
            OR vec_rsc_1_4_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_1_4_i_biwt_1 = '1' ) THEN
        vec_rsc_1_4_i_qa_d_bfwt_63_32 <= vec_rsc_1_4_i_qa_d(63 DOWNTO 32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_1_4_i_biwt = '1' ) THEN
        vec_rsc_1_4_i_qa_d_bfwt_31_0 <= vec_rsc_1_4_i_qa_d(31 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_1_4_i_oswt : IN STD_LOGIC;
    vec_rsc_1_4_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_1_4_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_4_i_biwt : OUT STD_LOGIC;
    vec_rsc_1_4_i_bdwt : OUT STD_LOGIC;
    vec_rsc_1_4_i_biwt_1 : OUT STD_LOGIC;
    vec_rsc_1_4_i_bdwt_2 : OUT STD_LOGIC;
    vec_rsc_1_4_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_1_4_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_1_4_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_4_i_dswt_pff : STD_LOGIC;

  SIGNAL VEC_LOOP_and_140_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_144_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_142_nl : STD_LOGIC;
BEGIN
  vec_rsc_1_4_i_bdwt <= vec_rsc_1_4_i_oswt AND core_wen;
  vec_rsc_1_4_i_biwt <= (NOT core_wten) AND vec_rsc_1_4_i_oswt;
  vec_rsc_1_4_i_bdwt_2 <= vec_rsc_1_4_i_oswt_1 AND core_wen;
  vec_rsc_1_4_i_biwt_1 <= (NOT core_wten) AND vec_rsc_1_4_i_oswt_1;
  VEC_LOOP_and_140_nl <= (vec_rsc_1_4_i_wea_d_core_psct(0)) AND vec_rsc_1_4_i_dswt_pff;
  vec_rsc_1_4_i_wea_d_core_sct <= STD_LOGIC_VECTOR'( '0' & VEC_LOOP_and_140_nl);
  vec_rsc_1_4_i_dswt_pff <= (NOT core_wten_pff) AND vec_rsc_1_4_i_oswt_pff;
  VEC_LOOP_and_144_nl <= (NOT core_wten_pff) AND vec_rsc_1_4_i_oswt_1_pff;
  vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND STD_LOGIC_VECTOR'( VEC_LOOP_and_144_nl & vec_rsc_1_4_i_dswt_pff);
  VEC_LOOP_and_142_nl <= (vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0))
      AND vec_rsc_1_4_i_dswt_pff;
  vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= STD_LOGIC_VECTOR'( '0'
      & VEC_LOOP_and_142_nl);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_1_3_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_3_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_3_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_3_i_biwt : IN STD_LOGIC;
    vec_rsc_1_3_i_bdwt : IN STD_LOGIC;
    vec_rsc_1_3_i_biwt_1 : IN STD_LOGIC;
    vec_rsc_1_3_i_bdwt_2 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_3_i_bcwt : STD_LOGIC;
  SIGNAL vec_rsc_1_3_i_bcwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_1_3_i_qa_d_bfwt_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_qa_d_bfwt_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL VEC_LOOP_mux_46_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_47_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  VEC_LOOP_mux_46_nl <= MUX_v_32_2_2((vec_rsc_1_3_i_qa_d(63 DOWNTO 32)), vec_rsc_1_3_i_qa_d_bfwt_63_32,
      vec_rsc_1_3_i_bcwt_1);
  VEC_LOOP_mux_47_nl <= MUX_v_32_2_2((vec_rsc_1_3_i_qa_d(31 DOWNTO 0)), vec_rsc_1_3_i_qa_d_bfwt_31_0,
      vec_rsc_1_3_i_bcwt);
  vec_rsc_1_3_i_qa_d_mxwt <= VEC_LOOP_mux_46_nl & VEC_LOOP_mux_47_nl;
  vec_rsc_1_3_i_da_d <= vec_rsc_1_3_i_da_d_core(31 DOWNTO 0);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        vec_rsc_1_3_i_bcwt <= '0';
        vec_rsc_1_3_i_bcwt_1 <= '0';
      ELSE
        vec_rsc_1_3_i_bcwt <= NOT((NOT(vec_rsc_1_3_i_bcwt OR vec_rsc_1_3_i_biwt))
            OR vec_rsc_1_3_i_bdwt);
        vec_rsc_1_3_i_bcwt_1 <= NOT((NOT(vec_rsc_1_3_i_bcwt_1 OR vec_rsc_1_3_i_biwt_1))
            OR vec_rsc_1_3_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_1_3_i_biwt_1 = '1' ) THEN
        vec_rsc_1_3_i_qa_d_bfwt_63_32 <= vec_rsc_1_3_i_qa_d(63 DOWNTO 32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_1_3_i_biwt = '1' ) THEN
        vec_rsc_1_3_i_qa_d_bfwt_31_0 <= vec_rsc_1_3_i_qa_d(31 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_1_3_i_oswt : IN STD_LOGIC;
    vec_rsc_1_3_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_1_3_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_3_i_biwt : OUT STD_LOGIC;
    vec_rsc_1_3_i_bdwt : OUT STD_LOGIC;
    vec_rsc_1_3_i_biwt_1 : OUT STD_LOGIC;
    vec_rsc_1_3_i_bdwt_2 : OUT STD_LOGIC;
    vec_rsc_1_3_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_1_3_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_1_3_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_3_i_dswt_pff : STD_LOGIC;

  SIGNAL VEC_LOOP_and_129_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_133_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_131_nl : STD_LOGIC;
BEGIN
  vec_rsc_1_3_i_bdwt <= vec_rsc_1_3_i_oswt AND core_wen;
  vec_rsc_1_3_i_biwt <= (NOT core_wten) AND vec_rsc_1_3_i_oswt;
  vec_rsc_1_3_i_bdwt_2 <= vec_rsc_1_3_i_oswt_1 AND core_wen;
  vec_rsc_1_3_i_biwt_1 <= (NOT core_wten) AND vec_rsc_1_3_i_oswt_1;
  VEC_LOOP_and_129_nl <= (vec_rsc_1_3_i_wea_d_core_psct(0)) AND vec_rsc_1_3_i_dswt_pff;
  vec_rsc_1_3_i_wea_d_core_sct <= STD_LOGIC_VECTOR'( '0' & VEC_LOOP_and_129_nl);
  vec_rsc_1_3_i_dswt_pff <= (NOT core_wten_pff) AND vec_rsc_1_3_i_oswt_pff;
  VEC_LOOP_and_133_nl <= (NOT core_wten_pff) AND vec_rsc_1_3_i_oswt_1_pff;
  vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND STD_LOGIC_VECTOR'( VEC_LOOP_and_133_nl & vec_rsc_1_3_i_dswt_pff);
  VEC_LOOP_and_131_nl <= (vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0))
      AND vec_rsc_1_3_i_dswt_pff;
  vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= STD_LOGIC_VECTOR'( '0'
      & VEC_LOOP_and_131_nl);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_1_2_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_2_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_2_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_2_i_biwt : IN STD_LOGIC;
    vec_rsc_1_2_i_bdwt : IN STD_LOGIC;
    vec_rsc_1_2_i_biwt_1 : IN STD_LOGIC;
    vec_rsc_1_2_i_bdwt_2 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_2_i_bcwt : STD_LOGIC;
  SIGNAL vec_rsc_1_2_i_bcwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_1_2_i_qa_d_bfwt_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_qa_d_bfwt_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL VEC_LOOP_mux_42_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_43_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  VEC_LOOP_mux_42_nl <= MUX_v_32_2_2((vec_rsc_1_2_i_qa_d(63 DOWNTO 32)), vec_rsc_1_2_i_qa_d_bfwt_63_32,
      vec_rsc_1_2_i_bcwt_1);
  VEC_LOOP_mux_43_nl <= MUX_v_32_2_2((vec_rsc_1_2_i_qa_d(31 DOWNTO 0)), vec_rsc_1_2_i_qa_d_bfwt_31_0,
      vec_rsc_1_2_i_bcwt);
  vec_rsc_1_2_i_qa_d_mxwt <= VEC_LOOP_mux_42_nl & VEC_LOOP_mux_43_nl;
  vec_rsc_1_2_i_da_d <= vec_rsc_1_2_i_da_d_core(31 DOWNTO 0);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        vec_rsc_1_2_i_bcwt <= '0';
        vec_rsc_1_2_i_bcwt_1 <= '0';
      ELSE
        vec_rsc_1_2_i_bcwt <= NOT((NOT(vec_rsc_1_2_i_bcwt OR vec_rsc_1_2_i_biwt))
            OR vec_rsc_1_2_i_bdwt);
        vec_rsc_1_2_i_bcwt_1 <= NOT((NOT(vec_rsc_1_2_i_bcwt_1 OR vec_rsc_1_2_i_biwt_1))
            OR vec_rsc_1_2_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_1_2_i_biwt_1 = '1' ) THEN
        vec_rsc_1_2_i_qa_d_bfwt_63_32 <= vec_rsc_1_2_i_qa_d(63 DOWNTO 32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_1_2_i_biwt = '1' ) THEN
        vec_rsc_1_2_i_qa_d_bfwt_31_0 <= vec_rsc_1_2_i_qa_d(31 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_1_2_i_oswt : IN STD_LOGIC;
    vec_rsc_1_2_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_1_2_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_2_i_biwt : OUT STD_LOGIC;
    vec_rsc_1_2_i_bdwt : OUT STD_LOGIC;
    vec_rsc_1_2_i_biwt_1 : OUT STD_LOGIC;
    vec_rsc_1_2_i_bdwt_2 : OUT STD_LOGIC;
    vec_rsc_1_2_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_1_2_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_1_2_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_2_i_dswt_pff : STD_LOGIC;

  SIGNAL VEC_LOOP_and_118_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_122_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_120_nl : STD_LOGIC;
BEGIN
  vec_rsc_1_2_i_bdwt <= vec_rsc_1_2_i_oswt AND core_wen;
  vec_rsc_1_2_i_biwt <= (NOT core_wten) AND vec_rsc_1_2_i_oswt;
  vec_rsc_1_2_i_bdwt_2 <= vec_rsc_1_2_i_oswt_1 AND core_wen;
  vec_rsc_1_2_i_biwt_1 <= (NOT core_wten) AND vec_rsc_1_2_i_oswt_1;
  VEC_LOOP_and_118_nl <= (vec_rsc_1_2_i_wea_d_core_psct(0)) AND vec_rsc_1_2_i_dswt_pff;
  vec_rsc_1_2_i_wea_d_core_sct <= STD_LOGIC_VECTOR'( '0' & VEC_LOOP_and_118_nl);
  vec_rsc_1_2_i_dswt_pff <= (NOT core_wten_pff) AND vec_rsc_1_2_i_oswt_pff;
  VEC_LOOP_and_122_nl <= (NOT core_wten_pff) AND vec_rsc_1_2_i_oswt_1_pff;
  vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND STD_LOGIC_VECTOR'( VEC_LOOP_and_122_nl & vec_rsc_1_2_i_dswt_pff);
  VEC_LOOP_and_120_nl <= (vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0))
      AND vec_rsc_1_2_i_dswt_pff;
  vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= STD_LOGIC_VECTOR'( '0'
      & VEC_LOOP_and_120_nl);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_1_1_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_1_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_1_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_1_i_biwt : IN STD_LOGIC;
    vec_rsc_1_1_i_bdwt : IN STD_LOGIC;
    vec_rsc_1_1_i_biwt_1 : IN STD_LOGIC;
    vec_rsc_1_1_i_bdwt_2 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_1_i_bcwt : STD_LOGIC;
  SIGNAL vec_rsc_1_1_i_bcwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_1_1_i_qa_d_bfwt_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_qa_d_bfwt_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL VEC_LOOP_mux_38_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_39_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  VEC_LOOP_mux_38_nl <= MUX_v_32_2_2((vec_rsc_1_1_i_qa_d(63 DOWNTO 32)), vec_rsc_1_1_i_qa_d_bfwt_63_32,
      vec_rsc_1_1_i_bcwt_1);
  VEC_LOOP_mux_39_nl <= MUX_v_32_2_2((vec_rsc_1_1_i_qa_d(31 DOWNTO 0)), vec_rsc_1_1_i_qa_d_bfwt_31_0,
      vec_rsc_1_1_i_bcwt);
  vec_rsc_1_1_i_qa_d_mxwt <= VEC_LOOP_mux_38_nl & VEC_LOOP_mux_39_nl;
  vec_rsc_1_1_i_da_d <= vec_rsc_1_1_i_da_d_core(31 DOWNTO 0);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        vec_rsc_1_1_i_bcwt <= '0';
        vec_rsc_1_1_i_bcwt_1 <= '0';
      ELSE
        vec_rsc_1_1_i_bcwt <= NOT((NOT(vec_rsc_1_1_i_bcwt OR vec_rsc_1_1_i_biwt))
            OR vec_rsc_1_1_i_bdwt);
        vec_rsc_1_1_i_bcwt_1 <= NOT((NOT(vec_rsc_1_1_i_bcwt_1 OR vec_rsc_1_1_i_biwt_1))
            OR vec_rsc_1_1_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_1_1_i_biwt_1 = '1' ) THEN
        vec_rsc_1_1_i_qa_d_bfwt_63_32 <= vec_rsc_1_1_i_qa_d(63 DOWNTO 32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_1_1_i_biwt = '1' ) THEN
        vec_rsc_1_1_i_qa_d_bfwt_31_0 <= vec_rsc_1_1_i_qa_d(31 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_1_1_i_oswt : IN STD_LOGIC;
    vec_rsc_1_1_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_1_1_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_1_i_biwt : OUT STD_LOGIC;
    vec_rsc_1_1_i_bdwt : OUT STD_LOGIC;
    vec_rsc_1_1_i_biwt_1 : OUT STD_LOGIC;
    vec_rsc_1_1_i_bdwt_2 : OUT STD_LOGIC;
    vec_rsc_1_1_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_1_1_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_1_1_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_1_i_dswt_pff : STD_LOGIC;

  SIGNAL VEC_LOOP_and_107_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_111_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_109_nl : STD_LOGIC;
BEGIN
  vec_rsc_1_1_i_bdwt <= vec_rsc_1_1_i_oswt AND core_wen;
  vec_rsc_1_1_i_biwt <= (NOT core_wten) AND vec_rsc_1_1_i_oswt;
  vec_rsc_1_1_i_bdwt_2 <= vec_rsc_1_1_i_oswt_1 AND core_wen;
  vec_rsc_1_1_i_biwt_1 <= (NOT core_wten) AND vec_rsc_1_1_i_oswt_1;
  VEC_LOOP_and_107_nl <= (vec_rsc_1_1_i_wea_d_core_psct(0)) AND vec_rsc_1_1_i_dswt_pff;
  vec_rsc_1_1_i_wea_d_core_sct <= STD_LOGIC_VECTOR'( '0' & VEC_LOOP_and_107_nl);
  vec_rsc_1_1_i_dswt_pff <= (NOT core_wten_pff) AND vec_rsc_1_1_i_oswt_pff;
  VEC_LOOP_and_111_nl <= (NOT core_wten_pff) AND vec_rsc_1_1_i_oswt_1_pff;
  vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND STD_LOGIC_VECTOR'( VEC_LOOP_and_111_nl & vec_rsc_1_1_i_dswt_pff);
  VEC_LOOP_and_109_nl <= (vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0))
      AND vec_rsc_1_1_i_dswt_pff;
  vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= STD_LOGIC_VECTOR'( '0'
      & VEC_LOOP_and_109_nl);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_1_0_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_0_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_0_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_0_i_biwt : IN STD_LOGIC;
    vec_rsc_1_0_i_bdwt : IN STD_LOGIC;
    vec_rsc_1_0_i_biwt_1 : IN STD_LOGIC;
    vec_rsc_1_0_i_bdwt_2 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_0_i_bcwt : STD_LOGIC;
  SIGNAL vec_rsc_1_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_1_0_i_qa_d_bfwt_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_qa_d_bfwt_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL VEC_LOOP_mux_34_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_35_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  VEC_LOOP_mux_34_nl <= MUX_v_32_2_2((vec_rsc_1_0_i_qa_d(63 DOWNTO 32)), vec_rsc_1_0_i_qa_d_bfwt_63_32,
      vec_rsc_1_0_i_bcwt_1);
  VEC_LOOP_mux_35_nl <= MUX_v_32_2_2((vec_rsc_1_0_i_qa_d(31 DOWNTO 0)), vec_rsc_1_0_i_qa_d_bfwt_31_0,
      vec_rsc_1_0_i_bcwt);
  vec_rsc_1_0_i_qa_d_mxwt <= VEC_LOOP_mux_34_nl & VEC_LOOP_mux_35_nl;
  vec_rsc_1_0_i_da_d <= vec_rsc_1_0_i_da_d_core(31 DOWNTO 0);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        vec_rsc_1_0_i_bcwt <= '0';
        vec_rsc_1_0_i_bcwt_1 <= '0';
      ELSE
        vec_rsc_1_0_i_bcwt <= NOT((NOT(vec_rsc_1_0_i_bcwt OR vec_rsc_1_0_i_biwt))
            OR vec_rsc_1_0_i_bdwt);
        vec_rsc_1_0_i_bcwt_1 <= NOT((NOT(vec_rsc_1_0_i_bcwt_1 OR vec_rsc_1_0_i_biwt_1))
            OR vec_rsc_1_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_1_0_i_biwt_1 = '1' ) THEN
        vec_rsc_1_0_i_qa_d_bfwt_63_32 <= vec_rsc_1_0_i_qa_d(63 DOWNTO 32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_1_0_i_biwt = '1' ) THEN
        vec_rsc_1_0_i_qa_d_bfwt_31_0 <= vec_rsc_1_0_i_qa_d(31 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_1_0_i_oswt : IN STD_LOGIC;
    vec_rsc_1_0_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_1_0_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_0_i_biwt : OUT STD_LOGIC;
    vec_rsc_1_0_i_bdwt : OUT STD_LOGIC;
    vec_rsc_1_0_i_biwt_1 : OUT STD_LOGIC;
    vec_rsc_1_0_i_bdwt_2 : OUT STD_LOGIC;
    vec_rsc_1_0_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_1_0_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_1_0_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_0_i_dswt_pff : STD_LOGIC;

  SIGNAL VEC_LOOP_and_96_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_100_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_98_nl : STD_LOGIC;
BEGIN
  vec_rsc_1_0_i_bdwt <= vec_rsc_1_0_i_oswt AND core_wen;
  vec_rsc_1_0_i_biwt <= (NOT core_wten) AND vec_rsc_1_0_i_oswt;
  vec_rsc_1_0_i_bdwt_2 <= vec_rsc_1_0_i_oswt_1 AND core_wen;
  vec_rsc_1_0_i_biwt_1 <= (NOT core_wten) AND vec_rsc_1_0_i_oswt_1;
  VEC_LOOP_and_96_nl <= (vec_rsc_1_0_i_wea_d_core_psct(0)) AND vec_rsc_1_0_i_dswt_pff;
  vec_rsc_1_0_i_wea_d_core_sct <= STD_LOGIC_VECTOR'( '0' & VEC_LOOP_and_96_nl);
  vec_rsc_1_0_i_dswt_pff <= (NOT core_wten_pff) AND vec_rsc_1_0_i_oswt_pff;
  VEC_LOOP_and_100_nl <= (NOT core_wten_pff) AND vec_rsc_1_0_i_oswt_1_pff;
  vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND STD_LOGIC_VECTOR'( VEC_LOOP_and_100_nl & vec_rsc_1_0_i_dswt_pff);
  VEC_LOOP_and_98_nl <= (vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0))
      AND vec_rsc_1_0_i_dswt_pff;
  vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= STD_LOGIC_VECTOR'( '0'
      & VEC_LOOP_and_98_nl);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_7_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_i_biwt : IN STD_LOGIC;
    vec_rsc_0_7_i_bdwt : IN STD_LOGIC;
    vec_rsc_0_7_i_biwt_1 : IN STD_LOGIC;
    vec_rsc_0_7_i_bdwt_2 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_7_i_bcwt : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_bcwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_qa_d_bfwt_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_qa_d_bfwt_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL VEC_LOOP_mux_30_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_31_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  VEC_LOOP_mux_30_nl <= MUX_v_32_2_2((vec_rsc_0_7_i_qa_d(63 DOWNTO 32)), vec_rsc_0_7_i_qa_d_bfwt_63_32,
      vec_rsc_0_7_i_bcwt_1);
  VEC_LOOP_mux_31_nl <= MUX_v_32_2_2((vec_rsc_0_7_i_qa_d(31 DOWNTO 0)), vec_rsc_0_7_i_qa_d_bfwt_31_0,
      vec_rsc_0_7_i_bcwt);
  vec_rsc_0_7_i_qa_d_mxwt <= VEC_LOOP_mux_30_nl & VEC_LOOP_mux_31_nl;
  vec_rsc_0_7_i_da_d <= vec_rsc_0_7_i_da_d_core(31 DOWNTO 0);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        vec_rsc_0_7_i_bcwt <= '0';
        vec_rsc_0_7_i_bcwt_1 <= '0';
      ELSE
        vec_rsc_0_7_i_bcwt <= NOT((NOT(vec_rsc_0_7_i_bcwt OR vec_rsc_0_7_i_biwt))
            OR vec_rsc_0_7_i_bdwt);
        vec_rsc_0_7_i_bcwt_1 <= NOT((NOT(vec_rsc_0_7_i_bcwt_1 OR vec_rsc_0_7_i_biwt_1))
            OR vec_rsc_0_7_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_0_7_i_biwt_1 = '1' ) THEN
        vec_rsc_0_7_i_qa_d_bfwt_63_32 <= vec_rsc_0_7_i_qa_d(63 DOWNTO 32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_0_7_i_biwt = '1' ) THEN
        vec_rsc_0_7_i_qa_d_bfwt_31_0 <= vec_rsc_0_7_i_qa_d(31 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_0_7_i_oswt : IN STD_LOGIC;
    vec_rsc_0_7_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_0_7_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_7_i_biwt : OUT STD_LOGIC;
    vec_rsc_0_7_i_bdwt : OUT STD_LOGIC;
    vec_rsc_0_7_i_biwt_1 : OUT STD_LOGIC;
    vec_rsc_0_7_i_bdwt_2 : OUT STD_LOGIC;
    vec_rsc_0_7_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_0_7_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_0_7_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_7_i_dswt_pff : STD_LOGIC;

  SIGNAL VEC_LOOP_and_85_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_89_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_87_nl : STD_LOGIC;
BEGIN
  vec_rsc_0_7_i_bdwt <= vec_rsc_0_7_i_oswt AND core_wen;
  vec_rsc_0_7_i_biwt <= (NOT core_wten) AND vec_rsc_0_7_i_oswt;
  vec_rsc_0_7_i_bdwt_2 <= vec_rsc_0_7_i_oswt_1 AND core_wen;
  vec_rsc_0_7_i_biwt_1 <= (NOT core_wten) AND vec_rsc_0_7_i_oswt_1;
  VEC_LOOP_and_85_nl <= (vec_rsc_0_7_i_wea_d_core_psct(0)) AND vec_rsc_0_7_i_dswt_pff;
  vec_rsc_0_7_i_wea_d_core_sct <= STD_LOGIC_VECTOR'( '0' & VEC_LOOP_and_85_nl);
  vec_rsc_0_7_i_dswt_pff <= (NOT core_wten_pff) AND vec_rsc_0_7_i_oswt_pff;
  VEC_LOOP_and_89_nl <= (NOT core_wten_pff) AND vec_rsc_0_7_i_oswt_1_pff;
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND STD_LOGIC_VECTOR'( VEC_LOOP_and_89_nl & vec_rsc_0_7_i_dswt_pff);
  VEC_LOOP_and_87_nl <= (vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0))
      AND vec_rsc_0_7_i_dswt_pff;
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= STD_LOGIC_VECTOR'( '0'
      & VEC_LOOP_and_87_nl);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_6_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_i_biwt : IN STD_LOGIC;
    vec_rsc_0_6_i_bdwt : IN STD_LOGIC;
    vec_rsc_0_6_i_biwt_1 : IN STD_LOGIC;
    vec_rsc_0_6_i_bdwt_2 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_6_i_bcwt : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_bcwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_qa_d_bfwt_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_qa_d_bfwt_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL VEC_LOOP_mux_26_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_27_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  VEC_LOOP_mux_26_nl <= MUX_v_32_2_2((vec_rsc_0_6_i_qa_d(63 DOWNTO 32)), vec_rsc_0_6_i_qa_d_bfwt_63_32,
      vec_rsc_0_6_i_bcwt_1);
  VEC_LOOP_mux_27_nl <= MUX_v_32_2_2((vec_rsc_0_6_i_qa_d(31 DOWNTO 0)), vec_rsc_0_6_i_qa_d_bfwt_31_0,
      vec_rsc_0_6_i_bcwt);
  vec_rsc_0_6_i_qa_d_mxwt <= VEC_LOOP_mux_26_nl & VEC_LOOP_mux_27_nl;
  vec_rsc_0_6_i_da_d <= vec_rsc_0_6_i_da_d_core(31 DOWNTO 0);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        vec_rsc_0_6_i_bcwt <= '0';
        vec_rsc_0_6_i_bcwt_1 <= '0';
      ELSE
        vec_rsc_0_6_i_bcwt <= NOT((NOT(vec_rsc_0_6_i_bcwt OR vec_rsc_0_6_i_biwt))
            OR vec_rsc_0_6_i_bdwt);
        vec_rsc_0_6_i_bcwt_1 <= NOT((NOT(vec_rsc_0_6_i_bcwt_1 OR vec_rsc_0_6_i_biwt_1))
            OR vec_rsc_0_6_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_0_6_i_biwt_1 = '1' ) THEN
        vec_rsc_0_6_i_qa_d_bfwt_63_32 <= vec_rsc_0_6_i_qa_d(63 DOWNTO 32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_0_6_i_biwt = '1' ) THEN
        vec_rsc_0_6_i_qa_d_bfwt_31_0 <= vec_rsc_0_6_i_qa_d(31 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_0_6_i_oswt : IN STD_LOGIC;
    vec_rsc_0_6_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_0_6_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_6_i_biwt : OUT STD_LOGIC;
    vec_rsc_0_6_i_bdwt : OUT STD_LOGIC;
    vec_rsc_0_6_i_biwt_1 : OUT STD_LOGIC;
    vec_rsc_0_6_i_bdwt_2 : OUT STD_LOGIC;
    vec_rsc_0_6_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_0_6_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_0_6_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_6_i_dswt_pff : STD_LOGIC;

  SIGNAL VEC_LOOP_and_74_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_78_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_76_nl : STD_LOGIC;
BEGIN
  vec_rsc_0_6_i_bdwt <= vec_rsc_0_6_i_oswt AND core_wen;
  vec_rsc_0_6_i_biwt <= (NOT core_wten) AND vec_rsc_0_6_i_oswt;
  vec_rsc_0_6_i_bdwt_2 <= vec_rsc_0_6_i_oswt_1 AND core_wen;
  vec_rsc_0_6_i_biwt_1 <= (NOT core_wten) AND vec_rsc_0_6_i_oswt_1;
  VEC_LOOP_and_74_nl <= (vec_rsc_0_6_i_wea_d_core_psct(0)) AND vec_rsc_0_6_i_dswt_pff;
  vec_rsc_0_6_i_wea_d_core_sct <= STD_LOGIC_VECTOR'( '0' & VEC_LOOP_and_74_nl);
  vec_rsc_0_6_i_dswt_pff <= (NOT core_wten_pff) AND vec_rsc_0_6_i_oswt_pff;
  VEC_LOOP_and_78_nl <= (NOT core_wten_pff) AND vec_rsc_0_6_i_oswt_1_pff;
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND STD_LOGIC_VECTOR'( VEC_LOOP_and_78_nl & vec_rsc_0_6_i_dswt_pff);
  VEC_LOOP_and_76_nl <= (vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0))
      AND vec_rsc_0_6_i_dswt_pff;
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= STD_LOGIC_VECTOR'( '0'
      & VEC_LOOP_and_76_nl);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_5_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_i_biwt : IN STD_LOGIC;
    vec_rsc_0_5_i_bdwt : IN STD_LOGIC;
    vec_rsc_0_5_i_biwt_1 : IN STD_LOGIC;
    vec_rsc_0_5_i_bdwt_2 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_5_i_bcwt : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_bcwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_qa_d_bfwt_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_qa_d_bfwt_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL VEC_LOOP_mux_22_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_23_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  VEC_LOOP_mux_22_nl <= MUX_v_32_2_2((vec_rsc_0_5_i_qa_d(63 DOWNTO 32)), vec_rsc_0_5_i_qa_d_bfwt_63_32,
      vec_rsc_0_5_i_bcwt_1);
  VEC_LOOP_mux_23_nl <= MUX_v_32_2_2((vec_rsc_0_5_i_qa_d(31 DOWNTO 0)), vec_rsc_0_5_i_qa_d_bfwt_31_0,
      vec_rsc_0_5_i_bcwt);
  vec_rsc_0_5_i_qa_d_mxwt <= VEC_LOOP_mux_22_nl & VEC_LOOP_mux_23_nl;
  vec_rsc_0_5_i_da_d <= vec_rsc_0_5_i_da_d_core(31 DOWNTO 0);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        vec_rsc_0_5_i_bcwt <= '0';
        vec_rsc_0_5_i_bcwt_1 <= '0';
      ELSE
        vec_rsc_0_5_i_bcwt <= NOT((NOT(vec_rsc_0_5_i_bcwt OR vec_rsc_0_5_i_biwt))
            OR vec_rsc_0_5_i_bdwt);
        vec_rsc_0_5_i_bcwt_1 <= NOT((NOT(vec_rsc_0_5_i_bcwt_1 OR vec_rsc_0_5_i_biwt_1))
            OR vec_rsc_0_5_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_0_5_i_biwt_1 = '1' ) THEN
        vec_rsc_0_5_i_qa_d_bfwt_63_32 <= vec_rsc_0_5_i_qa_d(63 DOWNTO 32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_0_5_i_biwt = '1' ) THEN
        vec_rsc_0_5_i_qa_d_bfwt_31_0 <= vec_rsc_0_5_i_qa_d(31 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_0_5_i_oswt : IN STD_LOGIC;
    vec_rsc_0_5_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_0_5_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_5_i_biwt : OUT STD_LOGIC;
    vec_rsc_0_5_i_bdwt : OUT STD_LOGIC;
    vec_rsc_0_5_i_biwt_1 : OUT STD_LOGIC;
    vec_rsc_0_5_i_bdwt_2 : OUT STD_LOGIC;
    vec_rsc_0_5_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_0_5_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_0_5_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_5_i_dswt_pff : STD_LOGIC;

  SIGNAL VEC_LOOP_and_63_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_67_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_65_nl : STD_LOGIC;
BEGIN
  vec_rsc_0_5_i_bdwt <= vec_rsc_0_5_i_oswt AND core_wen;
  vec_rsc_0_5_i_biwt <= (NOT core_wten) AND vec_rsc_0_5_i_oswt;
  vec_rsc_0_5_i_bdwt_2 <= vec_rsc_0_5_i_oswt_1 AND core_wen;
  vec_rsc_0_5_i_biwt_1 <= (NOT core_wten) AND vec_rsc_0_5_i_oswt_1;
  VEC_LOOP_and_63_nl <= (vec_rsc_0_5_i_wea_d_core_psct(0)) AND vec_rsc_0_5_i_dswt_pff;
  vec_rsc_0_5_i_wea_d_core_sct <= STD_LOGIC_VECTOR'( '0' & VEC_LOOP_and_63_nl);
  vec_rsc_0_5_i_dswt_pff <= (NOT core_wten_pff) AND vec_rsc_0_5_i_oswt_pff;
  VEC_LOOP_and_67_nl <= (NOT core_wten_pff) AND vec_rsc_0_5_i_oswt_1_pff;
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND STD_LOGIC_VECTOR'( VEC_LOOP_and_67_nl & vec_rsc_0_5_i_dswt_pff);
  VEC_LOOP_and_65_nl <= (vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0))
      AND vec_rsc_0_5_i_dswt_pff;
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= STD_LOGIC_VECTOR'( '0'
      & VEC_LOOP_and_65_nl);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_4_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_i_biwt : IN STD_LOGIC;
    vec_rsc_0_4_i_bdwt : IN STD_LOGIC;
    vec_rsc_0_4_i_biwt_1 : IN STD_LOGIC;
    vec_rsc_0_4_i_bdwt_2 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_4_i_bcwt : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_bcwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_qa_d_bfwt_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_qa_d_bfwt_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL VEC_LOOP_mux_18_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_19_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  VEC_LOOP_mux_18_nl <= MUX_v_32_2_2((vec_rsc_0_4_i_qa_d(63 DOWNTO 32)), vec_rsc_0_4_i_qa_d_bfwt_63_32,
      vec_rsc_0_4_i_bcwt_1);
  VEC_LOOP_mux_19_nl <= MUX_v_32_2_2((vec_rsc_0_4_i_qa_d(31 DOWNTO 0)), vec_rsc_0_4_i_qa_d_bfwt_31_0,
      vec_rsc_0_4_i_bcwt);
  vec_rsc_0_4_i_qa_d_mxwt <= VEC_LOOP_mux_18_nl & VEC_LOOP_mux_19_nl;
  vec_rsc_0_4_i_da_d <= vec_rsc_0_4_i_da_d_core(31 DOWNTO 0);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        vec_rsc_0_4_i_bcwt <= '0';
        vec_rsc_0_4_i_bcwt_1 <= '0';
      ELSE
        vec_rsc_0_4_i_bcwt <= NOT((NOT(vec_rsc_0_4_i_bcwt OR vec_rsc_0_4_i_biwt))
            OR vec_rsc_0_4_i_bdwt);
        vec_rsc_0_4_i_bcwt_1 <= NOT((NOT(vec_rsc_0_4_i_bcwt_1 OR vec_rsc_0_4_i_biwt_1))
            OR vec_rsc_0_4_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_0_4_i_biwt_1 = '1' ) THEN
        vec_rsc_0_4_i_qa_d_bfwt_63_32 <= vec_rsc_0_4_i_qa_d(63 DOWNTO 32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_0_4_i_biwt = '1' ) THEN
        vec_rsc_0_4_i_qa_d_bfwt_31_0 <= vec_rsc_0_4_i_qa_d(31 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_0_4_i_oswt : IN STD_LOGIC;
    vec_rsc_0_4_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_0_4_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_4_i_biwt : OUT STD_LOGIC;
    vec_rsc_0_4_i_bdwt : OUT STD_LOGIC;
    vec_rsc_0_4_i_biwt_1 : OUT STD_LOGIC;
    vec_rsc_0_4_i_bdwt_2 : OUT STD_LOGIC;
    vec_rsc_0_4_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_0_4_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_0_4_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_4_i_dswt_pff : STD_LOGIC;

  SIGNAL VEC_LOOP_and_52_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_56_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_54_nl : STD_LOGIC;
BEGIN
  vec_rsc_0_4_i_bdwt <= vec_rsc_0_4_i_oswt AND core_wen;
  vec_rsc_0_4_i_biwt <= (NOT core_wten) AND vec_rsc_0_4_i_oswt;
  vec_rsc_0_4_i_bdwt_2 <= vec_rsc_0_4_i_oswt_1 AND core_wen;
  vec_rsc_0_4_i_biwt_1 <= (NOT core_wten) AND vec_rsc_0_4_i_oswt_1;
  VEC_LOOP_and_52_nl <= (vec_rsc_0_4_i_wea_d_core_psct(0)) AND vec_rsc_0_4_i_dswt_pff;
  vec_rsc_0_4_i_wea_d_core_sct <= STD_LOGIC_VECTOR'( '0' & VEC_LOOP_and_52_nl);
  vec_rsc_0_4_i_dswt_pff <= (NOT core_wten_pff) AND vec_rsc_0_4_i_oswt_pff;
  VEC_LOOP_and_56_nl <= (NOT core_wten_pff) AND vec_rsc_0_4_i_oswt_1_pff;
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND STD_LOGIC_VECTOR'( VEC_LOOP_and_56_nl & vec_rsc_0_4_i_dswt_pff);
  VEC_LOOP_and_54_nl <= (vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0))
      AND vec_rsc_0_4_i_dswt_pff;
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= STD_LOGIC_VECTOR'( '0'
      & VEC_LOOP_and_54_nl);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_3_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_i_biwt : IN STD_LOGIC;
    vec_rsc_0_3_i_bdwt : IN STD_LOGIC;
    vec_rsc_0_3_i_biwt_1 : IN STD_LOGIC;
    vec_rsc_0_3_i_bdwt_2 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_3_i_bcwt : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_bcwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_qa_d_bfwt_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_qa_d_bfwt_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL VEC_LOOP_mux_14_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_15_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  VEC_LOOP_mux_14_nl <= MUX_v_32_2_2((vec_rsc_0_3_i_qa_d(63 DOWNTO 32)), vec_rsc_0_3_i_qa_d_bfwt_63_32,
      vec_rsc_0_3_i_bcwt_1);
  VEC_LOOP_mux_15_nl <= MUX_v_32_2_2((vec_rsc_0_3_i_qa_d(31 DOWNTO 0)), vec_rsc_0_3_i_qa_d_bfwt_31_0,
      vec_rsc_0_3_i_bcwt);
  vec_rsc_0_3_i_qa_d_mxwt <= VEC_LOOP_mux_14_nl & VEC_LOOP_mux_15_nl;
  vec_rsc_0_3_i_da_d <= vec_rsc_0_3_i_da_d_core(31 DOWNTO 0);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        vec_rsc_0_3_i_bcwt <= '0';
        vec_rsc_0_3_i_bcwt_1 <= '0';
      ELSE
        vec_rsc_0_3_i_bcwt <= NOT((NOT(vec_rsc_0_3_i_bcwt OR vec_rsc_0_3_i_biwt))
            OR vec_rsc_0_3_i_bdwt);
        vec_rsc_0_3_i_bcwt_1 <= NOT((NOT(vec_rsc_0_3_i_bcwt_1 OR vec_rsc_0_3_i_biwt_1))
            OR vec_rsc_0_3_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_0_3_i_biwt_1 = '1' ) THEN
        vec_rsc_0_3_i_qa_d_bfwt_63_32 <= vec_rsc_0_3_i_qa_d(63 DOWNTO 32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_0_3_i_biwt = '1' ) THEN
        vec_rsc_0_3_i_qa_d_bfwt_31_0 <= vec_rsc_0_3_i_qa_d(31 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_0_3_i_oswt : IN STD_LOGIC;
    vec_rsc_0_3_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_0_3_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_3_i_biwt : OUT STD_LOGIC;
    vec_rsc_0_3_i_bdwt : OUT STD_LOGIC;
    vec_rsc_0_3_i_biwt_1 : OUT STD_LOGIC;
    vec_rsc_0_3_i_bdwt_2 : OUT STD_LOGIC;
    vec_rsc_0_3_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_0_3_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_0_3_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_3_i_dswt_pff : STD_LOGIC;

  SIGNAL VEC_LOOP_and_41_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_45_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_43_nl : STD_LOGIC;
BEGIN
  vec_rsc_0_3_i_bdwt <= vec_rsc_0_3_i_oswt AND core_wen;
  vec_rsc_0_3_i_biwt <= (NOT core_wten) AND vec_rsc_0_3_i_oswt;
  vec_rsc_0_3_i_bdwt_2 <= vec_rsc_0_3_i_oswt_1 AND core_wen;
  vec_rsc_0_3_i_biwt_1 <= (NOT core_wten) AND vec_rsc_0_3_i_oswt_1;
  VEC_LOOP_and_41_nl <= (vec_rsc_0_3_i_wea_d_core_psct(0)) AND vec_rsc_0_3_i_dswt_pff;
  vec_rsc_0_3_i_wea_d_core_sct <= STD_LOGIC_VECTOR'( '0' & VEC_LOOP_and_41_nl);
  vec_rsc_0_3_i_dswt_pff <= (NOT core_wten_pff) AND vec_rsc_0_3_i_oswt_pff;
  VEC_LOOP_and_45_nl <= (NOT core_wten_pff) AND vec_rsc_0_3_i_oswt_1_pff;
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND STD_LOGIC_VECTOR'( VEC_LOOP_and_45_nl & vec_rsc_0_3_i_dswt_pff);
  VEC_LOOP_and_43_nl <= (vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0))
      AND vec_rsc_0_3_i_dswt_pff;
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= STD_LOGIC_VECTOR'( '0'
      & VEC_LOOP_and_43_nl);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_2_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_i_biwt : IN STD_LOGIC;
    vec_rsc_0_2_i_bdwt : IN STD_LOGIC;
    vec_rsc_0_2_i_biwt_1 : IN STD_LOGIC;
    vec_rsc_0_2_i_bdwt_2 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_2_i_bcwt : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_bcwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_qa_d_bfwt_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_qa_d_bfwt_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL VEC_LOOP_mux_10_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_11_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  VEC_LOOP_mux_10_nl <= MUX_v_32_2_2((vec_rsc_0_2_i_qa_d(63 DOWNTO 32)), vec_rsc_0_2_i_qa_d_bfwt_63_32,
      vec_rsc_0_2_i_bcwt_1);
  VEC_LOOP_mux_11_nl <= MUX_v_32_2_2((vec_rsc_0_2_i_qa_d(31 DOWNTO 0)), vec_rsc_0_2_i_qa_d_bfwt_31_0,
      vec_rsc_0_2_i_bcwt);
  vec_rsc_0_2_i_qa_d_mxwt <= VEC_LOOP_mux_10_nl & VEC_LOOP_mux_11_nl;
  vec_rsc_0_2_i_da_d <= vec_rsc_0_2_i_da_d_core(31 DOWNTO 0);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        vec_rsc_0_2_i_bcwt <= '0';
        vec_rsc_0_2_i_bcwt_1 <= '0';
      ELSE
        vec_rsc_0_2_i_bcwt <= NOT((NOT(vec_rsc_0_2_i_bcwt OR vec_rsc_0_2_i_biwt))
            OR vec_rsc_0_2_i_bdwt);
        vec_rsc_0_2_i_bcwt_1 <= NOT((NOT(vec_rsc_0_2_i_bcwt_1 OR vec_rsc_0_2_i_biwt_1))
            OR vec_rsc_0_2_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_0_2_i_biwt_1 = '1' ) THEN
        vec_rsc_0_2_i_qa_d_bfwt_63_32 <= vec_rsc_0_2_i_qa_d(63 DOWNTO 32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_0_2_i_biwt = '1' ) THEN
        vec_rsc_0_2_i_qa_d_bfwt_31_0 <= vec_rsc_0_2_i_qa_d(31 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_0_2_i_oswt : IN STD_LOGIC;
    vec_rsc_0_2_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_0_2_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_2_i_biwt : OUT STD_LOGIC;
    vec_rsc_0_2_i_bdwt : OUT STD_LOGIC;
    vec_rsc_0_2_i_biwt_1 : OUT STD_LOGIC;
    vec_rsc_0_2_i_bdwt_2 : OUT STD_LOGIC;
    vec_rsc_0_2_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_0_2_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_0_2_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_2_i_dswt_pff : STD_LOGIC;

  SIGNAL VEC_LOOP_and_30_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_34_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_32_nl : STD_LOGIC;
BEGIN
  vec_rsc_0_2_i_bdwt <= vec_rsc_0_2_i_oswt AND core_wen;
  vec_rsc_0_2_i_biwt <= (NOT core_wten) AND vec_rsc_0_2_i_oswt;
  vec_rsc_0_2_i_bdwt_2 <= vec_rsc_0_2_i_oswt_1 AND core_wen;
  vec_rsc_0_2_i_biwt_1 <= (NOT core_wten) AND vec_rsc_0_2_i_oswt_1;
  VEC_LOOP_and_30_nl <= (vec_rsc_0_2_i_wea_d_core_psct(0)) AND vec_rsc_0_2_i_dswt_pff;
  vec_rsc_0_2_i_wea_d_core_sct <= STD_LOGIC_VECTOR'( '0' & VEC_LOOP_and_30_nl);
  vec_rsc_0_2_i_dswt_pff <= (NOT core_wten_pff) AND vec_rsc_0_2_i_oswt_pff;
  VEC_LOOP_and_34_nl <= (NOT core_wten_pff) AND vec_rsc_0_2_i_oswt_1_pff;
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND STD_LOGIC_VECTOR'( VEC_LOOP_and_34_nl & vec_rsc_0_2_i_dswt_pff);
  VEC_LOOP_and_32_nl <= (vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0))
      AND vec_rsc_0_2_i_dswt_pff;
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= STD_LOGIC_VECTOR'( '0'
      & VEC_LOOP_and_32_nl);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_1_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_i_biwt : IN STD_LOGIC;
    vec_rsc_0_1_i_bdwt : IN STD_LOGIC;
    vec_rsc_0_1_i_biwt_1 : IN STD_LOGIC;
    vec_rsc_0_1_i_bdwt_2 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_1_i_bcwt : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_bcwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_qa_d_bfwt_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_qa_d_bfwt_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL VEC_LOOP_mux_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_7_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  VEC_LOOP_mux_6_nl <= MUX_v_32_2_2((vec_rsc_0_1_i_qa_d(63 DOWNTO 32)), vec_rsc_0_1_i_qa_d_bfwt_63_32,
      vec_rsc_0_1_i_bcwt_1);
  VEC_LOOP_mux_7_nl <= MUX_v_32_2_2((vec_rsc_0_1_i_qa_d(31 DOWNTO 0)), vec_rsc_0_1_i_qa_d_bfwt_31_0,
      vec_rsc_0_1_i_bcwt);
  vec_rsc_0_1_i_qa_d_mxwt <= VEC_LOOP_mux_6_nl & VEC_LOOP_mux_7_nl;
  vec_rsc_0_1_i_da_d <= vec_rsc_0_1_i_da_d_core(31 DOWNTO 0);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        vec_rsc_0_1_i_bcwt <= '0';
        vec_rsc_0_1_i_bcwt_1 <= '0';
      ELSE
        vec_rsc_0_1_i_bcwt <= NOT((NOT(vec_rsc_0_1_i_bcwt OR vec_rsc_0_1_i_biwt))
            OR vec_rsc_0_1_i_bdwt);
        vec_rsc_0_1_i_bcwt_1 <= NOT((NOT(vec_rsc_0_1_i_bcwt_1 OR vec_rsc_0_1_i_biwt_1))
            OR vec_rsc_0_1_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_0_1_i_biwt_1 = '1' ) THEN
        vec_rsc_0_1_i_qa_d_bfwt_63_32 <= vec_rsc_0_1_i_qa_d(63 DOWNTO 32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_0_1_i_biwt = '1' ) THEN
        vec_rsc_0_1_i_qa_d_bfwt_31_0 <= vec_rsc_0_1_i_qa_d(31 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_0_1_i_oswt : IN STD_LOGIC;
    vec_rsc_0_1_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_0_1_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_1_i_biwt : OUT STD_LOGIC;
    vec_rsc_0_1_i_bdwt : OUT STD_LOGIC;
    vec_rsc_0_1_i_biwt_1 : OUT STD_LOGIC;
    vec_rsc_0_1_i_bdwt_2 : OUT STD_LOGIC;
    vec_rsc_0_1_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_0_1_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_0_1_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_1_i_dswt_pff : STD_LOGIC;

  SIGNAL VEC_LOOP_and_19_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_23_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_21_nl : STD_LOGIC;
BEGIN
  vec_rsc_0_1_i_bdwt <= vec_rsc_0_1_i_oswt AND core_wen;
  vec_rsc_0_1_i_biwt <= (NOT core_wten) AND vec_rsc_0_1_i_oswt;
  vec_rsc_0_1_i_bdwt_2 <= vec_rsc_0_1_i_oswt_1 AND core_wen;
  vec_rsc_0_1_i_biwt_1 <= (NOT core_wten) AND vec_rsc_0_1_i_oswt_1;
  VEC_LOOP_and_19_nl <= (vec_rsc_0_1_i_wea_d_core_psct(0)) AND vec_rsc_0_1_i_dswt_pff;
  vec_rsc_0_1_i_wea_d_core_sct <= STD_LOGIC_VECTOR'( '0' & VEC_LOOP_and_19_nl);
  vec_rsc_0_1_i_dswt_pff <= (NOT core_wten_pff) AND vec_rsc_0_1_i_oswt_pff;
  VEC_LOOP_and_23_nl <= (NOT core_wten_pff) AND vec_rsc_0_1_i_oswt_1_pff;
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND STD_LOGIC_VECTOR'( VEC_LOOP_and_23_nl & vec_rsc_0_1_i_dswt_pff);
  VEC_LOOP_and_21_nl <= (vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0))
      AND vec_rsc_0_1_i_dswt_pff;
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= STD_LOGIC_VECTOR'( '0'
      & VEC_LOOP_and_21_nl);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_wait_dp IS
  PORT(
    ensig_cgo_iro : IN STD_LOGIC;
    ensig_cgo_iro_1 : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    ensig_cgo : IN STD_LOGIC;
    mult_cmp_ccs_ccore_en : OUT STD_LOGIC;
    ensig_cgo_1 : IN STD_LOGIC;
    modulo_sub_cmp_ccs_ccore_en : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_wait_dp IS
  -- Default Constants

BEGIN
  mult_cmp_ccs_ccore_en <= core_wen AND (ensig_cgo OR ensig_cgo_iro);
  modulo_sub_cmp_ccs_ccore_en <= core_wen AND (ensig_cgo_1 OR ensig_cgo_iro_1);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_0_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_biwt : IN STD_LOGIC;
    vec_rsc_0_0_i_bdwt : IN STD_LOGIC;
    vec_rsc_0_0_i_biwt_1 : IN STD_LOGIC;
    vec_rsc_0_0_i_bdwt_2 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_0_i_bcwt : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_qa_d_bfwt_63_32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_qa_d_bfwt_31_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL VEC_LOOP_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  VEC_LOOP_mux_2_nl <= MUX_v_32_2_2((vec_rsc_0_0_i_qa_d(63 DOWNTO 32)), vec_rsc_0_0_i_qa_d_bfwt_63_32,
      vec_rsc_0_0_i_bcwt_1);
  VEC_LOOP_mux_3_nl <= MUX_v_32_2_2((vec_rsc_0_0_i_qa_d(31 DOWNTO 0)), vec_rsc_0_0_i_qa_d_bfwt_31_0,
      vec_rsc_0_0_i_bcwt);
  vec_rsc_0_0_i_qa_d_mxwt <= VEC_LOOP_mux_2_nl & VEC_LOOP_mux_3_nl;
  vec_rsc_0_0_i_da_d <= vec_rsc_0_0_i_da_d_core(31 DOWNTO 0);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        vec_rsc_0_0_i_bcwt <= '0';
        vec_rsc_0_0_i_bcwt_1 <= '0';
      ELSE
        vec_rsc_0_0_i_bcwt <= NOT((NOT(vec_rsc_0_0_i_bcwt OR vec_rsc_0_0_i_biwt))
            OR vec_rsc_0_0_i_bdwt);
        vec_rsc_0_0_i_bcwt_1 <= NOT((NOT(vec_rsc_0_0_i_bcwt_1 OR vec_rsc_0_0_i_biwt_1))
            OR vec_rsc_0_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_0_0_i_biwt_1 = '1' ) THEN
        vec_rsc_0_0_i_qa_d_bfwt_63_32 <= vec_rsc_0_0_i_qa_d(63 DOWNTO 32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( vec_rsc_0_0_i_biwt = '1' ) THEN
        vec_rsc_0_0_i_qa_d_bfwt_31_0 <= vec_rsc_0_0_i_qa_d(31 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_0_0_i_oswt : IN STD_LOGIC;
    vec_rsc_0_0_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_0_0_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_0_i_biwt : OUT STD_LOGIC;
    vec_rsc_0_0_i_bdwt : OUT STD_LOGIC;
    vec_rsc_0_0_i_biwt_1 : OUT STD_LOGIC;
    vec_rsc_0_0_i_bdwt_2 : OUT STD_LOGIC;
    vec_rsc_0_0_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_0_0_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_0_0_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_0_i_dswt_pff : STD_LOGIC;

  SIGNAL VEC_LOOP_and_8_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_12_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_and_10_nl : STD_LOGIC;
BEGIN
  vec_rsc_0_0_i_bdwt <= vec_rsc_0_0_i_oswt AND core_wen;
  vec_rsc_0_0_i_biwt <= (NOT core_wten) AND vec_rsc_0_0_i_oswt;
  vec_rsc_0_0_i_bdwt_2 <= vec_rsc_0_0_i_oswt_1 AND core_wen;
  vec_rsc_0_0_i_biwt_1 <= (NOT core_wten) AND vec_rsc_0_0_i_oswt_1;
  VEC_LOOP_and_8_nl <= (vec_rsc_0_0_i_wea_d_core_psct(0)) AND vec_rsc_0_0_i_dswt_pff;
  vec_rsc_0_0_i_wea_d_core_sct <= STD_LOGIC_VECTOR'( '0' & VEC_LOOP_and_8_nl);
  vec_rsc_0_0_i_dswt_pff <= (NOT core_wten_pff) AND vec_rsc_0_0_i_oswt_pff;
  VEC_LOOP_and_12_nl <= (NOT core_wten_pff) AND vec_rsc_0_0_i_oswt_1_pff;
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND STD_LOGIC_VECTOR'( VEC_LOOP_and_12_nl & vec_rsc_0_0_i_dswt_pff);
  VEC_LOOP_and_10_nl <= (vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0))
      AND vec_rsc_0_0_i_dswt_pff;
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= STD_LOGIC_VECTOR'( '0'
      & VEC_LOOP_and_10_nl);
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_complete_rsci_complete_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_complete_rsci_complete_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    complete_rsci_oswt : IN STD_LOGIC;
    complete_rsci_wen_comp : OUT STD_LOGIC;
    complete_rsci_biwt : IN STD_LOGIC;
    complete_rsci_bdwt : IN STD_LOGIC;
    complete_rsci_bcwt : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_complete_rsci_complete_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_complete_rsci_complete_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL complete_rsci_bcwt_drv : STD_LOGIC;

BEGIN
  -- Output Reader Assignments
  complete_rsci_bcwt <= complete_rsci_bcwt_drv;

  complete_rsci_wen_comp <= (NOT complete_rsci_oswt) OR complete_rsci_biwt OR complete_rsci_bcwt_drv;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        complete_rsci_bcwt_drv <= '0';
      ELSE
        complete_rsci_bcwt_drv <= NOT((NOT(complete_rsci_bcwt_drv OR complete_rsci_biwt))
            OR complete_rsci_bdwt);
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_complete_rsci_complete_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_complete_rsci_complete_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    complete_rsci_oswt : IN STD_LOGIC;
    complete_rsci_biwt : OUT STD_LOGIC;
    complete_rsci_bdwt : OUT STD_LOGIC;
    complete_rsci_bcwt : IN STD_LOGIC;
    complete_rsci_ivld_core_sct : OUT STD_LOGIC;
    complete_rsci_irdy : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_complete_rsci_complete_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_complete_rsci_complete_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL complete_rsci_ogwt : STD_LOGIC;

BEGIN
  complete_rsci_bdwt <= complete_rsci_oswt AND core_wen;
  complete_rsci_biwt <= complete_rsci_ogwt AND complete_rsci_irdy;
  complete_rsci_ogwt <= complete_rsci_oswt AND (NOT complete_rsci_bcwt);
  complete_rsci_ivld_core_sct <= complete_rsci_ogwt;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_run_rsci_run_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_run_rsci_run_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    run_rsci_ivld_mxwt : OUT STD_LOGIC;
    run_rsci_ivld : IN STD_LOGIC;
    run_rsci_biwt : IN STD_LOGIC;
    run_rsci_bdwt : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_run_rsci_run_wait_dp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_run_rsci_run_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL run_rsci_bcwt : STD_LOGIC;
  SIGNAL run_rsci_ivld_bfwt : STD_LOGIC;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  run_rsci_ivld_mxwt <= MUX_s_1_2_2(run_rsci_ivld, run_rsci_ivld_bfwt, run_rsci_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        run_rsci_bcwt <= '0';
      ELSE
        run_rsci_bcwt <= NOT((NOT(run_rsci_bcwt OR run_rsci_biwt)) OR run_rsci_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( run_rsci_biwt = '1' ) THEN
        run_rsci_ivld_bfwt <= run_rsci_ivld;
      END IF;
    END IF;
  END PROCESS;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_run_rsci_run_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_run_rsci_run_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    run_rsci_oswt : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    run_rsci_biwt : OUT STD_LOGIC;
    run_rsci_bdwt : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_run_rsci_run_wait_ctrl;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_run_rsci_run_wait_ctrl IS
  -- Default Constants

BEGIN
  run_rsci_bdwt <= run_rsci_oswt AND core_wen;
  run_rsci_biwt <= (NOT core_wten) AND run_rsci_oswt;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_0_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_0_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_0_obj_twiddle_h_rsc_triosy_0_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_0_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_0_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_0_obj_twiddle_h_rsc_triosy_0_0_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_0_obj_twiddle_h_rsc_triosy_0_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_0_obj_iswt0 => twiddle_h_rsc_triosy_0_0_obj_iswt0,
      twiddle_h_rsc_triosy_0_0_obj_ld_core_sct => twiddle_h_rsc_triosy_0_0_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_1_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_1_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_1_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_1_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_1_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_1_obj_twiddle_h_rsc_triosy_0_1_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_1_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_1_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_1_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_1_obj_twiddle_h_rsc_triosy_0_1_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_1_obj_twiddle_h_rsc_triosy_0_1_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_1_obj_iswt0 => twiddle_h_rsc_triosy_0_1_obj_iswt0,
      twiddle_h_rsc_triosy_0_1_obj_ld_core_sct => twiddle_h_rsc_triosy_0_1_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_2_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_2_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_2_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_2_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_2_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_2_obj_twiddle_h_rsc_triosy_0_2_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_2_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_2_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_2_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_2_obj_twiddle_h_rsc_triosy_0_2_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_2_obj_twiddle_h_rsc_triosy_0_2_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_2_obj_iswt0 => twiddle_h_rsc_triosy_0_2_obj_iswt0,
      twiddle_h_rsc_triosy_0_2_obj_ld_core_sct => twiddle_h_rsc_triosy_0_2_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_3_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_3_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_3_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_3_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_3_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_3_obj_twiddle_h_rsc_triosy_0_3_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_3_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_3_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_3_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_3_obj_twiddle_h_rsc_triosy_0_3_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_3_obj_twiddle_h_rsc_triosy_0_3_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_3_obj_iswt0 => twiddle_h_rsc_triosy_0_3_obj_iswt0,
      twiddle_h_rsc_triosy_0_3_obj_ld_core_sct => twiddle_h_rsc_triosy_0_3_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_4_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_4_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_4_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_4_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_4_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_4_obj_twiddle_h_rsc_triosy_0_4_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_4_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_4_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_4_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_4_obj_twiddle_h_rsc_triosy_0_4_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_4_obj_twiddle_h_rsc_triosy_0_4_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_4_obj_iswt0 => twiddle_h_rsc_triosy_0_4_obj_iswt0,
      twiddle_h_rsc_triosy_0_4_obj_ld_core_sct => twiddle_h_rsc_triosy_0_4_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_5_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_5_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_5_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_5_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_5_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_5_obj_twiddle_h_rsc_triosy_0_5_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_5_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_5_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_5_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_5_obj_twiddle_h_rsc_triosy_0_5_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_5_obj_twiddle_h_rsc_triosy_0_5_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_5_obj_iswt0 => twiddle_h_rsc_triosy_0_5_obj_iswt0,
      twiddle_h_rsc_triosy_0_5_obj_ld_core_sct => twiddle_h_rsc_triosy_0_5_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_6_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_6_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_6_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_6_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_6_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_6_obj_twiddle_h_rsc_triosy_0_6_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_6_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_6_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_6_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_6_obj_twiddle_h_rsc_triosy_0_6_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_6_obj_twiddle_h_rsc_triosy_0_6_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_6_obj_iswt0 => twiddle_h_rsc_triosy_0_6_obj_iswt0,
      twiddle_h_rsc_triosy_0_6_obj_ld_core_sct => twiddle_h_rsc_triosy_0_6_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_7_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_7_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_7_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_7_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_7_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_7_obj_twiddle_h_rsc_triosy_0_7_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_7_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_7_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_7_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_7_obj_twiddle_h_rsc_triosy_0_7_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_7_obj_twiddle_h_rsc_triosy_0_7_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_7_obj_iswt0 => twiddle_h_rsc_triosy_0_7_obj_iswt0,
      twiddle_h_rsc_triosy_0_7_obj_ld_core_sct => twiddle_h_rsc_triosy_0_7_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_0_obj IS
  PORT(
    twiddle_h_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_0_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_1_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_0_obj_twiddle_h_rsc_triosy_1_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_1_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_1_0_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_1_0_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_0_obj_twiddle_h_rsc_triosy_1_0_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_0_obj_twiddle_h_rsc_triosy_1_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_1_0_obj_iswt0 => twiddle_h_rsc_triosy_1_0_obj_iswt0,
      twiddle_h_rsc_triosy_1_0_obj_ld_core_sct => twiddle_h_rsc_triosy_1_0_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_1_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_1_obj IS
  PORT(
    twiddle_h_rsc_triosy_1_1_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_1_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_1_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_1_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_1_1_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_1_obj_twiddle_h_rsc_triosy_1_1_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_1_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_1_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_1_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_1_1_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_1_1_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_1_obj_twiddle_h_rsc_triosy_1_1_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_1_obj_twiddle_h_rsc_triosy_1_1_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_1_1_obj_iswt0 => twiddle_h_rsc_triosy_1_1_obj_iswt0,
      twiddle_h_rsc_triosy_1_1_obj_ld_core_sct => twiddle_h_rsc_triosy_1_1_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_2_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_2_obj IS
  PORT(
    twiddle_h_rsc_triosy_1_2_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_2_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_2_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_2_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_1_2_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_2_obj_twiddle_h_rsc_triosy_1_2_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_2_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_2_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_1_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_1_2_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_1_2_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_2_obj_twiddle_h_rsc_triosy_1_2_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_2_obj_twiddle_h_rsc_triosy_1_2_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_1_2_obj_iswt0 => twiddle_h_rsc_triosy_1_2_obj_iswt0,
      twiddle_h_rsc_triosy_1_2_obj_ld_core_sct => twiddle_h_rsc_triosy_1_2_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_3_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_3_obj IS
  PORT(
    twiddle_h_rsc_triosy_1_3_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_3_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_3_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_3_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_1_3_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_3_obj_twiddle_h_rsc_triosy_1_3_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_3_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_3_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_1_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_1_3_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_1_3_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_3_obj_twiddle_h_rsc_triosy_1_3_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_3_obj_twiddle_h_rsc_triosy_1_3_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_1_3_obj_iswt0 => twiddle_h_rsc_triosy_1_3_obj_iswt0,
      twiddle_h_rsc_triosy_1_3_obj_ld_core_sct => twiddle_h_rsc_triosy_1_3_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_4_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_4_obj IS
  PORT(
    twiddle_h_rsc_triosy_1_4_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_4_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_4_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_4_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_1_4_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_4_obj_twiddle_h_rsc_triosy_1_4_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_4_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_4_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_1_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_1_4_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_1_4_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_4_obj_twiddle_h_rsc_triosy_1_4_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_4_obj_twiddle_h_rsc_triosy_1_4_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_1_4_obj_iswt0 => twiddle_h_rsc_triosy_1_4_obj_iswt0,
      twiddle_h_rsc_triosy_1_4_obj_ld_core_sct => twiddle_h_rsc_triosy_1_4_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_5_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_5_obj IS
  PORT(
    twiddle_h_rsc_triosy_1_5_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_5_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_5_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_5_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_1_5_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_5_obj_twiddle_h_rsc_triosy_1_5_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_5_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_5_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_1_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_1_5_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_1_5_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_5_obj_twiddle_h_rsc_triosy_1_5_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_5_obj_twiddle_h_rsc_triosy_1_5_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_1_5_obj_iswt0 => twiddle_h_rsc_triosy_1_5_obj_iswt0,
      twiddle_h_rsc_triosy_1_5_obj_ld_core_sct => twiddle_h_rsc_triosy_1_5_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_6_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_6_obj IS
  PORT(
    twiddle_h_rsc_triosy_1_6_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_6_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_6_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_6_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_1_6_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_6_obj_twiddle_h_rsc_triosy_1_6_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_6_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_6_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_1_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_1_6_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_1_6_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_6_obj_twiddle_h_rsc_triosy_1_6_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_6_obj_twiddle_h_rsc_triosy_1_6_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_1_6_obj_iswt0 => twiddle_h_rsc_triosy_1_6_obj_iswt0,
      twiddle_h_rsc_triosy_1_6_obj_ld_core_sct => twiddle_h_rsc_triosy_1_6_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_7_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_7_obj IS
  PORT(
    twiddle_h_rsc_triosy_1_7_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_1_7_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_7_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_7_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_1_7_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_7_obj_twiddle_h_rsc_triosy_1_7_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_7_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_7_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_1_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_1_7_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_1_7_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_7_obj_twiddle_h_rsc_triosy_1_7_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_7_obj_twiddle_h_rsc_triosy_1_7_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_1_7_obj_iswt0 => twiddle_h_rsc_triosy_1_7_obj_iswt0,
      twiddle_h_rsc_triosy_1_7_obj_ld_core_sct => twiddle_h_rsc_triosy_1_7_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_0_obj IS
  PORT(
    twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_0_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_0_obj_twiddle_rsc_triosy_0_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_0_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_0_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_0_obj_twiddle_rsc_triosy_0_0_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_0_obj_twiddle_rsc_triosy_0_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_0_obj_iswt0 => twiddle_rsc_triosy_0_0_obj_iswt0,
      twiddle_rsc_triosy_0_0_obj_ld_core_sct => twiddle_rsc_triosy_0_0_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_1_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_1_obj IS
  PORT(
    twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_1_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_1_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_1_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_1_obj_twiddle_rsc_triosy_0_1_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_1_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_1_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_1_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_1_obj_twiddle_rsc_triosy_0_1_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_1_obj_twiddle_rsc_triosy_0_1_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_1_obj_iswt0 => twiddle_rsc_triosy_0_1_obj_iswt0,
      twiddle_rsc_triosy_0_1_obj_ld_core_sct => twiddle_rsc_triosy_0_1_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_2_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_2_obj IS
  PORT(
    twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_2_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_2_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_2_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_2_obj_twiddle_rsc_triosy_0_2_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_2_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_2_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_2_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_2_obj_twiddle_rsc_triosy_0_2_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_2_obj_twiddle_rsc_triosy_0_2_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_2_obj_iswt0 => twiddle_rsc_triosy_0_2_obj_iswt0,
      twiddle_rsc_triosy_0_2_obj_ld_core_sct => twiddle_rsc_triosy_0_2_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_3_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_3_obj IS
  PORT(
    twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_3_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_3_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_3_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_3_obj_twiddle_rsc_triosy_0_3_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_3_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_3_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_3_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_3_obj_twiddle_rsc_triosy_0_3_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_3_obj_twiddle_rsc_triosy_0_3_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_3_obj_iswt0 => twiddle_rsc_triosy_0_3_obj_iswt0,
      twiddle_rsc_triosy_0_3_obj_ld_core_sct => twiddle_rsc_triosy_0_3_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_4_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_4_obj IS
  PORT(
    twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_4_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_4_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_4_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_4_obj_twiddle_rsc_triosy_0_4_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_4_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_4_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_4_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_4_obj_twiddle_rsc_triosy_0_4_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_4_obj_twiddle_rsc_triosy_0_4_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_4_obj_iswt0 => twiddle_rsc_triosy_0_4_obj_iswt0,
      twiddle_rsc_triosy_0_4_obj_ld_core_sct => twiddle_rsc_triosy_0_4_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_5_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_5_obj IS
  PORT(
    twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_5_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_5_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_5_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_5_obj_twiddle_rsc_triosy_0_5_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_5_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_5_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_5_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_5_obj_twiddle_rsc_triosy_0_5_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_5_obj_twiddle_rsc_triosy_0_5_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_5_obj_iswt0 => twiddle_rsc_triosy_0_5_obj_iswt0,
      twiddle_rsc_triosy_0_5_obj_ld_core_sct => twiddle_rsc_triosy_0_5_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_6_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_6_obj IS
  PORT(
    twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_6_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_6_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_6_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_6_obj_twiddle_rsc_triosy_0_6_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_6_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_6_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_6_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_6_obj_twiddle_rsc_triosy_0_6_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_6_obj_twiddle_rsc_triosy_0_6_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_6_obj_iswt0 => twiddle_rsc_triosy_0_6_obj_iswt0,
      twiddle_rsc_triosy_0_6_obj_ld_core_sct => twiddle_rsc_triosy_0_6_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_7_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_7_obj IS
  PORT(
    twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_7_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_7_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_7_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_7_obj_twiddle_rsc_triosy_0_7_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_7_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_7_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_7_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_7_obj_twiddle_rsc_triosy_0_7_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_7_obj_twiddle_rsc_triosy_0_7_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_7_obj_iswt0 => twiddle_rsc_triosy_0_7_obj_iswt0,
      twiddle_rsc_triosy_0_7_obj_ld_core_sct => twiddle_rsc_triosy_0_7_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_0_obj IS
  PORT(
    twiddle_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_0_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_1_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_0_obj_twiddle_rsc_triosy_1_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_1_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_1_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_1_0_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_1_0_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_0_obj_twiddle_rsc_triosy_1_0_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_0_obj_twiddle_rsc_triosy_1_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_1_0_obj_iswt0 => twiddle_rsc_triosy_1_0_obj_iswt0,
      twiddle_rsc_triosy_1_0_obj_ld_core_sct => twiddle_rsc_triosy_1_0_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_1_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_1_obj IS
  PORT(
    twiddle_rsc_triosy_1_1_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_1_1_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_1_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_1_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_1_1_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_1_obj_twiddle_rsc_triosy_1_1_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_1_1_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_1_1_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_1_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_1_1_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_1_1_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_1_obj_twiddle_rsc_triosy_1_1_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_1_obj_twiddle_rsc_triosy_1_1_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_1_1_obj_iswt0 => twiddle_rsc_triosy_1_1_obj_iswt0,
      twiddle_rsc_triosy_1_1_obj_ld_core_sct => twiddle_rsc_triosy_1_1_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_2_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_2_obj IS
  PORT(
    twiddle_rsc_triosy_1_2_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_1_2_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_2_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_2_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_1_2_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_2_obj_twiddle_rsc_triosy_1_2_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_1_2_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_1_2_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_1_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_1_2_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_1_2_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_2_obj_twiddle_rsc_triosy_1_2_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_2_obj_twiddle_rsc_triosy_1_2_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_1_2_obj_iswt0 => twiddle_rsc_triosy_1_2_obj_iswt0,
      twiddle_rsc_triosy_1_2_obj_ld_core_sct => twiddle_rsc_triosy_1_2_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_3_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_3_obj IS
  PORT(
    twiddle_rsc_triosy_1_3_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_1_3_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_3_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_3_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_1_3_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_3_obj_twiddle_rsc_triosy_1_3_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_1_3_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_1_3_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_1_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_1_3_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_1_3_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_3_obj_twiddle_rsc_triosy_1_3_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_3_obj_twiddle_rsc_triosy_1_3_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_1_3_obj_iswt0 => twiddle_rsc_triosy_1_3_obj_iswt0,
      twiddle_rsc_triosy_1_3_obj_ld_core_sct => twiddle_rsc_triosy_1_3_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_4_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_4_obj IS
  PORT(
    twiddle_rsc_triosy_1_4_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_1_4_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_4_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_4_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_1_4_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_4_obj_twiddle_rsc_triosy_1_4_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_1_4_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_1_4_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_1_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_1_4_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_1_4_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_4_obj_twiddle_rsc_triosy_1_4_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_4_obj_twiddle_rsc_triosy_1_4_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_1_4_obj_iswt0 => twiddle_rsc_triosy_1_4_obj_iswt0,
      twiddle_rsc_triosy_1_4_obj_ld_core_sct => twiddle_rsc_triosy_1_4_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_5_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_5_obj IS
  PORT(
    twiddle_rsc_triosy_1_5_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_1_5_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_5_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_5_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_1_5_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_5_obj_twiddle_rsc_triosy_1_5_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_1_5_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_1_5_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_1_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_1_5_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_1_5_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_5_obj_twiddle_rsc_triosy_1_5_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_5_obj_twiddle_rsc_triosy_1_5_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_1_5_obj_iswt0 => twiddle_rsc_triosy_1_5_obj_iswt0,
      twiddle_rsc_triosy_1_5_obj_ld_core_sct => twiddle_rsc_triosy_1_5_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_6_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_6_obj IS
  PORT(
    twiddle_rsc_triosy_1_6_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_1_6_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_6_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_6_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_1_6_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_6_obj_twiddle_rsc_triosy_1_6_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_1_6_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_1_6_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_1_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_1_6_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_1_6_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_6_obj_twiddle_rsc_triosy_1_6_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_6_obj_twiddle_rsc_triosy_1_6_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_1_6_obj_iswt0 => twiddle_rsc_triosy_1_6_obj_iswt0,
      twiddle_rsc_triosy_1_6_obj_ld_core_sct => twiddle_rsc_triosy_1_6_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_7_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_7_obj IS
  PORT(
    twiddle_rsc_triosy_1_7_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_1_7_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_7_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_7_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_1_7_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_7_obj_twiddle_rsc_triosy_1_7_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_1_7_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_1_7_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_1_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_1_7_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_1_7_lz
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_7_obj_twiddle_rsc_triosy_1_7_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_7_obj_twiddle_rsc_triosy_1_7_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_1_7_obj_iswt0 => twiddle_rsc_triosy_1_7_obj_iswt0,
      twiddle_rsc_triosy_1_7_obj_ld_core_sct => twiddle_rsc_triosy_1_7_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_r_rsc_triosy_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_r_rsc_triosy_obj IS
  PORT(
    r_rsc_triosy_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    r_rsc_triosy_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_r_rsc_triosy_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_r_rsc_triosy_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL r_rsc_triosy_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_r_rsc_triosy_obj_r_rsc_triosy_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      r_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
      r_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  r_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => r_rsc_triosy_obj_ld_core_sct,
      lz => r_rsc_triosy_lz
    );
  inPlaceNTT_DIF_precomp_core_r_rsc_triosy_obj_r_rsc_triosy_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_r_rsc_triosy_obj_r_rsc_triosy_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      r_rsc_triosy_obj_iswt0 => r_rsc_triosy_obj_iswt0,
      r_rsc_triosy_obj_ld_core_sct => r_rsc_triosy_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_p_rsc_triosy_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_p_rsc_triosy_obj IS
  PORT(
    p_rsc_triosy_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    p_rsc_triosy_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_p_rsc_triosy_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_p_rsc_triosy_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL p_rsc_triosy_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_p_rsc_triosy_obj_p_rsc_triosy_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      p_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
      p_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  p_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => p_rsc_triosy_obj_ld_core_sct,
      lz => p_rsc_triosy_lz
    );
  inPlaceNTT_DIF_precomp_core_p_rsc_triosy_obj_p_rsc_triosy_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_p_rsc_triosy_obj_p_rsc_triosy_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      p_rsc_triosy_obj_iswt0 => p_rsc_triosy_obj_iswt0,
      p_rsc_triosy_obj_ld_core_sct => p_rsc_triosy_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_0_obj IS
  PORT(
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_0_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_triosy_0_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_0_obj_vec_rsc_triosy_0_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC;
      vec_rsc_triosy_0_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  vec_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => vec_rsc_triosy_0_0_obj_ld_core_sct,
      lz => vec_rsc_triosy_0_0_lz
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_0_obj_vec_rsc_triosy_0_0_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_0_obj_vec_rsc_triosy_0_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      vec_rsc_triosy_0_0_obj_iswt0 => vec_rsc_triosy_0_0_obj_iswt0,
      vec_rsc_triosy_0_0_obj_ld_core_sct => vec_rsc_triosy_0_0_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_1_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_1_obj IS
  PORT(
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_1_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_1_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_triosy_0_1_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_1_obj_vec_rsc_triosy_0_1_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC;
      vec_rsc_triosy_0_1_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  vec_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => vec_rsc_triosy_0_1_obj_ld_core_sct,
      lz => vec_rsc_triosy_0_1_lz
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_1_obj_vec_rsc_triosy_0_1_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_1_obj_vec_rsc_triosy_0_1_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      vec_rsc_triosy_0_1_obj_iswt0 => vec_rsc_triosy_0_1_obj_iswt0,
      vec_rsc_triosy_0_1_obj_ld_core_sct => vec_rsc_triosy_0_1_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_2_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_2_obj IS
  PORT(
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_2_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_2_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_triosy_0_2_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_2_obj_vec_rsc_triosy_0_2_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC;
      vec_rsc_triosy_0_2_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  vec_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => vec_rsc_triosy_0_2_obj_ld_core_sct,
      lz => vec_rsc_triosy_0_2_lz
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_2_obj_vec_rsc_triosy_0_2_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_2_obj_vec_rsc_triosy_0_2_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      vec_rsc_triosy_0_2_obj_iswt0 => vec_rsc_triosy_0_2_obj_iswt0,
      vec_rsc_triosy_0_2_obj_ld_core_sct => vec_rsc_triosy_0_2_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_3_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_3_obj IS
  PORT(
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_3_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_3_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_triosy_0_3_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_3_obj_vec_rsc_triosy_0_3_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC;
      vec_rsc_triosy_0_3_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  vec_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => vec_rsc_triosy_0_3_obj_ld_core_sct,
      lz => vec_rsc_triosy_0_3_lz
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_3_obj_vec_rsc_triosy_0_3_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_3_obj_vec_rsc_triosy_0_3_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      vec_rsc_triosy_0_3_obj_iswt0 => vec_rsc_triosy_0_3_obj_iswt0,
      vec_rsc_triosy_0_3_obj_ld_core_sct => vec_rsc_triosy_0_3_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_4_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_4_obj IS
  PORT(
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_4_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_4_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_triosy_0_4_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_4_obj_vec_rsc_triosy_0_4_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC;
      vec_rsc_triosy_0_4_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  vec_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => vec_rsc_triosy_0_4_obj_ld_core_sct,
      lz => vec_rsc_triosy_0_4_lz
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_4_obj_vec_rsc_triosy_0_4_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_4_obj_vec_rsc_triosy_0_4_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      vec_rsc_triosy_0_4_obj_iswt0 => vec_rsc_triosy_0_4_obj_iswt0,
      vec_rsc_triosy_0_4_obj_ld_core_sct => vec_rsc_triosy_0_4_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_5_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_5_obj IS
  PORT(
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_5_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_5_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_triosy_0_5_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_5_obj_vec_rsc_triosy_0_5_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC;
      vec_rsc_triosy_0_5_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  vec_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => vec_rsc_triosy_0_5_obj_ld_core_sct,
      lz => vec_rsc_triosy_0_5_lz
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_5_obj_vec_rsc_triosy_0_5_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_5_obj_vec_rsc_triosy_0_5_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      vec_rsc_triosy_0_5_obj_iswt0 => vec_rsc_triosy_0_5_obj_iswt0,
      vec_rsc_triosy_0_5_obj_ld_core_sct => vec_rsc_triosy_0_5_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_6_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_6_obj IS
  PORT(
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_6_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_6_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_triosy_0_6_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_6_obj_vec_rsc_triosy_0_6_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC;
      vec_rsc_triosy_0_6_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  vec_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => vec_rsc_triosy_0_6_obj_ld_core_sct,
      lz => vec_rsc_triosy_0_6_lz
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_6_obj_vec_rsc_triosy_0_6_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_6_obj_vec_rsc_triosy_0_6_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      vec_rsc_triosy_0_6_obj_iswt0 => vec_rsc_triosy_0_6_obj_iswt0,
      vec_rsc_triosy_0_6_obj_ld_core_sct => vec_rsc_triosy_0_6_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_7_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_7_obj IS
  PORT(
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_7_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_7_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_triosy_0_7_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_7_obj_vec_rsc_triosy_0_7_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC;
      vec_rsc_triosy_0_7_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  vec_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => vec_rsc_triosy_0_7_obj_ld_core_sct,
      lz => vec_rsc_triosy_0_7_lz
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_7_obj_vec_rsc_triosy_0_7_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_7_obj_vec_rsc_triosy_0_7_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      vec_rsc_triosy_0_7_obj_iswt0 => vec_rsc_triosy_0_7_obj_iswt0,
      vec_rsc_triosy_0_7_obj_ld_core_sct => vec_rsc_triosy_0_7_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_0_obj IS
  PORT(
    vec_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_0_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_triosy_1_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_0_obj_vec_rsc_triosy_1_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC;
      vec_rsc_triosy_1_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  vec_rsc_triosy_1_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => vec_rsc_triosy_1_0_obj_ld_core_sct,
      lz => vec_rsc_triosy_1_0_lz
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_0_obj_vec_rsc_triosy_1_0_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_0_obj_vec_rsc_triosy_1_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      vec_rsc_triosy_1_0_obj_iswt0 => vec_rsc_triosy_1_0_obj_iswt0,
      vec_rsc_triosy_1_0_obj_ld_core_sct => vec_rsc_triosy_1_0_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_1_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_1_obj IS
  PORT(
    vec_rsc_triosy_1_1_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_1_1_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_1_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_1_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_triosy_1_1_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_1_obj_vec_rsc_triosy_1_1_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_1_1_obj_iswt0 : IN STD_LOGIC;
      vec_rsc_triosy_1_1_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  vec_rsc_triosy_1_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => vec_rsc_triosy_1_1_obj_ld_core_sct,
      lz => vec_rsc_triosy_1_1_lz
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_1_obj_vec_rsc_triosy_1_1_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_1_obj_vec_rsc_triosy_1_1_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      vec_rsc_triosy_1_1_obj_iswt0 => vec_rsc_triosy_1_1_obj_iswt0,
      vec_rsc_triosy_1_1_obj_ld_core_sct => vec_rsc_triosy_1_1_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_2_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_2_obj IS
  PORT(
    vec_rsc_triosy_1_2_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_1_2_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_2_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_2_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_triosy_1_2_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_2_obj_vec_rsc_triosy_1_2_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_1_2_obj_iswt0 : IN STD_LOGIC;
      vec_rsc_triosy_1_2_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  vec_rsc_triosy_1_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => vec_rsc_triosy_1_2_obj_ld_core_sct,
      lz => vec_rsc_triosy_1_2_lz
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_2_obj_vec_rsc_triosy_1_2_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_2_obj_vec_rsc_triosy_1_2_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      vec_rsc_triosy_1_2_obj_iswt0 => vec_rsc_triosy_1_2_obj_iswt0,
      vec_rsc_triosy_1_2_obj_ld_core_sct => vec_rsc_triosy_1_2_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_3_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_3_obj IS
  PORT(
    vec_rsc_triosy_1_3_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_1_3_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_3_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_3_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_triosy_1_3_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_3_obj_vec_rsc_triosy_1_3_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_1_3_obj_iswt0 : IN STD_LOGIC;
      vec_rsc_triosy_1_3_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  vec_rsc_triosy_1_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => vec_rsc_triosy_1_3_obj_ld_core_sct,
      lz => vec_rsc_triosy_1_3_lz
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_3_obj_vec_rsc_triosy_1_3_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_3_obj_vec_rsc_triosy_1_3_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      vec_rsc_triosy_1_3_obj_iswt0 => vec_rsc_triosy_1_3_obj_iswt0,
      vec_rsc_triosy_1_3_obj_ld_core_sct => vec_rsc_triosy_1_3_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_4_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_4_obj IS
  PORT(
    vec_rsc_triosy_1_4_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_1_4_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_4_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_4_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_triosy_1_4_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_4_obj_vec_rsc_triosy_1_4_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_1_4_obj_iswt0 : IN STD_LOGIC;
      vec_rsc_triosy_1_4_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  vec_rsc_triosy_1_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => vec_rsc_triosy_1_4_obj_ld_core_sct,
      lz => vec_rsc_triosy_1_4_lz
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_4_obj_vec_rsc_triosy_1_4_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_4_obj_vec_rsc_triosy_1_4_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      vec_rsc_triosy_1_4_obj_iswt0 => vec_rsc_triosy_1_4_obj_iswt0,
      vec_rsc_triosy_1_4_obj_ld_core_sct => vec_rsc_triosy_1_4_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_5_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_5_obj IS
  PORT(
    vec_rsc_triosy_1_5_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_1_5_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_5_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_5_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_triosy_1_5_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_5_obj_vec_rsc_triosy_1_5_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_1_5_obj_iswt0 : IN STD_LOGIC;
      vec_rsc_triosy_1_5_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  vec_rsc_triosy_1_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => vec_rsc_triosy_1_5_obj_ld_core_sct,
      lz => vec_rsc_triosy_1_5_lz
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_5_obj_vec_rsc_triosy_1_5_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_5_obj_vec_rsc_triosy_1_5_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      vec_rsc_triosy_1_5_obj_iswt0 => vec_rsc_triosy_1_5_obj_iswt0,
      vec_rsc_triosy_1_5_obj_ld_core_sct => vec_rsc_triosy_1_5_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_6_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_6_obj IS
  PORT(
    vec_rsc_triosy_1_6_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_1_6_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_6_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_6_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_triosy_1_6_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_6_obj_vec_rsc_triosy_1_6_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_1_6_obj_iswt0 : IN STD_LOGIC;
      vec_rsc_triosy_1_6_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  vec_rsc_triosy_1_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => vec_rsc_triosy_1_6_obj_ld_core_sct,
      lz => vec_rsc_triosy_1_6_lz
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_6_obj_vec_rsc_triosy_1_6_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_6_obj_vec_rsc_triosy_1_6_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      vec_rsc_triosy_1_6_obj_iswt0 => vec_rsc_triosy_1_6_obj_iswt0,
      vec_rsc_triosy_1_6_obj_ld_core_sct => vec_rsc_triosy_1_6_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_7_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_7_obj IS
  PORT(
    vec_rsc_triosy_1_7_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_triosy_1_7_obj_iswt0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_7_obj;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_7_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_triosy_1_7_obj_ld_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_7_obj_vec_rsc_triosy_1_7_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_1_7_obj_iswt0 : IN STD_LOGIC;
      vec_rsc_triosy_1_7_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  vec_rsc_triosy_1_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => vec_rsc_triosy_1_7_obj_ld_core_sct,
      lz => vec_rsc_triosy_1_7_lz
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_7_obj_vec_rsc_triosy_1_7_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_7_obj_vec_rsc_triosy_1_7_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      vec_rsc_triosy_1_7_obj_iswt0 => vec_rsc_triosy_1_7_obj_iswt0,
      vec_rsc_triosy_1_7_obj_ld_core_sct => vec_rsc_triosy_1_7_obj_ld_core_sct
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_1_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_1_7_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_1_7_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_7_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_1_7_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_7_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_1_7_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_1_7_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_1_7_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_1_7_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_1_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_7_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_7_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_1_7_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_dp_inst_twiddle_h_rsc_1_7_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_dp_inst_twiddle_h_rsc_1_7_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsc_1_7_i_oswt => twiddle_h_rsc_1_7_i_oswt,
      twiddle_h_rsc_1_7_i_biwt => twiddle_h_rsc_1_7_i_biwt,
      twiddle_h_rsc_1_7_i_bdwt => twiddle_h_rsc_1_7_i_bdwt,
      twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_h_rsc_1_7_i_oswt_pff => twiddle_h_rsc_1_7_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_dp_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_1_7_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_dp_inst_twiddle_h_rsc_1_7_i_qb_d,
      twiddle_h_rsc_1_7_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_dp_inst_twiddle_h_rsc_1_7_i_qb_d_mxwt,
      twiddle_h_rsc_1_7_i_biwt => twiddle_h_rsc_1_7_i_biwt,
      twiddle_h_rsc_1_7_i_bdwt => twiddle_h_rsc_1_7_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_dp_inst_twiddle_h_rsc_1_7_i_qb_d
      <= twiddle_h_rsc_1_7_i_qb_d;
  twiddle_h_rsc_1_7_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_twiddle_h_rsc_1_7_wait_dp_inst_twiddle_h_rsc_1_7_i_qb_d_mxwt;

  twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_1_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_1_6_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_1_6_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_6_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_1_6_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_6_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_1_6_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_1_6_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_1_6_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_1_6_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_1_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_6_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_6_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_1_6_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_dp_inst_twiddle_h_rsc_1_6_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_dp_inst_twiddle_h_rsc_1_6_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsc_1_6_i_oswt => twiddle_h_rsc_1_6_i_oswt,
      twiddle_h_rsc_1_6_i_biwt => twiddle_h_rsc_1_6_i_biwt,
      twiddle_h_rsc_1_6_i_bdwt => twiddle_h_rsc_1_6_i_bdwt,
      twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_h_rsc_1_6_i_oswt_pff => twiddle_h_rsc_1_6_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_dp_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_1_6_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_dp_inst_twiddle_h_rsc_1_6_i_qb_d,
      twiddle_h_rsc_1_6_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_dp_inst_twiddle_h_rsc_1_6_i_qb_d_mxwt,
      twiddle_h_rsc_1_6_i_biwt => twiddle_h_rsc_1_6_i_biwt,
      twiddle_h_rsc_1_6_i_bdwt => twiddle_h_rsc_1_6_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_dp_inst_twiddle_h_rsc_1_6_i_qb_d
      <= twiddle_h_rsc_1_6_i_qb_d;
  twiddle_h_rsc_1_6_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_twiddle_h_rsc_1_6_wait_dp_inst_twiddle_h_rsc_1_6_i_qb_d_mxwt;

  twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_1_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_1_5_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_1_5_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_5_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_1_5_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_5_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_1_5_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_1_5_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_1_5_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_1_5_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_1_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_5_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_5_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_1_5_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_dp_inst_twiddle_h_rsc_1_5_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_dp_inst_twiddle_h_rsc_1_5_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsc_1_5_i_oswt => twiddle_h_rsc_1_5_i_oswt,
      twiddle_h_rsc_1_5_i_biwt => twiddle_h_rsc_1_5_i_biwt,
      twiddle_h_rsc_1_5_i_bdwt => twiddle_h_rsc_1_5_i_bdwt,
      twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_h_rsc_1_5_i_oswt_pff => twiddle_h_rsc_1_5_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_dp_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_1_5_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_dp_inst_twiddle_h_rsc_1_5_i_qb_d,
      twiddle_h_rsc_1_5_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_dp_inst_twiddle_h_rsc_1_5_i_qb_d_mxwt,
      twiddle_h_rsc_1_5_i_biwt => twiddle_h_rsc_1_5_i_biwt,
      twiddle_h_rsc_1_5_i_bdwt => twiddle_h_rsc_1_5_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_dp_inst_twiddle_h_rsc_1_5_i_qb_d
      <= twiddle_h_rsc_1_5_i_qb_d;
  twiddle_h_rsc_1_5_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_twiddle_h_rsc_1_5_wait_dp_inst_twiddle_h_rsc_1_5_i_qb_d_mxwt;

  twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_1_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_1_4_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_1_4_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_4_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_1_4_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_4_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_1_4_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_1_4_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_1_4_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_1_4_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_1_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_4_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_4_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_1_4_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_dp_inst_twiddle_h_rsc_1_4_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_dp_inst_twiddle_h_rsc_1_4_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsc_1_4_i_oswt => twiddle_h_rsc_1_4_i_oswt,
      twiddle_h_rsc_1_4_i_biwt => twiddle_h_rsc_1_4_i_biwt,
      twiddle_h_rsc_1_4_i_bdwt => twiddle_h_rsc_1_4_i_bdwt,
      twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_h_rsc_1_4_i_oswt_pff => twiddle_h_rsc_1_4_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_dp_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_1_4_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_dp_inst_twiddle_h_rsc_1_4_i_qb_d,
      twiddle_h_rsc_1_4_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_dp_inst_twiddle_h_rsc_1_4_i_qb_d_mxwt,
      twiddle_h_rsc_1_4_i_biwt => twiddle_h_rsc_1_4_i_biwt,
      twiddle_h_rsc_1_4_i_bdwt => twiddle_h_rsc_1_4_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_dp_inst_twiddle_h_rsc_1_4_i_qb_d
      <= twiddle_h_rsc_1_4_i_qb_d;
  twiddle_h_rsc_1_4_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_twiddle_h_rsc_1_4_wait_dp_inst_twiddle_h_rsc_1_4_i_qb_d_mxwt;

  twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_1_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_1_3_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_1_3_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_3_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_1_3_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_3_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_1_3_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_1_3_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_1_3_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_1_3_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_1_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_3_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_3_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_1_3_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_dp_inst_twiddle_h_rsc_1_3_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_dp_inst_twiddle_h_rsc_1_3_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsc_1_3_i_oswt => twiddle_h_rsc_1_3_i_oswt,
      twiddle_h_rsc_1_3_i_biwt => twiddle_h_rsc_1_3_i_biwt,
      twiddle_h_rsc_1_3_i_bdwt => twiddle_h_rsc_1_3_i_bdwt,
      twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_h_rsc_1_3_i_oswt_pff => twiddle_h_rsc_1_3_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_dp_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_1_3_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_dp_inst_twiddle_h_rsc_1_3_i_qb_d,
      twiddle_h_rsc_1_3_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_dp_inst_twiddle_h_rsc_1_3_i_qb_d_mxwt,
      twiddle_h_rsc_1_3_i_biwt => twiddle_h_rsc_1_3_i_biwt,
      twiddle_h_rsc_1_3_i_bdwt => twiddle_h_rsc_1_3_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_dp_inst_twiddle_h_rsc_1_3_i_qb_d
      <= twiddle_h_rsc_1_3_i_qb_d;
  twiddle_h_rsc_1_3_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_twiddle_h_rsc_1_3_wait_dp_inst_twiddle_h_rsc_1_3_i_qb_d_mxwt;

  twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_1_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_1_2_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_1_2_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_2_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_1_2_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_2_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_1_2_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_1_2_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_1_2_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_1_2_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_1_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_2_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_2_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_1_2_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_dp_inst_twiddle_h_rsc_1_2_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_dp_inst_twiddle_h_rsc_1_2_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsc_1_2_i_oswt => twiddle_h_rsc_1_2_i_oswt,
      twiddle_h_rsc_1_2_i_biwt => twiddle_h_rsc_1_2_i_biwt,
      twiddle_h_rsc_1_2_i_bdwt => twiddle_h_rsc_1_2_i_bdwt,
      twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_h_rsc_1_2_i_oswt_pff => twiddle_h_rsc_1_2_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_dp_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_1_2_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_dp_inst_twiddle_h_rsc_1_2_i_qb_d,
      twiddle_h_rsc_1_2_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_dp_inst_twiddle_h_rsc_1_2_i_qb_d_mxwt,
      twiddle_h_rsc_1_2_i_biwt => twiddle_h_rsc_1_2_i_biwt,
      twiddle_h_rsc_1_2_i_bdwt => twiddle_h_rsc_1_2_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_dp_inst_twiddle_h_rsc_1_2_i_qb_d
      <= twiddle_h_rsc_1_2_i_qb_d;
  twiddle_h_rsc_1_2_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_twiddle_h_rsc_1_2_wait_dp_inst_twiddle_h_rsc_1_2_i_qb_d_mxwt;

  twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_1_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_1_1_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_1_1_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_1_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_1_1_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_1_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_1_1_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_1_1_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_1_1_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_1_1_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_1_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_1_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_1_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_1_1_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_dp_inst_twiddle_h_rsc_1_1_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_dp_inst_twiddle_h_rsc_1_1_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsc_1_1_i_oswt => twiddle_h_rsc_1_1_i_oswt,
      twiddle_h_rsc_1_1_i_biwt => twiddle_h_rsc_1_1_i_biwt,
      twiddle_h_rsc_1_1_i_bdwt => twiddle_h_rsc_1_1_i_bdwt,
      twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_h_rsc_1_1_i_oswt_pff => twiddle_h_rsc_1_1_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_dp_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_1_1_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_dp_inst_twiddle_h_rsc_1_1_i_qb_d,
      twiddle_h_rsc_1_1_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_dp_inst_twiddle_h_rsc_1_1_i_qb_d_mxwt,
      twiddle_h_rsc_1_1_i_biwt => twiddle_h_rsc_1_1_i_biwt,
      twiddle_h_rsc_1_1_i_bdwt => twiddle_h_rsc_1_1_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_dp_inst_twiddle_h_rsc_1_1_i_qb_d
      <= twiddle_h_rsc_1_1_i_qb_d;
  twiddle_h_rsc_1_1_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_twiddle_h_rsc_1_1_wait_dp_inst_twiddle_h_rsc_1_1_i_qb_d_mxwt;

  twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_1_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_1_0_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_1_0_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_0_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_1_0_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_0_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_1_0_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_1_0_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_1_0_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_1_0_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_1_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_0_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_0_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_1_0_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_dp_inst_twiddle_h_rsc_1_0_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_dp_inst_twiddle_h_rsc_1_0_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsc_1_0_i_oswt => twiddle_h_rsc_1_0_i_oswt,
      twiddle_h_rsc_1_0_i_biwt => twiddle_h_rsc_1_0_i_biwt,
      twiddle_h_rsc_1_0_i_bdwt => twiddle_h_rsc_1_0_i_bdwt,
      twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_h_rsc_1_0_i_oswt_pff => twiddle_h_rsc_1_0_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_dp_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_1_0_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_dp_inst_twiddle_h_rsc_1_0_i_qb_d,
      twiddle_h_rsc_1_0_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_dp_inst_twiddle_h_rsc_1_0_i_qb_d_mxwt,
      twiddle_h_rsc_1_0_i_biwt => twiddle_h_rsc_1_0_i_biwt,
      twiddle_h_rsc_1_0_i_bdwt => twiddle_h_rsc_1_0_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_dp_inst_twiddle_h_rsc_1_0_i_qb_d
      <= twiddle_h_rsc_1_0_i_qb_d;
  twiddle_h_rsc_1_0_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_twiddle_h_rsc_1_0_wait_dp_inst_twiddle_h_rsc_1_0_i_qb_d_mxwt;

  twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_7_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_7_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_7_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_7_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsc_0_7_i_oswt => twiddle_h_rsc_0_7_i_oswt,
      twiddle_h_rsc_0_7_i_biwt => twiddle_h_rsc_0_7_i_biwt,
      twiddle_h_rsc_0_7_i_bdwt => twiddle_h_rsc_0_7_i_bdwt,
      twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_h_rsc_0_7_i_oswt_pff => twiddle_h_rsc_0_7_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_dp_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_7_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_qb_d,
      twiddle_h_rsc_0_7_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_qb_d_mxwt,
      twiddle_h_rsc_0_7_i_biwt => twiddle_h_rsc_0_7_i_biwt,
      twiddle_h_rsc_0_7_i_bdwt => twiddle_h_rsc_0_7_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_qb_d
      <= twiddle_h_rsc_0_7_i_qb_d;
  twiddle_h_rsc_0_7_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_qb_d_mxwt;

  twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_6_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_6_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_6_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_6_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsc_0_6_i_oswt => twiddle_h_rsc_0_6_i_oswt,
      twiddle_h_rsc_0_6_i_biwt => twiddle_h_rsc_0_6_i_biwt,
      twiddle_h_rsc_0_6_i_bdwt => twiddle_h_rsc_0_6_i_bdwt,
      twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_h_rsc_0_6_i_oswt_pff => twiddle_h_rsc_0_6_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_dp_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_6_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_qb_d,
      twiddle_h_rsc_0_6_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_qb_d_mxwt,
      twiddle_h_rsc_0_6_i_biwt => twiddle_h_rsc_0_6_i_biwt,
      twiddle_h_rsc_0_6_i_bdwt => twiddle_h_rsc_0_6_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_qb_d
      <= twiddle_h_rsc_0_6_i_qb_d;
  twiddle_h_rsc_0_6_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_qb_d_mxwt;

  twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_5_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_5_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_5_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_5_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsc_0_5_i_oswt => twiddle_h_rsc_0_5_i_oswt,
      twiddle_h_rsc_0_5_i_biwt => twiddle_h_rsc_0_5_i_biwt,
      twiddle_h_rsc_0_5_i_bdwt => twiddle_h_rsc_0_5_i_bdwt,
      twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_h_rsc_0_5_i_oswt_pff => twiddle_h_rsc_0_5_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_dp_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_5_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_qb_d,
      twiddle_h_rsc_0_5_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_qb_d_mxwt,
      twiddle_h_rsc_0_5_i_biwt => twiddle_h_rsc_0_5_i_biwt,
      twiddle_h_rsc_0_5_i_bdwt => twiddle_h_rsc_0_5_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_qb_d
      <= twiddle_h_rsc_0_5_i_qb_d;
  twiddle_h_rsc_0_5_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_qb_d_mxwt;

  twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_4_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_4_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_4_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_4_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsc_0_4_i_oswt => twiddle_h_rsc_0_4_i_oswt,
      twiddle_h_rsc_0_4_i_biwt => twiddle_h_rsc_0_4_i_biwt,
      twiddle_h_rsc_0_4_i_bdwt => twiddle_h_rsc_0_4_i_bdwt,
      twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_h_rsc_0_4_i_oswt_pff => twiddle_h_rsc_0_4_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_dp_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_4_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_qb_d,
      twiddle_h_rsc_0_4_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_qb_d_mxwt,
      twiddle_h_rsc_0_4_i_biwt => twiddle_h_rsc_0_4_i_biwt,
      twiddle_h_rsc_0_4_i_bdwt => twiddle_h_rsc_0_4_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_qb_d
      <= twiddle_h_rsc_0_4_i_qb_d;
  twiddle_h_rsc_0_4_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_qb_d_mxwt;

  twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_3_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_3_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_3_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_3_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsc_0_3_i_oswt => twiddle_h_rsc_0_3_i_oswt,
      twiddle_h_rsc_0_3_i_biwt => twiddle_h_rsc_0_3_i_biwt,
      twiddle_h_rsc_0_3_i_bdwt => twiddle_h_rsc_0_3_i_bdwt,
      twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_h_rsc_0_3_i_oswt_pff => twiddle_h_rsc_0_3_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_dp_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_3_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_qb_d,
      twiddle_h_rsc_0_3_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_qb_d_mxwt,
      twiddle_h_rsc_0_3_i_biwt => twiddle_h_rsc_0_3_i_biwt,
      twiddle_h_rsc_0_3_i_bdwt => twiddle_h_rsc_0_3_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_qb_d
      <= twiddle_h_rsc_0_3_i_qb_d;
  twiddle_h_rsc_0_3_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_qb_d_mxwt;

  twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_2_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_2_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_2_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_2_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsc_0_2_i_oswt => twiddle_h_rsc_0_2_i_oswt,
      twiddle_h_rsc_0_2_i_biwt => twiddle_h_rsc_0_2_i_biwt,
      twiddle_h_rsc_0_2_i_bdwt => twiddle_h_rsc_0_2_i_bdwt,
      twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_h_rsc_0_2_i_oswt_pff => twiddle_h_rsc_0_2_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_dp_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_2_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_qb_d,
      twiddle_h_rsc_0_2_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_qb_d_mxwt,
      twiddle_h_rsc_0_2_i_biwt => twiddle_h_rsc_0_2_i_biwt,
      twiddle_h_rsc_0_2_i_bdwt => twiddle_h_rsc_0_2_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_qb_d
      <= twiddle_h_rsc_0_2_i_qb_d;
  twiddle_h_rsc_0_2_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_qb_d_mxwt;

  twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_1_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_1_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_1_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_1_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsc_0_1_i_oswt => twiddle_h_rsc_0_1_i_oswt,
      twiddle_h_rsc_0_1_i_biwt => twiddle_h_rsc_0_1_i_biwt,
      twiddle_h_rsc_0_1_i_bdwt => twiddle_h_rsc_0_1_i_bdwt,
      twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_h_rsc_0_1_i_oswt_pff => twiddle_h_rsc_0_1_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_dp_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_1_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_qb_d,
      twiddle_h_rsc_0_1_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_qb_d_mxwt,
      twiddle_h_rsc_0_1_i_biwt => twiddle_h_rsc_0_1_i_biwt,
      twiddle_h_rsc_0_1_i_bdwt => twiddle_h_rsc_0_1_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_qb_d
      <= twiddle_h_rsc_0_1_i_qb_d;
  twiddle_h_rsc_0_1_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_qb_d_mxwt;

  twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_0_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_0_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_0_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_0_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsc_0_0_i_oswt => twiddle_h_rsc_0_0_i_oswt,
      twiddle_h_rsc_0_0_i_biwt => twiddle_h_rsc_0_0_i_biwt,
      twiddle_h_rsc_0_0_i_bdwt => twiddle_h_rsc_0_0_i_bdwt,
      twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_h_rsc_0_0_i_oswt_pff => twiddle_h_rsc_0_0_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_dp_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_0_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_qb_d,
      twiddle_h_rsc_0_0_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_qb_d_mxwt,
      twiddle_h_rsc_0_0_i_biwt => twiddle_h_rsc_0_0_i_biwt,
      twiddle_h_rsc_0_0_i_bdwt => twiddle_h_rsc_0_0_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_qb_d
      <= twiddle_h_rsc_0_0_i_qb_d;
  twiddle_h_rsc_0_0_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_qb_d_mxwt;

  twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_1_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_1_7_i_oswt : IN STD_LOGIC;
    twiddle_rsc_1_7_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_7_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_1_7_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_7_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_1_7_i_oswt : IN STD_LOGIC;
      twiddle_rsc_1_7_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_1_7_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_rsc_1_7_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_1_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_7_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_7_i_biwt : IN STD_LOGIC;
      twiddle_rsc_1_7_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_dp_inst_twiddle_rsc_1_7_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_dp_inst_twiddle_rsc_1_7_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_1_7_i_oswt => twiddle_rsc_1_7_i_oswt,
      twiddle_rsc_1_7_i_biwt => twiddle_rsc_1_7_i_biwt,
      twiddle_rsc_1_7_i_bdwt => twiddle_rsc_1_7_i_bdwt,
      twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_rsc_1_7_i_oswt_pff => twiddle_rsc_1_7_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_dp_inst :
      inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_1_7_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_dp_inst_twiddle_rsc_1_7_i_qb_d,
      twiddle_rsc_1_7_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_dp_inst_twiddle_rsc_1_7_i_qb_d_mxwt,
      twiddle_rsc_1_7_i_biwt => twiddle_rsc_1_7_i_biwt,
      twiddle_rsc_1_7_i_bdwt => twiddle_rsc_1_7_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_dp_inst_twiddle_rsc_1_7_i_qb_d
      <= twiddle_rsc_1_7_i_qb_d;
  twiddle_rsc_1_7_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_twiddle_rsc_1_7_wait_dp_inst_twiddle_rsc_1_7_i_qb_d_mxwt;

  twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_1_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_1_6_i_oswt : IN STD_LOGIC;
    twiddle_rsc_1_6_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_6_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_1_6_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_6_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_1_6_i_oswt : IN STD_LOGIC;
      twiddle_rsc_1_6_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_1_6_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_rsc_1_6_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_1_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_6_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_6_i_biwt : IN STD_LOGIC;
      twiddle_rsc_1_6_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_dp_inst_twiddle_rsc_1_6_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_dp_inst_twiddle_rsc_1_6_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_1_6_i_oswt => twiddle_rsc_1_6_i_oswt,
      twiddle_rsc_1_6_i_biwt => twiddle_rsc_1_6_i_biwt,
      twiddle_rsc_1_6_i_bdwt => twiddle_rsc_1_6_i_bdwt,
      twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_rsc_1_6_i_oswt_pff => twiddle_rsc_1_6_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_dp_inst :
      inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_1_6_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_dp_inst_twiddle_rsc_1_6_i_qb_d,
      twiddle_rsc_1_6_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_dp_inst_twiddle_rsc_1_6_i_qb_d_mxwt,
      twiddle_rsc_1_6_i_biwt => twiddle_rsc_1_6_i_biwt,
      twiddle_rsc_1_6_i_bdwt => twiddle_rsc_1_6_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_dp_inst_twiddle_rsc_1_6_i_qb_d
      <= twiddle_rsc_1_6_i_qb_d;
  twiddle_rsc_1_6_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_twiddle_rsc_1_6_wait_dp_inst_twiddle_rsc_1_6_i_qb_d_mxwt;

  twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_1_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_1_5_i_oswt : IN STD_LOGIC;
    twiddle_rsc_1_5_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_5_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_1_5_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_5_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_1_5_i_oswt : IN STD_LOGIC;
      twiddle_rsc_1_5_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_1_5_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_rsc_1_5_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_1_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_5_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_5_i_biwt : IN STD_LOGIC;
      twiddle_rsc_1_5_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_dp_inst_twiddle_rsc_1_5_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_dp_inst_twiddle_rsc_1_5_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_1_5_i_oswt => twiddle_rsc_1_5_i_oswt,
      twiddle_rsc_1_5_i_biwt => twiddle_rsc_1_5_i_biwt,
      twiddle_rsc_1_5_i_bdwt => twiddle_rsc_1_5_i_bdwt,
      twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_rsc_1_5_i_oswt_pff => twiddle_rsc_1_5_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_dp_inst :
      inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_1_5_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_dp_inst_twiddle_rsc_1_5_i_qb_d,
      twiddle_rsc_1_5_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_dp_inst_twiddle_rsc_1_5_i_qb_d_mxwt,
      twiddle_rsc_1_5_i_biwt => twiddle_rsc_1_5_i_biwt,
      twiddle_rsc_1_5_i_bdwt => twiddle_rsc_1_5_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_dp_inst_twiddle_rsc_1_5_i_qb_d
      <= twiddle_rsc_1_5_i_qb_d;
  twiddle_rsc_1_5_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_twiddle_rsc_1_5_wait_dp_inst_twiddle_rsc_1_5_i_qb_d_mxwt;

  twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_1_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_1_4_i_oswt : IN STD_LOGIC;
    twiddle_rsc_1_4_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_4_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_1_4_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_4_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_1_4_i_oswt : IN STD_LOGIC;
      twiddle_rsc_1_4_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_1_4_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_rsc_1_4_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_1_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_4_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_4_i_biwt : IN STD_LOGIC;
      twiddle_rsc_1_4_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_dp_inst_twiddle_rsc_1_4_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_dp_inst_twiddle_rsc_1_4_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_1_4_i_oswt => twiddle_rsc_1_4_i_oswt,
      twiddle_rsc_1_4_i_biwt => twiddle_rsc_1_4_i_biwt,
      twiddle_rsc_1_4_i_bdwt => twiddle_rsc_1_4_i_bdwt,
      twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_rsc_1_4_i_oswt_pff => twiddle_rsc_1_4_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_dp_inst :
      inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_1_4_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_dp_inst_twiddle_rsc_1_4_i_qb_d,
      twiddle_rsc_1_4_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_dp_inst_twiddle_rsc_1_4_i_qb_d_mxwt,
      twiddle_rsc_1_4_i_biwt => twiddle_rsc_1_4_i_biwt,
      twiddle_rsc_1_4_i_bdwt => twiddle_rsc_1_4_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_dp_inst_twiddle_rsc_1_4_i_qb_d
      <= twiddle_rsc_1_4_i_qb_d;
  twiddle_rsc_1_4_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_twiddle_rsc_1_4_wait_dp_inst_twiddle_rsc_1_4_i_qb_d_mxwt;

  twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_1_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_1_3_i_oswt : IN STD_LOGIC;
    twiddle_rsc_1_3_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_3_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_1_3_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_3_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_1_3_i_oswt : IN STD_LOGIC;
      twiddle_rsc_1_3_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_1_3_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_rsc_1_3_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_1_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_3_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_3_i_biwt : IN STD_LOGIC;
      twiddle_rsc_1_3_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_dp_inst_twiddle_rsc_1_3_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_dp_inst_twiddle_rsc_1_3_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_1_3_i_oswt => twiddle_rsc_1_3_i_oswt,
      twiddle_rsc_1_3_i_biwt => twiddle_rsc_1_3_i_biwt,
      twiddle_rsc_1_3_i_bdwt => twiddle_rsc_1_3_i_bdwt,
      twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_rsc_1_3_i_oswt_pff => twiddle_rsc_1_3_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_dp_inst :
      inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_1_3_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_dp_inst_twiddle_rsc_1_3_i_qb_d,
      twiddle_rsc_1_3_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_dp_inst_twiddle_rsc_1_3_i_qb_d_mxwt,
      twiddle_rsc_1_3_i_biwt => twiddle_rsc_1_3_i_biwt,
      twiddle_rsc_1_3_i_bdwt => twiddle_rsc_1_3_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_dp_inst_twiddle_rsc_1_3_i_qb_d
      <= twiddle_rsc_1_3_i_qb_d;
  twiddle_rsc_1_3_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_twiddle_rsc_1_3_wait_dp_inst_twiddle_rsc_1_3_i_qb_d_mxwt;

  twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_1_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_1_2_i_oswt : IN STD_LOGIC;
    twiddle_rsc_1_2_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_2_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_1_2_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_2_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_1_2_i_oswt : IN STD_LOGIC;
      twiddle_rsc_1_2_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_1_2_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_rsc_1_2_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_1_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_2_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_2_i_biwt : IN STD_LOGIC;
      twiddle_rsc_1_2_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_dp_inst_twiddle_rsc_1_2_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_dp_inst_twiddle_rsc_1_2_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_1_2_i_oswt => twiddle_rsc_1_2_i_oswt,
      twiddle_rsc_1_2_i_biwt => twiddle_rsc_1_2_i_biwt,
      twiddle_rsc_1_2_i_bdwt => twiddle_rsc_1_2_i_bdwt,
      twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_rsc_1_2_i_oswt_pff => twiddle_rsc_1_2_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_dp_inst :
      inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_1_2_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_dp_inst_twiddle_rsc_1_2_i_qb_d,
      twiddle_rsc_1_2_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_dp_inst_twiddle_rsc_1_2_i_qb_d_mxwt,
      twiddle_rsc_1_2_i_biwt => twiddle_rsc_1_2_i_biwt,
      twiddle_rsc_1_2_i_bdwt => twiddle_rsc_1_2_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_dp_inst_twiddle_rsc_1_2_i_qb_d
      <= twiddle_rsc_1_2_i_qb_d;
  twiddle_rsc_1_2_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_twiddle_rsc_1_2_wait_dp_inst_twiddle_rsc_1_2_i_qb_d_mxwt;

  twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_1_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_1_1_i_oswt : IN STD_LOGIC;
    twiddle_rsc_1_1_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_1_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_1_1_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_1_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_1_1_i_oswt : IN STD_LOGIC;
      twiddle_rsc_1_1_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_1_1_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_rsc_1_1_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_1_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_1_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_1_i_biwt : IN STD_LOGIC;
      twiddle_rsc_1_1_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_dp_inst_twiddle_rsc_1_1_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_dp_inst_twiddle_rsc_1_1_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_1_1_i_oswt => twiddle_rsc_1_1_i_oswt,
      twiddle_rsc_1_1_i_biwt => twiddle_rsc_1_1_i_biwt,
      twiddle_rsc_1_1_i_bdwt => twiddle_rsc_1_1_i_bdwt,
      twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_rsc_1_1_i_oswt_pff => twiddle_rsc_1_1_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_dp_inst :
      inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_1_1_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_dp_inst_twiddle_rsc_1_1_i_qb_d,
      twiddle_rsc_1_1_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_dp_inst_twiddle_rsc_1_1_i_qb_d_mxwt,
      twiddle_rsc_1_1_i_biwt => twiddle_rsc_1_1_i_biwt,
      twiddle_rsc_1_1_i_bdwt => twiddle_rsc_1_1_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_dp_inst_twiddle_rsc_1_1_i_qb_d
      <= twiddle_rsc_1_1_i_qb_d;
  twiddle_rsc_1_1_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_twiddle_rsc_1_1_wait_dp_inst_twiddle_rsc_1_1_i_qb_d_mxwt;

  twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_1_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_1_0_i_oswt : IN STD_LOGIC;
    twiddle_rsc_1_0_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_0_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_1_0_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_0_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_1_0_i_oswt : IN STD_LOGIC;
      twiddle_rsc_1_0_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_1_0_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_rsc_1_0_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_1_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_0_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_0_i_biwt : IN STD_LOGIC;
      twiddle_rsc_1_0_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_dp_inst_twiddle_rsc_1_0_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_dp_inst_twiddle_rsc_1_0_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_1_0_i_oswt => twiddle_rsc_1_0_i_oswt,
      twiddle_rsc_1_0_i_biwt => twiddle_rsc_1_0_i_biwt,
      twiddle_rsc_1_0_i_bdwt => twiddle_rsc_1_0_i_bdwt,
      twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_rsc_1_0_i_oswt_pff => twiddle_rsc_1_0_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_dp_inst :
      inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_1_0_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_dp_inst_twiddle_rsc_1_0_i_qb_d,
      twiddle_rsc_1_0_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_dp_inst_twiddle_rsc_1_0_i_qb_d_mxwt,
      twiddle_rsc_1_0_i_biwt => twiddle_rsc_1_0_i_biwt,
      twiddle_rsc_1_0_i_bdwt => twiddle_rsc_1_0_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_dp_inst_twiddle_rsc_1_0_i_qb_d
      <= twiddle_rsc_1_0_i_qb_d;
  twiddle_rsc_1_0_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_twiddle_rsc_1_0_wait_dp_inst_twiddle_rsc_1_0_i_qb_d_mxwt;

  twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_0_7_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_7_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_7_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_7_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_0_7_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_7_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_7_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_7_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_7_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_7_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_7_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_0_7_i_oswt => twiddle_rsc_0_7_i_oswt,
      twiddle_rsc_0_7_i_biwt => twiddle_rsc_0_7_i_biwt,
      twiddle_rsc_0_7_i_bdwt => twiddle_rsc_0_7_i_bdwt,
      twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_rsc_0_7_i_oswt_pff => twiddle_rsc_0_7_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_dp_inst :
      inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_7_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_qb_d,
      twiddle_rsc_0_7_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_qb_d_mxwt,
      twiddle_rsc_0_7_i_biwt => twiddle_rsc_0_7_i_biwt,
      twiddle_rsc_0_7_i_bdwt => twiddle_rsc_0_7_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_qb_d
      <= twiddle_rsc_0_7_i_qb_d;
  twiddle_rsc_0_7_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_qb_d_mxwt;

  twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_0_6_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_6_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_6_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_6_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_0_6_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_6_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_6_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_6_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_6_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_6_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_6_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_0_6_i_oswt => twiddle_rsc_0_6_i_oswt,
      twiddle_rsc_0_6_i_biwt => twiddle_rsc_0_6_i_biwt,
      twiddle_rsc_0_6_i_bdwt => twiddle_rsc_0_6_i_bdwt,
      twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_rsc_0_6_i_oswt_pff => twiddle_rsc_0_6_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_dp_inst :
      inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_6_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_qb_d,
      twiddle_rsc_0_6_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_qb_d_mxwt,
      twiddle_rsc_0_6_i_biwt => twiddle_rsc_0_6_i_biwt,
      twiddle_rsc_0_6_i_bdwt => twiddle_rsc_0_6_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_qb_d
      <= twiddle_rsc_0_6_i_qb_d;
  twiddle_rsc_0_6_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_qb_d_mxwt;

  twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_0_5_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_5_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_5_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_5_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_0_5_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_5_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_5_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_5_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_5_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_5_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_5_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_0_5_i_oswt => twiddle_rsc_0_5_i_oswt,
      twiddle_rsc_0_5_i_biwt => twiddle_rsc_0_5_i_biwt,
      twiddle_rsc_0_5_i_bdwt => twiddle_rsc_0_5_i_bdwt,
      twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_rsc_0_5_i_oswt_pff => twiddle_rsc_0_5_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_dp_inst :
      inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_5_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_qb_d,
      twiddle_rsc_0_5_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_qb_d_mxwt,
      twiddle_rsc_0_5_i_biwt => twiddle_rsc_0_5_i_biwt,
      twiddle_rsc_0_5_i_bdwt => twiddle_rsc_0_5_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_qb_d
      <= twiddle_rsc_0_5_i_qb_d;
  twiddle_rsc_0_5_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_qb_d_mxwt;

  twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_0_4_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_4_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_4_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_4_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_0_4_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_4_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_4_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_4_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_4_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_4_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_4_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_0_4_i_oswt => twiddle_rsc_0_4_i_oswt,
      twiddle_rsc_0_4_i_biwt => twiddle_rsc_0_4_i_biwt,
      twiddle_rsc_0_4_i_bdwt => twiddle_rsc_0_4_i_bdwt,
      twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_rsc_0_4_i_oswt_pff => twiddle_rsc_0_4_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_dp_inst :
      inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_4_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_qb_d,
      twiddle_rsc_0_4_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_qb_d_mxwt,
      twiddle_rsc_0_4_i_biwt => twiddle_rsc_0_4_i_biwt,
      twiddle_rsc_0_4_i_bdwt => twiddle_rsc_0_4_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_qb_d
      <= twiddle_rsc_0_4_i_qb_d;
  twiddle_rsc_0_4_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_qb_d_mxwt;

  twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_0_3_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_3_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_3_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_3_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_0_3_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_3_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_3_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_3_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_3_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_3_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_3_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_0_3_i_oswt => twiddle_rsc_0_3_i_oswt,
      twiddle_rsc_0_3_i_biwt => twiddle_rsc_0_3_i_biwt,
      twiddle_rsc_0_3_i_bdwt => twiddle_rsc_0_3_i_bdwt,
      twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_rsc_0_3_i_oswt_pff => twiddle_rsc_0_3_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_dp_inst :
      inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_3_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_qb_d,
      twiddle_rsc_0_3_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_qb_d_mxwt,
      twiddle_rsc_0_3_i_biwt => twiddle_rsc_0_3_i_biwt,
      twiddle_rsc_0_3_i_bdwt => twiddle_rsc_0_3_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_qb_d
      <= twiddle_rsc_0_3_i_qb_d;
  twiddle_rsc_0_3_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_qb_d_mxwt;

  twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_0_2_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_2_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_2_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_2_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_0_2_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_2_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_2_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_2_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_2_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_2_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_2_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_0_2_i_oswt => twiddle_rsc_0_2_i_oswt,
      twiddle_rsc_0_2_i_biwt => twiddle_rsc_0_2_i_biwt,
      twiddle_rsc_0_2_i_bdwt => twiddle_rsc_0_2_i_bdwt,
      twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_rsc_0_2_i_oswt_pff => twiddle_rsc_0_2_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_dp_inst :
      inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_2_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_qb_d,
      twiddle_rsc_0_2_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_qb_d_mxwt,
      twiddle_rsc_0_2_i_biwt => twiddle_rsc_0_2_i_biwt,
      twiddle_rsc_0_2_i_bdwt => twiddle_rsc_0_2_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_qb_d
      <= twiddle_rsc_0_2_i_qb_d;
  twiddle_rsc_0_2_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_qb_d_mxwt;

  twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_0_1_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_1_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_1_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_1_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_0_1_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_1_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_1_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_1_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_1_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_1_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_1_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_0_1_i_oswt => twiddle_rsc_0_1_i_oswt,
      twiddle_rsc_0_1_i_biwt => twiddle_rsc_0_1_i_biwt,
      twiddle_rsc_0_1_i_bdwt => twiddle_rsc_0_1_i_bdwt,
      twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_rsc_0_1_i_oswt_pff => twiddle_rsc_0_1_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_dp_inst :
      inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_1_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_qb_d,
      twiddle_rsc_0_1_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_qb_d_mxwt,
      twiddle_rsc_0_1_i_biwt => twiddle_rsc_0_1_i_biwt,
      twiddle_rsc_0_1_i_bdwt => twiddle_rsc_0_1_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_qb_d
      <= twiddle_rsc_0_1_i_qb_d;
  twiddle_rsc_0_1_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_qb_d_mxwt;

  twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_0_0_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_0_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_i_oswt_pff : IN STD_LOGIC;
    core_wten_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_0_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_0_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_0_0_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_0_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_0_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_0_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_0_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_0_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_0_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_ctrl_inst
      : inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_0_0_i_oswt => twiddle_rsc_0_0_i_oswt,
      twiddle_rsc_0_0_i_biwt => twiddle_rsc_0_0_i_biwt,
      twiddle_rsc_0_0_i_bdwt => twiddle_rsc_0_0_i_bdwt,
      twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct => twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct,
      twiddle_rsc_0_0_i_oswt_pff => twiddle_rsc_0_0_i_oswt_pff,
      core_wten_pff => core_wten_pff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_dp_inst :
      inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_0_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_qb_d,
      twiddle_rsc_0_0_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_qb_d_mxwt,
      twiddle_rsc_0_0_i_biwt => twiddle_rsc_0_0_i_biwt,
      twiddle_rsc_0_0_i_bdwt => twiddle_rsc_0_0_i_bdwt
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_qb_d
      <= twiddle_rsc_0_0_i_qb_d;
  twiddle_rsc_0_0_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_qb_d_mxwt;

  twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_core_sct;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_1_7_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_7_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_1_7_i_oswt : IN STD_LOGIC;
    vec_rsc_1_7_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_1_7_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_7_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_7_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_1_7_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_1_7_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_7_i_biwt : STD_LOGIC;
  SIGNAL vec_rsc_1_7_i_bdwt : STD_LOGIC;
  SIGNAL vec_rsc_1_7_i_biwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_1_7_i_bdwt_2 : STD_LOGIC;
  SIGNAL vec_rsc_1_7_i_wea_d_core_sct : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_1_7_i_oswt : IN STD_LOGIC;
      vec_rsc_1_7_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_1_7_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_7_i_biwt : OUT STD_LOGIC;
      vec_rsc_1_7_i_bdwt : OUT STD_LOGIC;
      vec_rsc_1_7_i_biwt_1 : OUT STD_LOGIC;
      vec_rsc_1_7_i_bdwt_2 : OUT STD_LOGIC;
      vec_rsc_1_7_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_1_7_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_1_7_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_wea_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_1_7_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_7_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_7_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_7_i_biwt : IN STD_LOGIC;
      vec_rsc_1_7_i_bdwt : IN STD_LOGIC;
      vec_rsc_1_7_i_biwt_1 : IN STD_LOGIC;
      vec_rsc_1_7_i_bdwt_2 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp_inst_vec_rsc_1_7_i_da_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp_inst_vec_rsc_1_7_i_qa_d
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp_inst_vec_rsc_1_7_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp_inst_vec_rsc_1_7_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      vec_rsc_1_7_i_oswt => vec_rsc_1_7_i_oswt,
      vec_rsc_1_7_i_oswt_1 => vec_rsc_1_7_i_oswt_1,
      vec_rsc_1_7_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_wea_d_core_psct,
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      vec_rsc_1_7_i_biwt => vec_rsc_1_7_i_biwt,
      vec_rsc_1_7_i_bdwt => vec_rsc_1_7_i_bdwt,
      vec_rsc_1_7_i_biwt_1 => vec_rsc_1_7_i_biwt_1,
      vec_rsc_1_7_i_bdwt_2 => vec_rsc_1_7_i_bdwt_2,
      vec_rsc_1_7_i_wea_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_wea_d_core_sct,
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct,
      core_wten_pff => core_wten_pff,
      vec_rsc_1_7_i_oswt_pff => vec_rsc_1_7_i_oswt_pff,
      vec_rsc_1_7_i_oswt_1_pff => vec_rsc_1_7_i_oswt_1_pff
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_1_7_i_wea_d_core_psct(0)));
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0)));
  vec_rsc_1_7_i_wea_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_wea_d_core_sct;
  vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_ctrl_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;

  inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_1_7_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp_inst_vec_rsc_1_7_i_da_d,
      vec_rsc_1_7_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp_inst_vec_rsc_1_7_i_qa_d,
      vec_rsc_1_7_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp_inst_vec_rsc_1_7_i_da_d_core,
      vec_rsc_1_7_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp_inst_vec_rsc_1_7_i_qa_d_mxwt,
      vec_rsc_1_7_i_biwt => vec_rsc_1_7_i_biwt,
      vec_rsc_1_7_i_bdwt => vec_rsc_1_7_i_bdwt,
      vec_rsc_1_7_i_biwt_1 => vec_rsc_1_7_i_biwt_1,
      vec_rsc_1_7_i_bdwt_2 => vec_rsc_1_7_i_bdwt_2
    );
  vec_rsc_1_7_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp_inst_vec_rsc_1_7_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp_inst_vec_rsc_1_7_i_qa_d
      <= vec_rsc_1_7_i_qa_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp_inst_vec_rsc_1_7_i_da_d_core
      <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000") & (vec_rsc_1_7_i_da_d_core(31
      DOWNTO 0));
  vec_rsc_1_7_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_vec_rsc_1_7_wait_dp_inst_vec_rsc_1_7_i_qa_d_mxwt;

  vec_rsc_1_7_i_wea_d <= vec_rsc_1_7_i_wea_d_core_sct;
  vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;
  vec_rsc_1_7_i_da_d <= vec_rsc_1_7_i_da_d_reg;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_1_6_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_6_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_1_6_i_oswt : IN STD_LOGIC;
    vec_rsc_1_6_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_1_6_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_6_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_6_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_1_6_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_1_6_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_6_i_biwt : STD_LOGIC;
  SIGNAL vec_rsc_1_6_i_bdwt : STD_LOGIC;
  SIGNAL vec_rsc_1_6_i_biwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_1_6_i_bdwt_2 : STD_LOGIC;
  SIGNAL vec_rsc_1_6_i_wea_d_core_sct : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_1_6_i_oswt : IN STD_LOGIC;
      vec_rsc_1_6_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_1_6_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_6_i_biwt : OUT STD_LOGIC;
      vec_rsc_1_6_i_bdwt : OUT STD_LOGIC;
      vec_rsc_1_6_i_biwt_1 : OUT STD_LOGIC;
      vec_rsc_1_6_i_bdwt_2 : OUT STD_LOGIC;
      vec_rsc_1_6_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_1_6_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_1_6_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_wea_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_1_6_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_6_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_6_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_6_i_biwt : IN STD_LOGIC;
      vec_rsc_1_6_i_bdwt : IN STD_LOGIC;
      vec_rsc_1_6_i_biwt_1 : IN STD_LOGIC;
      vec_rsc_1_6_i_bdwt_2 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp_inst_vec_rsc_1_6_i_da_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp_inst_vec_rsc_1_6_i_qa_d
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp_inst_vec_rsc_1_6_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp_inst_vec_rsc_1_6_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      vec_rsc_1_6_i_oswt => vec_rsc_1_6_i_oswt,
      vec_rsc_1_6_i_oswt_1 => vec_rsc_1_6_i_oswt_1,
      vec_rsc_1_6_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_wea_d_core_psct,
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      vec_rsc_1_6_i_biwt => vec_rsc_1_6_i_biwt,
      vec_rsc_1_6_i_bdwt => vec_rsc_1_6_i_bdwt,
      vec_rsc_1_6_i_biwt_1 => vec_rsc_1_6_i_biwt_1,
      vec_rsc_1_6_i_bdwt_2 => vec_rsc_1_6_i_bdwt_2,
      vec_rsc_1_6_i_wea_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_wea_d_core_sct,
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct,
      core_wten_pff => core_wten_pff,
      vec_rsc_1_6_i_oswt_pff => vec_rsc_1_6_i_oswt_pff,
      vec_rsc_1_6_i_oswt_1_pff => vec_rsc_1_6_i_oswt_1_pff
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_1_6_i_wea_d_core_psct(0)));
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0)));
  vec_rsc_1_6_i_wea_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_wea_d_core_sct;
  vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_ctrl_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;

  inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_1_6_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp_inst_vec_rsc_1_6_i_da_d,
      vec_rsc_1_6_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp_inst_vec_rsc_1_6_i_qa_d,
      vec_rsc_1_6_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp_inst_vec_rsc_1_6_i_da_d_core,
      vec_rsc_1_6_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp_inst_vec_rsc_1_6_i_qa_d_mxwt,
      vec_rsc_1_6_i_biwt => vec_rsc_1_6_i_biwt,
      vec_rsc_1_6_i_bdwt => vec_rsc_1_6_i_bdwt,
      vec_rsc_1_6_i_biwt_1 => vec_rsc_1_6_i_biwt_1,
      vec_rsc_1_6_i_bdwt_2 => vec_rsc_1_6_i_bdwt_2
    );
  vec_rsc_1_6_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp_inst_vec_rsc_1_6_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp_inst_vec_rsc_1_6_i_qa_d
      <= vec_rsc_1_6_i_qa_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp_inst_vec_rsc_1_6_i_da_d_core
      <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000") & (vec_rsc_1_6_i_da_d_core(31
      DOWNTO 0));
  vec_rsc_1_6_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_vec_rsc_1_6_wait_dp_inst_vec_rsc_1_6_i_qa_d_mxwt;

  vec_rsc_1_6_i_wea_d <= vec_rsc_1_6_i_wea_d_core_sct;
  vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;
  vec_rsc_1_6_i_da_d <= vec_rsc_1_6_i_da_d_reg;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_1_5_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_5_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_1_5_i_oswt : IN STD_LOGIC;
    vec_rsc_1_5_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_1_5_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_5_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_5_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_1_5_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_1_5_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_5_i_biwt : STD_LOGIC;
  SIGNAL vec_rsc_1_5_i_bdwt : STD_LOGIC;
  SIGNAL vec_rsc_1_5_i_biwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_1_5_i_bdwt_2 : STD_LOGIC;
  SIGNAL vec_rsc_1_5_i_wea_d_core_sct : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_1_5_i_oswt : IN STD_LOGIC;
      vec_rsc_1_5_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_1_5_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_5_i_biwt : OUT STD_LOGIC;
      vec_rsc_1_5_i_bdwt : OUT STD_LOGIC;
      vec_rsc_1_5_i_biwt_1 : OUT STD_LOGIC;
      vec_rsc_1_5_i_bdwt_2 : OUT STD_LOGIC;
      vec_rsc_1_5_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_1_5_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_1_5_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_wea_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_1_5_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_5_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_5_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_5_i_biwt : IN STD_LOGIC;
      vec_rsc_1_5_i_bdwt : IN STD_LOGIC;
      vec_rsc_1_5_i_biwt_1 : IN STD_LOGIC;
      vec_rsc_1_5_i_bdwt_2 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp_inst_vec_rsc_1_5_i_da_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp_inst_vec_rsc_1_5_i_qa_d
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp_inst_vec_rsc_1_5_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp_inst_vec_rsc_1_5_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      vec_rsc_1_5_i_oswt => vec_rsc_1_5_i_oswt,
      vec_rsc_1_5_i_oswt_1 => vec_rsc_1_5_i_oswt_1,
      vec_rsc_1_5_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_wea_d_core_psct,
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      vec_rsc_1_5_i_biwt => vec_rsc_1_5_i_biwt,
      vec_rsc_1_5_i_bdwt => vec_rsc_1_5_i_bdwt,
      vec_rsc_1_5_i_biwt_1 => vec_rsc_1_5_i_biwt_1,
      vec_rsc_1_5_i_bdwt_2 => vec_rsc_1_5_i_bdwt_2,
      vec_rsc_1_5_i_wea_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_wea_d_core_sct,
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct,
      core_wten_pff => core_wten_pff,
      vec_rsc_1_5_i_oswt_pff => vec_rsc_1_5_i_oswt_pff,
      vec_rsc_1_5_i_oswt_1_pff => vec_rsc_1_5_i_oswt_1_pff
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_1_5_i_wea_d_core_psct(0)));
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0)));
  vec_rsc_1_5_i_wea_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_wea_d_core_sct;
  vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_ctrl_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;

  inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_1_5_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp_inst_vec_rsc_1_5_i_da_d,
      vec_rsc_1_5_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp_inst_vec_rsc_1_5_i_qa_d,
      vec_rsc_1_5_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp_inst_vec_rsc_1_5_i_da_d_core,
      vec_rsc_1_5_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp_inst_vec_rsc_1_5_i_qa_d_mxwt,
      vec_rsc_1_5_i_biwt => vec_rsc_1_5_i_biwt,
      vec_rsc_1_5_i_bdwt => vec_rsc_1_5_i_bdwt,
      vec_rsc_1_5_i_biwt_1 => vec_rsc_1_5_i_biwt_1,
      vec_rsc_1_5_i_bdwt_2 => vec_rsc_1_5_i_bdwt_2
    );
  vec_rsc_1_5_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp_inst_vec_rsc_1_5_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp_inst_vec_rsc_1_5_i_qa_d
      <= vec_rsc_1_5_i_qa_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp_inst_vec_rsc_1_5_i_da_d_core
      <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000") & (vec_rsc_1_5_i_da_d_core(31
      DOWNTO 0));
  vec_rsc_1_5_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_vec_rsc_1_5_wait_dp_inst_vec_rsc_1_5_i_qa_d_mxwt;

  vec_rsc_1_5_i_wea_d <= vec_rsc_1_5_i_wea_d_core_sct;
  vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;
  vec_rsc_1_5_i_da_d <= vec_rsc_1_5_i_da_d_reg;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_1_4_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_4_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_1_4_i_oswt : IN STD_LOGIC;
    vec_rsc_1_4_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_1_4_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_4_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_4_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_1_4_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_1_4_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_4_i_biwt : STD_LOGIC;
  SIGNAL vec_rsc_1_4_i_bdwt : STD_LOGIC;
  SIGNAL vec_rsc_1_4_i_biwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_1_4_i_bdwt_2 : STD_LOGIC;
  SIGNAL vec_rsc_1_4_i_wea_d_core_sct : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_1_4_i_oswt : IN STD_LOGIC;
      vec_rsc_1_4_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_1_4_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_4_i_biwt : OUT STD_LOGIC;
      vec_rsc_1_4_i_bdwt : OUT STD_LOGIC;
      vec_rsc_1_4_i_biwt_1 : OUT STD_LOGIC;
      vec_rsc_1_4_i_bdwt_2 : OUT STD_LOGIC;
      vec_rsc_1_4_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_1_4_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_1_4_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_wea_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_1_4_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_4_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_4_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_4_i_biwt : IN STD_LOGIC;
      vec_rsc_1_4_i_bdwt : IN STD_LOGIC;
      vec_rsc_1_4_i_biwt_1 : IN STD_LOGIC;
      vec_rsc_1_4_i_bdwt_2 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp_inst_vec_rsc_1_4_i_da_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp_inst_vec_rsc_1_4_i_qa_d
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp_inst_vec_rsc_1_4_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp_inst_vec_rsc_1_4_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      vec_rsc_1_4_i_oswt => vec_rsc_1_4_i_oswt,
      vec_rsc_1_4_i_oswt_1 => vec_rsc_1_4_i_oswt_1,
      vec_rsc_1_4_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_wea_d_core_psct,
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      vec_rsc_1_4_i_biwt => vec_rsc_1_4_i_biwt,
      vec_rsc_1_4_i_bdwt => vec_rsc_1_4_i_bdwt,
      vec_rsc_1_4_i_biwt_1 => vec_rsc_1_4_i_biwt_1,
      vec_rsc_1_4_i_bdwt_2 => vec_rsc_1_4_i_bdwt_2,
      vec_rsc_1_4_i_wea_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_wea_d_core_sct,
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct,
      core_wten_pff => core_wten_pff,
      vec_rsc_1_4_i_oswt_pff => vec_rsc_1_4_i_oswt_pff,
      vec_rsc_1_4_i_oswt_1_pff => vec_rsc_1_4_i_oswt_1_pff
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_1_4_i_wea_d_core_psct(0)));
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0)));
  vec_rsc_1_4_i_wea_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_wea_d_core_sct;
  vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_ctrl_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;

  inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_1_4_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp_inst_vec_rsc_1_4_i_da_d,
      vec_rsc_1_4_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp_inst_vec_rsc_1_4_i_qa_d,
      vec_rsc_1_4_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp_inst_vec_rsc_1_4_i_da_d_core,
      vec_rsc_1_4_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp_inst_vec_rsc_1_4_i_qa_d_mxwt,
      vec_rsc_1_4_i_biwt => vec_rsc_1_4_i_biwt,
      vec_rsc_1_4_i_bdwt => vec_rsc_1_4_i_bdwt,
      vec_rsc_1_4_i_biwt_1 => vec_rsc_1_4_i_biwt_1,
      vec_rsc_1_4_i_bdwt_2 => vec_rsc_1_4_i_bdwt_2
    );
  vec_rsc_1_4_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp_inst_vec_rsc_1_4_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp_inst_vec_rsc_1_4_i_qa_d
      <= vec_rsc_1_4_i_qa_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp_inst_vec_rsc_1_4_i_da_d_core
      <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000") & (vec_rsc_1_4_i_da_d_core(31
      DOWNTO 0));
  vec_rsc_1_4_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_vec_rsc_1_4_wait_dp_inst_vec_rsc_1_4_i_qa_d_mxwt;

  vec_rsc_1_4_i_wea_d <= vec_rsc_1_4_i_wea_d_core_sct;
  vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;
  vec_rsc_1_4_i_da_d <= vec_rsc_1_4_i_da_d_reg;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_1_3_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_3_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_1_3_i_oswt : IN STD_LOGIC;
    vec_rsc_1_3_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_1_3_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_3_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_3_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_1_3_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_1_3_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_3_i_biwt : STD_LOGIC;
  SIGNAL vec_rsc_1_3_i_bdwt : STD_LOGIC;
  SIGNAL vec_rsc_1_3_i_biwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_1_3_i_bdwt_2 : STD_LOGIC;
  SIGNAL vec_rsc_1_3_i_wea_d_core_sct : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_1_3_i_oswt : IN STD_LOGIC;
      vec_rsc_1_3_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_1_3_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_3_i_biwt : OUT STD_LOGIC;
      vec_rsc_1_3_i_bdwt : OUT STD_LOGIC;
      vec_rsc_1_3_i_biwt_1 : OUT STD_LOGIC;
      vec_rsc_1_3_i_bdwt_2 : OUT STD_LOGIC;
      vec_rsc_1_3_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_1_3_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_1_3_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_wea_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_1_3_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_3_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_3_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_3_i_biwt : IN STD_LOGIC;
      vec_rsc_1_3_i_bdwt : IN STD_LOGIC;
      vec_rsc_1_3_i_biwt_1 : IN STD_LOGIC;
      vec_rsc_1_3_i_bdwt_2 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp_inst_vec_rsc_1_3_i_da_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp_inst_vec_rsc_1_3_i_qa_d
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp_inst_vec_rsc_1_3_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp_inst_vec_rsc_1_3_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      vec_rsc_1_3_i_oswt => vec_rsc_1_3_i_oswt,
      vec_rsc_1_3_i_oswt_1 => vec_rsc_1_3_i_oswt_1,
      vec_rsc_1_3_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_wea_d_core_psct,
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      vec_rsc_1_3_i_biwt => vec_rsc_1_3_i_biwt,
      vec_rsc_1_3_i_bdwt => vec_rsc_1_3_i_bdwt,
      vec_rsc_1_3_i_biwt_1 => vec_rsc_1_3_i_biwt_1,
      vec_rsc_1_3_i_bdwt_2 => vec_rsc_1_3_i_bdwt_2,
      vec_rsc_1_3_i_wea_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_wea_d_core_sct,
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct,
      core_wten_pff => core_wten_pff,
      vec_rsc_1_3_i_oswt_pff => vec_rsc_1_3_i_oswt_pff,
      vec_rsc_1_3_i_oswt_1_pff => vec_rsc_1_3_i_oswt_1_pff
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_1_3_i_wea_d_core_psct(0)));
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0)));
  vec_rsc_1_3_i_wea_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_wea_d_core_sct;
  vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_ctrl_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;

  inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_1_3_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp_inst_vec_rsc_1_3_i_da_d,
      vec_rsc_1_3_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp_inst_vec_rsc_1_3_i_qa_d,
      vec_rsc_1_3_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp_inst_vec_rsc_1_3_i_da_d_core,
      vec_rsc_1_3_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp_inst_vec_rsc_1_3_i_qa_d_mxwt,
      vec_rsc_1_3_i_biwt => vec_rsc_1_3_i_biwt,
      vec_rsc_1_3_i_bdwt => vec_rsc_1_3_i_bdwt,
      vec_rsc_1_3_i_biwt_1 => vec_rsc_1_3_i_biwt_1,
      vec_rsc_1_3_i_bdwt_2 => vec_rsc_1_3_i_bdwt_2
    );
  vec_rsc_1_3_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp_inst_vec_rsc_1_3_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp_inst_vec_rsc_1_3_i_qa_d
      <= vec_rsc_1_3_i_qa_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp_inst_vec_rsc_1_3_i_da_d_core
      <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000") & (vec_rsc_1_3_i_da_d_core(31
      DOWNTO 0));
  vec_rsc_1_3_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_vec_rsc_1_3_wait_dp_inst_vec_rsc_1_3_i_qa_d_mxwt;

  vec_rsc_1_3_i_wea_d <= vec_rsc_1_3_i_wea_d_core_sct;
  vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;
  vec_rsc_1_3_i_da_d <= vec_rsc_1_3_i_da_d_reg;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_1_2_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_2_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_1_2_i_oswt : IN STD_LOGIC;
    vec_rsc_1_2_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_1_2_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_2_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_2_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_1_2_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_1_2_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_2_i_biwt : STD_LOGIC;
  SIGNAL vec_rsc_1_2_i_bdwt : STD_LOGIC;
  SIGNAL vec_rsc_1_2_i_biwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_1_2_i_bdwt_2 : STD_LOGIC;
  SIGNAL vec_rsc_1_2_i_wea_d_core_sct : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_1_2_i_oswt : IN STD_LOGIC;
      vec_rsc_1_2_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_1_2_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_2_i_biwt : OUT STD_LOGIC;
      vec_rsc_1_2_i_bdwt : OUT STD_LOGIC;
      vec_rsc_1_2_i_biwt_1 : OUT STD_LOGIC;
      vec_rsc_1_2_i_bdwt_2 : OUT STD_LOGIC;
      vec_rsc_1_2_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_1_2_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_1_2_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_wea_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_1_2_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_2_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_2_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_2_i_biwt : IN STD_LOGIC;
      vec_rsc_1_2_i_bdwt : IN STD_LOGIC;
      vec_rsc_1_2_i_biwt_1 : IN STD_LOGIC;
      vec_rsc_1_2_i_bdwt_2 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp_inst_vec_rsc_1_2_i_da_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp_inst_vec_rsc_1_2_i_qa_d
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp_inst_vec_rsc_1_2_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp_inst_vec_rsc_1_2_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      vec_rsc_1_2_i_oswt => vec_rsc_1_2_i_oswt,
      vec_rsc_1_2_i_oswt_1 => vec_rsc_1_2_i_oswt_1,
      vec_rsc_1_2_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_wea_d_core_psct,
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      vec_rsc_1_2_i_biwt => vec_rsc_1_2_i_biwt,
      vec_rsc_1_2_i_bdwt => vec_rsc_1_2_i_bdwt,
      vec_rsc_1_2_i_biwt_1 => vec_rsc_1_2_i_biwt_1,
      vec_rsc_1_2_i_bdwt_2 => vec_rsc_1_2_i_bdwt_2,
      vec_rsc_1_2_i_wea_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_wea_d_core_sct,
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct,
      core_wten_pff => core_wten_pff,
      vec_rsc_1_2_i_oswt_pff => vec_rsc_1_2_i_oswt_pff,
      vec_rsc_1_2_i_oswt_1_pff => vec_rsc_1_2_i_oswt_1_pff
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_1_2_i_wea_d_core_psct(0)));
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0)));
  vec_rsc_1_2_i_wea_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_wea_d_core_sct;
  vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_ctrl_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;

  inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_1_2_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp_inst_vec_rsc_1_2_i_da_d,
      vec_rsc_1_2_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp_inst_vec_rsc_1_2_i_qa_d,
      vec_rsc_1_2_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp_inst_vec_rsc_1_2_i_da_d_core,
      vec_rsc_1_2_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp_inst_vec_rsc_1_2_i_qa_d_mxwt,
      vec_rsc_1_2_i_biwt => vec_rsc_1_2_i_biwt,
      vec_rsc_1_2_i_bdwt => vec_rsc_1_2_i_bdwt,
      vec_rsc_1_2_i_biwt_1 => vec_rsc_1_2_i_biwt_1,
      vec_rsc_1_2_i_bdwt_2 => vec_rsc_1_2_i_bdwt_2
    );
  vec_rsc_1_2_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp_inst_vec_rsc_1_2_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp_inst_vec_rsc_1_2_i_qa_d
      <= vec_rsc_1_2_i_qa_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp_inst_vec_rsc_1_2_i_da_d_core
      <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000") & (vec_rsc_1_2_i_da_d_core(31
      DOWNTO 0));
  vec_rsc_1_2_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_vec_rsc_1_2_wait_dp_inst_vec_rsc_1_2_i_qa_d_mxwt;

  vec_rsc_1_2_i_wea_d <= vec_rsc_1_2_i_wea_d_core_sct;
  vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;
  vec_rsc_1_2_i_da_d <= vec_rsc_1_2_i_da_d_reg;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_1_1_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_1_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_1_1_i_oswt : IN STD_LOGIC;
    vec_rsc_1_1_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_1_1_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_1_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_1_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_1_1_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_1_1_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_1_i_biwt : STD_LOGIC;
  SIGNAL vec_rsc_1_1_i_bdwt : STD_LOGIC;
  SIGNAL vec_rsc_1_1_i_biwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_1_1_i_bdwt_2 : STD_LOGIC;
  SIGNAL vec_rsc_1_1_i_wea_d_core_sct : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_1_1_i_oswt : IN STD_LOGIC;
      vec_rsc_1_1_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_1_1_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_1_i_biwt : OUT STD_LOGIC;
      vec_rsc_1_1_i_bdwt : OUT STD_LOGIC;
      vec_rsc_1_1_i_biwt_1 : OUT STD_LOGIC;
      vec_rsc_1_1_i_bdwt_2 : OUT STD_LOGIC;
      vec_rsc_1_1_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_1_1_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_1_1_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_wea_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_1_1_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_1_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_1_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_1_i_biwt : IN STD_LOGIC;
      vec_rsc_1_1_i_bdwt : IN STD_LOGIC;
      vec_rsc_1_1_i_biwt_1 : IN STD_LOGIC;
      vec_rsc_1_1_i_bdwt_2 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp_inst_vec_rsc_1_1_i_da_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp_inst_vec_rsc_1_1_i_qa_d
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp_inst_vec_rsc_1_1_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp_inst_vec_rsc_1_1_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      vec_rsc_1_1_i_oswt => vec_rsc_1_1_i_oswt,
      vec_rsc_1_1_i_oswt_1 => vec_rsc_1_1_i_oswt_1,
      vec_rsc_1_1_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_wea_d_core_psct,
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      vec_rsc_1_1_i_biwt => vec_rsc_1_1_i_biwt,
      vec_rsc_1_1_i_bdwt => vec_rsc_1_1_i_bdwt,
      vec_rsc_1_1_i_biwt_1 => vec_rsc_1_1_i_biwt_1,
      vec_rsc_1_1_i_bdwt_2 => vec_rsc_1_1_i_bdwt_2,
      vec_rsc_1_1_i_wea_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_wea_d_core_sct,
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct,
      core_wten_pff => core_wten_pff,
      vec_rsc_1_1_i_oswt_pff => vec_rsc_1_1_i_oswt_pff,
      vec_rsc_1_1_i_oswt_1_pff => vec_rsc_1_1_i_oswt_1_pff
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_1_1_i_wea_d_core_psct(0)));
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0)));
  vec_rsc_1_1_i_wea_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_wea_d_core_sct;
  vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_ctrl_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;

  inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_1_1_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp_inst_vec_rsc_1_1_i_da_d,
      vec_rsc_1_1_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp_inst_vec_rsc_1_1_i_qa_d,
      vec_rsc_1_1_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp_inst_vec_rsc_1_1_i_da_d_core,
      vec_rsc_1_1_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp_inst_vec_rsc_1_1_i_qa_d_mxwt,
      vec_rsc_1_1_i_biwt => vec_rsc_1_1_i_biwt,
      vec_rsc_1_1_i_bdwt => vec_rsc_1_1_i_bdwt,
      vec_rsc_1_1_i_biwt_1 => vec_rsc_1_1_i_biwt_1,
      vec_rsc_1_1_i_bdwt_2 => vec_rsc_1_1_i_bdwt_2
    );
  vec_rsc_1_1_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp_inst_vec_rsc_1_1_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp_inst_vec_rsc_1_1_i_qa_d
      <= vec_rsc_1_1_i_qa_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp_inst_vec_rsc_1_1_i_da_d_core
      <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000") & (vec_rsc_1_1_i_da_d_core(31
      DOWNTO 0));
  vec_rsc_1_1_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_vec_rsc_1_1_wait_dp_inst_vec_rsc_1_1_i_qa_d_mxwt;

  vec_rsc_1_1_i_wea_d <= vec_rsc_1_1_i_wea_d_core_sct;
  vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;
  vec_rsc_1_1_i_da_d <= vec_rsc_1_1_i_da_d_reg;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_1_0_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_1_0_i_oswt : IN STD_LOGIC;
    vec_rsc_1_0_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_1_0_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_0_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_0_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_1_0_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_1_0_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_1_0_i_biwt : STD_LOGIC;
  SIGNAL vec_rsc_1_0_i_bdwt : STD_LOGIC;
  SIGNAL vec_rsc_1_0_i_biwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_1_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL vec_rsc_1_0_i_wea_d_core_sct : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_1_0_i_oswt : IN STD_LOGIC;
      vec_rsc_1_0_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_1_0_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_0_i_biwt : OUT STD_LOGIC;
      vec_rsc_1_0_i_bdwt : OUT STD_LOGIC;
      vec_rsc_1_0_i_biwt_1 : OUT STD_LOGIC;
      vec_rsc_1_0_i_bdwt_2 : OUT STD_LOGIC;
      vec_rsc_1_0_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_1_0_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_1_0_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_wea_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_1_0_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_0_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_0_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_0_i_biwt : IN STD_LOGIC;
      vec_rsc_1_0_i_bdwt : IN STD_LOGIC;
      vec_rsc_1_0_i_biwt_1 : IN STD_LOGIC;
      vec_rsc_1_0_i_bdwt_2 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp_inst_vec_rsc_1_0_i_da_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp_inst_vec_rsc_1_0_i_qa_d
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp_inst_vec_rsc_1_0_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp_inst_vec_rsc_1_0_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      vec_rsc_1_0_i_oswt => vec_rsc_1_0_i_oswt,
      vec_rsc_1_0_i_oswt_1 => vec_rsc_1_0_i_oswt_1,
      vec_rsc_1_0_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_wea_d_core_psct,
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      vec_rsc_1_0_i_biwt => vec_rsc_1_0_i_biwt,
      vec_rsc_1_0_i_bdwt => vec_rsc_1_0_i_bdwt,
      vec_rsc_1_0_i_biwt_1 => vec_rsc_1_0_i_biwt_1,
      vec_rsc_1_0_i_bdwt_2 => vec_rsc_1_0_i_bdwt_2,
      vec_rsc_1_0_i_wea_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_wea_d_core_sct,
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct,
      core_wten_pff => core_wten_pff,
      vec_rsc_1_0_i_oswt_pff => vec_rsc_1_0_i_oswt_pff,
      vec_rsc_1_0_i_oswt_1_pff => vec_rsc_1_0_i_oswt_1_pff
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_1_0_i_wea_d_core_psct(0)));
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0)));
  vec_rsc_1_0_i_wea_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_wea_d_core_sct;
  vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_ctrl_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;

  inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_1_0_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp_inst_vec_rsc_1_0_i_da_d,
      vec_rsc_1_0_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp_inst_vec_rsc_1_0_i_qa_d,
      vec_rsc_1_0_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp_inst_vec_rsc_1_0_i_da_d_core,
      vec_rsc_1_0_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp_inst_vec_rsc_1_0_i_qa_d_mxwt,
      vec_rsc_1_0_i_biwt => vec_rsc_1_0_i_biwt,
      vec_rsc_1_0_i_bdwt => vec_rsc_1_0_i_bdwt,
      vec_rsc_1_0_i_biwt_1 => vec_rsc_1_0_i_biwt_1,
      vec_rsc_1_0_i_bdwt_2 => vec_rsc_1_0_i_bdwt_2
    );
  vec_rsc_1_0_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp_inst_vec_rsc_1_0_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp_inst_vec_rsc_1_0_i_qa_d
      <= vec_rsc_1_0_i_qa_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp_inst_vec_rsc_1_0_i_da_d_core
      <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000") & (vec_rsc_1_0_i_da_d_core(31
      DOWNTO 0));
  vec_rsc_1_0_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_vec_rsc_1_0_wait_dp_inst_vec_rsc_1_0_i_qa_d_mxwt;

  vec_rsc_1_0_i_wea_d <= vec_rsc_1_0_i_wea_d_core_sct;
  vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;
  vec_rsc_1_0_i_da_d <= vec_rsc_1_0_i_da_d_reg;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_7_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_0_7_i_oswt : IN STD_LOGIC;
    vec_rsc_0_7_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_0_7_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_0_7_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_0_7_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_7_i_biwt : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_bdwt : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_biwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_bdwt_2 : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_wea_d_core_sct : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_0_7_i_oswt : IN STD_LOGIC;
      vec_rsc_0_7_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_0_7_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_7_i_biwt : OUT STD_LOGIC;
      vec_rsc_0_7_i_bdwt : OUT STD_LOGIC;
      vec_rsc_0_7_i_biwt_1 : OUT STD_LOGIC;
      vec_rsc_0_7_i_bdwt_2 : OUT STD_LOGIC;
      vec_rsc_0_7_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_0_7_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_0_7_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_wea_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_0_7_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_7_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_7_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_7_i_biwt : IN STD_LOGIC;
      vec_rsc_0_7_i_bdwt : IN STD_LOGIC;
      vec_rsc_0_7_i_biwt_1 : IN STD_LOGIC;
      vec_rsc_0_7_i_bdwt_2 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp_inst_vec_rsc_0_7_i_da_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp_inst_vec_rsc_0_7_i_qa_d
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp_inst_vec_rsc_0_7_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp_inst_vec_rsc_0_7_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      vec_rsc_0_7_i_oswt => vec_rsc_0_7_i_oswt,
      vec_rsc_0_7_i_oswt_1 => vec_rsc_0_7_i_oswt_1,
      vec_rsc_0_7_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_wea_d_core_psct,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      vec_rsc_0_7_i_biwt => vec_rsc_0_7_i_biwt,
      vec_rsc_0_7_i_bdwt => vec_rsc_0_7_i_bdwt,
      vec_rsc_0_7_i_biwt_1 => vec_rsc_0_7_i_biwt_1,
      vec_rsc_0_7_i_bdwt_2 => vec_rsc_0_7_i_bdwt_2,
      vec_rsc_0_7_i_wea_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_wea_d_core_sct,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct,
      core_wten_pff => core_wten_pff,
      vec_rsc_0_7_i_oswt_pff => vec_rsc_0_7_i_oswt_pff,
      vec_rsc_0_7_i_oswt_1_pff => vec_rsc_0_7_i_oswt_1_pff
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_0_7_i_wea_d_core_psct(0)));
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0)));
  vec_rsc_0_7_i_wea_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_wea_d_core_sct;
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_ctrl_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;

  inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_0_7_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp_inst_vec_rsc_0_7_i_da_d,
      vec_rsc_0_7_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp_inst_vec_rsc_0_7_i_qa_d,
      vec_rsc_0_7_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp_inst_vec_rsc_0_7_i_da_d_core,
      vec_rsc_0_7_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp_inst_vec_rsc_0_7_i_qa_d_mxwt,
      vec_rsc_0_7_i_biwt => vec_rsc_0_7_i_biwt,
      vec_rsc_0_7_i_bdwt => vec_rsc_0_7_i_bdwt,
      vec_rsc_0_7_i_biwt_1 => vec_rsc_0_7_i_biwt_1,
      vec_rsc_0_7_i_bdwt_2 => vec_rsc_0_7_i_bdwt_2
    );
  vec_rsc_0_7_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp_inst_vec_rsc_0_7_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp_inst_vec_rsc_0_7_i_qa_d
      <= vec_rsc_0_7_i_qa_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp_inst_vec_rsc_0_7_i_da_d_core
      <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000") & (vec_rsc_0_7_i_da_d_core(31
      DOWNTO 0));
  vec_rsc_0_7_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_vec_rsc_0_7_wait_dp_inst_vec_rsc_0_7_i_qa_d_mxwt;

  vec_rsc_0_7_i_wea_d <= vec_rsc_0_7_i_wea_d_core_sct;
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;
  vec_rsc_0_7_i_da_d <= vec_rsc_0_7_i_da_d_reg;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_6_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_0_6_i_oswt : IN STD_LOGIC;
    vec_rsc_0_6_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_0_6_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_0_6_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_0_6_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_6_i_biwt : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_bdwt : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_biwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_bdwt_2 : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_wea_d_core_sct : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_0_6_i_oswt : IN STD_LOGIC;
      vec_rsc_0_6_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_0_6_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_6_i_biwt : OUT STD_LOGIC;
      vec_rsc_0_6_i_bdwt : OUT STD_LOGIC;
      vec_rsc_0_6_i_biwt_1 : OUT STD_LOGIC;
      vec_rsc_0_6_i_bdwt_2 : OUT STD_LOGIC;
      vec_rsc_0_6_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_0_6_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_0_6_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_wea_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_0_6_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_6_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_6_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_6_i_biwt : IN STD_LOGIC;
      vec_rsc_0_6_i_bdwt : IN STD_LOGIC;
      vec_rsc_0_6_i_biwt_1 : IN STD_LOGIC;
      vec_rsc_0_6_i_bdwt_2 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp_inst_vec_rsc_0_6_i_da_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp_inst_vec_rsc_0_6_i_qa_d
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp_inst_vec_rsc_0_6_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp_inst_vec_rsc_0_6_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      vec_rsc_0_6_i_oswt => vec_rsc_0_6_i_oswt,
      vec_rsc_0_6_i_oswt_1 => vec_rsc_0_6_i_oswt_1,
      vec_rsc_0_6_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_wea_d_core_psct,
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      vec_rsc_0_6_i_biwt => vec_rsc_0_6_i_biwt,
      vec_rsc_0_6_i_bdwt => vec_rsc_0_6_i_bdwt,
      vec_rsc_0_6_i_biwt_1 => vec_rsc_0_6_i_biwt_1,
      vec_rsc_0_6_i_bdwt_2 => vec_rsc_0_6_i_bdwt_2,
      vec_rsc_0_6_i_wea_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_wea_d_core_sct,
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct,
      core_wten_pff => core_wten_pff,
      vec_rsc_0_6_i_oswt_pff => vec_rsc_0_6_i_oswt_pff,
      vec_rsc_0_6_i_oswt_1_pff => vec_rsc_0_6_i_oswt_1_pff
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_0_6_i_wea_d_core_psct(0)));
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0)));
  vec_rsc_0_6_i_wea_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_wea_d_core_sct;
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_ctrl_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;

  inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_0_6_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp_inst_vec_rsc_0_6_i_da_d,
      vec_rsc_0_6_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp_inst_vec_rsc_0_6_i_qa_d,
      vec_rsc_0_6_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp_inst_vec_rsc_0_6_i_da_d_core,
      vec_rsc_0_6_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp_inst_vec_rsc_0_6_i_qa_d_mxwt,
      vec_rsc_0_6_i_biwt => vec_rsc_0_6_i_biwt,
      vec_rsc_0_6_i_bdwt => vec_rsc_0_6_i_bdwt,
      vec_rsc_0_6_i_biwt_1 => vec_rsc_0_6_i_biwt_1,
      vec_rsc_0_6_i_bdwt_2 => vec_rsc_0_6_i_bdwt_2
    );
  vec_rsc_0_6_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp_inst_vec_rsc_0_6_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp_inst_vec_rsc_0_6_i_qa_d
      <= vec_rsc_0_6_i_qa_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp_inst_vec_rsc_0_6_i_da_d_core
      <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000") & (vec_rsc_0_6_i_da_d_core(31
      DOWNTO 0));
  vec_rsc_0_6_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_vec_rsc_0_6_wait_dp_inst_vec_rsc_0_6_i_qa_d_mxwt;

  vec_rsc_0_6_i_wea_d <= vec_rsc_0_6_i_wea_d_core_sct;
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;
  vec_rsc_0_6_i_da_d <= vec_rsc_0_6_i_da_d_reg;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_5_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_0_5_i_oswt : IN STD_LOGIC;
    vec_rsc_0_5_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_0_5_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_0_5_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_0_5_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_5_i_biwt : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_bdwt : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_biwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_bdwt_2 : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_wea_d_core_sct : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_0_5_i_oswt : IN STD_LOGIC;
      vec_rsc_0_5_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_0_5_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_5_i_biwt : OUT STD_LOGIC;
      vec_rsc_0_5_i_bdwt : OUT STD_LOGIC;
      vec_rsc_0_5_i_biwt_1 : OUT STD_LOGIC;
      vec_rsc_0_5_i_bdwt_2 : OUT STD_LOGIC;
      vec_rsc_0_5_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_0_5_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_0_5_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_wea_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_0_5_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_5_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_5_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_5_i_biwt : IN STD_LOGIC;
      vec_rsc_0_5_i_bdwt : IN STD_LOGIC;
      vec_rsc_0_5_i_biwt_1 : IN STD_LOGIC;
      vec_rsc_0_5_i_bdwt_2 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp_inst_vec_rsc_0_5_i_da_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp_inst_vec_rsc_0_5_i_qa_d
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp_inst_vec_rsc_0_5_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp_inst_vec_rsc_0_5_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      vec_rsc_0_5_i_oswt => vec_rsc_0_5_i_oswt,
      vec_rsc_0_5_i_oswt_1 => vec_rsc_0_5_i_oswt_1,
      vec_rsc_0_5_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_wea_d_core_psct,
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      vec_rsc_0_5_i_biwt => vec_rsc_0_5_i_biwt,
      vec_rsc_0_5_i_bdwt => vec_rsc_0_5_i_bdwt,
      vec_rsc_0_5_i_biwt_1 => vec_rsc_0_5_i_biwt_1,
      vec_rsc_0_5_i_bdwt_2 => vec_rsc_0_5_i_bdwt_2,
      vec_rsc_0_5_i_wea_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_wea_d_core_sct,
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct,
      core_wten_pff => core_wten_pff,
      vec_rsc_0_5_i_oswt_pff => vec_rsc_0_5_i_oswt_pff,
      vec_rsc_0_5_i_oswt_1_pff => vec_rsc_0_5_i_oswt_1_pff
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_0_5_i_wea_d_core_psct(0)));
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0)));
  vec_rsc_0_5_i_wea_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_wea_d_core_sct;
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_ctrl_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;

  inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_0_5_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp_inst_vec_rsc_0_5_i_da_d,
      vec_rsc_0_5_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp_inst_vec_rsc_0_5_i_qa_d,
      vec_rsc_0_5_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp_inst_vec_rsc_0_5_i_da_d_core,
      vec_rsc_0_5_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp_inst_vec_rsc_0_5_i_qa_d_mxwt,
      vec_rsc_0_5_i_biwt => vec_rsc_0_5_i_biwt,
      vec_rsc_0_5_i_bdwt => vec_rsc_0_5_i_bdwt,
      vec_rsc_0_5_i_biwt_1 => vec_rsc_0_5_i_biwt_1,
      vec_rsc_0_5_i_bdwt_2 => vec_rsc_0_5_i_bdwt_2
    );
  vec_rsc_0_5_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp_inst_vec_rsc_0_5_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp_inst_vec_rsc_0_5_i_qa_d
      <= vec_rsc_0_5_i_qa_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp_inst_vec_rsc_0_5_i_da_d_core
      <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000") & (vec_rsc_0_5_i_da_d_core(31
      DOWNTO 0));
  vec_rsc_0_5_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_vec_rsc_0_5_wait_dp_inst_vec_rsc_0_5_i_qa_d_mxwt;

  vec_rsc_0_5_i_wea_d <= vec_rsc_0_5_i_wea_d_core_sct;
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;
  vec_rsc_0_5_i_da_d <= vec_rsc_0_5_i_da_d_reg;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_4_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_0_4_i_oswt : IN STD_LOGIC;
    vec_rsc_0_4_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_0_4_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_0_4_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_0_4_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_4_i_biwt : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_bdwt : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_biwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_bdwt_2 : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_wea_d_core_sct : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_0_4_i_oswt : IN STD_LOGIC;
      vec_rsc_0_4_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_0_4_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_4_i_biwt : OUT STD_LOGIC;
      vec_rsc_0_4_i_bdwt : OUT STD_LOGIC;
      vec_rsc_0_4_i_biwt_1 : OUT STD_LOGIC;
      vec_rsc_0_4_i_bdwt_2 : OUT STD_LOGIC;
      vec_rsc_0_4_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_0_4_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_0_4_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_wea_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_0_4_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_4_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_4_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_4_i_biwt : IN STD_LOGIC;
      vec_rsc_0_4_i_bdwt : IN STD_LOGIC;
      vec_rsc_0_4_i_biwt_1 : IN STD_LOGIC;
      vec_rsc_0_4_i_bdwt_2 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp_inst_vec_rsc_0_4_i_da_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp_inst_vec_rsc_0_4_i_qa_d
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp_inst_vec_rsc_0_4_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp_inst_vec_rsc_0_4_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      vec_rsc_0_4_i_oswt => vec_rsc_0_4_i_oswt,
      vec_rsc_0_4_i_oswt_1 => vec_rsc_0_4_i_oswt_1,
      vec_rsc_0_4_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_wea_d_core_psct,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      vec_rsc_0_4_i_biwt => vec_rsc_0_4_i_biwt,
      vec_rsc_0_4_i_bdwt => vec_rsc_0_4_i_bdwt,
      vec_rsc_0_4_i_biwt_1 => vec_rsc_0_4_i_biwt_1,
      vec_rsc_0_4_i_bdwt_2 => vec_rsc_0_4_i_bdwt_2,
      vec_rsc_0_4_i_wea_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_wea_d_core_sct,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct,
      core_wten_pff => core_wten_pff,
      vec_rsc_0_4_i_oswt_pff => vec_rsc_0_4_i_oswt_pff,
      vec_rsc_0_4_i_oswt_1_pff => vec_rsc_0_4_i_oswt_1_pff
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_0_4_i_wea_d_core_psct(0)));
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0)));
  vec_rsc_0_4_i_wea_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_wea_d_core_sct;
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_ctrl_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;

  inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_0_4_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp_inst_vec_rsc_0_4_i_da_d,
      vec_rsc_0_4_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp_inst_vec_rsc_0_4_i_qa_d,
      vec_rsc_0_4_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp_inst_vec_rsc_0_4_i_da_d_core,
      vec_rsc_0_4_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp_inst_vec_rsc_0_4_i_qa_d_mxwt,
      vec_rsc_0_4_i_biwt => vec_rsc_0_4_i_biwt,
      vec_rsc_0_4_i_bdwt => vec_rsc_0_4_i_bdwt,
      vec_rsc_0_4_i_biwt_1 => vec_rsc_0_4_i_biwt_1,
      vec_rsc_0_4_i_bdwt_2 => vec_rsc_0_4_i_bdwt_2
    );
  vec_rsc_0_4_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp_inst_vec_rsc_0_4_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp_inst_vec_rsc_0_4_i_qa_d
      <= vec_rsc_0_4_i_qa_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp_inst_vec_rsc_0_4_i_da_d_core
      <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000") & (vec_rsc_0_4_i_da_d_core(31
      DOWNTO 0));
  vec_rsc_0_4_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_vec_rsc_0_4_wait_dp_inst_vec_rsc_0_4_i_qa_d_mxwt;

  vec_rsc_0_4_i_wea_d <= vec_rsc_0_4_i_wea_d_core_sct;
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;
  vec_rsc_0_4_i_da_d <= vec_rsc_0_4_i_da_d_reg;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_3_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_0_3_i_oswt : IN STD_LOGIC;
    vec_rsc_0_3_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_0_3_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_0_3_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_0_3_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_3_i_biwt : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_bdwt : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_biwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_bdwt_2 : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_wea_d_core_sct : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_0_3_i_oswt : IN STD_LOGIC;
      vec_rsc_0_3_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_0_3_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_3_i_biwt : OUT STD_LOGIC;
      vec_rsc_0_3_i_bdwt : OUT STD_LOGIC;
      vec_rsc_0_3_i_biwt_1 : OUT STD_LOGIC;
      vec_rsc_0_3_i_bdwt_2 : OUT STD_LOGIC;
      vec_rsc_0_3_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_0_3_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_0_3_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_wea_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_0_3_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_3_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_3_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_3_i_biwt : IN STD_LOGIC;
      vec_rsc_0_3_i_bdwt : IN STD_LOGIC;
      vec_rsc_0_3_i_biwt_1 : IN STD_LOGIC;
      vec_rsc_0_3_i_bdwt_2 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp_inst_vec_rsc_0_3_i_da_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp_inst_vec_rsc_0_3_i_qa_d
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp_inst_vec_rsc_0_3_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp_inst_vec_rsc_0_3_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      vec_rsc_0_3_i_oswt => vec_rsc_0_3_i_oswt,
      vec_rsc_0_3_i_oswt_1 => vec_rsc_0_3_i_oswt_1,
      vec_rsc_0_3_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_wea_d_core_psct,
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      vec_rsc_0_3_i_biwt => vec_rsc_0_3_i_biwt,
      vec_rsc_0_3_i_bdwt => vec_rsc_0_3_i_bdwt,
      vec_rsc_0_3_i_biwt_1 => vec_rsc_0_3_i_biwt_1,
      vec_rsc_0_3_i_bdwt_2 => vec_rsc_0_3_i_bdwt_2,
      vec_rsc_0_3_i_wea_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_wea_d_core_sct,
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct,
      core_wten_pff => core_wten_pff,
      vec_rsc_0_3_i_oswt_pff => vec_rsc_0_3_i_oswt_pff,
      vec_rsc_0_3_i_oswt_1_pff => vec_rsc_0_3_i_oswt_1_pff
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_0_3_i_wea_d_core_psct(0)));
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0)));
  vec_rsc_0_3_i_wea_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_wea_d_core_sct;
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_ctrl_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;

  inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_0_3_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp_inst_vec_rsc_0_3_i_da_d,
      vec_rsc_0_3_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp_inst_vec_rsc_0_3_i_qa_d,
      vec_rsc_0_3_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp_inst_vec_rsc_0_3_i_da_d_core,
      vec_rsc_0_3_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp_inst_vec_rsc_0_3_i_qa_d_mxwt,
      vec_rsc_0_3_i_biwt => vec_rsc_0_3_i_biwt,
      vec_rsc_0_3_i_bdwt => vec_rsc_0_3_i_bdwt,
      vec_rsc_0_3_i_biwt_1 => vec_rsc_0_3_i_biwt_1,
      vec_rsc_0_3_i_bdwt_2 => vec_rsc_0_3_i_bdwt_2
    );
  vec_rsc_0_3_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp_inst_vec_rsc_0_3_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp_inst_vec_rsc_0_3_i_qa_d
      <= vec_rsc_0_3_i_qa_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp_inst_vec_rsc_0_3_i_da_d_core
      <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000") & (vec_rsc_0_3_i_da_d_core(31
      DOWNTO 0));
  vec_rsc_0_3_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_vec_rsc_0_3_wait_dp_inst_vec_rsc_0_3_i_qa_d_mxwt;

  vec_rsc_0_3_i_wea_d <= vec_rsc_0_3_i_wea_d_core_sct;
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;
  vec_rsc_0_3_i_da_d <= vec_rsc_0_3_i_da_d_reg;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_2_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_0_2_i_oswt : IN STD_LOGIC;
    vec_rsc_0_2_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_0_2_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_0_2_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_0_2_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_2_i_biwt : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_bdwt : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_biwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_bdwt_2 : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_wea_d_core_sct : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_0_2_i_oswt : IN STD_LOGIC;
      vec_rsc_0_2_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_0_2_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_2_i_biwt : OUT STD_LOGIC;
      vec_rsc_0_2_i_bdwt : OUT STD_LOGIC;
      vec_rsc_0_2_i_biwt_1 : OUT STD_LOGIC;
      vec_rsc_0_2_i_bdwt_2 : OUT STD_LOGIC;
      vec_rsc_0_2_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_0_2_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_0_2_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_wea_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_0_2_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_2_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_2_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_2_i_biwt : IN STD_LOGIC;
      vec_rsc_0_2_i_bdwt : IN STD_LOGIC;
      vec_rsc_0_2_i_biwt_1 : IN STD_LOGIC;
      vec_rsc_0_2_i_bdwt_2 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp_inst_vec_rsc_0_2_i_da_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp_inst_vec_rsc_0_2_i_qa_d
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp_inst_vec_rsc_0_2_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp_inst_vec_rsc_0_2_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      vec_rsc_0_2_i_oswt => vec_rsc_0_2_i_oswt,
      vec_rsc_0_2_i_oswt_1 => vec_rsc_0_2_i_oswt_1,
      vec_rsc_0_2_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_wea_d_core_psct,
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      vec_rsc_0_2_i_biwt => vec_rsc_0_2_i_biwt,
      vec_rsc_0_2_i_bdwt => vec_rsc_0_2_i_bdwt,
      vec_rsc_0_2_i_biwt_1 => vec_rsc_0_2_i_biwt_1,
      vec_rsc_0_2_i_bdwt_2 => vec_rsc_0_2_i_bdwt_2,
      vec_rsc_0_2_i_wea_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_wea_d_core_sct,
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct,
      core_wten_pff => core_wten_pff,
      vec_rsc_0_2_i_oswt_pff => vec_rsc_0_2_i_oswt_pff,
      vec_rsc_0_2_i_oswt_1_pff => vec_rsc_0_2_i_oswt_1_pff
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_0_2_i_wea_d_core_psct(0)));
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0)));
  vec_rsc_0_2_i_wea_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_wea_d_core_sct;
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_ctrl_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;

  inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_0_2_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp_inst_vec_rsc_0_2_i_da_d,
      vec_rsc_0_2_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp_inst_vec_rsc_0_2_i_qa_d,
      vec_rsc_0_2_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp_inst_vec_rsc_0_2_i_da_d_core,
      vec_rsc_0_2_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp_inst_vec_rsc_0_2_i_qa_d_mxwt,
      vec_rsc_0_2_i_biwt => vec_rsc_0_2_i_biwt,
      vec_rsc_0_2_i_bdwt => vec_rsc_0_2_i_bdwt,
      vec_rsc_0_2_i_biwt_1 => vec_rsc_0_2_i_biwt_1,
      vec_rsc_0_2_i_bdwt_2 => vec_rsc_0_2_i_bdwt_2
    );
  vec_rsc_0_2_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp_inst_vec_rsc_0_2_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp_inst_vec_rsc_0_2_i_qa_d
      <= vec_rsc_0_2_i_qa_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp_inst_vec_rsc_0_2_i_da_d_core
      <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000") & (vec_rsc_0_2_i_da_d_core(31
      DOWNTO 0));
  vec_rsc_0_2_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_vec_rsc_0_2_wait_dp_inst_vec_rsc_0_2_i_qa_d_mxwt;

  vec_rsc_0_2_i_wea_d <= vec_rsc_0_2_i_wea_d_core_sct;
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;
  vec_rsc_0_2_i_da_d <= vec_rsc_0_2_i_da_d_reg;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_1_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_0_1_i_oswt : IN STD_LOGIC;
    vec_rsc_0_1_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_0_1_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_0_1_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_0_1_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_1_i_biwt : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_bdwt : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_biwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_bdwt_2 : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_wea_d_core_sct : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_0_1_i_oswt : IN STD_LOGIC;
      vec_rsc_0_1_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_0_1_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_1_i_biwt : OUT STD_LOGIC;
      vec_rsc_0_1_i_bdwt : OUT STD_LOGIC;
      vec_rsc_0_1_i_biwt_1 : OUT STD_LOGIC;
      vec_rsc_0_1_i_bdwt_2 : OUT STD_LOGIC;
      vec_rsc_0_1_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_0_1_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_0_1_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_wea_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_0_1_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_1_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_1_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_1_i_biwt : IN STD_LOGIC;
      vec_rsc_0_1_i_bdwt : IN STD_LOGIC;
      vec_rsc_0_1_i_biwt_1 : IN STD_LOGIC;
      vec_rsc_0_1_i_bdwt_2 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp_inst_vec_rsc_0_1_i_da_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp_inst_vec_rsc_0_1_i_qa_d
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp_inst_vec_rsc_0_1_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp_inst_vec_rsc_0_1_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      vec_rsc_0_1_i_oswt => vec_rsc_0_1_i_oswt,
      vec_rsc_0_1_i_oswt_1 => vec_rsc_0_1_i_oswt_1,
      vec_rsc_0_1_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_wea_d_core_psct,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      vec_rsc_0_1_i_biwt => vec_rsc_0_1_i_biwt,
      vec_rsc_0_1_i_bdwt => vec_rsc_0_1_i_bdwt,
      vec_rsc_0_1_i_biwt_1 => vec_rsc_0_1_i_biwt_1,
      vec_rsc_0_1_i_bdwt_2 => vec_rsc_0_1_i_bdwt_2,
      vec_rsc_0_1_i_wea_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_wea_d_core_sct,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct,
      core_wten_pff => core_wten_pff,
      vec_rsc_0_1_i_oswt_pff => vec_rsc_0_1_i_oswt_pff,
      vec_rsc_0_1_i_oswt_1_pff => vec_rsc_0_1_i_oswt_1_pff
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_0_1_i_wea_d_core_psct(0)));
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0)));
  vec_rsc_0_1_i_wea_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_wea_d_core_sct;
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_ctrl_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;

  inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_0_1_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp_inst_vec_rsc_0_1_i_da_d,
      vec_rsc_0_1_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp_inst_vec_rsc_0_1_i_qa_d,
      vec_rsc_0_1_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp_inst_vec_rsc_0_1_i_da_d_core,
      vec_rsc_0_1_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp_inst_vec_rsc_0_1_i_qa_d_mxwt,
      vec_rsc_0_1_i_biwt => vec_rsc_0_1_i_biwt,
      vec_rsc_0_1_i_bdwt => vec_rsc_0_1_i_bdwt,
      vec_rsc_0_1_i_biwt_1 => vec_rsc_0_1_i_biwt_1,
      vec_rsc_0_1_i_bdwt_2 => vec_rsc_0_1_i_bdwt_2
    );
  vec_rsc_0_1_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp_inst_vec_rsc_0_1_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp_inst_vec_rsc_0_1_i_qa_d
      <= vec_rsc_0_1_i_qa_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp_inst_vec_rsc_0_1_i_da_d_core
      <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000") & (vec_rsc_0_1_i_da_d_core(31
      DOWNTO 0));
  vec_rsc_0_1_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_vec_rsc_0_1_wait_dp_inst_vec_rsc_0_1_i_qa_d_mxwt;

  vec_rsc_0_1_i_wea_d <= vec_rsc_0_1_i_wea_d_core_sct;
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;
  vec_rsc_0_1_i_da_d <= vec_rsc_0_1_i_da_d_reg;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_0_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    vec_rsc_0_0_i_oswt : IN STD_LOGIC;
    vec_rsc_0_0_i_oswt_1 : IN STD_LOGIC;
    vec_rsc_0_0_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
        (1 DOWNTO 0);
    core_wten_pff : IN STD_LOGIC;
    vec_rsc_0_0_i_oswt_pff : IN STD_LOGIC;
    vec_rsc_0_0_i_oswt_1_pff : IN STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1 IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_0_i_biwt : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_bdwt : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_biwt_1 : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_wea_d_core_sct : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_0_0_i_oswt : IN STD_LOGIC;
      vec_rsc_0_0_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_0_0_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_0_i_biwt : OUT STD_LOGIC;
      vec_rsc_0_0_i_bdwt : OUT STD_LOGIC;
      vec_rsc_0_0_i_biwt_1 : OUT STD_LOGIC;
      vec_rsc_0_0_i_bdwt_2 : OUT STD_LOGIC;
      vec_rsc_0_0_i_wea_d_core_sct : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct : OUT STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_0_0_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_0_0_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_wea_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_0_0_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_biwt : IN STD_LOGIC;
      vec_rsc_0_0_i_bdwt : IN STD_LOGIC;
      vec_rsc_0_0_i_biwt_1 : IN STD_LOGIC;
      vec_rsc_0_0_i_bdwt_2 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp_inst_vec_rsc_0_0_i_da_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp_inst_vec_rsc_0_0_i_qa_d
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp_inst_vec_rsc_0_0_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp_inst_vec_rsc_0_0_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      vec_rsc_0_0_i_oswt => vec_rsc_0_0_i_oswt,
      vec_rsc_0_0_i_oswt_1 => vec_rsc_0_0_i_oswt_1,
      vec_rsc_0_0_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_wea_d_core_psct,
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      vec_rsc_0_0_i_biwt => vec_rsc_0_0_i_biwt,
      vec_rsc_0_0_i_bdwt => vec_rsc_0_0_i_bdwt,
      vec_rsc_0_0_i_biwt_1 => vec_rsc_0_0_i_biwt_1,
      vec_rsc_0_0_i_bdwt_2 => vec_rsc_0_0_i_bdwt_2,
      vec_rsc_0_0_i_wea_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_wea_d_core_sct,
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct,
      core_wten_pff => core_wten_pff,
      vec_rsc_0_0_i_oswt_pff => vec_rsc_0_0_i_oswt_pff,
      vec_rsc_0_0_i_oswt_1_pff => vec_rsc_0_0_i_oswt_1_pff
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_0_0_i_wea_d_core_psct(0)));
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & (vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct(0)));
  vec_rsc_0_0_i_wea_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_wea_d_core_sct;
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_ctrl_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;

  inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_0_0_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp_inst_vec_rsc_0_0_i_da_d,
      vec_rsc_0_0_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp_inst_vec_rsc_0_0_i_qa_d,
      vec_rsc_0_0_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp_inst_vec_rsc_0_0_i_da_d_core,
      vec_rsc_0_0_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp_inst_vec_rsc_0_0_i_qa_d_mxwt,
      vec_rsc_0_0_i_biwt => vec_rsc_0_0_i_biwt,
      vec_rsc_0_0_i_bdwt => vec_rsc_0_0_i_bdwt,
      vec_rsc_0_0_i_biwt_1 => vec_rsc_0_0_i_biwt_1,
      vec_rsc_0_0_i_bdwt_2 => vec_rsc_0_0_i_bdwt_2
    );
  vec_rsc_0_0_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp_inst_vec_rsc_0_0_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp_inst_vec_rsc_0_0_i_qa_d
      <= vec_rsc_0_0_i_qa_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp_inst_vec_rsc_0_0_i_da_d_core
      <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000") & (vec_rsc_0_0_i_da_d_core(31
      DOWNTO 0));
  vec_rsc_0_0_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_vec_rsc_0_0_wait_dp_inst_vec_rsc_0_0_i_qa_d_mxwt;

  vec_rsc_0_0_i_wea_d <= vec_rsc_0_0_i_wea_d_core_sct;
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_sct;
  vec_rsc_0_0_i_da_d <= vec_rsc_0_0_i_da_d_reg;
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_complete_rsci
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_complete_rsci IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    complete_rsc_rdy : IN STD_LOGIC;
    complete_rsc_vld : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    complete_rsci_oswt : IN STD_LOGIC;
    complete_rsci_wen_comp : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_complete_rsci;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_complete_rsci IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL complete_rsci_biwt : STD_LOGIC;
  SIGNAL complete_rsci_bdwt : STD_LOGIC;
  SIGNAL complete_rsci_bcwt : STD_LOGIC;
  SIGNAL complete_rsci_ivld_core_sct : STD_LOGIC;
  SIGNAL complete_rsci_irdy : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_complete_rsci_complete_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      complete_rsci_oswt : IN STD_LOGIC;
      complete_rsci_biwt : OUT STD_LOGIC;
      complete_rsci_bdwt : OUT STD_LOGIC;
      complete_rsci_bcwt : IN STD_LOGIC;
      complete_rsci_ivld_core_sct : OUT STD_LOGIC;
      complete_rsci_irdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_complete_rsci_complete_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      complete_rsci_oswt : IN STD_LOGIC;
      complete_rsci_wen_comp : OUT STD_LOGIC;
      complete_rsci_biwt : IN STD_LOGIC;
      complete_rsci_bdwt : IN STD_LOGIC;
      complete_rsci_bcwt : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  complete_rsci : work.ccs_sync_out_wait_pkg_v1.ccs_sync_out_wait_v1
    GENERIC MAP(
      rscid => 18
      )
    PORT MAP(
      vld => complete_rsc_vld,
      rdy => complete_rsc_rdy,
      ivld => complete_rsci_ivld_core_sct,
      irdy => complete_rsci_irdy
    );
  inPlaceNTT_DIF_precomp_core_complete_rsci_complete_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_complete_rsci_complete_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      complete_rsci_oswt => complete_rsci_oswt,
      complete_rsci_biwt => complete_rsci_biwt,
      complete_rsci_bdwt => complete_rsci_bdwt,
      complete_rsci_bcwt => complete_rsci_bcwt,
      complete_rsci_ivld_core_sct => complete_rsci_ivld_core_sct,
      complete_rsci_irdy => complete_rsci_irdy
    );
  inPlaceNTT_DIF_precomp_core_complete_rsci_complete_wait_dp_inst : inPlaceNTT_DIF_precomp_core_complete_rsci_complete_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      complete_rsci_oswt => complete_rsci_oswt,
      complete_rsci_wen_comp => complete_rsci_wen_comp,
      complete_rsci_biwt => complete_rsci_biwt,
      complete_rsci_bdwt => complete_rsci_bdwt,
      complete_rsci_bcwt => complete_rsci_bcwt
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core_run_rsci
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core_run_rsci IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    run_rsc_rdy : OUT STD_LOGIC;
    run_rsc_vld : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    run_rsci_oswt : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    run_rsci_ivld_mxwt : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp_core_run_rsci;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core_run_rsci IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL run_rsci_ivld : STD_LOGIC;
  SIGNAL run_rsci_biwt : STD_LOGIC;
  SIGNAL run_rsci_bdwt : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_run_rsci_run_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      run_rsci_oswt : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      run_rsci_biwt : OUT STD_LOGIC;
      run_rsci_bdwt : OUT STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_run_rsci_run_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      run_rsci_ivld_mxwt : OUT STD_LOGIC;
      run_rsci_ivld : IN STD_LOGIC;
      run_rsci_biwt : IN STD_LOGIC;
      run_rsci_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
BEGIN
  run_rsci : work.ccs_sync_in_wait_pkg_v1.ccs_sync_in_wait_v1
    GENERIC MAP(
      rscid => 12
      )
    PORT MAP(
      vld => run_rsc_vld,
      rdy => run_rsc_rdy,
      ivld => run_rsci_ivld,
      irdy => run_rsci_biwt
    );
  inPlaceNTT_DIF_precomp_core_run_rsci_run_wait_ctrl_inst : inPlaceNTT_DIF_precomp_core_run_rsci_run_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      run_rsci_oswt => run_rsci_oswt,
      core_wten => core_wten,
      run_rsci_biwt => run_rsci_biwt,
      run_rsci_bdwt => run_rsci_bdwt
    );
  inPlaceNTT_DIF_precomp_core_run_rsci_run_wait_dp_inst : inPlaceNTT_DIF_precomp_core_run_rsci_run_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      run_rsci_ivld_mxwt => run_rsci_ivld_mxwt,
      run_rsci_ivld => run_rsci_ivld,
      run_rsci_biwt => run_rsci_biwt,
      run_rsci_bdwt => run_rsci_bdwt
    );
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    run_rsc_rdy : OUT STD_LOGIC;
    run_rsc_vld : IN STD_LOGIC;
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    vec_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    vec_rsc_triosy_1_1_lz : OUT STD_LOGIC;
    vec_rsc_triosy_1_2_lz : OUT STD_LOGIC;
    vec_rsc_triosy_1_3_lz : OUT STD_LOGIC;
    vec_rsc_triosy_1_4_lz : OUT STD_LOGIC;
    vec_rsc_triosy_1_5_lz : OUT STD_LOGIC;
    vec_rsc_triosy_1_6_lz : OUT STD_LOGIC;
    vec_rsc_triosy_1_7_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_1_1_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_1_2_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_1_3_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_1_4_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_1_5_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_1_6_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_1_7_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_1_1_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_1_2_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_1_3_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_1_4_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_1_5_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_1_6_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_1_7_lz : OUT STD_LOGIC;
    complete_rsc_rdy : IN STD_LOGIC;
    complete_rsc_vld : OUT STD_LOGIC;
    vec_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    vec_rsc_0_0_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_1_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    vec_rsc_0_1_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_2_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    vec_rsc_0_2_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_3_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    vec_rsc_0_3_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_4_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    vec_rsc_0_4_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_5_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    vec_rsc_0_5_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_6_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    vec_rsc_0_6_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_7_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    vec_rsc_0_7_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_0_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    vec_rsc_1_0_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_1_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    vec_rsc_1_1_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_1_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_2_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    vec_rsc_1_2_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_2_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_3_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    vec_rsc_1_3_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_3_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_4_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    vec_rsc_1_4_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_4_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_5_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    vec_rsc_1_5_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_5_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_6_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    vec_rsc_1_6_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_6_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_7_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    vec_rsc_1_7_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_1_7_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    twiddle_rsc_0_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_1_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_1_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_1_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_1_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_1_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_1_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_1_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_1_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsc_1_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsc_1_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsc_1_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsc_1_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsc_1_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsc_1_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsc_1_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsc_1_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_0_i_adrb_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0)
  );
END inPlaceNTT_DIF_precomp_core;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL core_wten : STD_LOGIC;
  SIGNAL run_rsci_ivld_mxwt : STD_LOGIC;
  SIGNAL p_rsci_idat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL complete_rsci_wen_comp : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_qa_d_mxwt : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_qa_d_mxwt : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_qa_d_mxwt : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_qa_d_mxwt : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_qa_d_mxwt : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_qa_d_mxwt : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_qa_d_mxwt : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_qa_d_mxwt : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_qa_d_mxwt : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_qa_d_mxwt : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_qa_d_mxwt : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_qa_d_mxwt : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_qa_d_mxwt : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_qa_d_mxwt : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_qa_d_mxwt : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_qa_d_mxwt : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_0_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_1_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_2_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_3_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_4_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_5_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_6_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_7_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_0_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_1_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_2_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_3_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_4_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_5_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_6_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_7_i_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_cmp_return_rsc_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_cmp_ccs_ccore_en : STD_LOGIC;
  SIGNAL modulo_sub_cmp_return_rsc_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_cmp_ccs_ccore_en : STD_LOGIC;
  SIGNAL modulo_add_cmp_return_rsc_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL fsm_output : STD_LOGIC_VECTOR (21 DOWNTO 0);
  SIGNAL VEC_LOOP_acc_10_tmp : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL VEC_LOOP_acc_1_tmp : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL and_dcpl_7 : STD_LOGIC;
  SIGNAL and_dcpl_8 : STD_LOGIC;
  SIGNAL and_dcpl_13 : STD_LOGIC;
  SIGNAL and_dcpl_14 : STD_LOGIC;
  SIGNAL and_dcpl_19 : STD_LOGIC;
  SIGNAL and_dcpl_21 : STD_LOGIC;
  SIGNAL and_dcpl_23 : STD_LOGIC;
  SIGNAL and_dcpl_25 : STD_LOGIC;
  SIGNAL and_dcpl_27 : STD_LOGIC;
  SIGNAL and_dcpl_29 : STD_LOGIC;
  SIGNAL and_dcpl_31 : STD_LOGIC;
  SIGNAL and_dcpl_33 : STD_LOGIC;
  SIGNAL and_dcpl_35 : STD_LOGIC;
  SIGNAL and_dcpl_37 : STD_LOGIC;
  SIGNAL and_dcpl_39 : STD_LOGIC;
  SIGNAL and_dcpl_41 : STD_LOGIC;
  SIGNAL and_dcpl_43 : STD_LOGIC;
  SIGNAL and_dcpl_45 : STD_LOGIC;
  SIGNAL and_dcpl_47 : STD_LOGIC;
  SIGNAL and_dcpl_49 : STD_LOGIC;
  SIGNAL and_dcpl_63 : STD_LOGIC;
  SIGNAL and_dcpl_65 : STD_LOGIC;
  SIGNAL and_dcpl_67 : STD_LOGIC;
  SIGNAL and_dcpl_69 : STD_LOGIC;
  SIGNAL and_dcpl_83 : STD_LOGIC;
  SIGNAL and_dcpl_85 : STD_LOGIC;
  SIGNAL and_dcpl_87 : STD_LOGIC;
  SIGNAL and_dcpl_89 : STD_LOGIC;
  SIGNAL and_dcpl_103 : STD_LOGIC;
  SIGNAL and_dcpl_104 : STD_LOGIC;
  SIGNAL and_dcpl_106 : STD_LOGIC;
  SIGNAL and_dcpl_108 : STD_LOGIC;
  SIGNAL and_dcpl_110 : STD_LOGIC;
  SIGNAL and_dcpl_112 : STD_LOGIC;
  SIGNAL and_dcpl_117 : STD_LOGIC;
  SIGNAL and_dcpl_122 : STD_LOGIC;
  SIGNAL and_dcpl_129 : STD_LOGIC;
  SIGNAL and_dcpl_131 : STD_LOGIC;
  SIGNAL or_tmp_141 : STD_LOGIC;
  SIGNAL and_157_cse : STD_LOGIC;
  SIGNAL and_159_cse : STD_LOGIC;
  SIGNAL and_158_cse : STD_LOGIC;
  SIGNAL and_178_cse : STD_LOGIC;
  SIGNAL and_180_cse : STD_LOGIC;
  SIGNAL and_179_cse : STD_LOGIC;
  SIGNAL and_191_cse : STD_LOGIC;
  SIGNAL and_193_cse : STD_LOGIC;
  SIGNAL and_192_cse : STD_LOGIC;
  SIGNAL and_204_cse : STD_LOGIC;
  SIGNAL and_206_cse : STD_LOGIC;
  SIGNAL and_205_cse : STD_LOGIC;
  SIGNAL and_217_cse : STD_LOGIC;
  SIGNAL and_219_cse : STD_LOGIC;
  SIGNAL and_218_cse : STD_LOGIC;
  SIGNAL and_230_cse : STD_LOGIC;
  SIGNAL and_232_cse : STD_LOGIC;
  SIGNAL and_231_cse : STD_LOGIC;
  SIGNAL and_243_cse : STD_LOGIC;
  SIGNAL and_245_cse : STD_LOGIC;
  SIGNAL and_244_cse : STD_LOGIC;
  SIGNAL and_256_cse : STD_LOGIC;
  SIGNAL and_258_cse : STD_LOGIC;
  SIGNAL and_257_cse : STD_LOGIC;
  SIGNAL and_269_cse : STD_LOGIC;
  SIGNAL and_271_cse : STD_LOGIC;
  SIGNAL and_270_cse : STD_LOGIC;
  SIGNAL and_282_cse : STD_LOGIC;
  SIGNAL and_284_cse : STD_LOGIC;
  SIGNAL and_283_cse : STD_LOGIC;
  SIGNAL and_295_cse : STD_LOGIC;
  SIGNAL and_297_cse : STD_LOGIC;
  SIGNAL and_296_cse : STD_LOGIC;
  SIGNAL and_308_cse : STD_LOGIC;
  SIGNAL and_310_cse : STD_LOGIC;
  SIGNAL and_309_cse : STD_LOGIC;
  SIGNAL and_321_cse : STD_LOGIC;
  SIGNAL and_323_cse : STD_LOGIC;
  SIGNAL and_322_cse : STD_LOGIC;
  SIGNAL and_334_cse : STD_LOGIC;
  SIGNAL and_336_cse : STD_LOGIC;
  SIGNAL and_335_cse : STD_LOGIC;
  SIGNAL and_347_cse : STD_LOGIC;
  SIGNAL and_349_cse : STD_LOGIC;
  SIGNAL and_348_cse : STD_LOGIC;
  SIGNAL and_360_cse : STD_LOGIC;
  SIGNAL and_362_cse : STD_LOGIC;
  SIGNAL and_361_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_lshift_itm : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_psp_sva : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_twiddle_f_mul_cse_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_twiddle_f_nor_6_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_nor_3_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_nor_1_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_nor_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_k_10_0_sva_9_0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL VEC_LOOP_j_10_0_sva_1 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL VEC_LOOP_VEC_LOOP_and_10_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_acc_10_cse_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL reg_run_rsci_oswt_cse : STD_LOGIC;
  SIGNAL reg_complete_rsci_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_0_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_0_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_0_1_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_0_1_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_0_2_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_0_2_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_0_3_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_0_3_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_0_4_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_0_4_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_0_5_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_0_5_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_0_6_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_0_6_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_0_7_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_0_7_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_1_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_1_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_1_1_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_1_1_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_1_2_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_1_2_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_1_3_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_1_3_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_1_4_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_1_4_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_1_5_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_1_5_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_1_6_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_1_6_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_1_7_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_1_7_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_1_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_2_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_3_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_4_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_5_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_6_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_7_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_1_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_1_1_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_1_2_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_1_3_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_1_4_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_1_5_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_1_6_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_1_7_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_triosy_1_7_obj_iswt0_cse : STD_LOGIC;
  SIGNAL reg_ensig_cgo_cse : STD_LOGIC;
  SIGNAL reg_ensig_cgo_1_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_and_1_cse : STD_LOGIC;
  SIGNAL VEC_LOOP_and_cse : STD_LOGIC;
  SIGNAL VEC_LOOP_nor_9_cse : STD_LOGIC;
  SIGNAL VEC_LOOP_nor_2_cse : STD_LOGIC;
  SIGNAL VEC_LOOP_nor_19_cse : STD_LOGIC;
  SIGNAL VEC_LOOP_nor_12_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_help_and_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_help_and_1_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_help_and_2_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_help_and_3_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_help_and_4_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_help_and_5_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_help_and_6_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_help_and_7_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_help_and_8_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_help_and_9_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_help_and_10_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_help_and_11_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_help_and_12_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_help_and_13_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_help_and_14_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_help_and_15_cse : STD_LOGIC;
  SIGNAL VEC_LOOP_mux1h_rmff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL VEC_LOOP_mux_4_rmff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wea_d_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL or_21_rmff : STD_LOGIC;
  SIGNAL core_wten_iff : STD_LOGIC;
  SIGNAL or_15_rmff : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL and_161_rmff : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_wea_d_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL or_26_rmff : STD_LOGIC;
  SIGNAL or_24_rmff : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL and_182_rmff : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_wea_d_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL or_31_rmff : STD_LOGIC;
  SIGNAL or_29_rmff : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL and_195_rmff : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_wea_d_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL or_36_rmff : STD_LOGIC;
  SIGNAL or_34_rmff : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL and_208_rmff : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_wea_d_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL or_41_rmff : STD_LOGIC;
  SIGNAL or_39_rmff : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL and_221_rmff : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_wea_d_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL or_46_rmff : STD_LOGIC;
  SIGNAL or_44_rmff : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL and_234_rmff : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_wea_d_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL or_51_rmff : STD_LOGIC;
  SIGNAL or_49_rmff : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL and_247_rmff : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_wea_d_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL or_56_rmff : STD_LOGIC;
  SIGNAL or_54_rmff : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL and_260_rmff : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_wea_d_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL or_61_rmff : STD_LOGIC;
  SIGNAL or_59_rmff : STD_LOGIC;
  SIGNAL vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL and_273_rmff : STD_LOGIC;
  SIGNAL vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_wea_d_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL or_66_rmff : STD_LOGIC;
  SIGNAL or_64_rmff : STD_LOGIC;
  SIGNAL vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL and_286_rmff : STD_LOGIC;
  SIGNAL vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_wea_d_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL or_71_rmff : STD_LOGIC;
  SIGNAL or_69_rmff : STD_LOGIC;
  SIGNAL vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL and_299_rmff : STD_LOGIC;
  SIGNAL vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_wea_d_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL or_76_rmff : STD_LOGIC;
  SIGNAL or_74_rmff : STD_LOGIC;
  SIGNAL vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL and_312_rmff : STD_LOGIC;
  SIGNAL vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_wea_d_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL or_81_rmff : STD_LOGIC;
  SIGNAL or_79_rmff : STD_LOGIC;
  SIGNAL vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL and_325_rmff : STD_LOGIC;
  SIGNAL vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_wea_d_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL or_86_rmff : STD_LOGIC;
  SIGNAL or_84_rmff : STD_LOGIC;
  SIGNAL vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL and_338_rmff : STD_LOGIC;
  SIGNAL vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_wea_d_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL or_91_rmff : STD_LOGIC;
  SIGNAL or_89_rmff : STD_LOGIC;
  SIGNAL vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL and_351_rmff : STD_LOGIC;
  SIGNAL vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_da_d_reg : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_wea_d_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL or_96_rmff : STD_LOGIC;
  SIGNAL or_94_rmff : STD_LOGIC;
  SIGNAL vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL and_364_rmff : STD_LOGIC;
  SIGNAL vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg : STD_LOGIC_VECTOR (1
      DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL and_373_rmff : STD_LOGIC;
  SIGNAL twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL and_375_rmff : STD_LOGIC;
  SIGNAL twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL and_377_rmff : STD_LOGIC;
  SIGNAL twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL and_379_rmff : STD_LOGIC;
  SIGNAL twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL and_381_rmff : STD_LOGIC;
  SIGNAL twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL and_383_rmff : STD_LOGIC;
  SIGNAL twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL and_385_rmff : STD_LOGIC;
  SIGNAL twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL and_387_rmff : STD_LOGIC;
  SIGNAL twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL and_389_rmff : STD_LOGIC;
  SIGNAL twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL and_391_rmff : STD_LOGIC;
  SIGNAL twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL and_393_rmff : STD_LOGIC;
  SIGNAL twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL and_395_rmff : STD_LOGIC;
  SIGNAL twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL and_397_rmff : STD_LOGIC;
  SIGNAL twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL and_399_rmff : STD_LOGIC;
  SIGNAL twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL and_401_rmff : STD_LOGIC;
  SIGNAL twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL and_403_rmff : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL or_116_rmff : STD_LOGIC;
  SIGNAL or_118_rmff : STD_LOGIC;
  SIGNAL tmp_2_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_3_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_1_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL p_sva : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL STAGE_LOOP_i_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_twiddle_f_equal_tmp : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_equal_tmp_3 : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_equal_tmp_5 : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_equal_tmp_6 : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_equal_tmp_7 : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_equal_tmp_9 : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_equal_tmp_10 : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_equal_tmp_11 : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_equal_tmp_12 : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_equal_tmp_13 : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_equal_tmp_14 : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_equal_tmp_15 : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_nor_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_nor_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_nor_1_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_2_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_nor_3_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_4_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_5_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_6_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_nor_6_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_8_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_9_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_11_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_12_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_13_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_14_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_nor_1_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_nor_10_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_nor_11_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_17_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_nor_13_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_19_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_20_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_21_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_nor_16_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_23_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_24_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_25_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_26_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_27_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_28_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_29_itm : STD_LOGIC;
  SIGNAL STAGE_LOOP_i_3_0_sva_2 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_k_10_0_sva_2 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_twiddle_help_and_16_cse : STD_LOGIC;
  SIGNAL STAGE_LOOP_acc_itm_4_1 : STD_LOGIC;

  SIGNAL COMP_LOOP_k_not_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_twiddle_f_mux1h_1_nl : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_twiddle_f_not_7_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_10_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_1_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_3_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_7_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_15_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_16_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_18_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_VEC_LOOP_and_22_nl : STD_LOGIC;
  SIGNAL STAGE_LOOP_acc_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL p_rsci_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL p_rsci_idat_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT mult
    PORT (
      x_rsc_dat : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      y_rsc_dat : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      y_rsc_dat_1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      p_rsc_dat : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      return_rsc_z : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      ccs_ccore_start_rsc_dat : IN STD_LOGIC;
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_srst : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL mult_cmp_x_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_cmp_y_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_cmp_y_rsc_dat_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_cmp_p_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_cmp_return_rsc_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_cmp_ccs_ccore_start_rsc_dat : STD_LOGIC;

  COMPONENT modulo_sub
    PORT (
      base_rsc_dat : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      m_rsc_dat : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      return_rsc_z : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      ccs_ccore_start_rsc_dat : IN STD_LOGIC;
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_srst : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL modulo_sub_cmp_base_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_cmp_m_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_cmp_return_rsc_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_cmp_ccs_ccore_start_rsc_dat : STD_LOGIC;

  COMPONENT modulo_add
    PORT (
      base_rsc_dat : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      m_rsc_dat : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      return_rsc_z : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      ccs_ccore_start_rsc_dat : IN STD_LOGIC;
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_srst : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL modulo_add_cmp_base_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_cmp_m_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_cmp_return_rsc_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_cmp_ccs_ccore_start_rsc_dat : STD_LOGIC;

  SIGNAL COMP_LOOP_twiddle_f_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL COMP_LOOP_twiddle_f_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_twiddle_f_lshift_rg_z : STD_LOGIC_VECTOR (10 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_run_rsci
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      run_rsc_rdy : OUT STD_LOGIC;
      run_rsc_vld : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      run_rsci_oswt : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      run_rsci_ivld_mxwt : OUT STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_complete_rsci
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      complete_rsc_rdy : IN STD_LOGIC;
      complete_rsc_vld : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      complete_rsci_oswt : IN STD_LOGIC;
      complete_rsci_wen_comp : OUT STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_0_0_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_0_0_i_oswt : IN STD_LOGIC;
      vec_rsc_0_0_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_0_0_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_0_0_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_0_0_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_da_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR
      (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_oswt_1_pff
      : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_wait_dp
    PORT(
      ensig_cgo_iro : IN STD_LOGIC;
      ensig_cgo_iro_1 : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      ensig_cgo : IN STD_LOGIC;
      mult_cmp_ccs_ccore_en : OUT STD_LOGIC;
      ensig_cgo_1 : IN STD_LOGIC;
      modulo_sub_cmp_ccs_ccore_en : OUT STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_0_1_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_1_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_0_1_i_oswt : IN STD_LOGIC;
      vec_rsc_0_1_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_0_1_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_1_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_1_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_0_1_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_0_1_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_da_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR
      (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_oswt_1_pff
      : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_0_2_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_2_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_0_2_i_oswt : IN STD_LOGIC;
      vec_rsc_0_2_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_0_2_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_2_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_2_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_0_2_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_0_2_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_da_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR
      (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_oswt_1_pff
      : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_0_3_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_3_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_0_3_i_oswt : IN STD_LOGIC;
      vec_rsc_0_3_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_0_3_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_3_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_3_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_0_3_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_0_3_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_da_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR
      (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_oswt_1_pff
      : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_0_4_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_4_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_0_4_i_oswt : IN STD_LOGIC;
      vec_rsc_0_4_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_0_4_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_4_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_4_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_0_4_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_0_4_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_da_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR
      (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_oswt_1_pff
      : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_0_5_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_5_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_0_5_i_oswt : IN STD_LOGIC;
      vec_rsc_0_5_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_0_5_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_5_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_5_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_0_5_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_0_5_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_da_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR
      (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_oswt_1_pff
      : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_0_6_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_6_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_0_6_i_oswt : IN STD_LOGIC;
      vec_rsc_0_6_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_0_6_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_6_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_6_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_0_6_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_0_6_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_da_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR
      (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_oswt_1_pff
      : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_0_7_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_7_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_0_7_i_oswt : IN STD_LOGIC;
      vec_rsc_0_7_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_0_7_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_7_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_7_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_0_7_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_0_7_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_da_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR
      (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_oswt_1_pff
      : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_1_0_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_1_0_i_oswt : IN STD_LOGIC;
      vec_rsc_1_0_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_1_0_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_0_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_0_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_1_0_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_1_0_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_da_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_qa_d : STD_LOGIC_VECTOR
      (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_oswt_1_pff
      : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_1_1_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_1_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_1_1_i_oswt : IN STD_LOGIC;
      vec_rsc_1_1_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_1_1_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_1_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_1_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_1_1_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_1_1_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_da_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_qa_d : STD_LOGIC_VECTOR
      (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_oswt_1_pff
      : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_1_2_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_2_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_1_2_i_oswt : IN STD_LOGIC;
      vec_rsc_1_2_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_1_2_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_2_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_2_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_1_2_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_1_2_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_da_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_qa_d : STD_LOGIC_VECTOR
      (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_oswt_1_pff
      : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_1_3_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_3_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_1_3_i_oswt : IN STD_LOGIC;
      vec_rsc_1_3_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_1_3_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_3_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_3_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_1_3_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_1_3_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_da_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_qa_d : STD_LOGIC_VECTOR
      (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_oswt_1_pff
      : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_1_4_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_4_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_1_4_i_oswt : IN STD_LOGIC;
      vec_rsc_1_4_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_1_4_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_4_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_4_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_1_4_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_1_4_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_da_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_qa_d : STD_LOGIC_VECTOR
      (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_oswt_1_pff
      : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_1_5_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_5_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_1_5_i_oswt : IN STD_LOGIC;
      vec_rsc_1_5_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_1_5_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_5_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_5_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_1_5_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_1_5_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_da_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_qa_d : STD_LOGIC_VECTOR
      (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_oswt_1_pff
      : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_1_6_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_6_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_1_6_i_oswt : IN STD_LOGIC;
      vec_rsc_1_6_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_1_6_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_6_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_6_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_1_6_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_1_6_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_da_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_qa_d : STD_LOGIC_VECTOR
      (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_oswt_1_pff
      : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_1_7_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_7_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_1_7_i_oswt : IN STD_LOGIC;
      vec_rsc_1_7_i_oswt_1 : IN STD_LOGIC;
      vec_rsc_1_7_i_da_d_core : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_7_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_7_i_wea_d_core_psct : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct : IN STD_LOGIC_VECTOR
          (1 DOWNTO 0);
      core_wten_pff : IN STD_LOGIC;
      vec_rsc_1_7_i_oswt_pff : IN STD_LOGIC;
      vec_rsc_1_7_i_oswt_1_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_da_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_qa_d : STD_LOGIC_VECTOR
      (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_da_d_core
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_wea_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_oswt_1_pff
      : STD_LOGIC;

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_0_0_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_0_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_0_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_inst_twiddle_rsc_0_0_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_inst_twiddle_rsc_0_0_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_0_1_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_1_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_1_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_inst_twiddle_rsc_0_1_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_inst_twiddle_rsc_0_1_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_0_2_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_2_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_2_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_inst_twiddle_rsc_0_2_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_inst_twiddle_rsc_0_2_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_0_3_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_3_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_3_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_inst_twiddle_rsc_0_3_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_inst_twiddle_rsc_0_3_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_0_4_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_4_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_4_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_inst_twiddle_rsc_0_4_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_inst_twiddle_rsc_0_4_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_0_5_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_5_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_5_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_inst_twiddle_rsc_0_5_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_inst_twiddle_rsc_0_5_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_0_6_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_6_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_6_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_inst_twiddle_rsc_0_6_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_inst_twiddle_rsc_0_6_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_0_7_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_7_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_7_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_inst_twiddle_rsc_0_7_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_inst_twiddle_rsc_0_7_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_1_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_1_0_i_oswt : IN STD_LOGIC;
      twiddle_rsc_1_0_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_0_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_inst_twiddle_rsc_1_0_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_inst_twiddle_rsc_1_0_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_1_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_1_1_i_oswt : IN STD_LOGIC;
      twiddle_rsc_1_1_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_1_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_inst_twiddle_rsc_1_1_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_inst_twiddle_rsc_1_1_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_1_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_1_2_i_oswt : IN STD_LOGIC;
      twiddle_rsc_1_2_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_2_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_inst_twiddle_rsc_1_2_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_inst_twiddle_rsc_1_2_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_1_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_1_3_i_oswt : IN STD_LOGIC;
      twiddle_rsc_1_3_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_3_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_inst_twiddle_rsc_1_3_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_inst_twiddle_rsc_1_3_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_1_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_1_4_i_oswt : IN STD_LOGIC;
      twiddle_rsc_1_4_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_4_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_inst_twiddle_rsc_1_4_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_inst_twiddle_rsc_1_4_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_1_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_1_5_i_oswt : IN STD_LOGIC;
      twiddle_rsc_1_5_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_5_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_inst_twiddle_rsc_1_5_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_inst_twiddle_rsc_1_5_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_1_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_1_6_i_oswt : IN STD_LOGIC;
      twiddle_rsc_1_6_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_6_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_inst_twiddle_rsc_1_6_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_inst_twiddle_rsc_1_6_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_1_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_1_7_i_oswt : IN STD_LOGIC;
      twiddle_rsc_1_7_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_7_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_inst_twiddle_rsc_1_7_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_inst_twiddle_rsc_1_7_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_0_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_inst_twiddle_h_rsc_0_0_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_inst_twiddle_h_rsc_0_0_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_1_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_inst_twiddle_h_rsc_0_1_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_inst_twiddle_h_rsc_0_1_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_2_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_inst_twiddle_h_rsc_0_2_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_inst_twiddle_h_rsc_0_2_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_3_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_inst_twiddle_h_rsc_0_3_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_inst_twiddle_h_rsc_0_3_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_4_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_inst_twiddle_h_rsc_0_4_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_inst_twiddle_h_rsc_0_4_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_5_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_inst_twiddle_h_rsc_0_5_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_inst_twiddle_h_rsc_0_5_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_6_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_inst_twiddle_h_rsc_0_6_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_inst_twiddle_h_rsc_0_6_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_7_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_inst_twiddle_h_rsc_0_7_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_inst_twiddle_h_rsc_0_7_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_1_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_1_0_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_1_0_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_0_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_inst_twiddle_h_rsc_1_0_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_inst_twiddle_h_rsc_1_0_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_1_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_1_1_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_1_1_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_1_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_inst_twiddle_h_rsc_1_1_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_inst_twiddle_h_rsc_1_1_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_1_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_1_2_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_1_2_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_2_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_inst_twiddle_h_rsc_1_2_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_inst_twiddle_h_rsc_1_2_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_1_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_1_3_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_1_3_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_3_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_inst_twiddle_h_rsc_1_3_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_inst_twiddle_h_rsc_1_3_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_1_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_1_4_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_1_4_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_4_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_inst_twiddle_h_rsc_1_4_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_inst_twiddle_h_rsc_1_4_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_1_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_1_5_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_1_5_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_5_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_inst_twiddle_h_rsc_1_5_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_inst_twiddle_h_rsc_1_5_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_1_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_1_6_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_1_6_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_6_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_inst_twiddle_h_rsc_1_6_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_inst_twiddle_h_rsc_1_6_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_1_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_1_7_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_1_7_i_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_7_i_oswt_pff : IN STD_LOGIC;
      core_wten_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_inst_twiddle_h_rsc_1_7_i_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_inst_twiddle_h_rsc_1_7_i_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_7_obj
    PORT(
      vec_rsc_triosy_1_7_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_1_7_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_6_obj
    PORT(
      vec_rsc_triosy_1_6_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_1_6_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_5_obj
    PORT(
      vec_rsc_triosy_1_5_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_1_5_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_4_obj
    PORT(
      vec_rsc_triosy_1_4_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_1_4_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_3_obj
    PORT(
      vec_rsc_triosy_1_3_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_1_3_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_2_obj
    PORT(
      vec_rsc_triosy_1_2_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_1_2_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_1_obj
    PORT(
      vec_rsc_triosy_1_1_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_1_1_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_0_obj
    PORT(
      vec_rsc_triosy_1_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_7_obj
    PORT(
      vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_6_obj
    PORT(
      vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_5_obj
    PORT(
      vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_4_obj
    PORT(
      vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_3_obj
    PORT(
      vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_2_obj
    PORT(
      vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_1_obj
    PORT(
      vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_0_obj
    PORT(
      vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      vec_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_p_rsc_triosy_obj
    PORT(
      p_rsc_triosy_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      p_rsc_triosy_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_r_rsc_triosy_obj
    PORT(
      r_rsc_triosy_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      r_rsc_triosy_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_7_obj
    PORT(
      twiddle_rsc_triosy_1_7_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_1_7_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_6_obj
    PORT(
      twiddle_rsc_triosy_1_6_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_1_6_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_5_obj
    PORT(
      twiddle_rsc_triosy_1_5_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_1_5_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_4_obj
    PORT(
      twiddle_rsc_triosy_1_4_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_1_4_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_3_obj
    PORT(
      twiddle_rsc_triosy_1_3_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_1_3_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_2_obj
    PORT(
      twiddle_rsc_triosy_1_2_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_1_2_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_1_obj
    PORT(
      twiddle_rsc_triosy_1_1_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_1_1_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_0_obj
    PORT(
      twiddle_rsc_triosy_1_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_7_obj
    PORT(
      twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_6_obj
    PORT(
      twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_5_obj
    PORT(
      twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_4_obj
    PORT(
      twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_3_obj
    PORT(
      twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_2_obj
    PORT(
      twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_1_obj
    PORT(
      twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_0_obj
    PORT(
      twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_7_obj
    PORT(
      twiddle_h_rsc_triosy_1_7_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_7_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_6_obj
    PORT(
      twiddle_h_rsc_triosy_1_6_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_6_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_5_obj
    PORT(
      twiddle_h_rsc_triosy_1_5_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_5_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_4_obj
    PORT(
      twiddle_h_rsc_triosy_1_4_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_4_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_3_obj
    PORT(
      twiddle_h_rsc_triosy_1_3_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_3_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_2_obj
    PORT(
      twiddle_h_rsc_triosy_1_2_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_2_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_1_obj
    PORT(
      twiddle_h_rsc_triosy_1_1_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_1_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_0_obj
    PORT(
      twiddle_h_rsc_triosy_1_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_7_obj
    PORT(
      twiddle_h_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_6_obj
    PORT(
      twiddle_h_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_5_obj
    PORT(
      twiddle_h_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_4_obj
    PORT(
      twiddle_h_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_3_obj
    PORT(
      twiddle_h_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_2_obj
    PORT(
      twiddle_h_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_1_obj
    PORT(
      twiddle_h_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_0_obj
    PORT(
      twiddle_h_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_staller
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      core_wten : OUT STD_LOGIC;
      complete_rsci_wen_comp : IN STD_LOGIC;
      core_wten_pff : OUT STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_precomp_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      complete_rsci_wen_comp : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
      main_C_0_tr0 : IN STD_LOGIC;
      VEC_LOOP_C_11_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_4_tr0 : IN STD_LOGIC;
      STAGE_LOOP_C_1_tr0 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR
      (21 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_core_fsm_inst_main_C_0_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_precomp_core_core_fsm_inst_VEC_LOOP_C_11_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_precomp_core_core_fsm_inst_COMP_LOOP_C_4_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_precomp_core_core_fsm_inst_STAGE_LOOP_C_1_tr0 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_v_10_3_2(input_2 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(9 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(9 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_16_2(input_15 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(15 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_3_2(input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_10_2_2(input_0 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(9 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_4_2_2(input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION minimum(arg1,arg2:INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1<arg2)THEN
      RETURN arg1;
    ELSE
      RETURN arg2;
    END IF;
  END;

  FUNCTION maximum(arg1,arg2:INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1>arg2)THEN
      RETURN arg1;
    ELSE
      RETURN arg2;
    END IF;
  END;

  FUNCTION READSLICE_1_11(input_val:STD_LOGIC_VECTOR(10 DOWNTO 0);index:INTEGER)
  RETURN STD_LOGIC IS
    CONSTANT min_sat_index:INTEGER:= maximum( index, 0 );
    CONSTANT sat_index:INTEGER:= minimum( min_sat_index, 10);
  BEGIN
    RETURN input_val(sat_index);
  END;

BEGIN
  p_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 14,
      width => 32
      )
    PORT MAP(
      dat => p_rsci_dat,
      idat => p_rsci_idat_1
    );
  p_rsci_dat <= p_rsc_dat;
  p_rsci_idat <= p_rsci_idat_1;

  mult_cmp : mult
    PORT MAP(
      x_rsc_dat => mult_cmp_x_rsc_dat,
      y_rsc_dat => mult_cmp_y_rsc_dat,
      y_rsc_dat_1 => mult_cmp_y_rsc_dat_1,
      p_rsc_dat => mult_cmp_p_rsc_dat,
      return_rsc_z => mult_cmp_return_rsc_z_1,
      ccs_ccore_start_rsc_dat => mult_cmp_ccs_ccore_start_rsc_dat,
      ccs_ccore_clk => clk,
      ccs_ccore_srst => rst,
      ccs_ccore_en => mult_cmp_ccs_ccore_en
    );
  mult_cmp_x_rsc_dat <= modulo_sub_cmp_return_rsc_z;
  mult_cmp_y_rsc_dat <= tmp_2_lpi_3_dfm;
  mult_cmp_y_rsc_dat_1 <= tmp_3_lpi_3_dfm;
  mult_cmp_p_rsc_dat <= p_sva;
  mult_cmp_return_rsc_z <= mult_cmp_return_rsc_z_1;
  mult_cmp_ccs_ccore_start_rsc_dat <= fsm_output(9);

  modulo_sub_cmp : modulo_sub
    PORT MAP(
      base_rsc_dat => modulo_sub_cmp_base_rsc_dat,
      m_rsc_dat => modulo_sub_cmp_m_rsc_dat,
      return_rsc_z => modulo_sub_cmp_return_rsc_z_1,
      ccs_ccore_start_rsc_dat => modulo_sub_cmp_ccs_ccore_start_rsc_dat,
      ccs_ccore_clk => clk,
      ccs_ccore_srst => rst,
      ccs_ccore_en => modulo_sub_cmp_ccs_ccore_en
    );
  modulo_sub_cmp_base_rsc_dat <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_lpi_4_dfm)
      - UNSIGNED(tmp_1_lpi_4_dfm), 32));
  modulo_sub_cmp_m_rsc_dat <= p_sva;
  modulo_sub_cmp_return_rsc_z <= modulo_sub_cmp_return_rsc_z_1;
  modulo_sub_cmp_ccs_ccore_start_rsc_dat <= fsm_output(8);

  modulo_add_cmp : modulo_add
    PORT MAP(
      base_rsc_dat => modulo_add_cmp_base_rsc_dat,
      m_rsc_dat => modulo_add_cmp_m_rsc_dat,
      return_rsc_z => modulo_add_cmp_return_rsc_z_1,
      ccs_ccore_start_rsc_dat => modulo_add_cmp_ccs_ccore_start_rsc_dat,
      ccs_ccore_clk => clk,
      ccs_ccore_srst => rst,
      ccs_ccore_en => modulo_sub_cmp_ccs_ccore_en
    );
  modulo_add_cmp_base_rsc_dat <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_lpi_4_dfm)
      + UNSIGNED(tmp_1_lpi_4_dfm), 32));
  modulo_add_cmp_m_rsc_dat <= p_sva;
  modulo_add_cmp_return_rsc_z <= modulo_add_cmp_return_rsc_z_1;
  modulo_add_cmp_ccs_ccore_start_rsc_dat <= fsm_output(8);

  COMP_LOOP_twiddle_f_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_l_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 0,
      width_s => 4,
      width_z => 11
      )
    PORT MAP(
      a => COMP_LOOP_twiddle_f_lshift_rg_a,
      s => COMP_LOOP_twiddle_f_lshift_rg_s,
      z => COMP_LOOP_twiddle_f_lshift_rg_z
    );
  COMP_LOOP_twiddle_f_lshift_rg_a(0) <= '1';
  COMP_LOOP_twiddle_f_lshift_rg_s <= MUX_v_4_2_2(STAGE_LOOP_i_3_0_sva, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(NOT
      STAGE_LOOP_i_3_0_sva) + UNSIGNED'( "1011"), 4)), fsm_output(2));
  z_out <= COMP_LOOP_twiddle_f_lshift_rg_z;

  inPlaceNTT_DIF_precomp_core_run_rsci_inst : inPlaceNTT_DIF_precomp_core_run_rsci
    PORT MAP(
      clk => clk,
      rst => rst,
      run_rsc_rdy => run_rsc_rdy,
      run_rsc_vld => run_rsc_vld,
      core_wen => complete_rsci_wen_comp,
      run_rsci_oswt => reg_run_rsci_oswt_cse,
      core_wten => core_wten,
      run_rsci_ivld_mxwt => run_rsci_ivld_mxwt
    );
  inPlaceNTT_DIF_precomp_core_complete_rsci_inst : inPlaceNTT_DIF_precomp_core_complete_rsci
    PORT MAP(
      clk => clk,
      rst => rst,
      complete_rsc_rdy => complete_rsc_rdy,
      complete_rsc_vld => complete_rsc_vld,
      core_wen => complete_rsci_wen_comp,
      complete_rsci_oswt => reg_complete_rsci_oswt_cse,
      complete_rsci_wen_comp => complete_rsci_wen_comp
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_0_0_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_da_d,
      vec_rsc_0_0_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_qa_d,
      vec_rsc_0_0_i_wea_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_wea_d,
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      vec_rsc_0_0_i_oswt => reg_vec_rsc_0_0_i_oswt_cse,
      vec_rsc_0_0_i_oswt_1 => reg_vec_rsc_0_0_i_oswt_1_cse,
      vec_rsc_0_0_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_da_d_core,
      vec_rsc_0_0_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_qa_d_mxwt,
      vec_rsc_0_0_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_wea_d_core_psct,
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      core_wten_pff => core_wten_iff,
      vec_rsc_0_0_i_oswt_pff => or_15_rmff,
      vec_rsc_0_0_i_oswt_1_pff => inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_oswt_1_pff
    );
  vec_rsc_0_0_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_qa_d <= vec_rsc_0_0_i_qa_d;
  vec_rsc_0_0_i_wea_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_wea_d;
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_da_d_core <= STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000") & VEC_LOOP_mux_4_rmff;
  vec_rsc_0_0_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_qa_d_mxwt;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_21_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( and_161_rmff & and_158_cse);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_21_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_0_i_1_inst_vec_rsc_0_0_i_oswt_1_pff <= and_161_rmff;

  inPlaceNTT_DIF_precomp_core_wait_dp_inst : inPlaceNTT_DIF_precomp_core_wait_dp
    PORT MAP(
      ensig_cgo_iro => or_116_rmff,
      ensig_cgo_iro_1 => or_118_rmff,
      core_wen => complete_rsci_wen_comp,
      ensig_cgo => reg_ensig_cgo_cse,
      mult_cmp_ccs_ccore_en => mult_cmp_ccs_ccore_en,
      ensig_cgo_1 => reg_ensig_cgo_1_cse,
      modulo_sub_cmp_ccs_ccore_en => modulo_sub_cmp_ccs_ccore_en
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_0_1_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_da_d,
      vec_rsc_0_1_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_qa_d,
      vec_rsc_0_1_i_wea_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_wea_d,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      vec_rsc_0_1_i_oswt => reg_vec_rsc_0_1_i_oswt_cse,
      vec_rsc_0_1_i_oswt_1 => reg_vec_rsc_0_1_i_oswt_1_cse,
      vec_rsc_0_1_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_da_d_core,
      vec_rsc_0_1_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_qa_d_mxwt,
      vec_rsc_0_1_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_wea_d_core_psct,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      core_wten_pff => core_wten_iff,
      vec_rsc_0_1_i_oswt_pff => or_24_rmff,
      vec_rsc_0_1_i_oswt_1_pff => inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_oswt_1_pff
    );
  vec_rsc_0_1_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_qa_d <= vec_rsc_0_1_i_qa_d;
  vec_rsc_0_1_i_wea_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_wea_d;
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_da_d_core <= STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000") & VEC_LOOP_mux_4_rmff;
  vec_rsc_0_1_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_qa_d_mxwt;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_26_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( and_182_rmff & and_179_cse);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_26_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_1_i_1_inst_vec_rsc_0_1_i_oswt_1_pff <= and_182_rmff;

  inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_0_2_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_da_d,
      vec_rsc_0_2_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_qa_d,
      vec_rsc_0_2_i_wea_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_wea_d,
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      vec_rsc_0_2_i_oswt => reg_vec_rsc_0_2_i_oswt_cse,
      vec_rsc_0_2_i_oswt_1 => reg_vec_rsc_0_2_i_oswt_1_cse,
      vec_rsc_0_2_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_da_d_core,
      vec_rsc_0_2_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_qa_d_mxwt,
      vec_rsc_0_2_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_wea_d_core_psct,
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      core_wten_pff => core_wten_iff,
      vec_rsc_0_2_i_oswt_pff => or_29_rmff,
      vec_rsc_0_2_i_oswt_1_pff => inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_oswt_1_pff
    );
  vec_rsc_0_2_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_qa_d <= vec_rsc_0_2_i_qa_d;
  vec_rsc_0_2_i_wea_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_wea_d;
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_da_d_core <= STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000") & VEC_LOOP_mux_4_rmff;
  vec_rsc_0_2_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_qa_d_mxwt;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_31_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( and_195_rmff & and_192_cse);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_31_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_2_i_1_inst_vec_rsc_0_2_i_oswt_1_pff <= and_195_rmff;

  inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_0_3_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_da_d,
      vec_rsc_0_3_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_qa_d,
      vec_rsc_0_3_i_wea_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_wea_d,
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      vec_rsc_0_3_i_oswt => reg_vec_rsc_0_3_i_oswt_cse,
      vec_rsc_0_3_i_oswt_1 => reg_vec_rsc_0_3_i_oswt_1_cse,
      vec_rsc_0_3_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_da_d_core,
      vec_rsc_0_3_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_qa_d_mxwt,
      vec_rsc_0_3_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_wea_d_core_psct,
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      core_wten_pff => core_wten_iff,
      vec_rsc_0_3_i_oswt_pff => or_34_rmff,
      vec_rsc_0_3_i_oswt_1_pff => inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_oswt_1_pff
    );
  vec_rsc_0_3_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_qa_d <= vec_rsc_0_3_i_qa_d;
  vec_rsc_0_3_i_wea_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_wea_d;
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_da_d_core <= STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000") & VEC_LOOP_mux_4_rmff;
  vec_rsc_0_3_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_qa_d_mxwt;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_36_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( and_208_rmff & and_205_cse);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_36_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_3_i_1_inst_vec_rsc_0_3_i_oswt_1_pff <= and_208_rmff;

  inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_0_4_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_da_d,
      vec_rsc_0_4_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_qa_d,
      vec_rsc_0_4_i_wea_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_wea_d,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      vec_rsc_0_4_i_oswt => reg_vec_rsc_0_4_i_oswt_cse,
      vec_rsc_0_4_i_oswt_1 => reg_vec_rsc_0_4_i_oswt_1_cse,
      vec_rsc_0_4_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_da_d_core,
      vec_rsc_0_4_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_qa_d_mxwt,
      vec_rsc_0_4_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_wea_d_core_psct,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      core_wten_pff => core_wten_iff,
      vec_rsc_0_4_i_oswt_pff => or_39_rmff,
      vec_rsc_0_4_i_oswt_1_pff => inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_oswt_1_pff
    );
  vec_rsc_0_4_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_qa_d <= vec_rsc_0_4_i_qa_d;
  vec_rsc_0_4_i_wea_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_wea_d;
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_da_d_core <= STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000") & VEC_LOOP_mux_4_rmff;
  vec_rsc_0_4_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_qa_d_mxwt;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_41_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( and_221_rmff & and_218_cse);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_41_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_4_i_1_inst_vec_rsc_0_4_i_oswt_1_pff <= and_221_rmff;

  inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_0_5_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_da_d,
      vec_rsc_0_5_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_qa_d,
      vec_rsc_0_5_i_wea_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_wea_d,
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      vec_rsc_0_5_i_oswt => reg_vec_rsc_0_5_i_oswt_cse,
      vec_rsc_0_5_i_oswt_1 => reg_vec_rsc_0_5_i_oswt_1_cse,
      vec_rsc_0_5_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_da_d_core,
      vec_rsc_0_5_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_qa_d_mxwt,
      vec_rsc_0_5_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_wea_d_core_psct,
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      core_wten_pff => core_wten_iff,
      vec_rsc_0_5_i_oswt_pff => or_44_rmff,
      vec_rsc_0_5_i_oswt_1_pff => inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_oswt_1_pff
    );
  vec_rsc_0_5_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_qa_d <= vec_rsc_0_5_i_qa_d;
  vec_rsc_0_5_i_wea_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_wea_d;
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_da_d_core <= STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000") & VEC_LOOP_mux_4_rmff;
  vec_rsc_0_5_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_qa_d_mxwt;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_46_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( and_234_rmff & and_231_cse);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_46_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_5_i_1_inst_vec_rsc_0_5_i_oswt_1_pff <= and_234_rmff;

  inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_0_6_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_da_d,
      vec_rsc_0_6_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_qa_d,
      vec_rsc_0_6_i_wea_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_wea_d,
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      vec_rsc_0_6_i_oswt => reg_vec_rsc_0_6_i_oswt_cse,
      vec_rsc_0_6_i_oswt_1 => reg_vec_rsc_0_6_i_oswt_1_cse,
      vec_rsc_0_6_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_da_d_core,
      vec_rsc_0_6_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_qa_d_mxwt,
      vec_rsc_0_6_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_wea_d_core_psct,
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      core_wten_pff => core_wten_iff,
      vec_rsc_0_6_i_oswt_pff => or_49_rmff,
      vec_rsc_0_6_i_oswt_1_pff => inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_oswt_1_pff
    );
  vec_rsc_0_6_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_qa_d <= vec_rsc_0_6_i_qa_d;
  vec_rsc_0_6_i_wea_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_wea_d;
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_da_d_core <= STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000") & VEC_LOOP_mux_4_rmff;
  vec_rsc_0_6_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_qa_d_mxwt;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_51_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( and_247_rmff & and_244_cse);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_51_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_6_i_1_inst_vec_rsc_0_6_i_oswt_1_pff <= and_247_rmff;

  inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_0_7_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_da_d,
      vec_rsc_0_7_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_qa_d,
      vec_rsc_0_7_i_wea_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_wea_d,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      vec_rsc_0_7_i_oswt => reg_vec_rsc_0_7_i_oswt_cse,
      vec_rsc_0_7_i_oswt_1 => reg_vec_rsc_0_7_i_oswt_1_cse,
      vec_rsc_0_7_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_da_d_core,
      vec_rsc_0_7_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_qa_d_mxwt,
      vec_rsc_0_7_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_wea_d_core_psct,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      core_wten_pff => core_wten_iff,
      vec_rsc_0_7_i_oswt_pff => or_54_rmff,
      vec_rsc_0_7_i_oswt_1_pff => inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_oswt_1_pff
    );
  vec_rsc_0_7_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_qa_d <= vec_rsc_0_7_i_qa_d;
  vec_rsc_0_7_i_wea_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_wea_d;
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_da_d_core <= STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000") & VEC_LOOP_mux_4_rmff;
  vec_rsc_0_7_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_qa_d_mxwt;
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_56_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( and_260_rmff & and_257_cse);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_56_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_0_7_i_1_inst_vec_rsc_0_7_i_oswt_1_pff <= and_260_rmff;

  inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_1_0_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_da_d,
      vec_rsc_1_0_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_qa_d,
      vec_rsc_1_0_i_wea_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_wea_d,
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      vec_rsc_1_0_i_oswt => reg_vec_rsc_1_0_i_oswt_cse,
      vec_rsc_1_0_i_oswt_1 => reg_vec_rsc_1_0_i_oswt_1_cse,
      vec_rsc_1_0_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_da_d_core,
      vec_rsc_1_0_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_qa_d_mxwt,
      vec_rsc_1_0_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_wea_d_core_psct,
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      core_wten_pff => core_wten_iff,
      vec_rsc_1_0_i_oswt_pff => or_59_rmff,
      vec_rsc_1_0_i_oswt_1_pff => inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_oswt_1_pff
    );
  vec_rsc_1_0_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_qa_d <= vec_rsc_1_0_i_qa_d;
  vec_rsc_1_0_i_wea_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_wea_d;
  vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_da_d_core <= STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000") & VEC_LOOP_mux_4_rmff;
  vec_rsc_1_0_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_qa_d_mxwt;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_61_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( and_273_rmff & and_270_cse);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_61_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_0_i_1_inst_vec_rsc_1_0_i_oswt_1_pff <= and_273_rmff;

  inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_1_1_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_da_d,
      vec_rsc_1_1_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_qa_d,
      vec_rsc_1_1_i_wea_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_wea_d,
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      vec_rsc_1_1_i_oswt => reg_vec_rsc_1_1_i_oswt_cse,
      vec_rsc_1_1_i_oswt_1 => reg_vec_rsc_1_1_i_oswt_1_cse,
      vec_rsc_1_1_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_da_d_core,
      vec_rsc_1_1_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_qa_d_mxwt,
      vec_rsc_1_1_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_wea_d_core_psct,
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      core_wten_pff => core_wten_iff,
      vec_rsc_1_1_i_oswt_pff => or_64_rmff,
      vec_rsc_1_1_i_oswt_1_pff => inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_oswt_1_pff
    );
  vec_rsc_1_1_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_qa_d <= vec_rsc_1_1_i_qa_d;
  vec_rsc_1_1_i_wea_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_wea_d;
  vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_da_d_core <= STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000") & VEC_LOOP_mux_4_rmff;
  vec_rsc_1_1_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_qa_d_mxwt;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_66_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( and_286_rmff & and_283_cse);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_66_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_1_i_1_inst_vec_rsc_1_1_i_oswt_1_pff <= and_286_rmff;

  inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_1_2_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_da_d,
      vec_rsc_1_2_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_qa_d,
      vec_rsc_1_2_i_wea_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_wea_d,
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      vec_rsc_1_2_i_oswt => reg_vec_rsc_1_2_i_oswt_cse,
      vec_rsc_1_2_i_oswt_1 => reg_vec_rsc_1_2_i_oswt_1_cse,
      vec_rsc_1_2_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_da_d_core,
      vec_rsc_1_2_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_qa_d_mxwt,
      vec_rsc_1_2_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_wea_d_core_psct,
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      core_wten_pff => core_wten_iff,
      vec_rsc_1_2_i_oswt_pff => or_69_rmff,
      vec_rsc_1_2_i_oswt_1_pff => inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_oswt_1_pff
    );
  vec_rsc_1_2_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_qa_d <= vec_rsc_1_2_i_qa_d;
  vec_rsc_1_2_i_wea_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_wea_d;
  vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_da_d_core <= STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000") & VEC_LOOP_mux_4_rmff;
  vec_rsc_1_2_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_qa_d_mxwt;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_71_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( and_299_rmff & and_296_cse);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_71_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_2_i_1_inst_vec_rsc_1_2_i_oswt_1_pff <= and_299_rmff;

  inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_1_3_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_da_d,
      vec_rsc_1_3_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_qa_d,
      vec_rsc_1_3_i_wea_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_wea_d,
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      vec_rsc_1_3_i_oswt => reg_vec_rsc_1_3_i_oswt_cse,
      vec_rsc_1_3_i_oswt_1 => reg_vec_rsc_1_3_i_oswt_1_cse,
      vec_rsc_1_3_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_da_d_core,
      vec_rsc_1_3_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_qa_d_mxwt,
      vec_rsc_1_3_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_wea_d_core_psct,
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      core_wten_pff => core_wten_iff,
      vec_rsc_1_3_i_oswt_pff => or_74_rmff,
      vec_rsc_1_3_i_oswt_1_pff => inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_oswt_1_pff
    );
  vec_rsc_1_3_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_qa_d <= vec_rsc_1_3_i_qa_d;
  vec_rsc_1_3_i_wea_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_wea_d;
  vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_da_d_core <= STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000") & VEC_LOOP_mux_4_rmff;
  vec_rsc_1_3_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_qa_d_mxwt;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_76_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( and_312_rmff & and_309_cse);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_76_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_3_i_1_inst_vec_rsc_1_3_i_oswt_1_pff <= and_312_rmff;

  inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_1_4_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_da_d,
      vec_rsc_1_4_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_qa_d,
      vec_rsc_1_4_i_wea_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_wea_d,
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      vec_rsc_1_4_i_oswt => reg_vec_rsc_1_4_i_oswt_cse,
      vec_rsc_1_4_i_oswt_1 => reg_vec_rsc_1_4_i_oswt_1_cse,
      vec_rsc_1_4_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_da_d_core,
      vec_rsc_1_4_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_qa_d_mxwt,
      vec_rsc_1_4_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_wea_d_core_psct,
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      core_wten_pff => core_wten_iff,
      vec_rsc_1_4_i_oswt_pff => or_79_rmff,
      vec_rsc_1_4_i_oswt_1_pff => inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_oswt_1_pff
    );
  vec_rsc_1_4_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_qa_d <= vec_rsc_1_4_i_qa_d;
  vec_rsc_1_4_i_wea_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_wea_d;
  vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_da_d_core <= STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000") & VEC_LOOP_mux_4_rmff;
  vec_rsc_1_4_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_qa_d_mxwt;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_81_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( and_325_rmff & and_322_cse);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_81_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_4_i_1_inst_vec_rsc_1_4_i_oswt_1_pff <= and_325_rmff;

  inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_1_5_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_da_d,
      vec_rsc_1_5_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_qa_d,
      vec_rsc_1_5_i_wea_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_wea_d,
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      vec_rsc_1_5_i_oswt => reg_vec_rsc_1_5_i_oswt_cse,
      vec_rsc_1_5_i_oswt_1 => reg_vec_rsc_1_5_i_oswt_1_cse,
      vec_rsc_1_5_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_da_d_core,
      vec_rsc_1_5_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_qa_d_mxwt,
      vec_rsc_1_5_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_wea_d_core_psct,
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      core_wten_pff => core_wten_iff,
      vec_rsc_1_5_i_oswt_pff => or_84_rmff,
      vec_rsc_1_5_i_oswt_1_pff => inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_oswt_1_pff
    );
  vec_rsc_1_5_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_qa_d <= vec_rsc_1_5_i_qa_d;
  vec_rsc_1_5_i_wea_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_wea_d;
  vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_da_d_core <= STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000") & VEC_LOOP_mux_4_rmff;
  vec_rsc_1_5_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_qa_d_mxwt;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_86_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( and_338_rmff & and_335_cse);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_86_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_5_i_1_inst_vec_rsc_1_5_i_oswt_1_pff <= and_338_rmff;

  inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_1_6_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_da_d,
      vec_rsc_1_6_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_qa_d,
      vec_rsc_1_6_i_wea_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_wea_d,
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      vec_rsc_1_6_i_oswt => reg_vec_rsc_1_6_i_oswt_cse,
      vec_rsc_1_6_i_oswt_1 => reg_vec_rsc_1_6_i_oswt_1_cse,
      vec_rsc_1_6_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_da_d_core,
      vec_rsc_1_6_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_qa_d_mxwt,
      vec_rsc_1_6_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_wea_d_core_psct,
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      core_wten_pff => core_wten_iff,
      vec_rsc_1_6_i_oswt_pff => or_89_rmff,
      vec_rsc_1_6_i_oswt_1_pff => inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_oswt_1_pff
    );
  vec_rsc_1_6_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_qa_d <= vec_rsc_1_6_i_qa_d;
  vec_rsc_1_6_i_wea_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_wea_d;
  vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_da_d_core <= STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000") & VEC_LOOP_mux_4_rmff;
  vec_rsc_1_6_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_qa_d_mxwt;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_91_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( and_351_rmff & and_348_cse);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_91_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_6_i_1_inst_vec_rsc_1_6_i_oswt_1_pff <= and_351_rmff;

  inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_1_7_i_da_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_da_d,
      vec_rsc_1_7_i_qa_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_qa_d,
      vec_rsc_1_7_i_wea_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_wea_d,
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      vec_rsc_1_7_i_oswt => reg_vec_rsc_1_7_i_oswt_cse,
      vec_rsc_1_7_i_oswt_1 => reg_vec_rsc_1_7_i_oswt_1_cse,
      vec_rsc_1_7_i_da_d_core => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_da_d_core,
      vec_rsc_1_7_i_qa_d_mxwt => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_qa_d_mxwt,
      vec_rsc_1_7_i_wea_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_wea_d_core_psct,
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct,
      core_wten_pff => core_wten_iff,
      vec_rsc_1_7_i_oswt_pff => or_94_rmff,
      vec_rsc_1_7_i_oswt_1_pff => inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_oswt_1_pff
    );
  vec_rsc_1_7_i_da_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_da_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_qa_d <= vec_rsc_1_7_i_qa_d;
  vec_rsc_1_7_i_wea_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_wea_d;
  vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_da_d_core <= STD_LOGIC_VECTOR'(
      "00000000000000000000000000000000") & VEC_LOOP_mux_4_rmff;
  vec_rsc_1_7_i_qa_d_mxwt <= inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_qa_d_mxwt;
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_wea_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_96_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( and_364_rmff & and_361_cse);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_core_psct
      <= STD_LOGIC_VECTOR'( '0' & or_96_rmff);
  inPlaceNTT_DIF_precomp_core_vec_rsc_1_7_i_1_inst_vec_rsc_1_7_i_oswt_1_pff <= and_364_rmff;

  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_0_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_inst_twiddle_rsc_0_0_i_qb_d,
      twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_rsc_0_0_i_oswt => reg_twiddle_rsc_0_0_i_oswt_cse,
      twiddle_rsc_0_0_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_inst_twiddle_rsc_0_0_i_qb_d_mxwt,
      twiddle_rsc_0_0_i_oswt_pff => and_373_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_inst_twiddle_rsc_0_0_i_qb_d <=
      twiddle_rsc_0_0_i_qb_d;
  twiddle_rsc_0_0_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_0_i_1_inst_twiddle_rsc_0_0_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_1_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_inst_twiddle_rsc_0_1_i_qb_d,
      twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_rsc_0_1_i_oswt => reg_twiddle_rsc_0_1_i_oswt_cse,
      twiddle_rsc_0_1_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_inst_twiddle_rsc_0_1_i_qb_d_mxwt,
      twiddle_rsc_0_1_i_oswt_pff => and_375_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_inst_twiddle_rsc_0_1_i_qb_d <=
      twiddle_rsc_0_1_i_qb_d;
  twiddle_rsc_0_1_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_1_i_1_inst_twiddle_rsc_0_1_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_2_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_inst_twiddle_rsc_0_2_i_qb_d,
      twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_rsc_0_2_i_oswt => reg_twiddle_rsc_0_2_i_oswt_cse,
      twiddle_rsc_0_2_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_inst_twiddle_rsc_0_2_i_qb_d_mxwt,
      twiddle_rsc_0_2_i_oswt_pff => and_377_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_inst_twiddle_rsc_0_2_i_qb_d <=
      twiddle_rsc_0_2_i_qb_d;
  twiddle_rsc_0_2_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_2_i_1_inst_twiddle_rsc_0_2_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_3_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_inst_twiddle_rsc_0_3_i_qb_d,
      twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_rsc_0_3_i_oswt => reg_twiddle_rsc_0_3_i_oswt_cse,
      twiddle_rsc_0_3_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_inst_twiddle_rsc_0_3_i_qb_d_mxwt,
      twiddle_rsc_0_3_i_oswt_pff => and_379_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_inst_twiddle_rsc_0_3_i_qb_d <=
      twiddle_rsc_0_3_i_qb_d;
  twiddle_rsc_0_3_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_3_i_1_inst_twiddle_rsc_0_3_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_4_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_inst_twiddle_rsc_0_4_i_qb_d,
      twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_rsc_0_4_i_oswt => reg_twiddle_rsc_0_4_i_oswt_cse,
      twiddle_rsc_0_4_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_inst_twiddle_rsc_0_4_i_qb_d_mxwt,
      twiddle_rsc_0_4_i_oswt_pff => and_381_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_inst_twiddle_rsc_0_4_i_qb_d <=
      twiddle_rsc_0_4_i_qb_d;
  twiddle_rsc_0_4_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_4_i_1_inst_twiddle_rsc_0_4_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_5_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_inst_twiddle_rsc_0_5_i_qb_d,
      twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_rsc_0_5_i_oswt => reg_twiddle_rsc_0_5_i_oswt_cse,
      twiddle_rsc_0_5_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_inst_twiddle_rsc_0_5_i_qb_d_mxwt,
      twiddle_rsc_0_5_i_oswt_pff => and_383_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_inst_twiddle_rsc_0_5_i_qb_d <=
      twiddle_rsc_0_5_i_qb_d;
  twiddle_rsc_0_5_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_5_i_1_inst_twiddle_rsc_0_5_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_6_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_inst_twiddle_rsc_0_6_i_qb_d,
      twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_rsc_0_6_i_oswt => reg_twiddle_rsc_0_6_i_oswt_cse,
      twiddle_rsc_0_6_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_inst_twiddle_rsc_0_6_i_qb_d_mxwt,
      twiddle_rsc_0_6_i_oswt_pff => and_385_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_inst_twiddle_rsc_0_6_i_qb_d <=
      twiddle_rsc_0_6_i_qb_d;
  twiddle_rsc_0_6_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_6_i_1_inst_twiddle_rsc_0_6_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_7_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_inst_twiddle_rsc_0_7_i_qb_d,
      twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_rsc_0_7_i_oswt => reg_twiddle_rsc_0_7_i_oswt_cse,
      twiddle_rsc_0_7_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_inst_twiddle_rsc_0_7_i_qb_d_mxwt,
      twiddle_rsc_0_7_i_oswt_pff => and_387_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_inst_twiddle_rsc_0_7_i_qb_d <=
      twiddle_rsc_0_7_i_qb_d;
  twiddle_rsc_0_7_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_0_7_i_1_inst_twiddle_rsc_0_7_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_1_0_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_inst_twiddle_rsc_1_0_i_qb_d,
      twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_rsc_1_0_i_oswt => reg_twiddle_rsc_1_0_i_oswt_cse,
      twiddle_rsc_1_0_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_inst_twiddle_rsc_1_0_i_qb_d_mxwt,
      twiddle_rsc_1_0_i_oswt_pff => and_389_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_inst_twiddle_rsc_1_0_i_qb_d <=
      twiddle_rsc_1_0_i_qb_d;
  twiddle_rsc_1_0_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_0_i_1_inst_twiddle_rsc_1_0_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_1_1_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_inst_twiddle_rsc_1_1_i_qb_d,
      twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_rsc_1_1_i_oswt => reg_twiddle_rsc_1_1_i_oswt_cse,
      twiddle_rsc_1_1_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_inst_twiddle_rsc_1_1_i_qb_d_mxwt,
      twiddle_rsc_1_1_i_oswt_pff => and_391_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_inst_twiddle_rsc_1_1_i_qb_d <=
      twiddle_rsc_1_1_i_qb_d;
  twiddle_rsc_1_1_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_1_i_1_inst_twiddle_rsc_1_1_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_1_2_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_inst_twiddle_rsc_1_2_i_qb_d,
      twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_rsc_1_2_i_oswt => reg_twiddle_rsc_1_2_i_oswt_cse,
      twiddle_rsc_1_2_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_inst_twiddle_rsc_1_2_i_qb_d_mxwt,
      twiddle_rsc_1_2_i_oswt_pff => and_393_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_inst_twiddle_rsc_1_2_i_qb_d <=
      twiddle_rsc_1_2_i_qb_d;
  twiddle_rsc_1_2_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_2_i_1_inst_twiddle_rsc_1_2_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_1_3_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_inst_twiddle_rsc_1_3_i_qb_d,
      twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_rsc_1_3_i_oswt => reg_twiddle_rsc_1_3_i_oswt_cse,
      twiddle_rsc_1_3_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_inst_twiddle_rsc_1_3_i_qb_d_mxwt,
      twiddle_rsc_1_3_i_oswt_pff => and_395_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_inst_twiddle_rsc_1_3_i_qb_d <=
      twiddle_rsc_1_3_i_qb_d;
  twiddle_rsc_1_3_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_3_i_1_inst_twiddle_rsc_1_3_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_1_4_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_inst_twiddle_rsc_1_4_i_qb_d,
      twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_rsc_1_4_i_oswt => reg_twiddle_rsc_1_4_i_oswt_cse,
      twiddle_rsc_1_4_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_inst_twiddle_rsc_1_4_i_qb_d_mxwt,
      twiddle_rsc_1_4_i_oswt_pff => and_397_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_inst_twiddle_rsc_1_4_i_qb_d <=
      twiddle_rsc_1_4_i_qb_d;
  twiddle_rsc_1_4_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_4_i_1_inst_twiddle_rsc_1_4_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_1_5_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_inst_twiddle_rsc_1_5_i_qb_d,
      twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_rsc_1_5_i_oswt => reg_twiddle_rsc_1_5_i_oswt_cse,
      twiddle_rsc_1_5_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_inst_twiddle_rsc_1_5_i_qb_d_mxwt,
      twiddle_rsc_1_5_i_oswt_pff => and_399_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_inst_twiddle_rsc_1_5_i_qb_d <=
      twiddle_rsc_1_5_i_qb_d;
  twiddle_rsc_1_5_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_5_i_1_inst_twiddle_rsc_1_5_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_1_6_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_inst_twiddle_rsc_1_6_i_qb_d,
      twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_rsc_1_6_i_oswt => reg_twiddle_rsc_1_6_i_oswt_cse,
      twiddle_rsc_1_6_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_inst_twiddle_rsc_1_6_i_qb_d_mxwt,
      twiddle_rsc_1_6_i_oswt_pff => and_401_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_inst_twiddle_rsc_1_6_i_qb_d <=
      twiddle_rsc_1_6_i_qb_d;
  twiddle_rsc_1_6_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_6_i_1_inst_twiddle_rsc_1_6_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_1_7_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_inst_twiddle_rsc_1_7_i_qb_d,
      twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_rsc_1_7_i_oswt => reg_twiddle_rsc_1_7_i_oswt_cse,
      twiddle_rsc_1_7_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_inst_twiddle_rsc_1_7_i_qb_d_mxwt,
      twiddle_rsc_1_7_i_oswt_pff => and_403_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_inst_twiddle_rsc_1_7_i_qb_d <=
      twiddle_rsc_1_7_i_qb_d;
  twiddle_rsc_1_7_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_rsc_1_7_i_1_inst_twiddle_rsc_1_7_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_0_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_inst_twiddle_h_rsc_0_0_i_qb_d,
      twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_h_rsc_0_0_i_oswt => reg_twiddle_rsc_0_0_i_oswt_cse,
      twiddle_h_rsc_0_0_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_inst_twiddle_h_rsc_0_0_i_qb_d_mxwt,
      twiddle_h_rsc_0_0_i_oswt_pff => and_373_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_inst_twiddle_h_rsc_0_0_i_qb_d
      <= twiddle_h_rsc_0_0_i_qb_d;
  twiddle_h_rsc_0_0_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_0_i_1_inst_twiddle_h_rsc_0_0_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_1_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_inst_twiddle_h_rsc_0_1_i_qb_d,
      twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_h_rsc_0_1_i_oswt => reg_twiddle_rsc_0_1_i_oswt_cse,
      twiddle_h_rsc_0_1_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_inst_twiddle_h_rsc_0_1_i_qb_d_mxwt,
      twiddle_h_rsc_0_1_i_oswt_pff => and_375_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_inst_twiddle_h_rsc_0_1_i_qb_d
      <= twiddle_h_rsc_0_1_i_qb_d;
  twiddle_h_rsc_0_1_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_1_i_1_inst_twiddle_h_rsc_0_1_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_2_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_inst_twiddle_h_rsc_0_2_i_qb_d,
      twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_h_rsc_0_2_i_oswt => reg_twiddle_rsc_0_2_i_oswt_cse,
      twiddle_h_rsc_0_2_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_inst_twiddle_h_rsc_0_2_i_qb_d_mxwt,
      twiddle_h_rsc_0_2_i_oswt_pff => and_377_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_inst_twiddle_h_rsc_0_2_i_qb_d
      <= twiddle_h_rsc_0_2_i_qb_d;
  twiddle_h_rsc_0_2_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_2_i_1_inst_twiddle_h_rsc_0_2_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_3_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_inst_twiddle_h_rsc_0_3_i_qb_d,
      twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_h_rsc_0_3_i_oswt => reg_twiddle_rsc_0_3_i_oswt_cse,
      twiddle_h_rsc_0_3_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_inst_twiddle_h_rsc_0_3_i_qb_d_mxwt,
      twiddle_h_rsc_0_3_i_oswt_pff => and_379_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_inst_twiddle_h_rsc_0_3_i_qb_d
      <= twiddle_h_rsc_0_3_i_qb_d;
  twiddle_h_rsc_0_3_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_3_i_1_inst_twiddle_h_rsc_0_3_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_4_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_inst_twiddle_h_rsc_0_4_i_qb_d,
      twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_h_rsc_0_4_i_oswt => reg_twiddle_rsc_0_4_i_oswt_cse,
      twiddle_h_rsc_0_4_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_inst_twiddle_h_rsc_0_4_i_qb_d_mxwt,
      twiddle_h_rsc_0_4_i_oswt_pff => and_381_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_inst_twiddle_h_rsc_0_4_i_qb_d
      <= twiddle_h_rsc_0_4_i_qb_d;
  twiddle_h_rsc_0_4_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_4_i_1_inst_twiddle_h_rsc_0_4_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_5_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_inst_twiddle_h_rsc_0_5_i_qb_d,
      twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_h_rsc_0_5_i_oswt => reg_twiddle_rsc_0_5_i_oswt_cse,
      twiddle_h_rsc_0_5_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_inst_twiddle_h_rsc_0_5_i_qb_d_mxwt,
      twiddle_h_rsc_0_5_i_oswt_pff => and_383_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_inst_twiddle_h_rsc_0_5_i_qb_d
      <= twiddle_h_rsc_0_5_i_qb_d;
  twiddle_h_rsc_0_5_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_5_i_1_inst_twiddle_h_rsc_0_5_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_6_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_inst_twiddle_h_rsc_0_6_i_qb_d,
      twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_h_rsc_0_6_i_oswt => reg_twiddle_rsc_0_6_i_oswt_cse,
      twiddle_h_rsc_0_6_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_inst_twiddle_h_rsc_0_6_i_qb_d_mxwt,
      twiddle_h_rsc_0_6_i_oswt_pff => and_385_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_inst_twiddle_h_rsc_0_6_i_qb_d
      <= twiddle_h_rsc_0_6_i_qb_d;
  twiddle_h_rsc_0_6_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_6_i_1_inst_twiddle_h_rsc_0_6_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_7_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_inst_twiddle_h_rsc_0_7_i_qb_d,
      twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_h_rsc_0_7_i_oswt => reg_twiddle_rsc_0_7_i_oswt_cse,
      twiddle_h_rsc_0_7_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_inst_twiddle_h_rsc_0_7_i_qb_d_mxwt,
      twiddle_h_rsc_0_7_i_oswt_pff => and_387_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_inst_twiddle_h_rsc_0_7_i_qb_d
      <= twiddle_h_rsc_0_7_i_qb_d;
  twiddle_h_rsc_0_7_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_0_7_i_1_inst_twiddle_h_rsc_0_7_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_1_0_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_inst_twiddle_h_rsc_1_0_i_qb_d,
      twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_h_rsc_1_0_i_oswt => reg_twiddle_rsc_1_0_i_oswt_cse,
      twiddle_h_rsc_1_0_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_inst_twiddle_h_rsc_1_0_i_qb_d_mxwt,
      twiddle_h_rsc_1_0_i_oswt_pff => and_389_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_inst_twiddle_h_rsc_1_0_i_qb_d
      <= twiddle_h_rsc_1_0_i_qb_d;
  twiddle_h_rsc_1_0_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_0_i_1_inst_twiddle_h_rsc_1_0_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_1_1_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_inst_twiddle_h_rsc_1_1_i_qb_d,
      twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_h_rsc_1_1_i_oswt => reg_twiddle_rsc_1_1_i_oswt_cse,
      twiddle_h_rsc_1_1_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_inst_twiddle_h_rsc_1_1_i_qb_d_mxwt,
      twiddle_h_rsc_1_1_i_oswt_pff => and_391_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_inst_twiddle_h_rsc_1_1_i_qb_d
      <= twiddle_h_rsc_1_1_i_qb_d;
  twiddle_h_rsc_1_1_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_1_i_1_inst_twiddle_h_rsc_1_1_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_1_2_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_inst_twiddle_h_rsc_1_2_i_qb_d,
      twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_h_rsc_1_2_i_oswt => reg_twiddle_rsc_1_2_i_oswt_cse,
      twiddle_h_rsc_1_2_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_inst_twiddle_h_rsc_1_2_i_qb_d_mxwt,
      twiddle_h_rsc_1_2_i_oswt_pff => and_393_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_inst_twiddle_h_rsc_1_2_i_qb_d
      <= twiddle_h_rsc_1_2_i_qb_d;
  twiddle_h_rsc_1_2_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_2_i_1_inst_twiddle_h_rsc_1_2_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_1_3_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_inst_twiddle_h_rsc_1_3_i_qb_d,
      twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_h_rsc_1_3_i_oswt => reg_twiddle_rsc_1_3_i_oswt_cse,
      twiddle_h_rsc_1_3_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_inst_twiddle_h_rsc_1_3_i_qb_d_mxwt,
      twiddle_h_rsc_1_3_i_oswt_pff => and_395_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_inst_twiddle_h_rsc_1_3_i_qb_d
      <= twiddle_h_rsc_1_3_i_qb_d;
  twiddle_h_rsc_1_3_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_3_i_1_inst_twiddle_h_rsc_1_3_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_1_4_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_inst_twiddle_h_rsc_1_4_i_qb_d,
      twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_h_rsc_1_4_i_oswt => reg_twiddle_rsc_1_4_i_oswt_cse,
      twiddle_h_rsc_1_4_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_inst_twiddle_h_rsc_1_4_i_qb_d_mxwt,
      twiddle_h_rsc_1_4_i_oswt_pff => and_397_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_inst_twiddle_h_rsc_1_4_i_qb_d
      <= twiddle_h_rsc_1_4_i_qb_d;
  twiddle_h_rsc_1_4_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_4_i_1_inst_twiddle_h_rsc_1_4_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_1_5_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_inst_twiddle_h_rsc_1_5_i_qb_d,
      twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_h_rsc_1_5_i_oswt => reg_twiddle_rsc_1_5_i_oswt_cse,
      twiddle_h_rsc_1_5_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_inst_twiddle_h_rsc_1_5_i_qb_d_mxwt,
      twiddle_h_rsc_1_5_i_oswt_pff => and_399_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_inst_twiddle_h_rsc_1_5_i_qb_d
      <= twiddle_h_rsc_1_5_i_qb_d;
  twiddle_h_rsc_1_5_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_5_i_1_inst_twiddle_h_rsc_1_5_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_1_6_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_inst_twiddle_h_rsc_1_6_i_qb_d,
      twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_h_rsc_1_6_i_oswt => reg_twiddle_rsc_1_6_i_oswt_cse,
      twiddle_h_rsc_1_6_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_inst_twiddle_h_rsc_1_6_i_qb_d_mxwt,
      twiddle_h_rsc_1_6_i_oswt_pff => and_401_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_inst_twiddle_h_rsc_1_6_i_qb_d
      <= twiddle_h_rsc_1_6_i_qb_d;
  twiddle_h_rsc_1_6_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_6_i_1_inst_twiddle_h_rsc_1_6_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_1_7_i_qb_d => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_inst_twiddle_h_rsc_1_7_i_qb_d,
      twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => complete_rsci_wen_comp,
      core_wten => core_wten,
      twiddle_h_rsc_1_7_i_oswt => reg_twiddle_rsc_1_7_i_oswt_cse,
      twiddle_h_rsc_1_7_i_qb_d_mxwt => inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_inst_twiddle_h_rsc_1_7_i_qb_d_mxwt,
      twiddle_h_rsc_1_7_i_oswt_pff => and_403_rmff,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_inst_twiddle_h_rsc_1_7_i_qb_d
      <= twiddle_h_rsc_1_7_i_qb_d;
  twiddle_h_rsc_1_7_i_qb_d_mxwt <= inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_1_7_i_1_inst_twiddle_h_rsc_1_7_i_qb_d_mxwt;

  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_7_obj_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_7_obj
    PORT MAP(
      vec_rsc_triosy_1_7_lz => vec_rsc_triosy_1_7_lz,
      core_wten => core_wten,
      vec_rsc_triosy_1_7_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_6_obj_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_6_obj
    PORT MAP(
      vec_rsc_triosy_1_6_lz => vec_rsc_triosy_1_6_lz,
      core_wten => core_wten,
      vec_rsc_triosy_1_6_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_5_obj_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_5_obj
    PORT MAP(
      vec_rsc_triosy_1_5_lz => vec_rsc_triosy_1_5_lz,
      core_wten => core_wten,
      vec_rsc_triosy_1_5_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_4_obj_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_4_obj
    PORT MAP(
      vec_rsc_triosy_1_4_lz => vec_rsc_triosy_1_4_lz,
      core_wten => core_wten,
      vec_rsc_triosy_1_4_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_3_obj_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_3_obj
    PORT MAP(
      vec_rsc_triosy_1_3_lz => vec_rsc_triosy_1_3_lz,
      core_wten => core_wten,
      vec_rsc_triosy_1_3_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_2_obj_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_2_obj
    PORT MAP(
      vec_rsc_triosy_1_2_lz => vec_rsc_triosy_1_2_lz,
      core_wten => core_wten,
      vec_rsc_triosy_1_2_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_1_obj_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_1_obj
    PORT MAP(
      vec_rsc_triosy_1_1_lz => vec_rsc_triosy_1_1_lz,
      core_wten => core_wten,
      vec_rsc_triosy_1_1_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_0_obj_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_1_0_obj
    PORT MAP(
      vec_rsc_triosy_1_0_lz => vec_rsc_triosy_1_0_lz,
      core_wten => core_wten,
      vec_rsc_triosy_1_0_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_7_obj_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_7_obj
    PORT MAP(
      vec_rsc_triosy_0_7_lz => vec_rsc_triosy_0_7_lz,
      core_wten => core_wten,
      vec_rsc_triosy_0_7_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_6_obj_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_6_obj
    PORT MAP(
      vec_rsc_triosy_0_6_lz => vec_rsc_triosy_0_6_lz,
      core_wten => core_wten,
      vec_rsc_triosy_0_6_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_5_obj_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_5_obj
    PORT MAP(
      vec_rsc_triosy_0_5_lz => vec_rsc_triosy_0_5_lz,
      core_wten => core_wten,
      vec_rsc_triosy_0_5_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_4_obj_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_4_obj
    PORT MAP(
      vec_rsc_triosy_0_4_lz => vec_rsc_triosy_0_4_lz,
      core_wten => core_wten,
      vec_rsc_triosy_0_4_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_3_obj_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_3_obj
    PORT MAP(
      vec_rsc_triosy_0_3_lz => vec_rsc_triosy_0_3_lz,
      core_wten => core_wten,
      vec_rsc_triosy_0_3_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_2_obj_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_2_obj
    PORT MAP(
      vec_rsc_triosy_0_2_lz => vec_rsc_triosy_0_2_lz,
      core_wten => core_wten,
      vec_rsc_triosy_0_2_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_1_obj_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_1_obj
    PORT MAP(
      vec_rsc_triosy_0_1_lz => vec_rsc_triosy_0_1_lz,
      core_wten => core_wten,
      vec_rsc_triosy_0_1_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_0_obj_inst : inPlaceNTT_DIF_precomp_core_vec_rsc_triosy_0_0_obj
    PORT MAP(
      vec_rsc_triosy_0_0_lz => vec_rsc_triosy_0_0_lz,
      core_wten => core_wten,
      vec_rsc_triosy_0_0_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_p_rsc_triosy_obj_inst : inPlaceNTT_DIF_precomp_core_p_rsc_triosy_obj
    PORT MAP(
      p_rsc_triosy_lz => p_rsc_triosy_lz,
      core_wten => core_wten,
      p_rsc_triosy_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_r_rsc_triosy_obj_inst : inPlaceNTT_DIF_precomp_core_r_rsc_triosy_obj
    PORT MAP(
      r_rsc_triosy_lz => r_rsc_triosy_lz,
      core_wten => core_wten,
      r_rsc_triosy_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_7_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_7_obj
    PORT MAP(
      twiddle_rsc_triosy_1_7_lz => twiddle_rsc_triosy_1_7_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_1_7_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_6_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_6_obj
    PORT MAP(
      twiddle_rsc_triosy_1_6_lz => twiddle_rsc_triosy_1_6_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_1_6_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_5_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_5_obj
    PORT MAP(
      twiddle_rsc_triosy_1_5_lz => twiddle_rsc_triosy_1_5_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_1_5_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_4_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_4_obj
    PORT MAP(
      twiddle_rsc_triosy_1_4_lz => twiddle_rsc_triosy_1_4_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_1_4_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_3_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_3_obj
    PORT MAP(
      twiddle_rsc_triosy_1_3_lz => twiddle_rsc_triosy_1_3_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_1_3_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_2_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_2_obj
    PORT MAP(
      twiddle_rsc_triosy_1_2_lz => twiddle_rsc_triosy_1_2_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_1_2_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_1_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_1_obj
    PORT MAP(
      twiddle_rsc_triosy_1_1_lz => twiddle_rsc_triosy_1_1_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_1_1_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_0_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_1_0_obj
    PORT MAP(
      twiddle_rsc_triosy_1_0_lz => twiddle_rsc_triosy_1_0_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_1_0_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_7_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_7_obj
    PORT MAP(
      twiddle_rsc_triosy_0_7_lz => twiddle_rsc_triosy_0_7_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_7_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_6_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_6_obj
    PORT MAP(
      twiddle_rsc_triosy_0_6_lz => twiddle_rsc_triosy_0_6_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_6_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_5_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_5_obj
    PORT MAP(
      twiddle_rsc_triosy_0_5_lz => twiddle_rsc_triosy_0_5_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_5_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_4_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_4_obj
    PORT MAP(
      twiddle_rsc_triosy_0_4_lz => twiddle_rsc_triosy_0_4_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_4_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_3_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_3_obj
    PORT MAP(
      twiddle_rsc_triosy_0_3_lz => twiddle_rsc_triosy_0_3_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_3_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_2_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_2_obj
    PORT MAP(
      twiddle_rsc_triosy_0_2_lz => twiddle_rsc_triosy_0_2_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_2_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_1_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_1_obj
    PORT MAP(
      twiddle_rsc_triosy_0_1_lz => twiddle_rsc_triosy_0_1_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_1_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_0_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_rsc_triosy_0_0_obj
    PORT MAP(
      twiddle_rsc_triosy_0_0_lz => twiddle_rsc_triosy_0_0_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_0_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_7_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_7_obj
    PORT MAP(
      twiddle_h_rsc_triosy_1_7_lz => twiddle_h_rsc_triosy_1_7_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_1_7_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_6_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_6_obj
    PORT MAP(
      twiddle_h_rsc_triosy_1_6_lz => twiddle_h_rsc_triosy_1_6_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_1_6_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_5_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_5_obj
    PORT MAP(
      twiddle_h_rsc_triosy_1_5_lz => twiddle_h_rsc_triosy_1_5_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_1_5_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_4_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_4_obj
    PORT MAP(
      twiddle_h_rsc_triosy_1_4_lz => twiddle_h_rsc_triosy_1_4_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_1_4_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_3_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_3_obj
    PORT MAP(
      twiddle_h_rsc_triosy_1_3_lz => twiddle_h_rsc_triosy_1_3_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_1_3_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_2_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_2_obj
    PORT MAP(
      twiddle_h_rsc_triosy_1_2_lz => twiddle_h_rsc_triosy_1_2_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_1_2_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_1_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_1_obj
    PORT MAP(
      twiddle_h_rsc_triosy_1_1_lz => twiddle_h_rsc_triosy_1_1_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_1_1_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_0_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_1_0_obj
    PORT MAP(
      twiddle_h_rsc_triosy_1_0_lz => twiddle_h_rsc_triosy_1_0_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_1_0_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_7_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_7_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_7_lz => twiddle_h_rsc_triosy_0_7_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_7_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_6_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_6_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_6_lz => twiddle_h_rsc_triosy_0_6_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_6_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_5_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_5_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_5_lz => twiddle_h_rsc_triosy_0_5_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_5_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_4_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_4_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_4_lz => twiddle_h_rsc_triosy_0_4_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_4_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_3_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_3_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_3_lz => twiddle_h_rsc_triosy_0_3_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_3_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_2_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_2_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_2_lz => twiddle_h_rsc_triosy_0_2_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_2_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_1_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_1_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_1_lz => twiddle_h_rsc_triosy_0_1_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_1_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_0_obj_inst : inPlaceNTT_DIF_precomp_core_twiddle_h_rsc_triosy_0_0_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_0_lz => twiddle_h_rsc_triosy_0_0_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_0_obj_iswt0 => reg_vec_rsc_triosy_1_7_obj_iswt0_cse
    );
  inPlaceNTT_DIF_precomp_core_staller_inst : inPlaceNTT_DIF_precomp_core_staller
    PORT MAP(
      clk => clk,
      rst => rst,
      core_wten => core_wten,
      complete_rsci_wen_comp => complete_rsci_wen_comp,
      core_wten_pff => core_wten_iff
    );
  inPlaceNTT_DIF_precomp_core_core_fsm_inst : inPlaceNTT_DIF_precomp_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      complete_rsci_wen_comp => complete_rsci_wen_comp,
      fsm_output => inPlaceNTT_DIF_precomp_core_core_fsm_inst_fsm_output,
      main_C_0_tr0 => inPlaceNTT_DIF_precomp_core_core_fsm_inst_main_C_0_tr0,
      VEC_LOOP_C_11_tr0 => inPlaceNTT_DIF_precomp_core_core_fsm_inst_VEC_LOOP_C_11_tr0,
      COMP_LOOP_C_4_tr0 => inPlaceNTT_DIF_precomp_core_core_fsm_inst_COMP_LOOP_C_4_tr0,
      STAGE_LOOP_C_1_tr0 => inPlaceNTT_DIF_precomp_core_core_fsm_inst_STAGE_LOOP_C_1_tr0
    );
  fsm_output <= inPlaceNTT_DIF_precomp_core_core_fsm_inst_fsm_output;
  inPlaceNTT_DIF_precomp_core_core_fsm_inst_main_C_0_tr0 <= NOT VEC_LOOP_VEC_LOOP_and_10_itm;
  inPlaceNTT_DIF_precomp_core_core_fsm_inst_VEC_LOOP_C_11_tr0 <= VEC_LOOP_j_10_0_sva_1(10);
  inPlaceNTT_DIF_precomp_core_core_fsm_inst_COMP_LOOP_C_4_tr0 <= NOT (READSLICE_1_11(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(COMP_LOOP_k_10_0_sva_2)
      + SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10 DOWNTO 1)))) + SIGNED'( "00000000001"),
      11)), 10));
  inPlaceNTT_DIF_precomp_core_core_fsm_inst_STAGE_LOOP_C_1_tr0 <= NOT STAGE_LOOP_acc_itm_4_1;

  or_15_rmff <= and_157_cse OR and_158_cse OR and_159_cse;
  and_161_rmff <= VEC_LOOP_nor_12_cse AND VEC_LOOP_nor_19_cse AND (fsm_output(6));
  VEC_LOOP_mux1h_rmff <= MUX1HOT_v_6_3_2((VEC_LOOP_acc_1_tmp(8 DOWNTO 3)), (COMP_LOOP_twiddle_f_lshift_itm(8
      DOWNTO 3)), (VEC_LOOP_acc_10_cse_sva(8 DOWNTO 3)), STD_LOGIC_VECTOR'( (fsm_output(6))
      & (fsm_output(9)) & (fsm_output(16))));
  VEC_LOOP_mux_4_rmff <= MUX_v_32_2_2(modulo_add_cmp_return_rsc_z, mult_cmp_return_rsc_z,
      fsm_output(16));
  or_21_rmff <= and_157_cse OR and_159_cse;
  or_24_rmff <= and_178_cse OR and_179_cse OR and_180_cse;
  and_182_rmff <= VEC_LOOP_nor_12_cse AND and_dcpl_25 AND (fsm_output(6));
  or_26_rmff <= and_178_cse OR and_180_cse;
  or_29_rmff <= and_191_cse OR and_192_cse OR and_193_cse;
  and_195_rmff <= VEC_LOOP_nor_12_cse AND and_dcpl_33 AND (fsm_output(6));
  or_31_rmff <= and_191_cse OR and_193_cse;
  or_34_rmff <= and_204_cse OR and_205_cse OR and_206_cse;
  and_208_rmff <= VEC_LOOP_nor_12_cse AND and_dcpl_41 AND (fsm_output(6));
  or_36_rmff <= and_204_cse OR and_206_cse;
  or_39_rmff <= and_217_cse OR and_218_cse OR and_219_cse;
  and_221_rmff <= and_dcpl_49 AND VEC_LOOP_nor_19_cse AND (fsm_output(6));
  or_41_rmff <= and_217_cse OR and_219_cse;
  or_44_rmff <= and_230_cse OR and_231_cse OR and_232_cse;
  and_234_rmff <= and_dcpl_49 AND and_dcpl_25 AND (fsm_output(6));
  or_46_rmff <= and_230_cse OR and_232_cse;
  or_49_rmff <= and_243_cse OR and_244_cse OR and_245_cse;
  and_247_rmff <= and_dcpl_49 AND and_dcpl_33 AND (fsm_output(6));
  or_51_rmff <= and_243_cse OR and_245_cse;
  or_54_rmff <= and_256_cse OR and_257_cse OR and_258_cse;
  and_260_rmff <= and_dcpl_49 AND and_dcpl_41 AND (fsm_output(6));
  or_56_rmff <= and_256_cse OR and_258_cse;
  or_59_rmff <= and_269_cse OR and_270_cse OR and_271_cse;
  and_273_rmff <= and_dcpl_69 AND VEC_LOOP_nor_19_cse AND (fsm_output(6));
  or_61_rmff <= and_269_cse OR and_271_cse;
  or_64_rmff <= and_282_cse OR and_283_cse OR and_284_cse;
  and_286_rmff <= and_dcpl_69 AND and_dcpl_25 AND (fsm_output(6));
  or_66_rmff <= and_282_cse OR and_284_cse;
  or_69_rmff <= and_295_cse OR and_296_cse OR and_297_cse;
  and_299_rmff <= and_dcpl_69 AND and_dcpl_33 AND (fsm_output(6));
  or_71_rmff <= and_295_cse OR and_297_cse;
  or_74_rmff <= and_308_cse OR and_309_cse OR and_310_cse;
  and_312_rmff <= and_dcpl_69 AND and_dcpl_41 AND (fsm_output(6));
  or_76_rmff <= and_308_cse OR and_310_cse;
  or_79_rmff <= and_321_cse OR and_322_cse OR and_323_cse;
  and_325_rmff <= and_dcpl_89 AND VEC_LOOP_nor_19_cse AND (fsm_output(6));
  or_81_rmff <= and_321_cse OR and_323_cse;
  or_84_rmff <= and_334_cse OR and_335_cse OR and_336_cse;
  and_338_rmff <= and_dcpl_89 AND and_dcpl_25 AND (fsm_output(6));
  or_86_rmff <= and_334_cse OR and_336_cse;
  or_89_rmff <= and_347_cse OR and_348_cse OR and_349_cse;
  and_351_rmff <= and_dcpl_89 AND and_dcpl_33 AND (fsm_output(6));
  or_91_rmff <= and_347_cse OR and_349_cse;
  or_94_rmff <= and_360_cse OR and_361_cse OR and_362_cse;
  and_364_rmff <= and_dcpl_89 AND and_dcpl_41 AND (fsm_output(6));
  or_96_rmff <= and_360_cse OR and_362_cse;
  and_373_rmff <= and_dcpl_104 AND and_dcpl_103 AND (fsm_output(4));
  and_375_rmff <= and_dcpl_104 AND and_dcpl_106 AND (fsm_output(4));
  and_377_rmff <= and_dcpl_104 AND and_dcpl_108 AND (fsm_output(4));
  and_379_rmff <= and_dcpl_104 AND and_dcpl_110 AND (fsm_output(4));
  and_381_rmff <= and_dcpl_112 AND and_dcpl_103 AND (fsm_output(4));
  and_383_rmff <= and_dcpl_112 AND and_dcpl_106 AND (fsm_output(4));
  and_385_rmff <= and_dcpl_112 AND and_dcpl_108 AND (fsm_output(4));
  and_387_rmff <= and_dcpl_112 AND and_dcpl_110 AND (fsm_output(4));
  and_389_rmff <= and_dcpl_117 AND and_dcpl_103 AND (fsm_output(4));
  and_391_rmff <= and_dcpl_117 AND and_dcpl_106 AND (fsm_output(4));
  and_393_rmff <= and_dcpl_117 AND and_dcpl_108 AND (fsm_output(4));
  and_395_rmff <= and_dcpl_117 AND and_dcpl_110 AND (fsm_output(4));
  and_397_rmff <= and_dcpl_122 AND and_dcpl_103 AND (fsm_output(4));
  and_399_rmff <= and_dcpl_122 AND and_dcpl_106 AND (fsm_output(4));
  and_401_rmff <= and_dcpl_122 AND and_dcpl_108 AND (fsm_output(4));
  and_403_rmff <= and_dcpl_122 AND and_dcpl_110 AND (fsm_output(4));
  or_116_rmff <= CONV_SL_1_1(fsm_output(15 DOWNTO 9)/=STD_LOGIC_VECTOR'("0000000"));
  or_118_rmff <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("00"));
  COMP_LOOP_twiddle_f_and_1_cse <= complete_rsci_wen_comp AND (fsm_output(3));
  COMP_LOOP_twiddle_help_and_cse <= COMP_LOOP_twiddle_f_equal_tmp AND (NOT or_tmp_141);
  COMP_LOOP_twiddle_help_and_1_cse <= (COMP_LOOP_twiddle_f_mul_cse_sva(0)) AND COMP_LOOP_twiddle_f_nor_itm
      AND (NOT or_tmp_141);
  COMP_LOOP_twiddle_help_and_2_cse <= (COMP_LOOP_twiddle_f_mul_cse_sva(1)) AND COMP_LOOP_twiddle_f_nor_1_itm
      AND (NOT or_tmp_141);
  COMP_LOOP_twiddle_help_and_3_cse <= COMP_LOOP_twiddle_f_equal_tmp_3 AND (NOT or_tmp_141);
  COMP_LOOP_twiddle_help_and_4_cse <= (COMP_LOOP_twiddle_f_mul_cse_sva(2)) AND COMP_LOOP_twiddle_f_nor_3_itm
      AND (NOT or_tmp_141);
  COMP_LOOP_twiddle_help_and_5_cse <= COMP_LOOP_twiddle_f_equal_tmp_5 AND (NOT or_tmp_141);
  COMP_LOOP_twiddle_help_and_6_cse <= COMP_LOOP_twiddle_f_equal_tmp_6 AND (NOT or_tmp_141);
  COMP_LOOP_twiddle_help_and_7_cse <= COMP_LOOP_twiddle_f_equal_tmp_7 AND (NOT or_tmp_141);
  COMP_LOOP_twiddle_help_and_8_cse <= (COMP_LOOP_twiddle_f_mul_cse_sva(9)) AND COMP_LOOP_twiddle_f_nor_6_itm
      AND (NOT or_tmp_141);
  COMP_LOOP_twiddle_help_and_9_cse <= COMP_LOOP_twiddle_f_equal_tmp_9 AND (NOT or_tmp_141);
  COMP_LOOP_twiddle_help_and_10_cse <= COMP_LOOP_twiddle_f_equal_tmp_10 AND (NOT
      or_tmp_141);
  COMP_LOOP_twiddle_help_and_11_cse <= COMP_LOOP_twiddle_f_equal_tmp_11 AND (NOT
      or_tmp_141);
  COMP_LOOP_twiddle_help_and_12_cse <= COMP_LOOP_twiddle_f_equal_tmp_12 AND (NOT
      or_tmp_141);
  COMP_LOOP_twiddle_help_and_13_cse <= COMP_LOOP_twiddle_f_equal_tmp_13 AND (NOT
      or_tmp_141);
  COMP_LOOP_twiddle_help_and_14_cse <= COMP_LOOP_twiddle_f_equal_tmp_14 AND (NOT
      or_tmp_141);
  COMP_LOOP_twiddle_help_and_15_cse <= COMP_LOOP_twiddle_f_equal_tmp_15 AND (NOT
      or_tmp_141);
  COMP_LOOP_twiddle_help_and_16_cse <= complete_rsci_wen_comp AND (NOT or_tmp_141);
  VEC_LOOP_and_cse <= complete_rsci_wen_comp AND (fsm_output(6));
  VEC_LOOP_nor_12_cse <= NOT((VEC_LOOP_acc_10_tmp(9)) OR (VEC_LOOP_acc_10_tmp(2)));
  VEC_LOOP_nor_19_cse <= NOT(CONV_SL_1_1(VEC_LOOP_acc_10_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  VEC_LOOP_nor_2_cse <= NOT((VEC_LOOP_acc_1_tmp(9)) OR (VEC_LOOP_acc_1_tmp(2)));
  VEC_LOOP_nor_9_cse <= NOT(CONV_SL_1_1(VEC_LOOP_acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  STAGE_LOOP_i_3_0_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_LOOP_i_3_0_sva)
      + UNSIGNED'( "1111"), 4));
  VEC_LOOP_acc_1_tmp <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_twiddle_f_lshift_itm)
      + UNSIGNED(COMP_LOOP_k_10_0_sva_9_0), 10));
  COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'(
      UNSIGNED(COMP_LOOP_twiddle_f_lshift_itm) * UNSIGNED(COMP_LOOP_k_10_0_sva_9_0)),
      10));
  VEC_LOOP_acc_10_tmp <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_twiddle_f_lshift_itm)
      + UNSIGNED(COMP_LOOP_k_10_0_sva_9_0) + UNSIGNED(STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)), 10));
  COMP_LOOP_k_10_0_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_0_sva_9_0),
      10), 11) + UNSIGNED'( "00000000001"), 11));
  and_dcpl_7 <= NOT((COMP_LOOP_twiddle_f_lshift_itm(2)) OR (COMP_LOOP_twiddle_f_lshift_itm(9)));
  and_dcpl_8 <= NOT(CONV_SL_1_1(COMP_LOOP_twiddle_f_lshift_itm(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_13 <= NOT((VEC_LOOP_acc_10_cse_sva(2)) OR (VEC_LOOP_acc_10_cse_sva(9)));
  and_dcpl_14 <= NOT(CONV_SL_1_1(VEC_LOOP_acc_10_cse_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_19 <= CONV_SL_1_1(COMP_LOOP_twiddle_f_lshift_itm(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_21 <= CONV_SL_1_1(VEC_LOOP_acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_23 <= CONV_SL_1_1(VEC_LOOP_acc_10_cse_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_25 <= CONV_SL_1_1(VEC_LOOP_acc_10_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_27 <= CONV_SL_1_1(COMP_LOOP_twiddle_f_lshift_itm(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_29 <= CONV_SL_1_1(VEC_LOOP_acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_31 <= CONV_SL_1_1(VEC_LOOP_acc_10_cse_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_33 <= CONV_SL_1_1(VEC_LOOP_acc_10_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_35 <= CONV_SL_1_1(COMP_LOOP_twiddle_f_lshift_itm(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_37 <= CONV_SL_1_1(VEC_LOOP_acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_39 <= CONV_SL_1_1(VEC_LOOP_acc_10_cse_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_41 <= CONV_SL_1_1(VEC_LOOP_acc_10_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_43 <= (COMP_LOOP_twiddle_f_lshift_itm(2)) AND (NOT (COMP_LOOP_twiddle_f_lshift_itm(9)));
  and_dcpl_45 <= (NOT (VEC_LOOP_acc_1_tmp(9))) AND (VEC_LOOP_acc_1_tmp(2));
  and_dcpl_47 <= (VEC_LOOP_acc_10_cse_sva(2)) AND (NOT (VEC_LOOP_acc_10_cse_sva(9)));
  and_dcpl_49 <= (NOT (VEC_LOOP_acc_10_tmp(9))) AND (VEC_LOOP_acc_10_tmp(2));
  and_dcpl_63 <= (NOT (COMP_LOOP_twiddle_f_lshift_itm(2))) AND (COMP_LOOP_twiddle_f_lshift_itm(9));
  and_dcpl_65 <= (VEC_LOOP_acc_1_tmp(9)) AND (NOT (VEC_LOOP_acc_1_tmp(2)));
  and_dcpl_67 <= (NOT (VEC_LOOP_acc_10_cse_sva(2))) AND (VEC_LOOP_acc_10_cse_sva(9));
  and_dcpl_69 <= (VEC_LOOP_acc_10_tmp(9)) AND (NOT (VEC_LOOP_acc_10_tmp(2)));
  and_dcpl_83 <= (COMP_LOOP_twiddle_f_lshift_itm(2)) AND (COMP_LOOP_twiddle_f_lshift_itm(9));
  and_dcpl_85 <= (VEC_LOOP_acc_1_tmp(9)) AND (VEC_LOOP_acc_1_tmp(2));
  and_dcpl_87 <= (VEC_LOOP_acc_10_cse_sva(2)) AND (VEC_LOOP_acc_10_cse_sva(9));
  and_dcpl_89 <= (VEC_LOOP_acc_10_tmp(9)) AND (VEC_LOOP_acc_10_tmp(2));
  and_dcpl_103 <= NOT(CONV_SL_1_1(COMP_LOOP_twiddle_f_mul_cse_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_104 <= NOT((COMP_LOOP_twiddle_f_mul_cse_sva(9)) OR (COMP_LOOP_twiddle_f_mul_cse_sva(2)));
  and_dcpl_106 <= CONV_SL_1_1(COMP_LOOP_twiddle_f_mul_cse_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_108 <= CONV_SL_1_1(COMP_LOOP_twiddle_f_mul_cse_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_110 <= CONV_SL_1_1(COMP_LOOP_twiddle_f_mul_cse_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_112 <= (NOT (COMP_LOOP_twiddle_f_mul_cse_sva(9))) AND (COMP_LOOP_twiddle_f_mul_cse_sva(2));
  and_dcpl_117 <= (COMP_LOOP_twiddle_f_mul_cse_sva(9)) AND (NOT (COMP_LOOP_twiddle_f_mul_cse_sva(2)));
  and_dcpl_122 <= (COMP_LOOP_twiddle_f_mul_cse_sva(9)) AND (COMP_LOOP_twiddle_f_mul_cse_sva(2));
  and_dcpl_129 <= NOT((fsm_output(21)) OR (fsm_output(20)) OR (fsm_output(0)));
  and_dcpl_131 <= and_dcpl_129 AND (NOT (fsm_output(1))) AND (NOT (fsm_output(19)));
  and_157_cse <= and_dcpl_8 AND and_dcpl_7 AND (fsm_output(9));
  and_159_cse <= and_dcpl_14 AND and_dcpl_13 AND (fsm_output(16));
  and_158_cse <= VEC_LOOP_nor_2_cse AND VEC_LOOP_nor_9_cse AND (fsm_output(6));
  and_178_cse <= and_dcpl_19 AND and_dcpl_7 AND (fsm_output(9));
  and_180_cse <= and_dcpl_23 AND and_dcpl_13 AND (fsm_output(16));
  and_179_cse <= VEC_LOOP_nor_2_cse AND and_dcpl_21 AND (fsm_output(6));
  and_191_cse <= and_dcpl_27 AND and_dcpl_7 AND (fsm_output(9));
  and_193_cse <= and_dcpl_31 AND and_dcpl_13 AND (fsm_output(16));
  and_192_cse <= VEC_LOOP_nor_2_cse AND and_dcpl_29 AND (fsm_output(6));
  and_204_cse <= and_dcpl_35 AND and_dcpl_7 AND (fsm_output(9));
  and_206_cse <= and_dcpl_39 AND and_dcpl_13 AND (fsm_output(16));
  and_205_cse <= VEC_LOOP_nor_2_cse AND and_dcpl_37 AND (fsm_output(6));
  and_217_cse <= and_dcpl_8 AND and_dcpl_43 AND (fsm_output(9));
  and_219_cse <= and_dcpl_14 AND and_dcpl_47 AND (fsm_output(16));
  and_218_cse <= and_dcpl_45 AND VEC_LOOP_nor_9_cse AND (fsm_output(6));
  and_230_cse <= and_dcpl_19 AND and_dcpl_43 AND (fsm_output(9));
  and_232_cse <= and_dcpl_23 AND and_dcpl_47 AND (fsm_output(16));
  and_231_cse <= and_dcpl_45 AND and_dcpl_21 AND (fsm_output(6));
  and_243_cse <= and_dcpl_27 AND and_dcpl_43 AND (fsm_output(9));
  and_245_cse <= and_dcpl_31 AND and_dcpl_47 AND (fsm_output(16));
  and_244_cse <= and_dcpl_45 AND and_dcpl_29 AND (fsm_output(6));
  and_256_cse <= and_dcpl_35 AND and_dcpl_43 AND (fsm_output(9));
  and_258_cse <= and_dcpl_39 AND and_dcpl_47 AND (fsm_output(16));
  and_257_cse <= and_dcpl_45 AND and_dcpl_37 AND (fsm_output(6));
  and_269_cse <= and_dcpl_8 AND and_dcpl_63 AND (fsm_output(9));
  and_271_cse <= and_dcpl_14 AND and_dcpl_67 AND (fsm_output(16));
  and_270_cse <= and_dcpl_65 AND VEC_LOOP_nor_9_cse AND (fsm_output(6));
  and_282_cse <= and_dcpl_19 AND and_dcpl_63 AND (fsm_output(9));
  and_284_cse <= and_dcpl_23 AND and_dcpl_67 AND (fsm_output(16));
  and_283_cse <= and_dcpl_65 AND and_dcpl_21 AND (fsm_output(6));
  and_295_cse <= and_dcpl_27 AND and_dcpl_63 AND (fsm_output(9));
  and_297_cse <= and_dcpl_31 AND and_dcpl_67 AND (fsm_output(16));
  and_296_cse <= and_dcpl_65 AND and_dcpl_29 AND (fsm_output(6));
  and_308_cse <= and_dcpl_35 AND and_dcpl_63 AND (fsm_output(9));
  and_310_cse <= and_dcpl_39 AND and_dcpl_67 AND (fsm_output(16));
  and_309_cse <= and_dcpl_65 AND and_dcpl_37 AND (fsm_output(6));
  and_321_cse <= and_dcpl_8 AND and_dcpl_83 AND (fsm_output(9));
  and_323_cse <= and_dcpl_14 AND and_dcpl_87 AND (fsm_output(16));
  and_322_cse <= and_dcpl_85 AND VEC_LOOP_nor_9_cse AND (fsm_output(6));
  and_334_cse <= and_dcpl_19 AND and_dcpl_83 AND (fsm_output(9));
  and_336_cse <= and_dcpl_23 AND and_dcpl_87 AND (fsm_output(16));
  and_335_cse <= and_dcpl_85 AND and_dcpl_21 AND (fsm_output(6));
  and_347_cse <= and_dcpl_27 AND and_dcpl_83 AND (fsm_output(9));
  and_349_cse <= and_dcpl_31 AND and_dcpl_87 AND (fsm_output(16));
  and_348_cse <= and_dcpl_85 AND and_dcpl_29 AND (fsm_output(6));
  and_360_cse <= and_dcpl_35 AND and_dcpl_83 AND (fsm_output(9));
  and_362_cse <= and_dcpl_39 AND and_dcpl_87 AND (fsm_output(16));
  and_361_cse <= and_dcpl_85 AND and_dcpl_37 AND (fsm_output(6));
  or_tmp_141 <= NOT((fsm_output(18)) OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(2))
      OR (fsm_output(5)) OR (NOT and_dcpl_131));
  STAGE_LOOP_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT STAGE_LOOP_i_3_0_sva_2))
      + SIGNED'( "00001"), 5));
  STAGE_LOOP_acc_itm_4_1 <= STAGE_LOOP_acc_nl(4);
  vec_rsc_0_0_i_adra_d <= (VEC_LOOP_acc_10_tmp(8 DOWNTO 3)) & VEC_LOOP_mux1h_rmff;
  vec_rsc_0_0_i_wea_d <= vec_rsc_0_0_i_wea_d_reg;
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg;
  vec_rsc_0_1_i_adra_d <= (VEC_LOOP_acc_10_tmp(8 DOWNTO 3)) & VEC_LOOP_mux1h_rmff;
  vec_rsc_0_1_i_wea_d <= vec_rsc_0_1_i_wea_d_reg;
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg;
  vec_rsc_0_2_i_adra_d <= (VEC_LOOP_acc_10_tmp(8 DOWNTO 3)) & VEC_LOOP_mux1h_rmff;
  vec_rsc_0_2_i_wea_d <= vec_rsc_0_2_i_wea_d_reg;
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg;
  vec_rsc_0_3_i_adra_d <= (VEC_LOOP_acc_10_tmp(8 DOWNTO 3)) & VEC_LOOP_mux1h_rmff;
  vec_rsc_0_3_i_wea_d <= vec_rsc_0_3_i_wea_d_reg;
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg;
  vec_rsc_0_4_i_adra_d <= (VEC_LOOP_acc_10_tmp(8 DOWNTO 3)) & VEC_LOOP_mux1h_rmff;
  vec_rsc_0_4_i_wea_d <= vec_rsc_0_4_i_wea_d_reg;
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg;
  vec_rsc_0_5_i_adra_d <= (VEC_LOOP_acc_10_tmp(8 DOWNTO 3)) & VEC_LOOP_mux1h_rmff;
  vec_rsc_0_5_i_wea_d <= vec_rsc_0_5_i_wea_d_reg;
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg;
  vec_rsc_0_6_i_adra_d <= (VEC_LOOP_acc_10_tmp(8 DOWNTO 3)) & VEC_LOOP_mux1h_rmff;
  vec_rsc_0_6_i_wea_d <= vec_rsc_0_6_i_wea_d_reg;
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg;
  vec_rsc_0_7_i_adra_d <= (VEC_LOOP_acc_10_tmp(8 DOWNTO 3)) & VEC_LOOP_mux1h_rmff;
  vec_rsc_0_7_i_wea_d <= vec_rsc_0_7_i_wea_d_reg;
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg;
  vec_rsc_1_0_i_adra_d <= (VEC_LOOP_acc_10_tmp(8 DOWNTO 3)) & VEC_LOOP_mux1h_rmff;
  vec_rsc_1_0_i_wea_d <= vec_rsc_1_0_i_wea_d_reg;
  vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg;
  vec_rsc_1_1_i_adra_d <= (VEC_LOOP_acc_10_tmp(8 DOWNTO 3)) & VEC_LOOP_mux1h_rmff;
  vec_rsc_1_1_i_wea_d <= vec_rsc_1_1_i_wea_d_reg;
  vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg;
  vec_rsc_1_2_i_adra_d <= (VEC_LOOP_acc_10_tmp(8 DOWNTO 3)) & VEC_LOOP_mux1h_rmff;
  vec_rsc_1_2_i_wea_d <= vec_rsc_1_2_i_wea_d_reg;
  vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg;
  vec_rsc_1_3_i_adra_d <= (VEC_LOOP_acc_10_tmp(8 DOWNTO 3)) & VEC_LOOP_mux1h_rmff;
  vec_rsc_1_3_i_wea_d <= vec_rsc_1_3_i_wea_d_reg;
  vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg;
  vec_rsc_1_4_i_adra_d <= (VEC_LOOP_acc_10_tmp(8 DOWNTO 3)) & VEC_LOOP_mux1h_rmff;
  vec_rsc_1_4_i_wea_d <= vec_rsc_1_4_i_wea_d_reg;
  vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg;
  vec_rsc_1_5_i_adra_d <= (VEC_LOOP_acc_10_tmp(8 DOWNTO 3)) & VEC_LOOP_mux1h_rmff;
  vec_rsc_1_5_i_wea_d <= vec_rsc_1_5_i_wea_d_reg;
  vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg;
  vec_rsc_1_6_i_adra_d <= (VEC_LOOP_acc_10_tmp(8 DOWNTO 3)) & VEC_LOOP_mux1h_rmff;
  vec_rsc_1_6_i_wea_d <= vec_rsc_1_6_i_wea_d_reg;
  vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg;
  vec_rsc_1_7_i_adra_d <= (VEC_LOOP_acc_10_tmp(8 DOWNTO 3)) & VEC_LOOP_mux1h_rmff;
  vec_rsc_1_7_i_wea_d <= vec_rsc_1_7_i_wea_d_reg;
  vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d <= vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_reg;
  twiddle_rsc_0_0_i_adrb_d_pff <= COMP_LOOP_twiddle_f_mul_cse_sva(8 DOWNTO 3);
  twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d_reg;
  vec_rsc_0_0_i_da_d <= vec_rsc_0_0_i_da_d_reg;
  vec_rsc_0_1_i_da_d <= vec_rsc_0_1_i_da_d_reg;
  vec_rsc_0_2_i_da_d <= vec_rsc_0_2_i_da_d_reg;
  vec_rsc_0_3_i_da_d <= vec_rsc_0_3_i_da_d_reg;
  vec_rsc_0_4_i_da_d <= vec_rsc_0_4_i_da_d_reg;
  vec_rsc_0_5_i_da_d <= vec_rsc_0_5_i_da_d_reg;
  vec_rsc_0_6_i_da_d <= vec_rsc_0_6_i_da_d_reg;
  vec_rsc_0_7_i_da_d <= vec_rsc_0_7_i_da_d_reg;
  vec_rsc_1_0_i_da_d <= vec_rsc_1_0_i_da_d_reg;
  vec_rsc_1_1_i_da_d <= vec_rsc_1_1_i_da_d_reg;
  vec_rsc_1_2_i_da_d <= vec_rsc_1_2_i_da_d_reg;
  vec_rsc_1_3_i_da_d <= vec_rsc_1_3_i_da_d_reg;
  vec_rsc_1_4_i_da_d <= vec_rsc_1_4_i_da_d_reg;
  vec_rsc_1_5_i_da_d <= vec_rsc_1_5_i_da_d_reg;
  vec_rsc_1_6_i_da_d <= vec_rsc_1_6_i_da_d_reg;
  vec_rsc_1_7_i_da_d <= vec_rsc_1_7_i_da_d_reg;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( complete_rsci_wen_comp = '1' ) THEN
        tmp_lpi_4_dfm <= MUX1HOT_v_32_16_2((vec_rsc_0_0_i_qa_d_mxwt(31 DOWNTO 0)),
            (vec_rsc_0_1_i_qa_d_mxwt(31 DOWNTO 0)), (vec_rsc_0_2_i_qa_d_mxwt(31 DOWNTO
            0)), (vec_rsc_0_3_i_qa_d_mxwt(31 DOWNTO 0)), (vec_rsc_0_4_i_qa_d_mxwt(31
            DOWNTO 0)), (vec_rsc_0_5_i_qa_d_mxwt(31 DOWNTO 0)), (vec_rsc_0_6_i_qa_d_mxwt(31
            DOWNTO 0)), (vec_rsc_0_7_i_qa_d_mxwt(31 DOWNTO 0)), (vec_rsc_1_0_i_qa_d_mxwt(31
            DOWNTO 0)), (vec_rsc_1_1_i_qa_d_mxwt(31 DOWNTO 0)), (vec_rsc_1_2_i_qa_d_mxwt(31
            DOWNTO 0)), (vec_rsc_1_3_i_qa_d_mxwt(31 DOWNTO 0)), (vec_rsc_1_4_i_qa_d_mxwt(31
            DOWNTO 0)), (vec_rsc_1_5_i_qa_d_mxwt(31 DOWNTO 0)), (vec_rsc_1_6_i_qa_d_mxwt(31
            DOWNTO 0)), (vec_rsc_1_7_i_qa_d_mxwt(31 DOWNTO 0)), STD_LOGIC_VECTOR'(
            VEC_LOOP_VEC_LOOP_nor_itm & VEC_LOOP_VEC_LOOP_and_nl & VEC_LOOP_VEC_LOOP_and_1_nl
            & VEC_LOOP_VEC_LOOP_and_2_itm & VEC_LOOP_VEC_LOOP_and_3_nl & VEC_LOOP_VEC_LOOP_and_4_itm
            & VEC_LOOP_VEC_LOOP_and_5_itm & VEC_LOOP_VEC_LOOP_and_6_itm & VEC_LOOP_VEC_LOOP_and_7_nl
            & VEC_LOOP_VEC_LOOP_and_8_itm & VEC_LOOP_VEC_LOOP_and_9_itm & VEC_LOOP_VEC_LOOP_and_10_itm
            & VEC_LOOP_VEC_LOOP_and_11_itm & VEC_LOOP_VEC_LOOP_and_12_itm & VEC_LOOP_VEC_LOOP_and_13_itm
            & VEC_LOOP_VEC_LOOP_and_14_itm));
        tmp_1_lpi_4_dfm <= MUX1HOT_v_32_16_2((vec_rsc_0_0_i_qa_d_mxwt(63 DOWNTO 32)),
            (vec_rsc_0_1_i_qa_d_mxwt(63 DOWNTO 32)), (vec_rsc_0_2_i_qa_d_mxwt(63
            DOWNTO 32)), (vec_rsc_0_3_i_qa_d_mxwt(63 DOWNTO 32)), (vec_rsc_0_4_i_qa_d_mxwt(63
            DOWNTO 32)), (vec_rsc_0_5_i_qa_d_mxwt(63 DOWNTO 32)), (vec_rsc_0_6_i_qa_d_mxwt(63
            DOWNTO 32)), (vec_rsc_0_7_i_qa_d_mxwt(63 DOWNTO 32)), (vec_rsc_1_0_i_qa_d_mxwt(63
            DOWNTO 32)), (vec_rsc_1_1_i_qa_d_mxwt(63 DOWNTO 32)), (vec_rsc_1_2_i_qa_d_mxwt(63
            DOWNTO 32)), (vec_rsc_1_3_i_qa_d_mxwt(63 DOWNTO 32)), (vec_rsc_1_4_i_qa_d_mxwt(63
            DOWNTO 32)), (vec_rsc_1_5_i_qa_d_mxwt(63 DOWNTO 32)), (vec_rsc_1_6_i_qa_d_mxwt(63
            DOWNTO 32)), (vec_rsc_1_7_i_qa_d_mxwt(63 DOWNTO 32)), STD_LOGIC_VECTOR'(
            VEC_LOOP_VEC_LOOP_nor_1_itm & VEC_LOOP_VEC_LOOP_and_15_nl & VEC_LOOP_VEC_LOOP_and_16_nl
            & VEC_LOOP_VEC_LOOP_and_17_itm & VEC_LOOP_VEC_LOOP_and_18_nl & VEC_LOOP_VEC_LOOP_and_19_itm
            & VEC_LOOP_VEC_LOOP_and_20_itm & VEC_LOOP_VEC_LOOP_and_21_itm & VEC_LOOP_VEC_LOOP_and_22_nl
            & VEC_LOOP_VEC_LOOP_and_23_itm & VEC_LOOP_VEC_LOOP_and_24_itm & VEC_LOOP_VEC_LOOP_and_25_itm
            & VEC_LOOP_VEC_LOOP_and_26_itm & VEC_LOOP_VEC_LOOP_and_27_itm & VEC_LOOP_VEC_LOOP_and_28_itm
            & VEC_LOOP_VEC_LOOP_and_29_itm));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_run_rsci_oswt_cse <= '0';
        reg_complete_rsci_oswt_cse <= '0';
        reg_vec_rsc_0_0_i_oswt_cse <= '0';
        reg_vec_rsc_0_0_i_oswt_1_cse <= '0';
        reg_vec_rsc_0_1_i_oswt_cse <= '0';
        reg_vec_rsc_0_1_i_oswt_1_cse <= '0';
        reg_vec_rsc_0_2_i_oswt_cse <= '0';
        reg_vec_rsc_0_2_i_oswt_1_cse <= '0';
        reg_vec_rsc_0_3_i_oswt_cse <= '0';
        reg_vec_rsc_0_3_i_oswt_1_cse <= '0';
        reg_vec_rsc_0_4_i_oswt_cse <= '0';
        reg_vec_rsc_0_4_i_oswt_1_cse <= '0';
        reg_vec_rsc_0_5_i_oswt_cse <= '0';
        reg_vec_rsc_0_5_i_oswt_1_cse <= '0';
        reg_vec_rsc_0_6_i_oswt_cse <= '0';
        reg_vec_rsc_0_6_i_oswt_1_cse <= '0';
        reg_vec_rsc_0_7_i_oswt_cse <= '0';
        reg_vec_rsc_0_7_i_oswt_1_cse <= '0';
        reg_vec_rsc_1_0_i_oswt_cse <= '0';
        reg_vec_rsc_1_0_i_oswt_1_cse <= '0';
        reg_vec_rsc_1_1_i_oswt_cse <= '0';
        reg_vec_rsc_1_1_i_oswt_1_cse <= '0';
        reg_vec_rsc_1_2_i_oswt_cse <= '0';
        reg_vec_rsc_1_2_i_oswt_1_cse <= '0';
        reg_vec_rsc_1_3_i_oswt_cse <= '0';
        reg_vec_rsc_1_3_i_oswt_1_cse <= '0';
        reg_vec_rsc_1_4_i_oswt_cse <= '0';
        reg_vec_rsc_1_4_i_oswt_1_cse <= '0';
        reg_vec_rsc_1_5_i_oswt_cse <= '0';
        reg_vec_rsc_1_5_i_oswt_1_cse <= '0';
        reg_vec_rsc_1_6_i_oswt_cse <= '0';
        reg_vec_rsc_1_6_i_oswt_1_cse <= '0';
        reg_vec_rsc_1_7_i_oswt_cse <= '0';
        reg_vec_rsc_1_7_i_oswt_1_cse <= '0';
        reg_twiddle_rsc_0_0_i_oswt_cse <= '0';
        reg_twiddle_rsc_0_1_i_oswt_cse <= '0';
        reg_twiddle_rsc_0_2_i_oswt_cse <= '0';
        reg_twiddle_rsc_0_3_i_oswt_cse <= '0';
        reg_twiddle_rsc_0_4_i_oswt_cse <= '0';
        reg_twiddle_rsc_0_5_i_oswt_cse <= '0';
        reg_twiddle_rsc_0_6_i_oswt_cse <= '0';
        reg_twiddle_rsc_0_7_i_oswt_cse <= '0';
        reg_twiddle_rsc_1_0_i_oswt_cse <= '0';
        reg_twiddle_rsc_1_1_i_oswt_cse <= '0';
        reg_twiddle_rsc_1_2_i_oswt_cse <= '0';
        reg_twiddle_rsc_1_3_i_oswt_cse <= '0';
        reg_twiddle_rsc_1_4_i_oswt_cse <= '0';
        reg_twiddle_rsc_1_5_i_oswt_cse <= '0';
        reg_twiddle_rsc_1_6_i_oswt_cse <= '0';
        reg_twiddle_rsc_1_7_i_oswt_cse <= '0';
        reg_vec_rsc_triosy_1_7_obj_iswt0_cse <= '0';
        reg_ensig_cgo_cse <= '0';
        reg_ensig_cgo_1_cse <= '0';
        VEC_LOOP_VEC_LOOP_nor_1_itm <= '0';
        VEC_LOOP_nor_10_itm <= '0';
        VEC_LOOP_nor_11_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_17_itm <= '0';
        VEC_LOOP_nor_13_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_19_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_20_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_21_itm <= '0';
        VEC_LOOP_nor_16_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_23_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_24_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_25_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_26_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_27_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_28_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_29_itm <= '0';
        VEC_LOOP_VEC_LOOP_nor_itm <= '0';
        VEC_LOOP_nor_itm <= '0';
        VEC_LOOP_nor_1_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_2_itm <= '0';
        VEC_LOOP_nor_3_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_4_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_5_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_6_itm <= '0';
        VEC_LOOP_nor_6_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_8_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_9_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_11_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_12_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_13_itm <= '0';
        VEC_LOOP_VEC_LOOP_and_14_itm <= '0';
      ELSIF ( complete_rsci_wen_comp = '1' ) THEN
        reg_run_rsci_oswt_cse <= fsm_output(0);
        reg_complete_rsci_oswt_cse <= (NOT STAGE_LOOP_acc_itm_4_1) AND (fsm_output(19));
        reg_vec_rsc_0_0_i_oswt_cse <= or_15_rmff;
        reg_vec_rsc_0_0_i_oswt_1_cse <= and_161_rmff;
        reg_vec_rsc_0_1_i_oswt_cse <= or_24_rmff;
        reg_vec_rsc_0_1_i_oswt_1_cse <= and_182_rmff;
        reg_vec_rsc_0_2_i_oswt_cse <= or_29_rmff;
        reg_vec_rsc_0_2_i_oswt_1_cse <= and_195_rmff;
        reg_vec_rsc_0_3_i_oswt_cse <= or_34_rmff;
        reg_vec_rsc_0_3_i_oswt_1_cse <= and_208_rmff;
        reg_vec_rsc_0_4_i_oswt_cse <= or_39_rmff;
        reg_vec_rsc_0_4_i_oswt_1_cse <= and_221_rmff;
        reg_vec_rsc_0_5_i_oswt_cse <= or_44_rmff;
        reg_vec_rsc_0_5_i_oswt_1_cse <= and_234_rmff;
        reg_vec_rsc_0_6_i_oswt_cse <= or_49_rmff;
        reg_vec_rsc_0_6_i_oswt_1_cse <= and_247_rmff;
        reg_vec_rsc_0_7_i_oswt_cse <= or_54_rmff;
        reg_vec_rsc_0_7_i_oswt_1_cse <= and_260_rmff;
        reg_vec_rsc_1_0_i_oswt_cse <= or_59_rmff;
        reg_vec_rsc_1_0_i_oswt_1_cse <= and_273_rmff;
        reg_vec_rsc_1_1_i_oswt_cse <= or_64_rmff;
        reg_vec_rsc_1_1_i_oswt_1_cse <= and_286_rmff;
        reg_vec_rsc_1_2_i_oswt_cse <= or_69_rmff;
        reg_vec_rsc_1_2_i_oswt_1_cse <= and_299_rmff;
        reg_vec_rsc_1_3_i_oswt_cse <= or_74_rmff;
        reg_vec_rsc_1_3_i_oswt_1_cse <= and_312_rmff;
        reg_vec_rsc_1_4_i_oswt_cse <= or_79_rmff;
        reg_vec_rsc_1_4_i_oswt_1_cse <= and_325_rmff;
        reg_vec_rsc_1_5_i_oswt_cse <= or_84_rmff;
        reg_vec_rsc_1_5_i_oswt_1_cse <= and_338_rmff;
        reg_vec_rsc_1_6_i_oswt_cse <= or_89_rmff;
        reg_vec_rsc_1_6_i_oswt_1_cse <= and_351_rmff;
        reg_vec_rsc_1_7_i_oswt_cse <= or_94_rmff;
        reg_vec_rsc_1_7_i_oswt_1_cse <= and_364_rmff;
        reg_twiddle_rsc_0_0_i_oswt_cse <= and_373_rmff;
        reg_twiddle_rsc_0_1_i_oswt_cse <= and_375_rmff;
        reg_twiddle_rsc_0_2_i_oswt_cse <= and_377_rmff;
        reg_twiddle_rsc_0_3_i_oswt_cse <= and_379_rmff;
        reg_twiddle_rsc_0_4_i_oswt_cse <= and_381_rmff;
        reg_twiddle_rsc_0_5_i_oswt_cse <= and_383_rmff;
        reg_twiddle_rsc_0_6_i_oswt_cse <= and_385_rmff;
        reg_twiddle_rsc_0_7_i_oswt_cse <= and_387_rmff;
        reg_twiddle_rsc_1_0_i_oswt_cse <= and_389_rmff;
        reg_twiddle_rsc_1_1_i_oswt_cse <= and_391_rmff;
        reg_twiddle_rsc_1_2_i_oswt_cse <= and_393_rmff;
        reg_twiddle_rsc_1_3_i_oswt_cse <= and_395_rmff;
        reg_twiddle_rsc_1_4_i_oswt_cse <= and_397_rmff;
        reg_twiddle_rsc_1_5_i_oswt_cse <= and_399_rmff;
        reg_twiddle_rsc_1_6_i_oswt_cse <= and_401_rmff;
        reg_twiddle_rsc_1_7_i_oswt_cse <= and_403_rmff;
        reg_vec_rsc_triosy_1_7_obj_iswt0_cse <= fsm_output(20);
        reg_ensig_cgo_cse <= or_116_rmff;
        reg_ensig_cgo_1_cse <= or_118_rmff;
        VEC_LOOP_VEC_LOOP_nor_1_itm <= NOT((VEC_LOOP_acc_10_tmp(9)) OR (VEC_LOOP_acc_10_tmp(2))
            OR (VEC_LOOP_acc_10_tmp(1)) OR (VEC_LOOP_acc_10_tmp(0)));
        VEC_LOOP_nor_10_itm <= NOT((VEC_LOOP_acc_10_tmp(9)) OR (VEC_LOOP_acc_10_tmp(2))
            OR (VEC_LOOP_acc_10_tmp(1)));
        VEC_LOOP_nor_11_itm <= NOT((VEC_LOOP_acc_10_tmp(9)) OR (VEC_LOOP_acc_10_tmp(2))
            OR (VEC_LOOP_acc_10_tmp(0)));
        VEC_LOOP_VEC_LOOP_and_17_itm <= CONV_SL_1_1(VEC_LOOP_acc_10_tmp(1 DOWNTO
            0)=STD_LOGIC_VECTOR'("11")) AND VEC_LOOP_nor_12_cse;
        VEC_LOOP_nor_13_itm <= NOT((VEC_LOOP_acc_10_tmp(9)) OR (VEC_LOOP_acc_10_tmp(1))
            OR (VEC_LOOP_acc_10_tmp(0)));
        VEC_LOOP_VEC_LOOP_and_19_itm <= (VEC_LOOP_acc_10_tmp(2)) AND (VEC_LOOP_acc_10_tmp(0))
            AND (NOT((VEC_LOOP_acc_10_tmp(9)) OR (VEC_LOOP_acc_10_tmp(1))));
        VEC_LOOP_VEC_LOOP_and_20_itm <= (VEC_LOOP_acc_10_tmp(2)) AND (VEC_LOOP_acc_10_tmp(1))
            AND (NOT((VEC_LOOP_acc_10_tmp(9)) OR (VEC_LOOP_acc_10_tmp(0))));
        VEC_LOOP_VEC_LOOP_and_21_itm <= (VEC_LOOP_acc_10_tmp(2)) AND (VEC_LOOP_acc_10_tmp(1))
            AND (VEC_LOOP_acc_10_tmp(0)) AND (NOT (VEC_LOOP_acc_10_tmp(9)));
        VEC_LOOP_nor_16_itm <= NOT(CONV_SL_1_1(VEC_LOOP_acc_10_tmp(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        VEC_LOOP_VEC_LOOP_and_23_itm <= (VEC_LOOP_acc_10_tmp(9)) AND (VEC_LOOP_acc_10_tmp(0))
            AND (NOT(CONV_SL_1_1(VEC_LOOP_acc_10_tmp(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))));
        VEC_LOOP_VEC_LOOP_and_24_itm <= (VEC_LOOP_acc_10_tmp(9)) AND (VEC_LOOP_acc_10_tmp(1))
            AND (NOT((VEC_LOOP_acc_10_tmp(2)) OR (VEC_LOOP_acc_10_tmp(0))));
        VEC_LOOP_VEC_LOOP_and_25_itm <= (VEC_LOOP_acc_10_tmp(9)) AND (VEC_LOOP_acc_10_tmp(1))
            AND (VEC_LOOP_acc_10_tmp(0)) AND (NOT (VEC_LOOP_acc_10_tmp(2)));
        VEC_LOOP_VEC_LOOP_and_26_itm <= (VEC_LOOP_acc_10_tmp(9)) AND (VEC_LOOP_acc_10_tmp(2))
            AND VEC_LOOP_nor_19_cse;
        VEC_LOOP_VEC_LOOP_and_27_itm <= (VEC_LOOP_acc_10_tmp(9)) AND (VEC_LOOP_acc_10_tmp(2))
            AND (VEC_LOOP_acc_10_tmp(0)) AND (NOT (VEC_LOOP_acc_10_tmp(1)));
        VEC_LOOP_VEC_LOOP_and_28_itm <= (VEC_LOOP_acc_10_tmp(9)) AND (VEC_LOOP_acc_10_tmp(2))
            AND (VEC_LOOP_acc_10_tmp(1)) AND (NOT (VEC_LOOP_acc_10_tmp(0)));
        VEC_LOOP_VEC_LOOP_and_29_itm <= (VEC_LOOP_acc_10_tmp(9)) AND (VEC_LOOP_acc_10_tmp(2))
            AND (VEC_LOOP_acc_10_tmp(1)) AND (VEC_LOOP_acc_10_tmp(0));
        VEC_LOOP_VEC_LOOP_nor_itm <= NOT((VEC_LOOP_acc_1_tmp(9)) OR (VEC_LOOP_acc_1_tmp(2))
            OR (VEC_LOOP_acc_1_tmp(1)) OR (VEC_LOOP_acc_1_tmp(0)));
        VEC_LOOP_nor_itm <= NOT((VEC_LOOP_acc_1_tmp(9)) OR (VEC_LOOP_acc_1_tmp(2))
            OR (VEC_LOOP_acc_1_tmp(1)));
        VEC_LOOP_nor_1_itm <= NOT((VEC_LOOP_acc_1_tmp(9)) OR (VEC_LOOP_acc_1_tmp(2))
            OR (VEC_LOOP_acc_1_tmp(0)));
        VEC_LOOP_VEC_LOOP_and_2_itm <= CONV_SL_1_1(VEC_LOOP_acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
            AND VEC_LOOP_nor_2_cse;
        VEC_LOOP_nor_3_itm <= NOT((VEC_LOOP_acc_1_tmp(9)) OR (VEC_LOOP_acc_1_tmp(1))
            OR (VEC_LOOP_acc_1_tmp(0)));
        VEC_LOOP_VEC_LOOP_and_4_itm <= (VEC_LOOP_acc_1_tmp(2)) AND (VEC_LOOP_acc_1_tmp(0))
            AND (NOT((VEC_LOOP_acc_1_tmp(9)) OR (VEC_LOOP_acc_1_tmp(1))));
        VEC_LOOP_VEC_LOOP_and_5_itm <= (VEC_LOOP_acc_1_tmp(2)) AND (VEC_LOOP_acc_1_tmp(1))
            AND (NOT((VEC_LOOP_acc_1_tmp(9)) OR (VEC_LOOP_acc_1_tmp(0))));
        VEC_LOOP_VEC_LOOP_and_6_itm <= (VEC_LOOP_acc_1_tmp(2)) AND (VEC_LOOP_acc_1_tmp(1))
            AND (VEC_LOOP_acc_1_tmp(0)) AND (NOT (VEC_LOOP_acc_1_tmp(9)));
        VEC_LOOP_nor_6_itm <= NOT(CONV_SL_1_1(VEC_LOOP_acc_1_tmp(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        VEC_LOOP_VEC_LOOP_and_8_itm <= (VEC_LOOP_acc_1_tmp(9)) AND (VEC_LOOP_acc_1_tmp(0))
            AND (NOT(CONV_SL_1_1(VEC_LOOP_acc_1_tmp(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))));
        VEC_LOOP_VEC_LOOP_and_9_itm <= (VEC_LOOP_acc_1_tmp(9)) AND (VEC_LOOP_acc_1_tmp(1))
            AND (NOT((VEC_LOOP_acc_1_tmp(2)) OR (VEC_LOOP_acc_1_tmp(0))));
        VEC_LOOP_VEC_LOOP_and_11_itm <= (VEC_LOOP_acc_1_tmp(9)) AND (VEC_LOOP_acc_1_tmp(2))
            AND VEC_LOOP_nor_9_cse;
        VEC_LOOP_VEC_LOOP_and_12_itm <= (VEC_LOOP_acc_1_tmp(9)) AND (VEC_LOOP_acc_1_tmp(2))
            AND (VEC_LOOP_acc_1_tmp(0)) AND (NOT (VEC_LOOP_acc_1_tmp(1)));
        VEC_LOOP_VEC_LOOP_and_13_itm <= (VEC_LOOP_acc_1_tmp(9)) AND (VEC_LOOP_acc_1_tmp(2))
            AND (VEC_LOOP_acc_1_tmp(1)) AND (NOT (VEC_LOOP_acc_1_tmp(0)));
        VEC_LOOP_VEC_LOOP_and_14_itm <= (VEC_LOOP_acc_1_tmp(9)) AND (VEC_LOOP_acc_1_tmp(2))
            AND (VEC_LOOP_acc_1_tmp(1)) AND (VEC_LOOP_acc_1_tmp(0));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (complete_rsci_wen_comp AND ((fsm_output(19)) OR (fsm_output(0)))) = '1'
          ) THEN
        STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'( "1010"), STAGE_LOOP_i_3_0_sva_2,
            fsm_output(19));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (complete_rsci_wen_comp AND (NOT and_dcpl_129)) = '1' ) THEN
        p_sva <= p_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (complete_rsci_wen_comp AND (NOT and_dcpl_131)) = '1' ) THEN
        STAGE_LOOP_lshift_psp_sva <= z_out;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (complete_rsci_wen_comp AND ((fsm_output(1)) OR (fsm_output(18)))) = '1'
          ) THEN
        COMP_LOOP_k_10_0_sva_9_0 <= MUX_v_10_2_2(STD_LOGIC_VECTOR'("0000000000"),
            (COMP_LOOP_k_10_0_sva_2(9 DOWNTO 0)), COMP_LOOP_k_not_1_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_twiddle_f_lshift_itm <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (((fsm_output(17)) OR (fsm_output(6)) OR (fsm_output(2)) OR (fsm_output(5)))
          AND complete_rsci_wen_comp) = '1' ) THEN
        COMP_LOOP_twiddle_f_lshift_itm <= MUX_v_10_2_2(STD_LOGIC_VECTOR'("0000000000"),
            COMP_LOOP_twiddle_f_mux1h_1_nl, COMP_LOOP_twiddle_f_not_7_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_twiddle_f_mul_cse_sva <= STD_LOGIC_VECTOR'( "0000000000");
        COMP_LOOP_twiddle_f_equal_tmp <= '0';
        COMP_LOOP_twiddle_f_equal_tmp_3 <= '0';
        COMP_LOOP_twiddle_f_equal_tmp_5 <= '0';
        COMP_LOOP_twiddle_f_equal_tmp_6 <= '0';
        COMP_LOOP_twiddle_f_equal_tmp_7 <= '0';
        COMP_LOOP_twiddle_f_equal_tmp_9 <= '0';
        COMP_LOOP_twiddle_f_equal_tmp_10 <= '0';
        COMP_LOOP_twiddle_f_equal_tmp_11 <= '0';
        COMP_LOOP_twiddle_f_equal_tmp_12 <= '0';
        COMP_LOOP_twiddle_f_equal_tmp_13 <= '0';
        COMP_LOOP_twiddle_f_equal_tmp_14 <= '0';
        COMP_LOOP_twiddle_f_equal_tmp_15 <= '0';
        COMP_LOOP_twiddle_f_nor_6_itm <= '0';
        COMP_LOOP_twiddle_f_nor_3_itm <= '0';
        COMP_LOOP_twiddle_f_nor_1_itm <= '0';
        COMP_LOOP_twiddle_f_nor_itm <= '0';
      ELSIF ( COMP_LOOP_twiddle_f_and_1_cse = '1' ) THEN
        COMP_LOOP_twiddle_f_mul_cse_sva <= COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0;
        COMP_LOOP_twiddle_f_equal_tmp <= NOT((COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(9))
            OR (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(2)) OR (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(1))
            OR (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(0)));
        COMP_LOOP_twiddle_f_equal_tmp_3 <= (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(1))
            AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(0)) AND (NOT((COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(9))
            OR (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(2))));
        COMP_LOOP_twiddle_f_equal_tmp_5 <= (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(2))
            AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(0)) AND (NOT((COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(9))
            OR (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(1))));
        COMP_LOOP_twiddle_f_equal_tmp_6 <= (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(2))
            AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(1)) AND (NOT((COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(9))
            OR (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(0))));
        COMP_LOOP_twiddle_f_equal_tmp_7 <= (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(2))
            AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(1)) AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(0))
            AND (NOT (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(9)));
        COMP_LOOP_twiddle_f_equal_tmp_9 <= (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(9))
            AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(0)) AND (NOT(CONV_SL_1_1(COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(2
            DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))));
        COMP_LOOP_twiddle_f_equal_tmp_10 <= (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(9))
            AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(1)) AND (NOT((COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(2))
            OR (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(0))));
        COMP_LOOP_twiddle_f_equal_tmp_11 <= (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(9))
            AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(1)) AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(0))
            AND (NOT (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(2)));
        COMP_LOOP_twiddle_f_equal_tmp_12 <= (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(9))
            AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(2)) AND (NOT(CONV_SL_1_1(COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(1
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))));
        COMP_LOOP_twiddle_f_equal_tmp_13 <= (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(9))
            AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(2)) AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(0))
            AND (NOT (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(1)));
        COMP_LOOP_twiddle_f_equal_tmp_14 <= (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(9))
            AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(2)) AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(1))
            AND (NOT (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(0)));
        COMP_LOOP_twiddle_f_equal_tmp_15 <= (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(9))
            AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(2)) AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(1))
            AND (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(0));
        COMP_LOOP_twiddle_f_nor_6_itm <= NOT(CONV_SL_1_1(COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_twiddle_f_nor_3_itm <= NOT((COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(9))
            OR (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(1)) OR (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(0)));
        COMP_LOOP_twiddle_f_nor_1_itm <= NOT((COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(9))
            OR (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(2)) OR (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(0)));
        COMP_LOOP_twiddle_f_nor_itm <= NOT((COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(9))
            OR (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(2)) OR (COMP_LOOP_twiddle_f_mul_cse_sva_mx0w0(1)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_twiddle_help_and_16_cse = '1' ) THEN
        tmp_3_lpi_3_dfm <= MUX1HOT_v_32_16_2(twiddle_h_rsc_0_0_i_qb_d_mxwt, twiddle_h_rsc_0_1_i_qb_d_mxwt,
            twiddle_h_rsc_0_2_i_qb_d_mxwt, twiddle_h_rsc_0_3_i_qb_d_mxwt, twiddle_h_rsc_0_4_i_qb_d_mxwt,
            twiddle_h_rsc_0_5_i_qb_d_mxwt, twiddle_h_rsc_0_6_i_qb_d_mxwt, twiddle_h_rsc_0_7_i_qb_d_mxwt,
            twiddle_h_rsc_1_0_i_qb_d_mxwt, twiddle_h_rsc_1_1_i_qb_d_mxwt, twiddle_h_rsc_1_2_i_qb_d_mxwt,
            twiddle_h_rsc_1_3_i_qb_d_mxwt, twiddle_h_rsc_1_4_i_qb_d_mxwt, twiddle_h_rsc_1_5_i_qb_d_mxwt,
            twiddle_h_rsc_1_6_i_qb_d_mxwt, twiddle_h_rsc_1_7_i_qb_d_mxwt, STD_LOGIC_VECTOR'(
            COMP_LOOP_twiddle_help_and_cse & COMP_LOOP_twiddle_help_and_1_cse & COMP_LOOP_twiddle_help_and_2_cse
            & COMP_LOOP_twiddle_help_and_3_cse & COMP_LOOP_twiddle_help_and_4_cse
            & COMP_LOOP_twiddle_help_and_5_cse & COMP_LOOP_twiddle_help_and_6_cse
            & COMP_LOOP_twiddle_help_and_7_cse & COMP_LOOP_twiddle_help_and_8_cse
            & COMP_LOOP_twiddle_help_and_9_cse & COMP_LOOP_twiddle_help_and_10_cse
            & COMP_LOOP_twiddle_help_and_11_cse & COMP_LOOP_twiddle_help_and_12_cse
            & COMP_LOOP_twiddle_help_and_13_cse & COMP_LOOP_twiddle_help_and_14_cse
            & COMP_LOOP_twiddle_help_and_15_cse));
        tmp_2_lpi_3_dfm <= MUX1HOT_v_32_16_2(twiddle_rsc_0_0_i_qb_d_mxwt, twiddle_rsc_0_1_i_qb_d_mxwt,
            twiddle_rsc_0_2_i_qb_d_mxwt, twiddle_rsc_0_3_i_qb_d_mxwt, twiddle_rsc_0_4_i_qb_d_mxwt,
            twiddle_rsc_0_5_i_qb_d_mxwt, twiddle_rsc_0_6_i_qb_d_mxwt, twiddle_rsc_0_7_i_qb_d_mxwt,
            twiddle_rsc_1_0_i_qb_d_mxwt, twiddle_rsc_1_1_i_qb_d_mxwt, twiddle_rsc_1_2_i_qb_d_mxwt,
            twiddle_rsc_1_3_i_qb_d_mxwt, twiddle_rsc_1_4_i_qb_d_mxwt, twiddle_rsc_1_5_i_qb_d_mxwt,
            twiddle_rsc_1_6_i_qb_d_mxwt, twiddle_rsc_1_7_i_qb_d_mxwt, STD_LOGIC_VECTOR'(
            COMP_LOOP_twiddle_help_and_cse & COMP_LOOP_twiddle_help_and_1_cse & COMP_LOOP_twiddle_help_and_2_cse
            & COMP_LOOP_twiddle_help_and_3_cse & COMP_LOOP_twiddle_help_and_4_cse
            & COMP_LOOP_twiddle_help_and_5_cse & COMP_LOOP_twiddle_help_and_6_cse
            & COMP_LOOP_twiddle_help_and_7_cse & COMP_LOOP_twiddle_help_and_8_cse
            & COMP_LOOP_twiddle_help_and_9_cse & COMP_LOOP_twiddle_help_and_10_cse
            & COMP_LOOP_twiddle_help_and_11_cse & COMP_LOOP_twiddle_help_and_12_cse
            & COMP_LOOP_twiddle_help_and_13_cse & COMP_LOOP_twiddle_help_and_14_cse
            & COMP_LOOP_twiddle_help_and_15_cse));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        VEC_LOOP_acc_10_cse_sva <= STD_LOGIC_VECTOR'( "0000000000");
        VEC_LOOP_j_10_0_sva_1 <= STD_LOGIC_VECTOR'( "00000000000");
      ELSIF ( VEC_LOOP_and_cse = '1' ) THEN
        VEC_LOOP_acc_10_cse_sva <= VEC_LOOP_acc_10_tmp;
        VEC_LOOP_j_10_0_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_twiddle_f_lshift_itm),
            10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva), 11));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        VEC_LOOP_VEC_LOOP_and_10_itm <= '0';
      ELSIF ( (complete_rsci_wen_comp AND ((fsm_output(20)) OR (fsm_output(6))))
          = '1' ) THEN
        VEC_LOOP_VEC_LOOP_and_10_itm <= MUX_s_1_2_2(VEC_LOOP_VEC_LOOP_and_10_nl,
            run_rsci_ivld_mxwt, fsm_output(20));
      END IF;
    END IF;
  END PROCESS;
  VEC_LOOP_VEC_LOOP_and_nl <= (COMP_LOOP_twiddle_f_lshift_itm(0)) AND VEC_LOOP_nor_itm;
  VEC_LOOP_VEC_LOOP_and_1_nl <= (COMP_LOOP_twiddle_f_lshift_itm(1)) AND VEC_LOOP_nor_1_itm;
  VEC_LOOP_VEC_LOOP_and_3_nl <= (COMP_LOOP_twiddle_f_lshift_itm(2)) AND VEC_LOOP_nor_3_itm;
  VEC_LOOP_VEC_LOOP_and_7_nl <= (COMP_LOOP_twiddle_f_lshift_itm(9)) AND VEC_LOOP_nor_6_itm;
  VEC_LOOP_VEC_LOOP_and_15_nl <= (VEC_LOOP_acc_10_cse_sva(0)) AND VEC_LOOP_nor_10_itm;
  VEC_LOOP_VEC_LOOP_and_16_nl <= (VEC_LOOP_acc_10_cse_sva(1)) AND VEC_LOOP_nor_11_itm;
  VEC_LOOP_VEC_LOOP_and_18_nl <= (VEC_LOOP_acc_10_cse_sva(2)) AND VEC_LOOP_nor_13_itm;
  VEC_LOOP_VEC_LOOP_and_22_nl <= (VEC_LOOP_acc_10_cse_sva(9)) AND VEC_LOOP_nor_16_itm;
  COMP_LOOP_k_not_1_nl <= NOT (fsm_output(1));
  COMP_LOOP_twiddle_f_mux1h_1_nl <= MUX1HOT_v_10_3_2((z_out(9 DOWNTO 0)), VEC_LOOP_acc_1_tmp,
      (VEC_LOOP_j_10_0_sva_1(9 DOWNTO 0)), STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6))
      & (fsm_output(17))));
  COMP_LOOP_twiddle_f_not_7_nl <= NOT (fsm_output(5));
  VEC_LOOP_VEC_LOOP_and_10_nl <= (VEC_LOOP_acc_1_tmp(9)) AND (VEC_LOOP_acc_1_tmp(1))
      AND (VEC_LOOP_acc_1_tmp(0)) AND (NOT (VEC_LOOP_acc_1_tmp(2)));
END v5;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_precomp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_sync_in_wait_pkg_v1.ALL;
USE work.ccs_sync_out_wait_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_precomp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    run_rsc_rdy : OUT STD_LOGIC;
    run_rsc_vld : IN STD_LOGIC;
    vec_rsc_0_0_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_0_wea : OUT STD_LOGIC;
    vec_rsc_0_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_0_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_0_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_0_web : OUT STD_LOGIC;
    vec_rsc_0_0_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_0_1_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_1_wea : OUT STD_LOGIC;
    vec_rsc_0_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_1_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_1_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_1_web : OUT STD_LOGIC;
    vec_rsc_0_1_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_0_2_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_2_wea : OUT STD_LOGIC;
    vec_rsc_0_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_2_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_2_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_2_web : OUT STD_LOGIC;
    vec_rsc_0_2_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_0_3_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_3_wea : OUT STD_LOGIC;
    vec_rsc_0_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_3_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_3_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_3_web : OUT STD_LOGIC;
    vec_rsc_0_3_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_0_4_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_4_wea : OUT STD_LOGIC;
    vec_rsc_0_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_4_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_4_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_4_web : OUT STD_LOGIC;
    vec_rsc_0_4_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_0_5_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_5_wea : OUT STD_LOGIC;
    vec_rsc_0_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_5_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_5_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_5_web : OUT STD_LOGIC;
    vec_rsc_0_5_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_0_6_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_6_wea : OUT STD_LOGIC;
    vec_rsc_0_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_6_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_6_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_6_web : OUT STD_LOGIC;
    vec_rsc_0_6_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_0_7_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_7_wea : OUT STD_LOGIC;
    vec_rsc_0_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_7_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_7_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_0_7_web : OUT STD_LOGIC;
    vec_rsc_0_7_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    vec_rsc_1_0_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_1_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_0_wea : OUT STD_LOGIC;
    vec_rsc_1_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_0_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_1_0_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_0_web : OUT STD_LOGIC;
    vec_rsc_1_0_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    vec_rsc_1_1_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_1_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_1_wea : OUT STD_LOGIC;
    vec_rsc_1_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_1_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_1_1_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_1_web : OUT STD_LOGIC;
    vec_rsc_1_1_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_triosy_1_1_lz : OUT STD_LOGIC;
    vec_rsc_1_2_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_1_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_2_wea : OUT STD_LOGIC;
    vec_rsc_1_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_2_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_1_2_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_2_web : OUT STD_LOGIC;
    vec_rsc_1_2_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_triosy_1_2_lz : OUT STD_LOGIC;
    vec_rsc_1_3_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_1_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_3_wea : OUT STD_LOGIC;
    vec_rsc_1_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_3_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_1_3_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_3_web : OUT STD_LOGIC;
    vec_rsc_1_3_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_triosy_1_3_lz : OUT STD_LOGIC;
    vec_rsc_1_4_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_1_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_4_wea : OUT STD_LOGIC;
    vec_rsc_1_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_4_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_1_4_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_4_web : OUT STD_LOGIC;
    vec_rsc_1_4_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_triosy_1_4_lz : OUT STD_LOGIC;
    vec_rsc_1_5_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_1_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_5_wea : OUT STD_LOGIC;
    vec_rsc_1_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_5_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_1_5_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_5_web : OUT STD_LOGIC;
    vec_rsc_1_5_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_triosy_1_5_lz : OUT STD_LOGIC;
    vec_rsc_1_6_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_1_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_6_wea : OUT STD_LOGIC;
    vec_rsc_1_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_6_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_1_6_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_6_web : OUT STD_LOGIC;
    vec_rsc_1_6_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_triosy_1_6_lz : OUT STD_LOGIC;
    vec_rsc_1_7_adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_1_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_7_wea : OUT STD_LOGIC;
    vec_rsc_1_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_7_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_1_7_db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_1_7_web : OUT STD_LOGIC;
    vec_rsc_1_7_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    vec_rsc_triosy_1_7_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsc_0_0_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_0_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_rsc_0_1_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_1_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_rsc_0_2_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_2_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_rsc_0_3_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_3_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_rsc_0_4_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_4_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_rsc_0_5_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_5_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_rsc_0_6_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_6_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_rsc_0_7_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_7_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_rsc_1_0_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_1_0_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    twiddle_rsc_1_1_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_1_1_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_1_1_lz : OUT STD_LOGIC;
    twiddle_rsc_1_2_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_1_2_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_1_2_lz : OUT STD_LOGIC;
    twiddle_rsc_1_3_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_1_3_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_1_3_lz : OUT STD_LOGIC;
    twiddle_rsc_1_4_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_1_4_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_1_4_lz : OUT STD_LOGIC;
    twiddle_rsc_1_5_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_1_5_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_1_5_lz : OUT STD_LOGIC;
    twiddle_rsc_1_6_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_1_6_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_1_6_lz : OUT STD_LOGIC;
    twiddle_rsc_1_7_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_1_7_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_1_7_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_0_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_1_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_2_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_3_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_4_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_5_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_6_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_7_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_h_rsc_1_0_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_1_0_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    twiddle_h_rsc_1_1_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_1_1_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_1_1_lz : OUT STD_LOGIC;
    twiddle_h_rsc_1_2_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_1_2_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_1_2_lz : OUT STD_LOGIC;
    twiddle_h_rsc_1_3_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_1_3_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_1_3_lz : OUT STD_LOGIC;
    twiddle_h_rsc_1_4_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_1_4_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_1_4_lz : OUT STD_LOGIC;
    twiddle_h_rsc_1_5_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_1_5_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_1_5_lz : OUT STD_LOGIC;
    twiddle_h_rsc_1_6_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_1_6_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_1_6_lz : OUT STD_LOGIC;
    twiddle_h_rsc_1_7_adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_1_7_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_1_7_lz : OUT STD_LOGIC;
    complete_rsc_rdy : IN STD_LOGIC;
    complete_rsc_vld : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_precomp;

ARCHITECTURE v5 OF inPlaceNTT_DIF_precomp IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_0_i_adra_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_1_i_adra_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_2_i_adra_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_3_i_adra_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_4_i_adra_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_5_i_adra_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_6_i_adra_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_7_i_adra_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL twiddle_rsc_0_0_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_1_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_2_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_3_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_4_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_5_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_6_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_7_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_1_0_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_1_1_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_1_2_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_1_3_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_1_4_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_1_5_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_1_6_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_1_7_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_0_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_1_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_2_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_3_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_4_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_5_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_6_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_7_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_0_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_1_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_2_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_3_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_4_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_5_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_6_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsc_1_7_i_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_0_i_adrb_d_iff : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_22_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_adra_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_23_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_1_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_adra_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_24_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_2_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_adra_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_25_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_3_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_adra_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_26_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_4_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_adra_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_27_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_5_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_adra_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_28_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_6_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_adra_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_29_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_7_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_adra_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_30_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL vec_rsc_1_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_adra_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_31_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL vec_rsc_1_1_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_adra_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_32_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL vec_rsc_1_2_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_adra_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_33_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL vec_rsc_1_3_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_adra_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_34_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL vec_rsc_1_4_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_adra_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_35_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL vec_rsc_1_5_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_adra_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_36_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL vec_rsc_1_6_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_adra_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_37_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL vec_rsc_1_7_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_adra : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_adra_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_da_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_38_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_39_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_1_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_40_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_2_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_41_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_3_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_42_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_4_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_43_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_5_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_44_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_6_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_45_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_7_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_46_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_1_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_0_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_1_0_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_1_0_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_47_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_1_1_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_1_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_1_1_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_1_1_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_48_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_1_2_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_2_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_1_2_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_1_2_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_49_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_1_3_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_3_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_1_3_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_1_3_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_50_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_1_4_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_4_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_1_4_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_1_4_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_51_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_1_5_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_5_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_1_5_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_1_5_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_52_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_1_6_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_6_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_1_6_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_1_6_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_53_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_1_7_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_1_7_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_1_7_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_1_7_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_54_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_55_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_1_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_56_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_2_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_57_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_3_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_58_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_4_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_59_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_5_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_60_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_6_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_61_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_0_7_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_62_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_1_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_0_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_0_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_0_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_63_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_1_1_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_1_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_1_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_1_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_64_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_1_2_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_2_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_2_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_2_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_65_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_1_3_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_3_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_3_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_3_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_66_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_1_4_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_4_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_4_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_4_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_67_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_1_5_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_5_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_5_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_5_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_68_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_1_6_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_6_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_6_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_6_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_69_6_32_64_64_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsc_1_7_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_7_i_adrb : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_7_i_adrb_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_1_7_i_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_precomp_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      run_rsc_rdy : OUT STD_LOGIC;
      run_rsc_vld : IN STD_LOGIC;
      vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      vec_rsc_triosy_1_0_lz : OUT STD_LOGIC;
      vec_rsc_triosy_1_1_lz : OUT STD_LOGIC;
      vec_rsc_triosy_1_2_lz : OUT STD_LOGIC;
      vec_rsc_triosy_1_3_lz : OUT STD_LOGIC;
      vec_rsc_triosy_1_4_lz : OUT STD_LOGIC;
      vec_rsc_triosy_1_5_lz : OUT STD_LOGIC;
      vec_rsc_triosy_1_6_lz : OUT STD_LOGIC;
      vec_rsc_triosy_1_7_lz : OUT STD_LOGIC;
      p_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      p_rsc_triosy_lz : OUT STD_LOGIC;
      r_rsc_triosy_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_1_0_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_1_1_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_1_2_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_1_3_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_1_4_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_1_5_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_1_6_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_1_7_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_1_0_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_1_1_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_1_2_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_1_3_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_1_4_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_1_5_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_1_6_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_1_7_lz : OUT STD_LOGIC;
      complete_rsc_rdy : IN STD_LOGIC;
      complete_rsc_vld : OUT STD_LOGIC;
      vec_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      vec_rsc_0_0_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_1_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      vec_rsc_0_1_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_1_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_2_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      vec_rsc_0_2_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_2_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_3_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      vec_rsc_0_3_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_3_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_4_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      vec_rsc_0_4_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_4_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_5_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      vec_rsc_0_5_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_5_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_6_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      vec_rsc_0_6_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_6_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_7_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      vec_rsc_0_7_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_7_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_0_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      vec_rsc_1_0_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_1_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      vec_rsc_1_1_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_1_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_2_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      vec_rsc_1_2_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_2_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_3_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      vec_rsc_1_3_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_3_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_4_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      vec_rsc_1_4_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_4_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_5_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      vec_rsc_1_5_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_5_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_6_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      vec_rsc_1_6_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_6_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_7_i_adra_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      vec_rsc_1_7_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      vec_rsc_1_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_1_7_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      twiddle_rsc_0_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_1_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_1_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_1_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_1_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_1_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_1_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_1_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_1_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsc_1_0_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsc_1_1_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsc_1_2_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsc_1_3_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsc_1_4_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsc_1_5_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsc_1_6_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsc_1_7_i_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_0_i_adrb_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_p_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_adra_d : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_da_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_qa_d : STD_LOGIC_VECTOR (63
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_adra_d : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_da_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_qa_d : STD_LOGIC_VECTOR (63
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_adra_d : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_da_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_qa_d : STD_LOGIC_VECTOR (63
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_adra_d : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_da_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_qa_d : STD_LOGIC_VECTOR (63
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_adra_d : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_da_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_qa_d : STD_LOGIC_VECTOR (63
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_adra_d : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_da_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_qa_d : STD_LOGIC_VECTOR (63
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_adra_d : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_da_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_qa_d : STD_LOGIC_VECTOR (63
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_adra_d : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_da_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_qa_d : STD_LOGIC_VECTOR (63
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_wea_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d
      : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_0_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_1_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_2_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_3_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_4_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_5_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_6_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_7_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_0_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_1_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_2_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_3_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_4_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_5_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_6_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_7_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_0_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_1_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_2_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_3_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_4_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_5_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_6_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_7_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_0_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_1_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_2_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_3_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_4_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_5_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_6_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_7_i_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_0_i_adrb_d_pff : STD_LOGIC_VECTOR
      (5 DOWNTO 0);

BEGIN
  vec_rsc_0_0_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_22_6_32_64_64_32_1_gen
    PORT MAP(
      qb => vec_rsc_0_0_i_qb,
      web => vec_rsc_0_0_web,
      db => vec_rsc_0_0_i_db,
      adrb => vec_rsc_0_0_i_adrb,
      qa => vec_rsc_0_0_i_qa,
      wea => vec_rsc_0_0_wea,
      da => vec_rsc_0_0_i_da,
      adra => vec_rsc_0_0_i_adra,
      adra_d => vec_rsc_0_0_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => vec_rsc_0_0_i_da_d_1,
      qa_d => vec_rsc_0_0_i_qa_d_1,
      wea_d => vec_rsc_0_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  vec_rsc_0_0_i_qb <= vec_rsc_0_0_qb;
  vec_rsc_0_0_db <= vec_rsc_0_0_i_db;
  vec_rsc_0_0_adrb <= vec_rsc_0_0_i_adrb;
  vec_rsc_0_0_i_qa <= vec_rsc_0_0_qa;
  vec_rsc_0_0_da <= vec_rsc_0_0_i_da;
  vec_rsc_0_0_adra <= vec_rsc_0_0_i_adra;
  vec_rsc_0_0_i_adra_d_1 <= vec_rsc_0_0_i_adra_d;
  vec_rsc_0_0_i_da_d_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000")
      & vec_rsc_0_0_i_da_d;
  vec_rsc_0_0_i_qa_d <= vec_rsc_0_0_i_qa_d_1;
  vec_rsc_0_0_i_wea_d_1 <= vec_rsc_0_0_i_wea_d;
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  vec_rsc_0_1_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_23_6_32_64_64_32_1_gen
    PORT MAP(
      qb => vec_rsc_0_1_i_qb,
      web => vec_rsc_0_1_web,
      db => vec_rsc_0_1_i_db,
      adrb => vec_rsc_0_1_i_adrb,
      qa => vec_rsc_0_1_i_qa,
      wea => vec_rsc_0_1_wea,
      da => vec_rsc_0_1_i_da,
      adra => vec_rsc_0_1_i_adra,
      adra_d => vec_rsc_0_1_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => vec_rsc_0_1_i_da_d_1,
      qa_d => vec_rsc_0_1_i_qa_d_1,
      wea_d => vec_rsc_0_1_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  vec_rsc_0_1_i_qb <= vec_rsc_0_1_qb;
  vec_rsc_0_1_db <= vec_rsc_0_1_i_db;
  vec_rsc_0_1_adrb <= vec_rsc_0_1_i_adrb;
  vec_rsc_0_1_i_qa <= vec_rsc_0_1_qa;
  vec_rsc_0_1_da <= vec_rsc_0_1_i_da;
  vec_rsc_0_1_adra <= vec_rsc_0_1_i_adra;
  vec_rsc_0_1_i_adra_d_1 <= vec_rsc_0_1_i_adra_d;
  vec_rsc_0_1_i_da_d_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000")
      & vec_rsc_0_1_i_da_d;
  vec_rsc_0_1_i_qa_d <= vec_rsc_0_1_i_qa_d_1;
  vec_rsc_0_1_i_wea_d_1 <= vec_rsc_0_1_i_wea_d;
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  vec_rsc_0_2_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_24_6_32_64_64_32_1_gen
    PORT MAP(
      qb => vec_rsc_0_2_i_qb,
      web => vec_rsc_0_2_web,
      db => vec_rsc_0_2_i_db,
      adrb => vec_rsc_0_2_i_adrb,
      qa => vec_rsc_0_2_i_qa,
      wea => vec_rsc_0_2_wea,
      da => vec_rsc_0_2_i_da,
      adra => vec_rsc_0_2_i_adra,
      adra_d => vec_rsc_0_2_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => vec_rsc_0_2_i_da_d_1,
      qa_d => vec_rsc_0_2_i_qa_d_1,
      wea_d => vec_rsc_0_2_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  vec_rsc_0_2_i_qb <= vec_rsc_0_2_qb;
  vec_rsc_0_2_db <= vec_rsc_0_2_i_db;
  vec_rsc_0_2_adrb <= vec_rsc_0_2_i_adrb;
  vec_rsc_0_2_i_qa <= vec_rsc_0_2_qa;
  vec_rsc_0_2_da <= vec_rsc_0_2_i_da;
  vec_rsc_0_2_adra <= vec_rsc_0_2_i_adra;
  vec_rsc_0_2_i_adra_d_1 <= vec_rsc_0_2_i_adra_d;
  vec_rsc_0_2_i_da_d_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000")
      & vec_rsc_0_2_i_da_d;
  vec_rsc_0_2_i_qa_d <= vec_rsc_0_2_i_qa_d_1;
  vec_rsc_0_2_i_wea_d_1 <= vec_rsc_0_2_i_wea_d;
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  vec_rsc_0_3_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_25_6_32_64_64_32_1_gen
    PORT MAP(
      qb => vec_rsc_0_3_i_qb,
      web => vec_rsc_0_3_web,
      db => vec_rsc_0_3_i_db,
      adrb => vec_rsc_0_3_i_adrb,
      qa => vec_rsc_0_3_i_qa,
      wea => vec_rsc_0_3_wea,
      da => vec_rsc_0_3_i_da,
      adra => vec_rsc_0_3_i_adra,
      adra_d => vec_rsc_0_3_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => vec_rsc_0_3_i_da_d_1,
      qa_d => vec_rsc_0_3_i_qa_d_1,
      wea_d => vec_rsc_0_3_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  vec_rsc_0_3_i_qb <= vec_rsc_0_3_qb;
  vec_rsc_0_3_db <= vec_rsc_0_3_i_db;
  vec_rsc_0_3_adrb <= vec_rsc_0_3_i_adrb;
  vec_rsc_0_3_i_qa <= vec_rsc_0_3_qa;
  vec_rsc_0_3_da <= vec_rsc_0_3_i_da;
  vec_rsc_0_3_adra <= vec_rsc_0_3_i_adra;
  vec_rsc_0_3_i_adra_d_1 <= vec_rsc_0_3_i_adra_d;
  vec_rsc_0_3_i_da_d_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000")
      & vec_rsc_0_3_i_da_d;
  vec_rsc_0_3_i_qa_d <= vec_rsc_0_3_i_qa_d_1;
  vec_rsc_0_3_i_wea_d_1 <= vec_rsc_0_3_i_wea_d;
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  vec_rsc_0_4_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_26_6_32_64_64_32_1_gen
    PORT MAP(
      qb => vec_rsc_0_4_i_qb,
      web => vec_rsc_0_4_web,
      db => vec_rsc_0_4_i_db,
      adrb => vec_rsc_0_4_i_adrb,
      qa => vec_rsc_0_4_i_qa,
      wea => vec_rsc_0_4_wea,
      da => vec_rsc_0_4_i_da,
      adra => vec_rsc_0_4_i_adra,
      adra_d => vec_rsc_0_4_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => vec_rsc_0_4_i_da_d_1,
      qa_d => vec_rsc_0_4_i_qa_d_1,
      wea_d => vec_rsc_0_4_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  vec_rsc_0_4_i_qb <= vec_rsc_0_4_qb;
  vec_rsc_0_4_db <= vec_rsc_0_4_i_db;
  vec_rsc_0_4_adrb <= vec_rsc_0_4_i_adrb;
  vec_rsc_0_4_i_qa <= vec_rsc_0_4_qa;
  vec_rsc_0_4_da <= vec_rsc_0_4_i_da;
  vec_rsc_0_4_adra <= vec_rsc_0_4_i_adra;
  vec_rsc_0_4_i_adra_d_1 <= vec_rsc_0_4_i_adra_d;
  vec_rsc_0_4_i_da_d_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000")
      & vec_rsc_0_4_i_da_d;
  vec_rsc_0_4_i_qa_d <= vec_rsc_0_4_i_qa_d_1;
  vec_rsc_0_4_i_wea_d_1 <= vec_rsc_0_4_i_wea_d;
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  vec_rsc_0_5_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_27_6_32_64_64_32_1_gen
    PORT MAP(
      qb => vec_rsc_0_5_i_qb,
      web => vec_rsc_0_5_web,
      db => vec_rsc_0_5_i_db,
      adrb => vec_rsc_0_5_i_adrb,
      qa => vec_rsc_0_5_i_qa,
      wea => vec_rsc_0_5_wea,
      da => vec_rsc_0_5_i_da,
      adra => vec_rsc_0_5_i_adra,
      adra_d => vec_rsc_0_5_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => vec_rsc_0_5_i_da_d_1,
      qa_d => vec_rsc_0_5_i_qa_d_1,
      wea_d => vec_rsc_0_5_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  vec_rsc_0_5_i_qb <= vec_rsc_0_5_qb;
  vec_rsc_0_5_db <= vec_rsc_0_5_i_db;
  vec_rsc_0_5_adrb <= vec_rsc_0_5_i_adrb;
  vec_rsc_0_5_i_qa <= vec_rsc_0_5_qa;
  vec_rsc_0_5_da <= vec_rsc_0_5_i_da;
  vec_rsc_0_5_adra <= vec_rsc_0_5_i_adra;
  vec_rsc_0_5_i_adra_d_1 <= vec_rsc_0_5_i_adra_d;
  vec_rsc_0_5_i_da_d_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000")
      & vec_rsc_0_5_i_da_d;
  vec_rsc_0_5_i_qa_d <= vec_rsc_0_5_i_qa_d_1;
  vec_rsc_0_5_i_wea_d_1 <= vec_rsc_0_5_i_wea_d;
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  vec_rsc_0_6_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_28_6_32_64_64_32_1_gen
    PORT MAP(
      qb => vec_rsc_0_6_i_qb,
      web => vec_rsc_0_6_web,
      db => vec_rsc_0_6_i_db,
      adrb => vec_rsc_0_6_i_adrb,
      qa => vec_rsc_0_6_i_qa,
      wea => vec_rsc_0_6_wea,
      da => vec_rsc_0_6_i_da,
      adra => vec_rsc_0_6_i_adra,
      adra_d => vec_rsc_0_6_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => vec_rsc_0_6_i_da_d_1,
      qa_d => vec_rsc_0_6_i_qa_d_1,
      wea_d => vec_rsc_0_6_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  vec_rsc_0_6_i_qb <= vec_rsc_0_6_qb;
  vec_rsc_0_6_db <= vec_rsc_0_6_i_db;
  vec_rsc_0_6_adrb <= vec_rsc_0_6_i_adrb;
  vec_rsc_0_6_i_qa <= vec_rsc_0_6_qa;
  vec_rsc_0_6_da <= vec_rsc_0_6_i_da;
  vec_rsc_0_6_adra <= vec_rsc_0_6_i_adra;
  vec_rsc_0_6_i_adra_d_1 <= vec_rsc_0_6_i_adra_d;
  vec_rsc_0_6_i_da_d_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000")
      & vec_rsc_0_6_i_da_d;
  vec_rsc_0_6_i_qa_d <= vec_rsc_0_6_i_qa_d_1;
  vec_rsc_0_6_i_wea_d_1 <= vec_rsc_0_6_i_wea_d;
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  vec_rsc_0_7_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_29_6_32_64_64_32_1_gen
    PORT MAP(
      qb => vec_rsc_0_7_i_qb,
      web => vec_rsc_0_7_web,
      db => vec_rsc_0_7_i_db,
      adrb => vec_rsc_0_7_i_adrb,
      qa => vec_rsc_0_7_i_qa,
      wea => vec_rsc_0_7_wea,
      da => vec_rsc_0_7_i_da,
      adra => vec_rsc_0_7_i_adra,
      adra_d => vec_rsc_0_7_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => vec_rsc_0_7_i_da_d_1,
      qa_d => vec_rsc_0_7_i_qa_d_1,
      wea_d => vec_rsc_0_7_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  vec_rsc_0_7_i_qb <= vec_rsc_0_7_qb;
  vec_rsc_0_7_db <= vec_rsc_0_7_i_db;
  vec_rsc_0_7_adrb <= vec_rsc_0_7_i_adrb;
  vec_rsc_0_7_i_qa <= vec_rsc_0_7_qa;
  vec_rsc_0_7_da <= vec_rsc_0_7_i_da;
  vec_rsc_0_7_adra <= vec_rsc_0_7_i_adra;
  vec_rsc_0_7_i_adra_d_1 <= vec_rsc_0_7_i_adra_d;
  vec_rsc_0_7_i_da_d_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000")
      & vec_rsc_0_7_i_da_d;
  vec_rsc_0_7_i_qa_d <= vec_rsc_0_7_i_qa_d_1;
  vec_rsc_0_7_i_wea_d_1 <= vec_rsc_0_7_i_wea_d;
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  vec_rsc_1_0_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_30_6_32_64_64_32_1_gen
    PORT MAP(
      qb => vec_rsc_1_0_i_qb,
      web => vec_rsc_1_0_web,
      db => vec_rsc_1_0_i_db,
      adrb => vec_rsc_1_0_i_adrb,
      qa => vec_rsc_1_0_i_qa,
      wea => vec_rsc_1_0_wea,
      da => vec_rsc_1_0_i_da,
      adra => vec_rsc_1_0_i_adra,
      adra_d => vec_rsc_1_0_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => vec_rsc_1_0_i_da_d_1,
      qa_d => vec_rsc_1_0_i_qa_d_1,
      wea_d => vec_rsc_1_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  vec_rsc_1_0_i_qb <= vec_rsc_1_0_qb;
  vec_rsc_1_0_db <= vec_rsc_1_0_i_db;
  vec_rsc_1_0_adrb <= vec_rsc_1_0_i_adrb;
  vec_rsc_1_0_i_qa <= vec_rsc_1_0_qa;
  vec_rsc_1_0_da <= vec_rsc_1_0_i_da;
  vec_rsc_1_0_adra <= vec_rsc_1_0_i_adra;
  vec_rsc_1_0_i_adra_d_1 <= vec_rsc_1_0_i_adra_d;
  vec_rsc_1_0_i_da_d_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000")
      & vec_rsc_1_0_i_da_d;
  vec_rsc_1_0_i_qa_d <= vec_rsc_1_0_i_qa_d_1;
  vec_rsc_1_0_i_wea_d_1 <= vec_rsc_1_0_i_wea_d;
  vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  vec_rsc_1_1_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_31_6_32_64_64_32_1_gen
    PORT MAP(
      qb => vec_rsc_1_1_i_qb,
      web => vec_rsc_1_1_web,
      db => vec_rsc_1_1_i_db,
      adrb => vec_rsc_1_1_i_adrb,
      qa => vec_rsc_1_1_i_qa,
      wea => vec_rsc_1_1_wea,
      da => vec_rsc_1_1_i_da,
      adra => vec_rsc_1_1_i_adra,
      adra_d => vec_rsc_1_1_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => vec_rsc_1_1_i_da_d_1,
      qa_d => vec_rsc_1_1_i_qa_d_1,
      wea_d => vec_rsc_1_1_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  vec_rsc_1_1_i_qb <= vec_rsc_1_1_qb;
  vec_rsc_1_1_db <= vec_rsc_1_1_i_db;
  vec_rsc_1_1_adrb <= vec_rsc_1_1_i_adrb;
  vec_rsc_1_1_i_qa <= vec_rsc_1_1_qa;
  vec_rsc_1_1_da <= vec_rsc_1_1_i_da;
  vec_rsc_1_1_adra <= vec_rsc_1_1_i_adra;
  vec_rsc_1_1_i_adra_d_1 <= vec_rsc_1_1_i_adra_d;
  vec_rsc_1_1_i_da_d_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000")
      & vec_rsc_1_1_i_da_d;
  vec_rsc_1_1_i_qa_d <= vec_rsc_1_1_i_qa_d_1;
  vec_rsc_1_1_i_wea_d_1 <= vec_rsc_1_1_i_wea_d;
  vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  vec_rsc_1_2_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_32_6_32_64_64_32_1_gen
    PORT MAP(
      qb => vec_rsc_1_2_i_qb,
      web => vec_rsc_1_2_web,
      db => vec_rsc_1_2_i_db,
      adrb => vec_rsc_1_2_i_adrb,
      qa => vec_rsc_1_2_i_qa,
      wea => vec_rsc_1_2_wea,
      da => vec_rsc_1_2_i_da,
      adra => vec_rsc_1_2_i_adra,
      adra_d => vec_rsc_1_2_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => vec_rsc_1_2_i_da_d_1,
      qa_d => vec_rsc_1_2_i_qa_d_1,
      wea_d => vec_rsc_1_2_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  vec_rsc_1_2_i_qb <= vec_rsc_1_2_qb;
  vec_rsc_1_2_db <= vec_rsc_1_2_i_db;
  vec_rsc_1_2_adrb <= vec_rsc_1_2_i_adrb;
  vec_rsc_1_2_i_qa <= vec_rsc_1_2_qa;
  vec_rsc_1_2_da <= vec_rsc_1_2_i_da;
  vec_rsc_1_2_adra <= vec_rsc_1_2_i_adra;
  vec_rsc_1_2_i_adra_d_1 <= vec_rsc_1_2_i_adra_d;
  vec_rsc_1_2_i_da_d_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000")
      & vec_rsc_1_2_i_da_d;
  vec_rsc_1_2_i_qa_d <= vec_rsc_1_2_i_qa_d_1;
  vec_rsc_1_2_i_wea_d_1 <= vec_rsc_1_2_i_wea_d;
  vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  vec_rsc_1_3_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_33_6_32_64_64_32_1_gen
    PORT MAP(
      qb => vec_rsc_1_3_i_qb,
      web => vec_rsc_1_3_web,
      db => vec_rsc_1_3_i_db,
      adrb => vec_rsc_1_3_i_adrb,
      qa => vec_rsc_1_3_i_qa,
      wea => vec_rsc_1_3_wea,
      da => vec_rsc_1_3_i_da,
      adra => vec_rsc_1_3_i_adra,
      adra_d => vec_rsc_1_3_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => vec_rsc_1_3_i_da_d_1,
      qa_d => vec_rsc_1_3_i_qa_d_1,
      wea_d => vec_rsc_1_3_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  vec_rsc_1_3_i_qb <= vec_rsc_1_3_qb;
  vec_rsc_1_3_db <= vec_rsc_1_3_i_db;
  vec_rsc_1_3_adrb <= vec_rsc_1_3_i_adrb;
  vec_rsc_1_3_i_qa <= vec_rsc_1_3_qa;
  vec_rsc_1_3_da <= vec_rsc_1_3_i_da;
  vec_rsc_1_3_adra <= vec_rsc_1_3_i_adra;
  vec_rsc_1_3_i_adra_d_1 <= vec_rsc_1_3_i_adra_d;
  vec_rsc_1_3_i_da_d_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000")
      & vec_rsc_1_3_i_da_d;
  vec_rsc_1_3_i_qa_d <= vec_rsc_1_3_i_qa_d_1;
  vec_rsc_1_3_i_wea_d_1 <= vec_rsc_1_3_i_wea_d;
  vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  vec_rsc_1_4_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_34_6_32_64_64_32_1_gen
    PORT MAP(
      qb => vec_rsc_1_4_i_qb,
      web => vec_rsc_1_4_web,
      db => vec_rsc_1_4_i_db,
      adrb => vec_rsc_1_4_i_adrb,
      qa => vec_rsc_1_4_i_qa,
      wea => vec_rsc_1_4_wea,
      da => vec_rsc_1_4_i_da,
      adra => vec_rsc_1_4_i_adra,
      adra_d => vec_rsc_1_4_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => vec_rsc_1_4_i_da_d_1,
      qa_d => vec_rsc_1_4_i_qa_d_1,
      wea_d => vec_rsc_1_4_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  vec_rsc_1_4_i_qb <= vec_rsc_1_4_qb;
  vec_rsc_1_4_db <= vec_rsc_1_4_i_db;
  vec_rsc_1_4_adrb <= vec_rsc_1_4_i_adrb;
  vec_rsc_1_4_i_qa <= vec_rsc_1_4_qa;
  vec_rsc_1_4_da <= vec_rsc_1_4_i_da;
  vec_rsc_1_4_adra <= vec_rsc_1_4_i_adra;
  vec_rsc_1_4_i_adra_d_1 <= vec_rsc_1_4_i_adra_d;
  vec_rsc_1_4_i_da_d_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000")
      & vec_rsc_1_4_i_da_d;
  vec_rsc_1_4_i_qa_d <= vec_rsc_1_4_i_qa_d_1;
  vec_rsc_1_4_i_wea_d_1 <= vec_rsc_1_4_i_wea_d;
  vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  vec_rsc_1_5_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_35_6_32_64_64_32_1_gen
    PORT MAP(
      qb => vec_rsc_1_5_i_qb,
      web => vec_rsc_1_5_web,
      db => vec_rsc_1_5_i_db,
      adrb => vec_rsc_1_5_i_adrb,
      qa => vec_rsc_1_5_i_qa,
      wea => vec_rsc_1_5_wea,
      da => vec_rsc_1_5_i_da,
      adra => vec_rsc_1_5_i_adra,
      adra_d => vec_rsc_1_5_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => vec_rsc_1_5_i_da_d_1,
      qa_d => vec_rsc_1_5_i_qa_d_1,
      wea_d => vec_rsc_1_5_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  vec_rsc_1_5_i_qb <= vec_rsc_1_5_qb;
  vec_rsc_1_5_db <= vec_rsc_1_5_i_db;
  vec_rsc_1_5_adrb <= vec_rsc_1_5_i_adrb;
  vec_rsc_1_5_i_qa <= vec_rsc_1_5_qa;
  vec_rsc_1_5_da <= vec_rsc_1_5_i_da;
  vec_rsc_1_5_adra <= vec_rsc_1_5_i_adra;
  vec_rsc_1_5_i_adra_d_1 <= vec_rsc_1_5_i_adra_d;
  vec_rsc_1_5_i_da_d_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000")
      & vec_rsc_1_5_i_da_d;
  vec_rsc_1_5_i_qa_d <= vec_rsc_1_5_i_qa_d_1;
  vec_rsc_1_5_i_wea_d_1 <= vec_rsc_1_5_i_wea_d;
  vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  vec_rsc_1_6_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_36_6_32_64_64_32_1_gen
    PORT MAP(
      qb => vec_rsc_1_6_i_qb,
      web => vec_rsc_1_6_web,
      db => vec_rsc_1_6_i_db,
      adrb => vec_rsc_1_6_i_adrb,
      qa => vec_rsc_1_6_i_qa,
      wea => vec_rsc_1_6_wea,
      da => vec_rsc_1_6_i_da,
      adra => vec_rsc_1_6_i_adra,
      adra_d => vec_rsc_1_6_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => vec_rsc_1_6_i_da_d_1,
      qa_d => vec_rsc_1_6_i_qa_d_1,
      wea_d => vec_rsc_1_6_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  vec_rsc_1_6_i_qb <= vec_rsc_1_6_qb;
  vec_rsc_1_6_db <= vec_rsc_1_6_i_db;
  vec_rsc_1_6_adrb <= vec_rsc_1_6_i_adrb;
  vec_rsc_1_6_i_qa <= vec_rsc_1_6_qa;
  vec_rsc_1_6_da <= vec_rsc_1_6_i_da;
  vec_rsc_1_6_adra <= vec_rsc_1_6_i_adra;
  vec_rsc_1_6_i_adra_d_1 <= vec_rsc_1_6_i_adra_d;
  vec_rsc_1_6_i_da_d_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000")
      & vec_rsc_1_6_i_da_d;
  vec_rsc_1_6_i_qa_d <= vec_rsc_1_6_i_qa_d_1;
  vec_rsc_1_6_i_wea_d_1 <= vec_rsc_1_6_i_wea_d;
  vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  vec_rsc_1_7_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_37_6_32_64_64_32_1_gen
    PORT MAP(
      qb => vec_rsc_1_7_i_qb,
      web => vec_rsc_1_7_web,
      db => vec_rsc_1_7_i_db,
      adrb => vec_rsc_1_7_i_adrb,
      qa => vec_rsc_1_7_i_qa,
      wea => vec_rsc_1_7_wea,
      da => vec_rsc_1_7_i_da,
      adra => vec_rsc_1_7_i_adra,
      adra_d => vec_rsc_1_7_i_adra_d_1,
      clka => clk,
      clka_en => '1',
      da_d => vec_rsc_1_7_i_da_d_1,
      qa_d => vec_rsc_1_7_i_qa_d_1,
      wea_d => vec_rsc_1_7_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  vec_rsc_1_7_i_qb <= vec_rsc_1_7_qb;
  vec_rsc_1_7_db <= vec_rsc_1_7_i_db;
  vec_rsc_1_7_adrb <= vec_rsc_1_7_i_adrb;
  vec_rsc_1_7_i_qa <= vec_rsc_1_7_qa;
  vec_rsc_1_7_da <= vec_rsc_1_7_i_da;
  vec_rsc_1_7_adra <= vec_rsc_1_7_i_adra;
  vec_rsc_1_7_i_adra_d_1 <= vec_rsc_1_7_i_adra_d;
  vec_rsc_1_7_i_da_d_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000")
      & vec_rsc_1_7_i_da_d;
  vec_rsc_1_7_i_qa_d <= vec_rsc_1_7_i_qa_d_1;
  vec_rsc_1_7_i_wea_d_1 <= vec_rsc_1_7_i_wea_d;
  vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  twiddle_rsc_0_0_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_38_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_0_i_qb,
      adrb => twiddle_rsc_0_0_i_adrb,
      adrb_d => twiddle_rsc_0_0_i_adrb_d,
      qb_d => twiddle_rsc_0_0_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_0_i_qb <= twiddle_rsc_0_0_qb;
  twiddle_rsc_0_0_adrb <= twiddle_rsc_0_0_i_adrb;
  twiddle_rsc_0_0_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_rsc_0_0_i_qb_d <= twiddle_rsc_0_0_i_qb_d_1;

  twiddle_rsc_0_1_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_39_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_1_i_qb,
      adrb => twiddle_rsc_0_1_i_adrb,
      adrb_d => twiddle_rsc_0_1_i_adrb_d,
      qb_d => twiddle_rsc_0_1_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_1_i_qb <= twiddle_rsc_0_1_qb;
  twiddle_rsc_0_1_adrb <= twiddle_rsc_0_1_i_adrb;
  twiddle_rsc_0_1_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_rsc_0_1_i_qb_d <= twiddle_rsc_0_1_i_qb_d_1;

  twiddle_rsc_0_2_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_40_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_2_i_qb,
      adrb => twiddle_rsc_0_2_i_adrb,
      adrb_d => twiddle_rsc_0_2_i_adrb_d,
      qb_d => twiddle_rsc_0_2_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_2_i_qb <= twiddle_rsc_0_2_qb;
  twiddle_rsc_0_2_adrb <= twiddle_rsc_0_2_i_adrb;
  twiddle_rsc_0_2_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_rsc_0_2_i_qb_d <= twiddle_rsc_0_2_i_qb_d_1;

  twiddle_rsc_0_3_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_41_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_3_i_qb,
      adrb => twiddle_rsc_0_3_i_adrb,
      adrb_d => twiddle_rsc_0_3_i_adrb_d,
      qb_d => twiddle_rsc_0_3_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_3_i_qb <= twiddle_rsc_0_3_qb;
  twiddle_rsc_0_3_adrb <= twiddle_rsc_0_3_i_adrb;
  twiddle_rsc_0_3_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_rsc_0_3_i_qb_d <= twiddle_rsc_0_3_i_qb_d_1;

  twiddle_rsc_0_4_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_42_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_4_i_qb,
      adrb => twiddle_rsc_0_4_i_adrb,
      adrb_d => twiddle_rsc_0_4_i_adrb_d,
      qb_d => twiddle_rsc_0_4_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_4_i_qb <= twiddle_rsc_0_4_qb;
  twiddle_rsc_0_4_adrb <= twiddle_rsc_0_4_i_adrb;
  twiddle_rsc_0_4_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_rsc_0_4_i_qb_d <= twiddle_rsc_0_4_i_qb_d_1;

  twiddle_rsc_0_5_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_43_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_5_i_qb,
      adrb => twiddle_rsc_0_5_i_adrb,
      adrb_d => twiddle_rsc_0_5_i_adrb_d,
      qb_d => twiddle_rsc_0_5_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_5_i_qb <= twiddle_rsc_0_5_qb;
  twiddle_rsc_0_5_adrb <= twiddle_rsc_0_5_i_adrb;
  twiddle_rsc_0_5_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_rsc_0_5_i_qb_d <= twiddle_rsc_0_5_i_qb_d_1;

  twiddle_rsc_0_6_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_44_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_6_i_qb,
      adrb => twiddle_rsc_0_6_i_adrb,
      adrb_d => twiddle_rsc_0_6_i_adrb_d,
      qb_d => twiddle_rsc_0_6_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_6_i_qb <= twiddle_rsc_0_6_qb;
  twiddle_rsc_0_6_adrb <= twiddle_rsc_0_6_i_adrb;
  twiddle_rsc_0_6_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_rsc_0_6_i_qb_d <= twiddle_rsc_0_6_i_qb_d_1;

  twiddle_rsc_0_7_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_45_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_0_7_i_qb,
      adrb => twiddle_rsc_0_7_i_adrb,
      adrb_d => twiddle_rsc_0_7_i_adrb_d,
      qb_d => twiddle_rsc_0_7_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_7_i_qb <= twiddle_rsc_0_7_qb;
  twiddle_rsc_0_7_adrb <= twiddle_rsc_0_7_i_adrb;
  twiddle_rsc_0_7_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_rsc_0_7_i_qb_d <= twiddle_rsc_0_7_i_qb_d_1;

  twiddle_rsc_1_0_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_46_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_1_0_i_qb,
      adrb => twiddle_rsc_1_0_i_adrb,
      adrb_d => twiddle_rsc_1_0_i_adrb_d,
      qb_d => twiddle_rsc_1_0_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_1_0_i_qb <= twiddle_rsc_1_0_qb;
  twiddle_rsc_1_0_adrb <= twiddle_rsc_1_0_i_adrb;
  twiddle_rsc_1_0_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_rsc_1_0_i_qb_d <= twiddle_rsc_1_0_i_qb_d_1;

  twiddle_rsc_1_1_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_47_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_1_1_i_qb,
      adrb => twiddle_rsc_1_1_i_adrb,
      adrb_d => twiddle_rsc_1_1_i_adrb_d,
      qb_d => twiddle_rsc_1_1_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_1_1_i_qb <= twiddle_rsc_1_1_qb;
  twiddle_rsc_1_1_adrb <= twiddle_rsc_1_1_i_adrb;
  twiddle_rsc_1_1_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_rsc_1_1_i_qb_d <= twiddle_rsc_1_1_i_qb_d_1;

  twiddle_rsc_1_2_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_48_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_1_2_i_qb,
      adrb => twiddle_rsc_1_2_i_adrb,
      adrb_d => twiddle_rsc_1_2_i_adrb_d,
      qb_d => twiddle_rsc_1_2_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_1_2_i_qb <= twiddle_rsc_1_2_qb;
  twiddle_rsc_1_2_adrb <= twiddle_rsc_1_2_i_adrb;
  twiddle_rsc_1_2_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_rsc_1_2_i_qb_d <= twiddle_rsc_1_2_i_qb_d_1;

  twiddle_rsc_1_3_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_49_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_1_3_i_qb,
      adrb => twiddle_rsc_1_3_i_adrb,
      adrb_d => twiddle_rsc_1_3_i_adrb_d,
      qb_d => twiddle_rsc_1_3_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_1_3_i_qb <= twiddle_rsc_1_3_qb;
  twiddle_rsc_1_3_adrb <= twiddle_rsc_1_3_i_adrb;
  twiddle_rsc_1_3_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_rsc_1_3_i_qb_d <= twiddle_rsc_1_3_i_qb_d_1;

  twiddle_rsc_1_4_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_50_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_1_4_i_qb,
      adrb => twiddle_rsc_1_4_i_adrb,
      adrb_d => twiddle_rsc_1_4_i_adrb_d,
      qb_d => twiddle_rsc_1_4_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_1_4_i_qb <= twiddle_rsc_1_4_qb;
  twiddle_rsc_1_4_adrb <= twiddle_rsc_1_4_i_adrb;
  twiddle_rsc_1_4_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_rsc_1_4_i_qb_d <= twiddle_rsc_1_4_i_qb_d_1;

  twiddle_rsc_1_5_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_51_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_1_5_i_qb,
      adrb => twiddle_rsc_1_5_i_adrb,
      adrb_d => twiddle_rsc_1_5_i_adrb_d,
      qb_d => twiddle_rsc_1_5_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_1_5_i_qb <= twiddle_rsc_1_5_qb;
  twiddle_rsc_1_5_adrb <= twiddle_rsc_1_5_i_adrb;
  twiddle_rsc_1_5_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_rsc_1_5_i_qb_d <= twiddle_rsc_1_5_i_qb_d_1;

  twiddle_rsc_1_6_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_52_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_1_6_i_qb,
      adrb => twiddle_rsc_1_6_i_adrb,
      adrb_d => twiddle_rsc_1_6_i_adrb_d,
      qb_d => twiddle_rsc_1_6_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_1_6_i_qb <= twiddle_rsc_1_6_qb;
  twiddle_rsc_1_6_adrb <= twiddle_rsc_1_6_i_adrb;
  twiddle_rsc_1_6_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_rsc_1_6_i_qb_d <= twiddle_rsc_1_6_i_qb_d_1;

  twiddle_rsc_1_7_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_53_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_rsc_1_7_i_qb,
      adrb => twiddle_rsc_1_7_i_adrb,
      adrb_d => twiddle_rsc_1_7_i_adrb_d,
      qb_d => twiddle_rsc_1_7_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_1_7_i_qb <= twiddle_rsc_1_7_qb;
  twiddle_rsc_1_7_adrb <= twiddle_rsc_1_7_i_adrb;
  twiddle_rsc_1_7_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_rsc_1_7_i_qb_d <= twiddle_rsc_1_7_i_qb_d_1;

  twiddle_h_rsc_0_0_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_54_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_0_i_qb,
      adrb => twiddle_h_rsc_0_0_i_adrb,
      adrb_d => twiddle_h_rsc_0_0_i_adrb_d,
      qb_d => twiddle_h_rsc_0_0_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsc_0_0_i_qb <= twiddle_h_rsc_0_0_qb;
  twiddle_h_rsc_0_0_adrb <= twiddle_h_rsc_0_0_i_adrb;
  twiddle_h_rsc_0_0_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_h_rsc_0_0_i_qb_d <= twiddle_h_rsc_0_0_i_qb_d_1;

  twiddle_h_rsc_0_1_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_55_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_1_i_qb,
      adrb => twiddle_h_rsc_0_1_i_adrb,
      adrb_d => twiddle_h_rsc_0_1_i_adrb_d,
      qb_d => twiddle_h_rsc_0_1_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsc_0_1_i_qb <= twiddle_h_rsc_0_1_qb;
  twiddle_h_rsc_0_1_adrb <= twiddle_h_rsc_0_1_i_adrb;
  twiddle_h_rsc_0_1_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_h_rsc_0_1_i_qb_d <= twiddle_h_rsc_0_1_i_qb_d_1;

  twiddle_h_rsc_0_2_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_56_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_2_i_qb,
      adrb => twiddle_h_rsc_0_2_i_adrb,
      adrb_d => twiddle_h_rsc_0_2_i_adrb_d,
      qb_d => twiddle_h_rsc_0_2_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsc_0_2_i_qb <= twiddle_h_rsc_0_2_qb;
  twiddle_h_rsc_0_2_adrb <= twiddle_h_rsc_0_2_i_adrb;
  twiddle_h_rsc_0_2_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_h_rsc_0_2_i_qb_d <= twiddle_h_rsc_0_2_i_qb_d_1;

  twiddle_h_rsc_0_3_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_57_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_3_i_qb,
      adrb => twiddle_h_rsc_0_3_i_adrb,
      adrb_d => twiddle_h_rsc_0_3_i_adrb_d,
      qb_d => twiddle_h_rsc_0_3_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsc_0_3_i_qb <= twiddle_h_rsc_0_3_qb;
  twiddle_h_rsc_0_3_adrb <= twiddle_h_rsc_0_3_i_adrb;
  twiddle_h_rsc_0_3_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_h_rsc_0_3_i_qb_d <= twiddle_h_rsc_0_3_i_qb_d_1;

  twiddle_h_rsc_0_4_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_58_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_4_i_qb,
      adrb => twiddle_h_rsc_0_4_i_adrb,
      adrb_d => twiddle_h_rsc_0_4_i_adrb_d,
      qb_d => twiddle_h_rsc_0_4_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsc_0_4_i_qb <= twiddle_h_rsc_0_4_qb;
  twiddle_h_rsc_0_4_adrb <= twiddle_h_rsc_0_4_i_adrb;
  twiddle_h_rsc_0_4_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_h_rsc_0_4_i_qb_d <= twiddle_h_rsc_0_4_i_qb_d_1;

  twiddle_h_rsc_0_5_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_59_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_5_i_qb,
      adrb => twiddle_h_rsc_0_5_i_adrb,
      adrb_d => twiddle_h_rsc_0_5_i_adrb_d,
      qb_d => twiddle_h_rsc_0_5_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsc_0_5_i_qb <= twiddle_h_rsc_0_5_qb;
  twiddle_h_rsc_0_5_adrb <= twiddle_h_rsc_0_5_i_adrb;
  twiddle_h_rsc_0_5_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_h_rsc_0_5_i_qb_d <= twiddle_h_rsc_0_5_i_qb_d_1;

  twiddle_h_rsc_0_6_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_60_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_6_i_qb,
      adrb => twiddle_h_rsc_0_6_i_adrb,
      adrb_d => twiddle_h_rsc_0_6_i_adrb_d,
      qb_d => twiddle_h_rsc_0_6_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsc_0_6_i_qb <= twiddle_h_rsc_0_6_qb;
  twiddle_h_rsc_0_6_adrb <= twiddle_h_rsc_0_6_i_adrb;
  twiddle_h_rsc_0_6_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_h_rsc_0_6_i_qb_d <= twiddle_h_rsc_0_6_i_qb_d_1;

  twiddle_h_rsc_0_7_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_61_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_0_7_i_qb,
      adrb => twiddle_h_rsc_0_7_i_adrb,
      adrb_d => twiddle_h_rsc_0_7_i_adrb_d,
      qb_d => twiddle_h_rsc_0_7_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsc_0_7_i_qb <= twiddle_h_rsc_0_7_qb;
  twiddle_h_rsc_0_7_adrb <= twiddle_h_rsc_0_7_i_adrb;
  twiddle_h_rsc_0_7_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_h_rsc_0_7_i_qb_d <= twiddle_h_rsc_0_7_i_qb_d_1;

  twiddle_h_rsc_1_0_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_62_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_1_0_i_qb,
      adrb => twiddle_h_rsc_1_0_i_adrb,
      adrb_d => twiddle_h_rsc_1_0_i_adrb_d,
      qb_d => twiddle_h_rsc_1_0_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsc_1_0_i_qb <= twiddle_h_rsc_1_0_qb;
  twiddle_h_rsc_1_0_adrb <= twiddle_h_rsc_1_0_i_adrb;
  twiddle_h_rsc_1_0_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_h_rsc_1_0_i_qb_d <= twiddle_h_rsc_1_0_i_qb_d_1;

  twiddle_h_rsc_1_1_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_63_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_1_1_i_qb,
      adrb => twiddle_h_rsc_1_1_i_adrb,
      adrb_d => twiddle_h_rsc_1_1_i_adrb_d,
      qb_d => twiddle_h_rsc_1_1_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsc_1_1_i_qb <= twiddle_h_rsc_1_1_qb;
  twiddle_h_rsc_1_1_adrb <= twiddle_h_rsc_1_1_i_adrb;
  twiddle_h_rsc_1_1_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_h_rsc_1_1_i_qb_d <= twiddle_h_rsc_1_1_i_qb_d_1;

  twiddle_h_rsc_1_2_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_64_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_1_2_i_qb,
      adrb => twiddle_h_rsc_1_2_i_adrb,
      adrb_d => twiddle_h_rsc_1_2_i_adrb_d,
      qb_d => twiddle_h_rsc_1_2_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsc_1_2_i_qb <= twiddle_h_rsc_1_2_qb;
  twiddle_h_rsc_1_2_adrb <= twiddle_h_rsc_1_2_i_adrb;
  twiddle_h_rsc_1_2_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_h_rsc_1_2_i_qb_d <= twiddle_h_rsc_1_2_i_qb_d_1;

  twiddle_h_rsc_1_3_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_65_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_1_3_i_qb,
      adrb => twiddle_h_rsc_1_3_i_adrb,
      adrb_d => twiddle_h_rsc_1_3_i_adrb_d,
      qb_d => twiddle_h_rsc_1_3_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsc_1_3_i_qb <= twiddle_h_rsc_1_3_qb;
  twiddle_h_rsc_1_3_adrb <= twiddle_h_rsc_1_3_i_adrb;
  twiddle_h_rsc_1_3_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_h_rsc_1_3_i_qb_d <= twiddle_h_rsc_1_3_i_qb_d_1;

  twiddle_h_rsc_1_4_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_66_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_1_4_i_qb,
      adrb => twiddle_h_rsc_1_4_i_adrb,
      adrb_d => twiddle_h_rsc_1_4_i_adrb_d,
      qb_d => twiddle_h_rsc_1_4_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsc_1_4_i_qb <= twiddle_h_rsc_1_4_qb;
  twiddle_h_rsc_1_4_adrb <= twiddle_h_rsc_1_4_i_adrb;
  twiddle_h_rsc_1_4_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_h_rsc_1_4_i_qb_d <= twiddle_h_rsc_1_4_i_qb_d_1;

  twiddle_h_rsc_1_5_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_67_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_1_5_i_qb,
      adrb => twiddle_h_rsc_1_5_i_adrb,
      adrb_d => twiddle_h_rsc_1_5_i_adrb_d,
      qb_d => twiddle_h_rsc_1_5_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsc_1_5_i_qb <= twiddle_h_rsc_1_5_qb;
  twiddle_h_rsc_1_5_adrb <= twiddle_h_rsc_1_5_i_adrb;
  twiddle_h_rsc_1_5_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_h_rsc_1_5_i_qb_d <= twiddle_h_rsc_1_5_i_qb_d_1;

  twiddle_h_rsc_1_6_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_68_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_1_6_i_qb,
      adrb => twiddle_h_rsc_1_6_i_adrb,
      adrb_d => twiddle_h_rsc_1_6_i_adrb_d,
      qb_d => twiddle_h_rsc_1_6_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsc_1_6_i_qb <= twiddle_h_rsc_1_6_qb;
  twiddle_h_rsc_1_6_adrb <= twiddle_h_rsc_1_6_i_adrb;
  twiddle_h_rsc_1_6_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_h_rsc_1_6_i_qb_d <= twiddle_h_rsc_1_6_i_qb_d_1;

  twiddle_h_rsc_1_7_i : inPlaceNTT_DIF_precomp_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rport_69_6_32_64_64_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsc_1_7_i_qb,
      adrb => twiddle_h_rsc_1_7_i_adrb,
      adrb_d => twiddle_h_rsc_1_7_i_adrb_d,
      qb_d => twiddle_h_rsc_1_7_i_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsc_1_7_i_qb <= twiddle_h_rsc_1_7_qb;
  twiddle_h_rsc_1_7_adrb <= twiddle_h_rsc_1_7_i_adrb;
  twiddle_h_rsc_1_7_i_adrb_d <= twiddle_rsc_0_0_i_adrb_d_iff;
  twiddle_h_rsc_1_7_i_qb_d <= twiddle_h_rsc_1_7_i_qb_d_1;

  inPlaceNTT_DIF_precomp_core_inst : inPlaceNTT_DIF_precomp_core
    PORT MAP(
      clk => clk,
      rst => rst,
      run_rsc_rdy => run_rsc_rdy,
      run_rsc_vld => run_rsc_vld,
      vec_rsc_triosy_0_0_lz => vec_rsc_triosy_0_0_lz,
      vec_rsc_triosy_0_1_lz => vec_rsc_triosy_0_1_lz,
      vec_rsc_triosy_0_2_lz => vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz => vec_rsc_triosy_0_3_lz,
      vec_rsc_triosy_0_4_lz => vec_rsc_triosy_0_4_lz,
      vec_rsc_triosy_0_5_lz => vec_rsc_triosy_0_5_lz,
      vec_rsc_triosy_0_6_lz => vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz => vec_rsc_triosy_0_7_lz,
      vec_rsc_triosy_1_0_lz => vec_rsc_triosy_1_0_lz,
      vec_rsc_triosy_1_1_lz => vec_rsc_triosy_1_1_lz,
      vec_rsc_triosy_1_2_lz => vec_rsc_triosy_1_2_lz,
      vec_rsc_triosy_1_3_lz => vec_rsc_triosy_1_3_lz,
      vec_rsc_triosy_1_4_lz => vec_rsc_triosy_1_4_lz,
      vec_rsc_triosy_1_5_lz => vec_rsc_triosy_1_5_lz,
      vec_rsc_triosy_1_6_lz => vec_rsc_triosy_1_6_lz,
      vec_rsc_triosy_1_7_lz => vec_rsc_triosy_1_7_lz,
      p_rsc_dat => inPlaceNTT_DIF_precomp_core_inst_p_rsc_dat,
      p_rsc_triosy_lz => p_rsc_triosy_lz,
      r_rsc_triosy_lz => r_rsc_triosy_lz,
      twiddle_rsc_triosy_0_0_lz => twiddle_rsc_triosy_0_0_lz,
      twiddle_rsc_triosy_0_1_lz => twiddle_rsc_triosy_0_1_lz,
      twiddle_rsc_triosy_0_2_lz => twiddle_rsc_triosy_0_2_lz,
      twiddle_rsc_triosy_0_3_lz => twiddle_rsc_triosy_0_3_lz,
      twiddle_rsc_triosy_0_4_lz => twiddle_rsc_triosy_0_4_lz,
      twiddle_rsc_triosy_0_5_lz => twiddle_rsc_triosy_0_5_lz,
      twiddle_rsc_triosy_0_6_lz => twiddle_rsc_triosy_0_6_lz,
      twiddle_rsc_triosy_0_7_lz => twiddle_rsc_triosy_0_7_lz,
      twiddle_rsc_triosy_1_0_lz => twiddle_rsc_triosy_1_0_lz,
      twiddle_rsc_triosy_1_1_lz => twiddle_rsc_triosy_1_1_lz,
      twiddle_rsc_triosy_1_2_lz => twiddle_rsc_triosy_1_2_lz,
      twiddle_rsc_triosy_1_3_lz => twiddle_rsc_triosy_1_3_lz,
      twiddle_rsc_triosy_1_4_lz => twiddle_rsc_triosy_1_4_lz,
      twiddle_rsc_triosy_1_5_lz => twiddle_rsc_triosy_1_5_lz,
      twiddle_rsc_triosy_1_6_lz => twiddle_rsc_triosy_1_6_lz,
      twiddle_rsc_triosy_1_7_lz => twiddle_rsc_triosy_1_7_lz,
      twiddle_h_rsc_triosy_0_0_lz => twiddle_h_rsc_triosy_0_0_lz,
      twiddle_h_rsc_triosy_0_1_lz => twiddle_h_rsc_triosy_0_1_lz,
      twiddle_h_rsc_triosy_0_2_lz => twiddle_h_rsc_triosy_0_2_lz,
      twiddle_h_rsc_triosy_0_3_lz => twiddle_h_rsc_triosy_0_3_lz,
      twiddle_h_rsc_triosy_0_4_lz => twiddle_h_rsc_triosy_0_4_lz,
      twiddle_h_rsc_triosy_0_5_lz => twiddle_h_rsc_triosy_0_5_lz,
      twiddle_h_rsc_triosy_0_6_lz => twiddle_h_rsc_triosy_0_6_lz,
      twiddle_h_rsc_triosy_0_7_lz => twiddle_h_rsc_triosy_0_7_lz,
      twiddle_h_rsc_triosy_1_0_lz => twiddle_h_rsc_triosy_1_0_lz,
      twiddle_h_rsc_triosy_1_1_lz => twiddle_h_rsc_triosy_1_1_lz,
      twiddle_h_rsc_triosy_1_2_lz => twiddle_h_rsc_triosy_1_2_lz,
      twiddle_h_rsc_triosy_1_3_lz => twiddle_h_rsc_triosy_1_3_lz,
      twiddle_h_rsc_triosy_1_4_lz => twiddle_h_rsc_triosy_1_4_lz,
      twiddle_h_rsc_triosy_1_5_lz => twiddle_h_rsc_triosy_1_5_lz,
      twiddle_h_rsc_triosy_1_6_lz => twiddle_h_rsc_triosy_1_6_lz,
      twiddle_h_rsc_triosy_1_7_lz => twiddle_h_rsc_triosy_1_7_lz,
      complete_rsc_rdy => complete_rsc_rdy,
      complete_rsc_vld => complete_rsc_vld,
      vec_rsc_0_0_i_adra_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_adra_d,
      vec_rsc_0_0_i_da_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_da_d,
      vec_rsc_0_0_i_qa_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_qa_d,
      vec_rsc_0_0_i_wea_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_wea_d,
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      vec_rsc_0_1_i_adra_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_adra_d,
      vec_rsc_0_1_i_da_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_da_d,
      vec_rsc_0_1_i_qa_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_qa_d,
      vec_rsc_0_1_i_wea_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_wea_d,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      vec_rsc_0_2_i_adra_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_adra_d,
      vec_rsc_0_2_i_da_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_da_d,
      vec_rsc_0_2_i_qa_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_qa_d,
      vec_rsc_0_2_i_wea_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_wea_d,
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      vec_rsc_0_3_i_adra_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_adra_d,
      vec_rsc_0_3_i_da_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_da_d,
      vec_rsc_0_3_i_qa_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_qa_d,
      vec_rsc_0_3_i_wea_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_wea_d,
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      vec_rsc_0_4_i_adra_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_adra_d,
      vec_rsc_0_4_i_da_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_da_d,
      vec_rsc_0_4_i_qa_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_qa_d,
      vec_rsc_0_4_i_wea_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_wea_d,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      vec_rsc_0_5_i_adra_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_adra_d,
      vec_rsc_0_5_i_da_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_da_d,
      vec_rsc_0_5_i_qa_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_qa_d,
      vec_rsc_0_5_i_wea_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_wea_d,
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      vec_rsc_0_6_i_adra_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_adra_d,
      vec_rsc_0_6_i_da_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_da_d,
      vec_rsc_0_6_i_qa_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_qa_d,
      vec_rsc_0_6_i_wea_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_wea_d,
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      vec_rsc_0_7_i_adra_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_adra_d,
      vec_rsc_0_7_i_da_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_da_d,
      vec_rsc_0_7_i_qa_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_qa_d,
      vec_rsc_0_7_i_wea_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_wea_d,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      vec_rsc_1_0_i_adra_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_adra_d,
      vec_rsc_1_0_i_da_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_da_d,
      vec_rsc_1_0_i_qa_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_qa_d,
      vec_rsc_1_0_i_wea_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_wea_d,
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      vec_rsc_1_1_i_adra_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_adra_d,
      vec_rsc_1_1_i_da_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_da_d,
      vec_rsc_1_1_i_qa_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_qa_d,
      vec_rsc_1_1_i_wea_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_wea_d,
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      vec_rsc_1_2_i_adra_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_adra_d,
      vec_rsc_1_2_i_da_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_da_d,
      vec_rsc_1_2_i_qa_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_qa_d,
      vec_rsc_1_2_i_wea_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_wea_d,
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      vec_rsc_1_3_i_adra_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_adra_d,
      vec_rsc_1_3_i_da_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_da_d,
      vec_rsc_1_3_i_qa_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_qa_d,
      vec_rsc_1_3_i_wea_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_wea_d,
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      vec_rsc_1_4_i_adra_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_adra_d,
      vec_rsc_1_4_i_da_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_da_d,
      vec_rsc_1_4_i_qa_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_qa_d,
      vec_rsc_1_4_i_wea_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_wea_d,
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      vec_rsc_1_5_i_adra_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_adra_d,
      vec_rsc_1_5_i_da_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_da_d,
      vec_rsc_1_5_i_qa_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_qa_d,
      vec_rsc_1_5_i_wea_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_wea_d,
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      vec_rsc_1_6_i_adra_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_adra_d,
      vec_rsc_1_6_i_da_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_da_d,
      vec_rsc_1_6_i_qa_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_qa_d,
      vec_rsc_1_6_i_wea_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_wea_d,
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      vec_rsc_1_7_i_adra_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_adra_d,
      vec_rsc_1_7_i_da_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_da_d,
      vec_rsc_1_7_i_qa_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_qa_d,
      vec_rsc_1_7_i_wea_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_wea_d,
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d => inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      twiddle_rsc_0_0_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_0_i_qb_d,
      twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_1_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_1_i_qb_d,
      twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_2_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_2_i_qb_d,
      twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_3_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_3_i_qb_d,
      twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_4_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_4_i_qb_d,
      twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_5_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_5_i_qb_d,
      twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_6_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_6_i_qb_d,
      twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_7_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_7_i_qb_d,
      twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_1_0_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_0_i_qb_d,
      twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_1_1_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_1_i_qb_d,
      twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_1_2_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_2_i_qb_d,
      twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_1_3_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_3_i_qb_d,
      twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_1_4_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_4_i_qb_d,
      twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_1_5_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_5_i_qb_d,
      twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_1_6_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_6_i_qb_d,
      twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_1_7_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_7_i_qb_d,
      twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_0_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_0_i_qb_d,
      twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_0_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_1_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_1_i_qb_d,
      twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_1_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_2_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_2_i_qb_d,
      twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_2_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_3_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_3_i_qb_d,
      twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_3_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_4_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_4_i_qb_d,
      twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_4_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_5_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_5_i_qb_d,
      twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_5_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_6_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_6_i_qb_d,
      twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_6_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_7_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_7_i_qb_d,
      twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_0_7_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_1_0_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_0_i_qb_d,
      twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_0_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_1_1_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_1_i_qb_d,
      twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_1_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_1_2_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_2_i_qb_d,
      twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_2_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_1_3_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_3_i_qb_d,
      twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_3_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_1_4_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_4_i_qb_d,
      twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_4_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_1_5_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_5_i_qb_d,
      twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_5_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_1_6_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_6_i_qb_d,
      twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_6_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_1_7_i_qb_d => inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_7_i_qb_d,
      twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsc_1_7_i_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_0_i_adrb_d_pff => inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_0_i_adrb_d_pff
    );
  inPlaceNTT_DIF_precomp_core_inst_p_rsc_dat <= p_rsc_dat;
  vec_rsc_0_0_i_adra_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_adra_d;
  vec_rsc_0_0_i_da_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_da_d;
  inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_qa_d <= vec_rsc_0_0_i_qa_d;
  vec_rsc_0_0_i_wea_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_wea_d;
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  vec_rsc_0_1_i_adra_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_adra_d;
  vec_rsc_0_1_i_da_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_da_d;
  inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_qa_d <= vec_rsc_0_1_i_qa_d;
  vec_rsc_0_1_i_wea_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_wea_d;
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  vec_rsc_0_2_i_adra_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_adra_d;
  vec_rsc_0_2_i_da_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_da_d;
  inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_qa_d <= vec_rsc_0_2_i_qa_d;
  vec_rsc_0_2_i_wea_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_wea_d;
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_2_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  vec_rsc_0_3_i_adra_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_adra_d;
  vec_rsc_0_3_i_da_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_da_d;
  inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_qa_d <= vec_rsc_0_3_i_qa_d;
  vec_rsc_0_3_i_wea_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_wea_d;
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_3_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  vec_rsc_0_4_i_adra_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_adra_d;
  vec_rsc_0_4_i_da_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_da_d;
  inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_qa_d <= vec_rsc_0_4_i_qa_d;
  vec_rsc_0_4_i_wea_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_wea_d;
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_4_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  vec_rsc_0_5_i_adra_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_adra_d;
  vec_rsc_0_5_i_da_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_da_d;
  inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_qa_d <= vec_rsc_0_5_i_qa_d;
  vec_rsc_0_5_i_wea_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_wea_d;
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_5_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  vec_rsc_0_6_i_adra_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_adra_d;
  vec_rsc_0_6_i_da_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_da_d;
  inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_qa_d <= vec_rsc_0_6_i_qa_d;
  vec_rsc_0_6_i_wea_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_wea_d;
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_6_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  vec_rsc_0_7_i_adra_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_adra_d;
  vec_rsc_0_7_i_da_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_da_d;
  inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_qa_d <= vec_rsc_0_7_i_qa_d;
  vec_rsc_0_7_i_wea_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_wea_d;
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_0_7_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  vec_rsc_1_0_i_adra_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_adra_d;
  vec_rsc_1_0_i_da_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_da_d;
  inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_qa_d <= vec_rsc_1_0_i_qa_d;
  vec_rsc_1_0_i_wea_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_wea_d;
  vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  vec_rsc_1_1_i_adra_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_adra_d;
  vec_rsc_1_1_i_da_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_da_d;
  inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_qa_d <= vec_rsc_1_1_i_qa_d;
  vec_rsc_1_1_i_wea_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_wea_d;
  vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_1_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  vec_rsc_1_2_i_adra_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_adra_d;
  vec_rsc_1_2_i_da_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_da_d;
  inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_qa_d <= vec_rsc_1_2_i_qa_d;
  vec_rsc_1_2_i_wea_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_wea_d;
  vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_2_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  vec_rsc_1_3_i_adra_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_adra_d;
  vec_rsc_1_3_i_da_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_da_d;
  inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_qa_d <= vec_rsc_1_3_i_qa_d;
  vec_rsc_1_3_i_wea_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_wea_d;
  vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_3_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  vec_rsc_1_4_i_adra_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_adra_d;
  vec_rsc_1_4_i_da_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_da_d;
  inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_qa_d <= vec_rsc_1_4_i_qa_d;
  vec_rsc_1_4_i_wea_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_wea_d;
  vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_4_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  vec_rsc_1_5_i_adra_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_adra_d;
  vec_rsc_1_5_i_da_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_da_d;
  inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_qa_d <= vec_rsc_1_5_i_qa_d;
  vec_rsc_1_5_i_wea_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_wea_d;
  vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_5_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  vec_rsc_1_6_i_adra_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_adra_d;
  vec_rsc_1_6_i_da_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_da_d;
  inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_qa_d <= vec_rsc_1_6_i_qa_d;
  vec_rsc_1_6_i_wea_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_wea_d;
  vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_6_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  vec_rsc_1_7_i_adra_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_adra_d;
  vec_rsc_1_7_i_da_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_da_d;
  inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_qa_d <= vec_rsc_1_7_i_qa_d;
  vec_rsc_1_7_i_wea_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_wea_d;
  vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d <= inPlaceNTT_DIF_precomp_core_inst_vec_rsc_1_7_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_0_i_qb_d <= twiddle_rsc_0_0_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_1_i_qb_d <= twiddle_rsc_0_1_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_2_i_qb_d <= twiddle_rsc_0_2_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_3_i_qb_d <= twiddle_rsc_0_3_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_4_i_qb_d <= twiddle_rsc_0_4_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_5_i_qb_d <= twiddle_rsc_0_5_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_6_i_qb_d <= twiddle_rsc_0_6_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_7_i_qb_d <= twiddle_rsc_0_7_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_0_i_qb_d <= twiddle_rsc_1_0_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_1_i_qb_d <= twiddle_rsc_1_1_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_2_i_qb_d <= twiddle_rsc_1_2_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_3_i_qb_d <= twiddle_rsc_1_3_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_4_i_qb_d <= twiddle_rsc_1_4_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_5_i_qb_d <= twiddle_rsc_1_5_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_6_i_qb_d <= twiddle_rsc_1_6_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_1_7_i_qb_d <= twiddle_rsc_1_7_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_0_i_qb_d <= twiddle_h_rsc_0_0_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_1_i_qb_d <= twiddle_h_rsc_0_1_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_2_i_qb_d <= twiddle_h_rsc_0_2_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_3_i_qb_d <= twiddle_h_rsc_0_3_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_4_i_qb_d <= twiddle_h_rsc_0_4_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_5_i_qb_d <= twiddle_h_rsc_0_5_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_6_i_qb_d <= twiddle_h_rsc_0_6_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_0_7_i_qb_d <= twiddle_h_rsc_0_7_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_0_i_qb_d <= twiddle_h_rsc_1_0_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_1_i_qb_d <= twiddle_h_rsc_1_1_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_2_i_qb_d <= twiddle_h_rsc_1_2_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_3_i_qb_d <= twiddle_h_rsc_1_3_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_4_i_qb_d <= twiddle_h_rsc_1_4_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_5_i_qb_d <= twiddle_h_rsc_1_5_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_6_i_qb_d <= twiddle_h_rsc_1_6_i_qb_d;
  inPlaceNTT_DIF_precomp_core_inst_twiddle_h_rsc_1_7_i_qb_d <= twiddle_h_rsc_1_7_i_qb_d;
  twiddle_rsc_0_0_i_adrb_d_iff <= inPlaceNTT_DIF_precomp_core_inst_twiddle_rsc_0_0_i_adrb_d_pff;

END v5;



