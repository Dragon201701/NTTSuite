
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.v 
module mgc_rem(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_b-1:0] z;  
   reg  [width_b-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  rem_s(a,b,z);
	else
          rem_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> ../td_ccore_solutions/modulo_dev_bb61c76201db0c9669a47462bb7d006361ff_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Tue Jul 20 15:24:30 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    modulo_dev_core
// ------------------------------------------------------------------


module modulo_dev_core (
  base_rsc_dat, m_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [63:0] base_rsc_dat;
  input [63:0] m_rsc_dat;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [63:0] base_rsci_idat;
  wire [63:0] m_rsci_idat;
  reg [63:0] return_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire [64:0] rem_13_cmp_z;
  wire [64:0] rem_13_cmp_1_z;
  wire [64:0] rem_13_cmp_2_z;
  wire [64:0] rem_13_cmp_3_z;
  wire [64:0] rem_13_cmp_4_z;
  wire [64:0] rem_13_cmp_5_z;
  wire [64:0] rem_13_cmp_6_z;
  wire [64:0] rem_13_cmp_7_z;
  wire [64:0] rem_13_cmp_8_z;
  wire [64:0] rem_13_cmp_9_z;
  wire [64:0] rem_13_cmp_10_z;
  wire [64:0] rem_13_cmp_11_z;
  reg [63:0] rem_13_cmp_b_63_0;
  reg [63:0] rem_13_cmp_1_b_63_0;
  reg [63:0] rem_13_cmp_2_b_63_0;
  reg [63:0] rem_13_cmp_3_b_63_0;
  reg [63:0] rem_13_cmp_4_b_63_0;
  reg [63:0] rem_13_cmp_5_b_63_0;
  reg [63:0] rem_13_cmp_6_b_63_0;
  reg [63:0] rem_13_cmp_7_b_63_0;
  reg [63:0] rem_13_cmp_8_b_63_0;
  reg [63:0] rem_13_cmp_9_b_63_0;
  reg [63:0] rem_13_cmp_10_b_63_0;
  reg [63:0] rem_13_cmp_11_b_63_0;
  reg [63:0] rem_13_cmp_a_63_0;
  reg [63:0] rem_13_cmp_1_a_63_0;
  reg [63:0] rem_13_cmp_2_a_63_0;
  reg [63:0] rem_13_cmp_3_a_63_0;
  reg [63:0] rem_13_cmp_4_a_63_0;
  reg [63:0] rem_13_cmp_5_a_63_0;
  reg [63:0] rem_13_cmp_6_a_63_0;
  reg [63:0] rem_13_cmp_7_a_63_0;
  reg [63:0] rem_13_cmp_8_a_63_0;
  reg [63:0] rem_13_cmp_9_a_63_0;
  reg [63:0] rem_13_cmp_10_a_63_0;
  reg [63:0] rem_13_cmp_11_a_63_0;
  wire [1:0] acc_tmp;
  wire [2:0] nl_acc_tmp;
  wire [3:0] acc_1_tmp;
  wire [4:0] nl_acc_1_tmp;
  wire and_dcpl_1;
  wire and_dcpl_2;
  wire and_dcpl_3;
  wire and_dcpl_4;
  wire and_dcpl_6;
  wire and_dcpl_8;
  wire and_dcpl_9;
  wire and_dcpl_11;
  wire and_dcpl_13;
  wire and_dcpl_18;
  wire and_dcpl_23;
  wire and_dcpl_28;
  wire and_dcpl_29;
  wire and_dcpl_30;
  wire and_dcpl_31;
  wire and_dcpl_33;
  wire and_dcpl_35;
  wire and_dcpl_36;
  wire and_dcpl_38;
  wire and_dcpl_40;
  wire and_dcpl_45;
  wire and_dcpl_50;
  wire and_dcpl_55;
  wire and_dcpl_56;
  wire and_dcpl_57;
  wire and_dcpl_58;
  wire and_dcpl_60;
  wire and_dcpl_62;
  wire and_dcpl_63;
  wire and_dcpl_65;
  wire and_dcpl_67;
  wire and_dcpl_72;
  wire and_dcpl_77;
  wire and_dcpl_82;
  wire and_dcpl_83;
  wire and_dcpl_84;
  wire and_dcpl_85;
  wire and_dcpl_87;
  wire and_dcpl_89;
  wire and_dcpl_90;
  wire and_dcpl_92;
  wire and_dcpl_94;
  wire and_dcpl_99;
  wire and_dcpl_104;
  wire and_dcpl_109;
  wire and_dcpl_110;
  wire and_dcpl_111;
  wire and_dcpl_112;
  wire and_dcpl_114;
  wire and_dcpl_115;
  wire and_dcpl_117;
  wire and_dcpl_119;
  wire and_dcpl_121;
  wire and_dcpl_126;
  wire and_dcpl_129;
  wire and_dcpl_136;
  wire and_dcpl_137;
  wire and_dcpl_138;
  wire and_dcpl_139;
  wire and_dcpl_141;
  wire and_dcpl_143;
  wire and_dcpl_144;
  wire and_dcpl_146;
  wire and_dcpl_148;
  wire and_dcpl_153;
  wire and_dcpl_158;
  wire and_dcpl_163;
  wire and_dcpl_164;
  wire and_dcpl_165;
  wire and_dcpl_166;
  wire and_dcpl_168;
  wire and_dcpl_170;
  wire and_dcpl_171;
  wire and_dcpl_173;
  wire and_dcpl_175;
  wire and_dcpl_180;
  wire and_dcpl_185;
  wire and_dcpl_190;
  wire and_dcpl_191;
  wire and_dcpl_192;
  wire and_dcpl_193;
  wire and_dcpl_195;
  wire and_dcpl_197;
  wire and_dcpl_198;
  wire and_dcpl_200;
  wire and_dcpl_202;
  wire and_dcpl_207;
  wire and_dcpl_212;
  wire and_dcpl_217;
  wire and_dcpl_218;
  wire and_dcpl_219;
  wire and_dcpl_220;
  wire and_dcpl_222;
  wire and_dcpl_224;
  wire and_dcpl_225;
  wire and_dcpl_227;
  wire and_dcpl_229;
  wire and_dcpl_234;
  wire and_dcpl_239;
  wire and_dcpl_244;
  wire and_dcpl_245;
  wire and_dcpl_246;
  wire and_dcpl_247;
  wire and_dcpl_249;
  wire and_dcpl_251;
  wire and_dcpl_252;
  wire and_dcpl_254;
  wire and_dcpl_256;
  wire and_dcpl_261;
  wire and_dcpl_266;
  wire and_dcpl_271;
  wire and_dcpl_272;
  wire and_dcpl_274;
  wire and_dcpl_276;
  wire and_dcpl_278;
  wire and_dcpl_280;
  wire and_dcpl_285;
  wire and_dcpl_291;
  wire and_dcpl_292;
  wire and_dcpl_293;
  wire and_dcpl_294;
  wire and_dcpl_295;
  wire and_dcpl_296;
  wire and_dcpl_298;
  wire not_tmp_54;
  wire or_tmp_2;
  wire and_dcpl_300;
  wire and_dcpl_301;
  wire and_dcpl_302;
  wire and_dcpl_304;
  wire and_tmp;
  wire and_dcpl_306;
  wire and_dcpl_307;
  wire and_dcpl_308;
  wire and_dcpl_310;
  wire and_tmp_2;
  wire and_dcpl_312;
  wire and_dcpl_313;
  wire and_dcpl_314;
  wire and_dcpl_316;
  wire and_tmp_5;
  wire and_dcpl_318;
  wire and_tmp_9;
  wire and_dcpl_324;
  wire and_tmp_13;
  wire and_dcpl_330;
  wire mux_tmp_19;
  wire and_tmp_17;
  wire and_dcpl_336;
  wire mux_tmp_22;
  wire mux_tmp_23;
  wire and_tmp_21;
  wire and_dcpl_342;
  wire mux_tmp_26;
  wire mux_tmp_27;
  wire mux_tmp_28;
  wire and_tmp_25;
  wire and_dcpl_348;
  wire and_tmp_35;
  wire and_dcpl_355;
  wire and_dcpl_356;
  wire and_dcpl_358;
  wire or_tmp_80;
  wire and_dcpl_360;
  wire and_dcpl_362;
  wire mux_tmp_32;
  wire and_dcpl_364;
  wire and_dcpl_366;
  wire mux_tmp_34;
  wire mux_tmp_35;
  wire and_dcpl_368;
  wire and_dcpl_370;
  wire mux_tmp_37;
  wire mux_tmp_38;
  wire mux_tmp_39;
  wire and_dcpl_372;
  wire mux_tmp_41;
  wire mux_tmp_42;
  wire mux_tmp_43;
  wire mux_tmp_44;
  wire and_dcpl_376;
  wire mux_tmp_46;
  wire mux_tmp_47;
  wire mux_tmp_48;
  wire mux_tmp_49;
  wire mux_tmp_50;
  wire and_dcpl_379;
  wire mux_tmp_52;
  wire mux_tmp_53;
  wire mux_tmp_54;
  wire mux_tmp_55;
  wire mux_tmp_56;
  wire mux_tmp_57;
  wire and_dcpl_382;
  wire mux_tmp_59;
  wire mux_tmp_60;
  wire mux_tmp_61;
  wire mux_tmp_62;
  wire mux_tmp_63;
  wire mux_tmp_64;
  wire mux_tmp_65;
  wire and_dcpl_385;
  wire mux_tmp_67;
  wire mux_tmp_68;
  wire mux_tmp_69;
  wire mux_tmp_70;
  wire mux_tmp_71;
  wire mux_tmp_72;
  wire mux_tmp_73;
  wire mux_tmp_74;
  wire and_dcpl_388;
  wire and_tmp_44;
  wire mux_tmp_76;
  wire and_dcpl_393;
  wire and_dcpl_394;
  wire and_dcpl_395;
  wire or_tmp_185;
  wire and_dcpl_397;
  wire and_dcpl_398;
  wire and_tmp_45;
  wire and_dcpl_400;
  wire and_dcpl_401;
  wire and_tmp_47;
  wire and_dcpl_403;
  wire and_dcpl_404;
  wire and_tmp_50;
  wire and_dcpl_406;
  wire and_tmp_54;
  wire and_dcpl_409;
  wire and_tmp_58;
  wire and_dcpl_413;
  wire mux_tmp_84;
  wire and_tmp_62;
  wire and_dcpl_417;
  wire mux_tmp_87;
  wire mux_tmp_88;
  wire and_tmp_66;
  wire and_dcpl_421;
  wire mux_tmp_91;
  wire mux_tmp_92;
  wire mux_tmp_93;
  wire and_tmp_70;
  wire and_dcpl_425;
  wire and_tmp_80;
  wire and_dcpl_430;
  wire and_dcpl_431;
  wire or_tmp_263;
  wire and_dcpl_433;
  wire mux_tmp_97;
  wire and_dcpl_435;
  wire mux_tmp_99;
  wire mux_tmp_100;
  wire and_dcpl_437;
  wire mux_tmp_102;
  wire mux_tmp_103;
  wire mux_tmp_104;
  wire and_dcpl_439;
  wire mux_tmp_106;
  wire mux_tmp_107;
  wire mux_tmp_108;
  wire mux_tmp_109;
  wire and_dcpl_442;
  wire mux_tmp_111;
  wire mux_tmp_112;
  wire mux_tmp_113;
  wire mux_tmp_114;
  wire mux_tmp_115;
  wire and_dcpl_445;
  wire mux_tmp_117;
  wire mux_tmp_118;
  wire mux_tmp_119;
  wire mux_tmp_120;
  wire mux_tmp_121;
  wire mux_tmp_122;
  wire and_dcpl_448;
  wire mux_tmp_124;
  wire mux_tmp_125;
  wire mux_tmp_126;
  wire mux_tmp_127;
  wire mux_tmp_128;
  wire mux_tmp_129;
  wire mux_tmp_130;
  wire and_dcpl_451;
  wire mux_tmp_132;
  wire mux_tmp_133;
  wire mux_tmp_134;
  wire mux_tmp_135;
  wire mux_tmp_136;
  wire mux_tmp_137;
  wire mux_tmp_138;
  wire mux_tmp_139;
  wire and_dcpl_454;
  wire and_tmp_89;
  wire mux_tmp_141;
  wire and_dcpl_460;
  wire and_dcpl_461;
  wire and_dcpl_462;
  wire and_dcpl_463;
  wire not_tmp_332;
  wire or_tmp_368;
  wire and_dcpl_465;
  wire and_dcpl_466;
  wire and_dcpl_467;
  wire and_tmp_90;
  wire and_dcpl_469;
  wire and_dcpl_470;
  wire and_dcpl_471;
  wire and_tmp_92;
  wire and_dcpl_473;
  wire and_dcpl_474;
  wire and_dcpl_475;
  wire and_tmp_95;
  wire and_dcpl_477;
  wire and_tmp_99;
  wire and_dcpl_480;
  wire and_tmp_103;
  wire and_dcpl_483;
  wire mux_tmp_149;
  wire and_tmp_107;
  wire and_dcpl_486;
  wire mux_tmp_152;
  wire mux_tmp_153;
  wire and_tmp_111;
  wire and_dcpl_489;
  wire mux_tmp_156;
  wire mux_tmp_157;
  wire mux_tmp_158;
  wire and_tmp_115;
  wire and_dcpl_492;
  wire and_tmp_125;
  wire and_dcpl_498;
  wire or_tmp_446;
  wire and_dcpl_500;
  wire mux_tmp_162;
  wire and_dcpl_502;
  wire mux_tmp_164;
  wire mux_tmp_165;
  wire and_dcpl_504;
  wire mux_tmp_167;
  wire mux_tmp_168;
  wire mux_tmp_169;
  wire and_dcpl_506;
  wire mux_tmp_171;
  wire mux_tmp_172;
  wire mux_tmp_173;
  wire mux_tmp_174;
  wire and_dcpl_508;
  wire mux_tmp_176;
  wire mux_tmp_177;
  wire mux_tmp_178;
  wire mux_tmp_179;
  wire mux_tmp_180;
  wire and_dcpl_510;
  wire mux_tmp_182;
  wire mux_tmp_183;
  wire mux_tmp_184;
  wire mux_tmp_185;
  wire mux_tmp_186;
  wire mux_tmp_187;
  wire and_dcpl_512;
  wire mux_tmp_189;
  wire mux_tmp_190;
  wire mux_tmp_191;
  wire mux_tmp_192;
  wire mux_tmp_193;
  wire mux_tmp_194;
  wire mux_tmp_195;
  wire and_dcpl_514;
  wire mux_tmp_197;
  wire mux_tmp_198;
  wire mux_tmp_199;
  wire mux_tmp_200;
  wire mux_tmp_201;
  wire mux_tmp_202;
  wire mux_tmp_203;
  wire mux_tmp_204;
  wire and_dcpl_516;
  wire and_tmp_134;
  wire mux_tmp_206;
  wire and_dcpl_520;
  wire and_dcpl_521;
  wire or_tmp_551;
  wire and_dcpl_523;
  wire and_dcpl_524;
  wire and_tmp_135;
  wire and_dcpl_526;
  wire and_dcpl_527;
  wire and_tmp_137;
  wire and_dcpl_529;
  wire and_dcpl_530;
  wire and_tmp_140;
  wire and_dcpl_532;
  wire and_tmp_144;
  wire and_dcpl_534;
  wire and_tmp_148;
  wire and_dcpl_536;
  wire mux_tmp_214;
  wire and_tmp_152;
  wire and_dcpl_538;
  wire mux_tmp_217;
  wire mux_tmp_218;
  wire and_tmp_156;
  wire and_dcpl_540;
  wire mux_tmp_221;
  wire mux_tmp_222;
  wire mux_tmp_223;
  wire and_tmp_160;
  wire and_dcpl_542;
  wire and_tmp_170;
  wire and_dcpl_546;
  wire or_tmp_629;
  wire and_dcpl_548;
  wire mux_tmp_227;
  wire and_dcpl_550;
  wire mux_tmp_229;
  wire mux_tmp_230;
  wire and_dcpl_552;
  wire mux_tmp_232;
  wire mux_tmp_233;
  wire mux_tmp_234;
  wire and_dcpl_554;
  wire mux_tmp_236;
  wire mux_tmp_237;
  wire mux_tmp_238;
  wire mux_tmp_239;
  wire and_dcpl_556;
  wire mux_tmp_241;
  wire mux_tmp_242;
  wire mux_tmp_243;
  wire mux_tmp_244;
  wire mux_tmp_245;
  wire and_dcpl_558;
  wire mux_tmp_247;
  wire mux_tmp_248;
  wire mux_tmp_249;
  wire mux_tmp_250;
  wire mux_tmp_251;
  wire mux_tmp_252;
  wire and_dcpl_560;
  wire mux_tmp_254;
  wire mux_tmp_255;
  wire mux_tmp_256;
  wire mux_tmp_257;
  wire mux_tmp_258;
  wire mux_tmp_259;
  wire mux_tmp_260;
  wire and_dcpl_562;
  wire mux_tmp_262;
  wire mux_tmp_263;
  wire mux_tmp_264;
  wire mux_tmp_265;
  wire mux_tmp_266;
  wire mux_tmp_267;
  wire mux_tmp_268;
  wire mux_tmp_269;
  wire and_dcpl_564;
  wire and_tmp_179;
  wire mux_tmp_271;
  wire and_dcpl_568;
  wire and_dcpl_569;
  wire and_dcpl_570;
  wire and_dcpl_571;
  wire or_tmp_733;
  wire and_dcpl_573;
  wire and_dcpl_574;
  wire and_dcpl_575;
  wire and_tmp_180;
  wire and_dcpl_577;
  wire and_dcpl_578;
  wire and_dcpl_579;
  wire and_tmp_182;
  wire and_dcpl_581;
  wire and_dcpl_582;
  wire and_dcpl_583;
  wire and_tmp_185;
  wire and_dcpl_585;
  wire and_tmp_189;
  wire and_dcpl_589;
  wire and_tmp_193;
  wire and_dcpl_593;
  wire mux_tmp_279;
  wire and_tmp_197;
  wire and_dcpl_597;
  wire mux_tmp_282;
  wire mux_tmp_283;
  wire and_tmp_201;
  wire and_dcpl_601;
  wire mux_tmp_286;
  wire mux_tmp_287;
  wire mux_tmp_288;
  wire and_tmp_205;
  wire and_dcpl_605;
  wire or_tmp_808;
  wire mux_tmp_291;
  wire mux_tmp_292;
  wire mux_tmp_293;
  wire mux_tmp_294;
  wire mux_tmp_295;
  wire mux_tmp_296;
  wire mux_tmp_297;
  wire mux_tmp_298;
  wire and_tmp_206;
  wire and_dcpl_610;
  wire or_tmp_820;
  wire and_dcpl_612;
  wire mux_tmp_301;
  wire and_dcpl_614;
  wire mux_tmp_303;
  wire mux_tmp_304;
  wire and_dcpl_616;
  wire mux_tmp_306;
  wire mux_tmp_307;
  wire mux_tmp_308;
  wire and_dcpl_618;
  wire mux_tmp_310;
  wire mux_tmp_311;
  wire mux_tmp_312;
  wire mux_tmp_313;
  wire and_dcpl_622;
  wire mux_tmp_315;
  wire mux_tmp_316;
  wire mux_tmp_317;
  wire mux_tmp_318;
  wire mux_tmp_319;
  wire and_dcpl_625;
  wire mux_tmp_321;
  wire mux_tmp_322;
  wire mux_tmp_323;
  wire mux_tmp_324;
  wire mux_tmp_325;
  wire mux_tmp_326;
  wire and_dcpl_628;
  wire mux_tmp_328;
  wire mux_tmp_329;
  wire mux_tmp_330;
  wire mux_tmp_331;
  wire mux_tmp_332;
  wire mux_tmp_333;
  wire mux_tmp_334;
  wire and_dcpl_631;
  wire mux_tmp_336;
  wire mux_tmp_337;
  wire mux_tmp_338;
  wire mux_tmp_339;
  wire mux_tmp_340;
  wire mux_tmp_341;
  wire mux_tmp_342;
  wire mux_tmp_343;
  wire and_dcpl_634;
  wire or_tmp_921;
  wire mux_tmp_345;
  wire mux_tmp_346;
  wire mux_tmp_347;
  wire mux_tmp_348;
  wire mux_tmp_349;
  wire mux_tmp_350;
  wire mux_tmp_351;
  wire mux_tmp_352;
  wire mux_tmp_353;
  wire mux_tmp_354;
  wire and_dcpl_638;
  wire and_dcpl_639;
  wire or_tmp_934;
  wire and_dcpl_641;
  wire and_dcpl_642;
  wire and_tmp_207;
  wire and_dcpl_644;
  wire and_dcpl_645;
  wire and_tmp_209;
  wire and_dcpl_647;
  wire and_dcpl_648;
  wire and_tmp_212;
  wire and_dcpl_650;
  wire and_tmp_216;
  wire and_dcpl_653;
  wire and_tmp_220;
  wire and_dcpl_657;
  wire mux_tmp_362;
  wire and_tmp_224;
  wire and_dcpl_661;
  wire mux_tmp_365;
  wire mux_tmp_366;
  wire and_tmp_228;
  wire and_dcpl_665;
  wire mux_tmp_369;
  wire mux_tmp_370;
  wire mux_tmp_371;
  wire and_tmp_232;
  wire and_dcpl_669;
  wire or_tmp_1009;
  wire mux_tmp_374;
  wire mux_tmp_375;
  wire mux_tmp_376;
  wire mux_tmp_377;
  wire mux_tmp_378;
  wire mux_tmp_379;
  wire mux_tmp_380;
  wire mux_tmp_381;
  wire and_tmp_233;
  wire and_dcpl_673;
  wire or_tmp_1021;
  wire and_dcpl_675;
  wire mux_tmp_384;
  wire and_dcpl_677;
  wire mux_tmp_386;
  wire mux_tmp_387;
  wire and_dcpl_679;
  wire mux_tmp_389;
  wire mux_tmp_390;
  wire mux_tmp_391;
  wire and_dcpl_681;
  wire mux_tmp_393;
  wire mux_tmp_394;
  wire mux_tmp_395;
  wire mux_tmp_396;
  wire and_dcpl_684;
  wire mux_tmp_398;
  wire mux_tmp_399;
  wire mux_tmp_400;
  wire mux_tmp_401;
  wire mux_tmp_402;
  wire and_dcpl_687;
  wire mux_tmp_404;
  wire mux_tmp_405;
  wire mux_tmp_406;
  wire mux_tmp_407;
  wire mux_tmp_408;
  wire mux_tmp_409;
  wire and_dcpl_690;
  wire mux_tmp_411;
  wire mux_tmp_412;
  wire mux_tmp_413;
  wire mux_tmp_414;
  wire mux_tmp_415;
  wire mux_tmp_416;
  wire mux_tmp_417;
  wire and_dcpl_693;
  wire mux_tmp_419;
  wire mux_tmp_420;
  wire mux_tmp_421;
  wire mux_tmp_422;
  wire mux_tmp_423;
  wire mux_tmp_424;
  wire mux_tmp_425;
  wire mux_tmp_426;
  wire and_dcpl_696;
  wire or_tmp_1122;
  wire mux_tmp_428;
  wire mux_tmp_429;
  wire mux_tmp_430;
  wire mux_tmp_431;
  wire mux_tmp_432;
  wire mux_tmp_433;
  wire mux_tmp_434;
  wire mux_tmp_435;
  wire mux_tmp_436;
  wire mux_tmp_437;
  reg [1:0] rem_12cyc_st_10_1_0;
  reg [1:0] rem_12cyc_st_10_3_2;
  reg [1:0] rem_12cyc_st_9_1_0;
  reg [1:0] rem_12cyc_st_9_3_2;
  reg [1:0] rem_12cyc_st_8_1_0;
  reg [1:0] rem_12cyc_st_8_3_2;
  reg [1:0] rem_12cyc_st_7_1_0;
  reg [1:0] rem_12cyc_st_7_3_2;
  reg [1:0] rem_12cyc_st_6_1_0;
  reg [1:0] rem_12cyc_st_6_3_2;
  reg [1:0] rem_12cyc_st_5_1_0;
  reg [1:0] rem_12cyc_st_5_3_2;
  reg [1:0] rem_12cyc_st_4_1_0;
  reg [1:0] rem_12cyc_st_4_3_2;
  reg [1:0] rem_12cyc_st_3_1_0;
  reg [1:0] rem_12cyc_st_3_3_2;
  reg [1:0] rem_12cyc_st_2_1_0;
  reg [1:0] rem_12cyc_st_2_3_2;
  reg [1:0] rem_12cyc_1_0;
  reg [1:0] rem_12cyc_3_2;
  reg [1:0] rem_12cyc_st_12_3_2;
  reg [63:0] result_sva_duc;
  reg [1:0] rem_12cyc_st_12_1_0;
  reg asn_itm_12;
  reg main_stage_0_13;
  reg main_stage_0_3;
  reg asn_itm_1;
  reg main_stage_0_2;
  reg main_stage_0_4;
  reg asn_itm_2;
  reg main_stage_0_5;
  reg asn_itm_3;
  reg main_stage_0_6;
  reg asn_itm_4;
  reg asn_itm_5;
  reg main_stage_0_8;
  reg asn_itm_7;
  reg main_stage_0_9;
  reg asn_itm_8;
  reg main_stage_0_10;
  reg asn_itm_9;
  reg main_stage_0_7;
  reg asn_itm_6;
  reg main_stage_0_11;
  reg asn_itm_10;
  wire and_1173_cse;
  wire and_1175_cse;
  wire and_1177_cse;
  wire and_1179_cse;
  wire and_1181_cse;
  wire and_1183_cse;
  wire and_1185_cse;
  wire and_1187_cse;
  wire and_1189_cse;
  wire and_1191_cse;
  wire and_1193_cse;
  wire and_1195_cse;
  wire and_1197_cse;
  wire or_1_cse;
  wire or_6_cse;
  wire or_10_cse;
  wire or_15_cse;
  wire or_21_cse;
  wire or_28_cse;
  wire or_37_cse;
  wire or_48_cse;
  wire or_83_cse;
  wire nand_276_cse;
  wire or_88_cse;
  wire nand_274_cse;
  wire or_93_cse;
  wire nand_271_cse;
  wire or_100_cse;
  wire nand_267_cse;
  wire or_109_cse;
  wire or_120_cse;
  wire or_133_cse;
  wire or_148_cse;
  wire or_190_cse;
  wire or_195_cse;
  wire or_199_cse;
  wire or_204_cse;
  wire or_210_cse;
  wire or_217_cse;
  wire or_226_cse;
  wire or_237_cse;
  wire or_270_cse;
  wire or_275_cse;
  wire or_280_cse;
  wire or_287_cse;
  wire or_296_cse;
  wire or_307_cse;
  wire or_320_cse;
  wire or_335_cse;
  wire nand_281_cse;
  wire or_377_cse;
  wire or_382_cse;
  wire or_386_cse;
  wire or_391_cse;
  wire or_397_cse;
  wire nand_215_cse;
  wire or_404_cse;
  wire nand_212_cse;
  wire or_413_cse;
  wire nand_208_cse;
  wire or_424_cse;
  wire or_458_cse;
  wire or_463_cse;
  wire nand_198_cse;
  wire or_468_cse;
  wire or_475_cse;
  wire nand_189_cse;
  wire or_484_cse;
  wire or_495_cse;
  wire or_508_cse;
  wire nand_203_cse;
  wire or_523_cse;
  wire nand_250_cse;
  wire or_564_cse;
  wire or_569_cse;
  wire or_573_cse;
  wire or_578_cse;
  wire or_584_cse;
  wire or_591_cse;
  wire or_600_cse;
  wire or_611_cse;
  wire or_643_cse;
  wire or_648_cse;
  wire or_653_cse;
  wire or_660_cse;
  wire or_669_cse;
  wire or_680_cse;
  wire or_693_cse;
  wire or_708_cse;
  wire or_748_cse;
  wire or_753_cse;
  wire or_757_cse;
  wire or_762_cse;
  wire or_768_cse;
  wire or_775_cse;
  wire or_784_cse;
  wire or_795_cse;
  wire or_837_cse;
  wire nand_84_cse;
  wire or_842_cse;
  wire or_847_cse;
  wire nand_79_cse;
  wire or_854_cse;
  wire or_863_cse;
  wire or_874_cse;
  wire or_887_cse;
  wire or_902_cse;
  wire or_952_cse;
  wire or_957_cse;
  wire or_961_cse;
  wire or_966_cse;
  wire or_972_cse;
  wire or_979_cse;
  wire or_988_cse;
  wire or_999_cse;
  wire nand_57_cse;
  wire or_1045_cse;
  wire or_1050_cse;
  wire or_1057_cse;
  wire or_1066_cse;
  wire nand_36_cse;
  wire nand_29_cse;
  wire nand_21_cse;
  wire nand_222_cse;
  wire nand_223_cse;
  reg main_stage_0_12;
  reg [63:0] m_buf_sva_1;
  reg [63:0] m_buf_sva_2;
  reg [63:0] m_buf_sva_3;
  reg [63:0] m_buf_sva_4;
  reg [63:0] m_buf_sva_5;
  reg [63:0] m_buf_sva_6;
  reg [63:0] m_buf_sva_7;
  reg [63:0] m_buf_sva_8;
  reg [63:0] m_buf_sva_9;
  reg [63:0] m_buf_sva_10;
  reg [63:0] m_buf_sva_11;
  reg [63:0] m_buf_sva_12;
  reg asn_itm_11;
  reg [63:0] mut_2_63_0;
  reg [63:0] mut_3_63_0;
  reg [63:0] mut_4_63_0;
  reg [63:0] mut_5_63_0;
  reg [63:0] mut_6_63_0;
  reg [63:0] mut_7_63_0;
  reg [63:0] mut_8_63_0;
  reg [63:0] mut_9_63_0;
  reg [63:0] mut_10_63_0;
  reg [63:0] mut_11_63_0;
  reg [63:0] mut_1_2_63_0;
  reg [63:0] mut_1_3_63_0;
  reg [63:0] mut_1_4_63_0;
  reg [63:0] mut_1_5_63_0;
  reg [63:0] mut_1_6_63_0;
  reg [63:0] mut_1_7_63_0;
  reg [63:0] mut_1_8_63_0;
  reg [63:0] mut_1_9_63_0;
  reg [63:0] mut_1_10_63_0;
  reg [63:0] mut_1_11_63_0;
  reg [63:0] mut_2_2_63_0;
  reg [63:0] mut_2_3_63_0;
  reg [63:0] mut_2_4_63_0;
  reg [63:0] mut_2_5_63_0;
  reg [63:0] mut_2_6_63_0;
  reg [63:0] mut_2_7_63_0;
  reg [63:0] mut_2_8_63_0;
  reg [63:0] mut_2_9_63_0;
  reg [63:0] mut_2_10_63_0;
  reg [63:0] mut_2_11_63_0;
  reg [63:0] mut_3_2_63_0;
  reg [63:0] mut_3_3_63_0;
  reg [63:0] mut_3_4_63_0;
  reg [63:0] mut_3_5_63_0;
  reg [63:0] mut_3_6_63_0;
  reg [63:0] mut_3_7_63_0;
  reg [63:0] mut_3_8_63_0;
  reg [63:0] mut_3_9_63_0;
  reg [63:0] mut_3_10_63_0;
  reg [63:0] mut_3_11_63_0;
  reg [63:0] mut_4_2_63_0;
  reg [63:0] mut_4_3_63_0;
  reg [63:0] mut_4_4_63_0;
  reg [63:0] mut_4_5_63_0;
  reg [63:0] mut_4_6_63_0;
  reg [63:0] mut_4_7_63_0;
  reg [63:0] mut_4_8_63_0;
  reg [63:0] mut_4_9_63_0;
  reg [63:0] mut_4_10_63_0;
  reg [63:0] mut_4_11_63_0;
  reg [63:0] mut_5_2_63_0;
  reg [63:0] mut_5_3_63_0;
  reg [63:0] mut_5_4_63_0;
  reg [63:0] mut_5_5_63_0;
  reg [63:0] mut_5_6_63_0;
  reg [63:0] mut_5_7_63_0;
  reg [63:0] mut_5_8_63_0;
  reg [63:0] mut_5_9_63_0;
  reg [63:0] mut_5_10_63_0;
  reg [63:0] mut_5_11_63_0;
  reg [63:0] mut_6_2_63_0;
  reg [63:0] mut_6_3_63_0;
  reg [63:0] mut_6_4_63_0;
  reg [63:0] mut_6_5_63_0;
  reg [63:0] mut_6_6_63_0;
  reg [63:0] mut_6_7_63_0;
  reg [63:0] mut_6_8_63_0;
  reg [63:0] mut_6_9_63_0;
  reg [63:0] mut_6_10_63_0;
  reg [63:0] mut_6_11_63_0;
  reg [63:0] mut_7_2_63_0;
  reg [63:0] mut_7_3_63_0;
  reg [63:0] mut_7_4_63_0;
  reg [63:0] mut_7_5_63_0;
  reg [63:0] mut_7_6_63_0;
  reg [63:0] mut_7_7_63_0;
  reg [63:0] mut_7_8_63_0;
  reg [63:0] mut_7_9_63_0;
  reg [63:0] mut_7_10_63_0;
  reg [63:0] mut_7_11_63_0;
  reg [63:0] mut_8_2_63_0;
  reg [63:0] mut_8_3_63_0;
  reg [63:0] mut_8_4_63_0;
  reg [63:0] mut_8_5_63_0;
  reg [63:0] mut_8_6_63_0;
  reg [63:0] mut_8_7_63_0;
  reg [63:0] mut_8_8_63_0;
  reg [63:0] mut_8_9_63_0;
  reg [63:0] mut_8_10_63_0;
  reg [63:0] mut_8_11_63_0;
  reg [63:0] mut_9_2_63_0;
  reg [63:0] mut_9_3_63_0;
  reg [63:0] mut_9_4_63_0;
  reg [63:0] mut_9_5_63_0;
  reg [63:0] mut_9_6_63_0;
  reg [63:0] mut_9_7_63_0;
  reg [63:0] mut_9_8_63_0;
  reg [63:0] mut_9_9_63_0;
  reg [63:0] mut_9_10_63_0;
  reg [63:0] mut_9_11_63_0;
  reg [63:0] mut_10_2_63_0;
  reg [63:0] mut_10_3_63_0;
  reg [63:0] mut_10_4_63_0;
  reg [63:0] mut_10_5_63_0;
  reg [63:0] mut_10_6_63_0;
  reg [63:0] mut_10_7_63_0;
  reg [63:0] mut_10_8_63_0;
  reg [63:0] mut_10_9_63_0;
  reg [63:0] mut_10_10_63_0;
  reg [63:0] mut_10_11_63_0;
  reg [63:0] mut_11_2_63_0;
  reg [63:0] mut_11_3_63_0;
  reg [63:0] mut_11_4_63_0;
  reg [63:0] mut_11_5_63_0;
  reg [63:0] mut_11_6_63_0;
  reg [63:0] mut_11_7_63_0;
  reg [63:0] mut_11_8_63_0;
  reg [63:0] mut_11_9_63_0;
  reg [63:0] mut_11_10_63_0;
  reg [63:0] mut_11_11_63_0;
  reg [63:0] mut_12_2_63_0;
  reg [63:0] mut_12_3_63_0;
  reg [63:0] mut_12_4_63_0;
  reg [63:0] mut_12_5_63_0;
  reg [63:0] mut_12_6_63_0;
  reg [63:0] mut_12_7_63_0;
  reg [63:0] mut_12_8_63_0;
  reg [63:0] mut_12_9_63_0;
  reg [63:0] mut_12_10_63_0;
  reg [63:0] mut_12_11_63_0;
  reg [63:0] mut_13_2_63_0;
  reg [63:0] mut_13_3_63_0;
  reg [63:0] mut_13_4_63_0;
  reg [63:0] mut_13_5_63_0;
  reg [63:0] mut_13_6_63_0;
  reg [63:0] mut_13_7_63_0;
  reg [63:0] mut_13_8_63_0;
  reg [63:0] mut_13_9_63_0;
  reg [63:0] mut_13_10_63_0;
  reg [63:0] mut_13_11_63_0;
  reg [63:0] mut_14_2_63_0;
  reg [63:0] mut_14_3_63_0;
  reg [63:0] mut_14_4_63_0;
  reg [63:0] mut_14_5_63_0;
  reg [63:0] mut_14_6_63_0;
  reg [63:0] mut_14_7_63_0;
  reg [63:0] mut_14_8_63_0;
  reg [63:0] mut_14_9_63_0;
  reg [63:0] mut_14_10_63_0;
  reg [63:0] mut_14_11_63_0;
  reg [63:0] mut_15_2_63_0;
  reg [63:0] mut_15_3_63_0;
  reg [63:0] mut_15_4_63_0;
  reg [63:0] mut_15_5_63_0;
  reg [63:0] mut_15_6_63_0;
  reg [63:0] mut_15_7_63_0;
  reg [63:0] mut_15_8_63_0;
  reg [63:0] mut_15_9_63_0;
  reg [63:0] mut_15_10_63_0;
  reg [63:0] mut_15_11_63_0;
  reg [63:0] mut_16_2_63_0;
  reg [63:0] mut_16_3_63_0;
  reg [63:0] mut_16_4_63_0;
  reg [63:0] mut_16_5_63_0;
  reg [63:0] mut_16_6_63_0;
  reg [63:0] mut_16_7_63_0;
  reg [63:0] mut_16_8_63_0;
  reg [63:0] mut_16_9_63_0;
  reg [63:0] mut_16_10_63_0;
  reg [63:0] mut_16_11_63_0;
  reg [63:0] mut_17_2_63_0;
  reg [63:0] mut_17_3_63_0;
  reg [63:0] mut_17_4_63_0;
  reg [63:0] mut_17_5_63_0;
  reg [63:0] mut_17_6_63_0;
  reg [63:0] mut_17_7_63_0;
  reg [63:0] mut_17_8_63_0;
  reg [63:0] mut_17_9_63_0;
  reg [63:0] mut_17_10_63_0;
  reg [63:0] mut_17_11_63_0;
  reg [63:0] mut_18_2_63_0;
  reg [63:0] mut_18_3_63_0;
  reg [63:0] mut_18_4_63_0;
  reg [63:0] mut_18_5_63_0;
  reg [63:0] mut_18_6_63_0;
  reg [63:0] mut_18_7_63_0;
  reg [63:0] mut_18_8_63_0;
  reg [63:0] mut_18_9_63_0;
  reg [63:0] mut_18_10_63_0;
  reg [63:0] mut_18_11_63_0;
  reg [63:0] mut_19_2_63_0;
  reg [63:0] mut_19_3_63_0;
  reg [63:0] mut_19_4_63_0;
  reg [63:0] mut_19_5_63_0;
  reg [63:0] mut_19_6_63_0;
  reg [63:0] mut_19_7_63_0;
  reg [63:0] mut_19_8_63_0;
  reg [63:0] mut_19_9_63_0;
  reg [63:0] mut_19_10_63_0;
  reg [63:0] mut_19_11_63_0;
  reg [63:0] mut_20_2_63_0;
  reg [63:0] mut_20_3_63_0;
  reg [63:0] mut_20_4_63_0;
  reg [63:0] mut_20_5_63_0;
  reg [63:0] mut_20_6_63_0;
  reg [63:0] mut_20_7_63_0;
  reg [63:0] mut_20_8_63_0;
  reg [63:0] mut_20_9_63_0;
  reg [63:0] mut_20_10_63_0;
  reg [63:0] mut_20_11_63_0;
  reg [63:0] mut_21_2_63_0;
  reg [63:0] mut_21_3_63_0;
  reg [63:0] mut_21_4_63_0;
  reg [63:0] mut_21_5_63_0;
  reg [63:0] mut_21_6_63_0;
  reg [63:0] mut_21_7_63_0;
  reg [63:0] mut_21_8_63_0;
  reg [63:0] mut_21_9_63_0;
  reg [63:0] mut_21_10_63_0;
  reg [63:0] mut_21_11_63_0;
  reg [63:0] mut_22_2_63_0;
  reg [63:0] mut_22_3_63_0;
  reg [63:0] mut_22_4_63_0;
  reg [63:0] mut_22_5_63_0;
  reg [63:0] mut_22_6_63_0;
  reg [63:0] mut_22_7_63_0;
  reg [63:0] mut_22_8_63_0;
  reg [63:0] mut_22_9_63_0;
  reg [63:0] mut_22_10_63_0;
  reg [63:0] mut_22_11_63_0;
  reg [63:0] mut_23_2_63_0;
  reg [63:0] mut_23_3_63_0;
  reg [63:0] mut_23_4_63_0;
  reg [63:0] mut_23_5_63_0;
  reg [63:0] mut_23_6_63_0;
  reg [63:0] mut_23_7_63_0;
  reg [63:0] mut_23_8_63_0;
  reg [63:0] mut_23_9_63_0;
  reg [63:0] mut_23_10_63_0;
  reg [63:0] mut_23_11_63_0;
  reg [1:0] rem_12cyc_st_11_3_2;
  reg [1:0] rem_12cyc_st_11_1_0;
  wire [63:0] result_sva_duc_mx0;
  wire and_1203_cse;
  wire and_1205_cse;
  wire and_1207_cse;
  wire and_1209_cse;
  wire and_1211_cse;
  wire and_1213_cse;
  wire and_1215_cse;
  wire and_1217_cse;
  wire and_1219_cse;
  wire and_1221_cse;
  wire and_1223_cse;
  wire and_1225_cse;
  wire and_1227_cse;
  wire and_1229_cse;
  wire and_1231_cse;
  wire and_1233_cse;
  wire and_1235_cse;
  wire and_1237_cse;
  wire and_1239_cse;
  wire and_1241_cse;
  wire and_1243_cse;
  wire and_1245_cse;
  wire and_1247_cse;
  wire and_1249_cse;
  wire and_1251_cse;
  wire and_1253_cse;
  wire and_1255_cse;
  wire and_1257_cse;
  wire and_1259_cse;
  wire and_1261_cse;
  wire and_1263_cse;
  wire and_1265_cse;
  wire and_1267_cse;
  wire and_1269_cse;
  wire and_1271_cse;
  wire and_1273_cse;
  wire and_1275_cse;
  wire and_1277_cse;
  wire and_1279_cse;
  wire and_1281_cse;
  wire and_1283_cse;
  wire and_1285_cse;
  wire and_1287_cse;
  wire and_1289_cse;
  wire and_1291_cse;
  wire and_1293_cse;
  wire and_1295_cse;
  wire and_1297_cse;
  wire and_1299_cse;
  wire and_1301_cse;
  wire and_1303_cse;
  wire and_1305_cse;
  wire and_1307_cse;
  wire and_1309_cse;
  wire and_1311_cse;
  wire and_1313_cse;
  wire and_1315_cse;
  wire and_1317_cse;
  wire and_1319_cse;
  wire and_1321_cse;
  wire and_1323_cse;
  wire and_1325_cse;
  wire and_1327_cse;
  wire and_1329_cse;
  wire and_1331_cse;
  wire and_1333_cse;
  wire and_1335_cse;
  wire and_1337_cse;
  wire and_1339_cse;
  wire and_1341_cse;
  wire and_1343_cse;
  wire and_1345_cse;
  wire and_1347_cse;
  wire and_1349_cse;
  wire and_1351_cse;
  wire and_1353_cse;
  wire and_1355_cse;
  wire and_1357_cse;
  wire and_1359_cse;
  wire and_1361_cse;
  wire and_1363_cse;
  wire and_1365_cse;
  wire and_1367_cse;
  wire and_1369_cse;
  wire and_1371_cse;
  wire and_1373_cse;
  wire and_1375_cse;
  wire and_1377_cse;
  wire and_1379_cse;
  wire and_1381_cse;
  wire and_1383_cse;
  wire and_1385_cse;
  wire and_1387_cse;
  wire and_1389_cse;
  wire and_1391_cse;
  wire and_1393_cse;
  wire and_1395_cse;
  wire and_1397_cse;
  wire and_1399_cse;
  wire and_1401_cse;
  wire and_1403_cse;
  wire and_1405_cse;
  wire and_1407_cse;
  wire and_1409_cse;
  wire and_1411_cse;
  wire and_1413_cse;
  wire and_1415_cse;
  wire and_1417_cse;
  wire and_1419_cse;
  wire and_1421_cse;
  wire and_1423_cse;
  wire and_1425_cse;
  wire and_1427_cse;
  wire and_1429_cse;
  wire and_1431_cse;
  wire and_1433_cse;
  wire and_1435_cse;
  wire and_1437_cse;
  wire and_1439_cse;
  wire and_1441_cse;
  wire and_1443_cse;
  wire and_1445_cse;
  wire and_1447_cse;
  wire and_1449_cse;
  wire and_1451_cse;
  wire and_1453_cse;
  wire and_1455_cse;
  wire and_1457_cse;
  wire and_1459_cse;
  wire and_1461_cse;
  wire and_1463_cse;

  wire[63:0] qelse_acc_nl;
  wire[64:0] nl_qelse_acc_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] mux_12_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] mux_7_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] mux_3_nl;
  wire[0:0] mux_2_nl;
  wire[0:0] and_273_nl;
  wire[0:0] and_275_nl;
  wire[0:0] and_277_nl;
  wire[0:0] and_279_nl;
  wire[0:0] and_281_nl;
  wire[0:0] and_282_nl;
  wire[0:0] and_283_nl;
  wire[0:0] and_284_nl;
  wire[0:0] and_286_nl;
  wire[0:0] and_287_nl;
  wire[0:0] and_288_nl;
  wire[0:0] and_289_nl;
  wire[0:0] and_290_nl;
  wire[0:0] xor_nl;
  wire[0:0] nor_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] nor_518_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] nor_517_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] nor_516_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] nor_515_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] nor_514_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] nor_512_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] nor_513_nl;
  wire[0:0] nor_509_nl;
  wire[0:0] mux_22_nl;
  wire[0:0] nor_510_nl;
  wire[0:0] mux_23_nl;
  wire[0:0] nor_511_nl;
  wire[0:0] nor_505_nl;
  wire[0:0] nor_506_nl;
  wire[0:0] mux_26_nl;
  wire[0:0] nor_507_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] nor_508_nl;
  wire[0:0] nor_500_nl;
  wire[0:0] or_61_nl;
  wire[0:0] nor_501_nl;
  wire[0:0] nor_502_nl;
  wire[0:0] mux_31_nl;
  wire[0:0] nor_503_nl;
  wire[0:0] mux_32_nl;
  wire[0:0] nor_504_nl;
  wire[0:0] mux_33_nl;
  wire[0:0] nor_499_nl;
  wire[0:0] and_1168_nl;
  wire[0:0] mux_35_nl;
  wire[0:0] nor_498_nl;
  wire[0:0] and_1166_nl;
  wire[0:0] and_1167_nl;
  wire[0:0] mux_38_nl;
  wire[0:0] nor_497_nl;
  wire[0:0] and_1163_nl;
  wire[0:0] and_1164_nl;
  wire[0:0] and_1165_nl;
  wire[0:0] mux_42_nl;
  wire[0:0] nor_496_nl;
  wire[0:0] and_1159_nl;
  wire[0:0] and_1160_nl;
  wire[0:0] and_1161_nl;
  wire[0:0] and_1162_nl;
  wire[0:0] mux_47_nl;
  wire[0:0] nor_495_nl;
  wire[0:0] nor_493_nl;
  wire[0:0] and_1155_nl;
  wire[0:0] and_1156_nl;
  wire[0:0] and_1157_nl;
  wire[0:0] and_1158_nl;
  wire[0:0] mux_53_nl;
  wire[0:0] nor_494_nl;
  wire[0:0] nor_490_nl;
  wire[0:0] nor_491_nl;
  wire[0:0] and_1151_nl;
  wire[0:0] and_1152_nl;
  wire[0:0] and_1153_nl;
  wire[0:0] and_1154_nl;
  wire[0:0] mux_60_nl;
  wire[0:0] nor_492_nl;
  wire[0:0] nor_486_nl;
  wire[0:0] nor_487_nl;
  wire[0:0] nor_488_nl;
  wire[0:0] and_1147_nl;
  wire[0:0] and_1148_nl;
  wire[0:0] and_1149_nl;
  wire[0:0] and_1150_nl;
  wire[0:0] mux_68_nl;
  wire[0:0] nor_489_nl;
  wire[0:0] nor_481_nl;
  wire[0:0] or_165_nl;
  wire[0:0] nor_482_nl;
  wire[0:0] nor_483_nl;
  wire[0:0] nor_484_nl;
  wire[0:0] and_1143_nl;
  wire[0:0] and_1144_nl;
  wire[0:0] and_1145_nl;
  wire[0:0] and_1146_nl;
  wire[0:0] mux_77_nl;
  wire[0:0] nor_485_nl;
  wire[0:0] nor_480_nl;
  wire[0:0] or_175_nl;
  wire[0:0] mux_79_nl;
  wire[0:0] nor_479_nl;
  wire[0:0] mux_80_nl;
  wire[0:0] nor_478_nl;
  wire[0:0] mux_81_nl;
  wire[0:0] nor_477_nl;
  wire[0:0] mux_82_nl;
  wire[0:0] nor_476_nl;
  wire[0:0] mux_83_nl;
  wire[0:0] nor_475_nl;
  wire[0:0] mux_84_nl;
  wire[0:0] nor_473_nl;
  wire[0:0] mux_85_nl;
  wire[0:0] nor_474_nl;
  wire[0:0] nor_470_nl;
  wire[0:0] mux_87_nl;
  wire[0:0] nor_471_nl;
  wire[0:0] mux_88_nl;
  wire[0:0] nor_472_nl;
  wire[0:0] nor_466_nl;
  wire[0:0] nor_467_nl;
  wire[0:0] mux_91_nl;
  wire[0:0] nor_468_nl;
  wire[0:0] mux_92_nl;
  wire[0:0] nor_469_nl;
  wire[0:0] nor_461_nl;
  wire[0:0] or_250_nl;
  wire[0:0] nor_462_nl;
  wire[0:0] nor_463_nl;
  wire[0:0] mux_96_nl;
  wire[0:0] nor_464_nl;
  wire[0:0] mux_97_nl;
  wire[0:0] nor_465_nl;
  wire[0:0] mux_98_nl;
  wire[0:0] nor_460_nl;
  wire[0:0] and_1142_nl;
  wire[0:0] mux_100_nl;
  wire[0:0] nor_459_nl;
  wire[0:0] and_1140_nl;
  wire[0:0] and_1141_nl;
  wire[0:0] mux_103_nl;
  wire[0:0] nor_458_nl;
  wire[0:0] and_1137_nl;
  wire[0:0] and_1138_nl;
  wire[0:0] and_1139_nl;
  wire[0:0] mux_107_nl;
  wire[0:0] nor_457_nl;
  wire[0:0] and_1133_nl;
  wire[0:0] and_1134_nl;
  wire[0:0] and_1135_nl;
  wire[0:0] and_1136_nl;
  wire[0:0] mux_112_nl;
  wire[0:0] nor_456_nl;
  wire[0:0] nor_454_nl;
  wire[0:0] and_1129_nl;
  wire[0:0] and_1130_nl;
  wire[0:0] and_1131_nl;
  wire[0:0] and_1132_nl;
  wire[0:0] mux_118_nl;
  wire[0:0] nor_455_nl;
  wire[0:0] nor_451_nl;
  wire[0:0] nor_452_nl;
  wire[0:0] and_1125_nl;
  wire[0:0] and_1126_nl;
  wire[0:0] and_1127_nl;
  wire[0:0] and_1128_nl;
  wire[0:0] mux_125_nl;
  wire[0:0] nor_453_nl;
  wire[0:0] nor_447_nl;
  wire[0:0] nor_448_nl;
  wire[0:0] nor_449_nl;
  wire[0:0] and_1121_nl;
  wire[0:0] and_1122_nl;
  wire[0:0] and_1123_nl;
  wire[0:0] and_1124_nl;
  wire[0:0] mux_133_nl;
  wire[0:0] nor_450_nl;
  wire[0:0] nor_442_nl;
  wire[0:0] or_352_nl;
  wire[0:0] nor_443_nl;
  wire[0:0] nor_444_nl;
  wire[0:0] nor_445_nl;
  wire[0:0] and_1117_nl;
  wire[0:0] and_1118_nl;
  wire[0:0] and_1119_nl;
  wire[0:0] and_1120_nl;
  wire[0:0] mux_142_nl;
  wire[0:0] nor_446_nl;
  wire[0:0] and_1116_nl;
  wire[0:0] or_362_nl;
  wire[0:0] mux_144_nl;
  wire[0:0] and_1172_nl;
  wire[0:0] mux_145_nl;
  wire[0:0] and_1114_nl;
  wire[0:0] mux_146_nl;
  wire[0:0] and_1113_nl;
  wire[0:0] mux_147_nl;
  wire[0:0] and_1112_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] and_1111_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] and_1109_nl;
  wire[0:0] mux_150_nl;
  wire[0:0] and_1110_nl;
  wire[0:0] and_1106_nl;
  wire[0:0] mux_152_nl;
  wire[0:0] and_1107_nl;
  wire[0:0] mux_153_nl;
  wire[0:0] and_1108_nl;
  wire[0:0] and_1102_nl;
  wire[0:0] and_1103_nl;
  wire[0:0] mux_156_nl;
  wire[0:0] and_1104_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] and_1105_nl;
  wire[0:0] and_1097_nl;
  wire[0:0] or_437_nl;
  wire[0:0] and_1098_nl;
  wire[0:0] and_1099_nl;
  wire[0:0] mux_161_nl;
  wire[0:0] and_1100_nl;
  wire[0:0] mux_162_nl;
  wire[0:0] and_1101_nl;
  wire[0:0] mux_163_nl;
  wire[0:0] and_1171_nl;
  wire[0:0] and_1094_nl;
  wire[0:0] mux_165_nl;
  wire[0:0] and_1095_nl;
  wire[0:0] and_1091_nl;
  wire[0:0] and_1092_nl;
  wire[0:0] mux_168_nl;
  wire[0:0] and_1093_nl;
  wire[0:0] and_1087_nl;
  wire[0:0] and_1088_nl;
  wire[0:0] and_1089_nl;
  wire[0:0] mux_172_nl;
  wire[0:0] and_1090_nl;
  wire[0:0] and_1082_nl;
  wire[0:0] and_1083_nl;
  wire[0:0] and_1084_nl;
  wire[0:0] and_1085_nl;
  wire[0:0] mux_177_nl;
  wire[0:0] and_1086_nl;
  wire[0:0] and_1076_nl;
  wire[0:0] and_1077_nl;
  wire[0:0] and_1078_nl;
  wire[0:0] and_1079_nl;
  wire[0:0] and_1080_nl;
  wire[0:0] mux_183_nl;
  wire[0:0] and_1081_nl;
  wire[0:0] and_1069_nl;
  wire[0:0] and_1070_nl;
  wire[0:0] and_1071_nl;
  wire[0:0] and_1072_nl;
  wire[0:0] and_1073_nl;
  wire[0:0] and_1074_nl;
  wire[0:0] mux_190_nl;
  wire[0:0] and_1075_nl;
  wire[0:0] and_1061_nl;
  wire[0:0] and_1062_nl;
  wire[0:0] and_1063_nl;
  wire[0:0] and_1064_nl;
  wire[0:0] and_1065_nl;
  wire[0:0] and_1066_nl;
  wire[0:0] and_1067_nl;
  wire[0:0] mux_198_nl;
  wire[0:0] and_1068_nl;
  wire[0:0] and_1052_nl;
  wire[0:0] or_540_nl;
  wire[0:0] and_1053_nl;
  wire[0:0] and_1054_nl;
  wire[0:0] and_1055_nl;
  wire[0:0] and_1056_nl;
  wire[0:0] and_1057_nl;
  wire[0:0] and_1058_nl;
  wire[0:0] and_1059_nl;
  wire[0:0] mux_207_nl;
  wire[0:0] and_1060_nl;
  wire[0:0] nor_439_nl;
  wire[0:0] or_550_nl;
  wire[0:0] mux_209_nl;
  wire[0:0] and_1170_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] and_1050_nl;
  wire[0:0] mux_211_nl;
  wire[0:0] and_1049_nl;
  wire[0:0] mux_212_nl;
  wire[0:0] and_1048_nl;
  wire[0:0] mux_213_nl;
  wire[0:0] and_1047_nl;
  wire[0:0] mux_214_nl;
  wire[0:0] and_1045_nl;
  wire[0:0] mux_215_nl;
  wire[0:0] and_1046_nl;
  wire[0:0] and_1042_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] and_1043_nl;
  wire[0:0] mux_218_nl;
  wire[0:0] and_1044_nl;
  wire[0:0] and_1038_nl;
  wire[0:0] and_1039_nl;
  wire[0:0] mux_221_nl;
  wire[0:0] and_1040_nl;
  wire[0:0] mux_222_nl;
  wire[0:0] and_1041_nl;
  wire[0:0] and_1033_nl;
  wire[0:0] or_624_nl;
  wire[0:0] and_1034_nl;
  wire[0:0] and_1035_nl;
  wire[0:0] mux_226_nl;
  wire[0:0] and_1036_nl;
  wire[0:0] mux_227_nl;
  wire[0:0] and_1037_nl;
  wire[0:0] mux_228_nl;
  wire[0:0] and_1169_nl;
  wire[0:0] and_1030_nl;
  wire[0:0] mux_230_nl;
  wire[0:0] and_1031_nl;
  wire[0:0] and_1027_nl;
  wire[0:0] and_1028_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] and_1029_nl;
  wire[0:0] and_1023_nl;
  wire[0:0] and_1024_nl;
  wire[0:0] and_1025_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] and_1026_nl;
  wire[0:0] and_1018_nl;
  wire[0:0] and_1019_nl;
  wire[0:0] and_1020_nl;
  wire[0:0] and_1021_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] and_1022_nl;
  wire[0:0] and_1012_nl;
  wire[0:0] and_1013_nl;
  wire[0:0] and_1014_nl;
  wire[0:0] and_1015_nl;
  wire[0:0] and_1016_nl;
  wire[0:0] mux_248_nl;
  wire[0:0] and_1017_nl;
  wire[0:0] and_1005_nl;
  wire[0:0] and_1006_nl;
  wire[0:0] and_1007_nl;
  wire[0:0] and_1008_nl;
  wire[0:0] and_1009_nl;
  wire[0:0] and_1010_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] and_1011_nl;
  wire[0:0] and_997_nl;
  wire[0:0] and_998_nl;
  wire[0:0] and_999_nl;
  wire[0:0] and_1000_nl;
  wire[0:0] and_1001_nl;
  wire[0:0] and_1002_nl;
  wire[0:0] and_1003_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] and_1004_nl;
  wire[0:0] and_988_nl;
  wire[0:0] or_725_nl;
  wire[0:0] and_989_nl;
  wire[0:0] and_990_nl;
  wire[0:0] and_991_nl;
  wire[0:0] and_992_nl;
  wire[0:0] and_993_nl;
  wire[0:0] and_994_nl;
  wire[0:0] and_995_nl;
  wire[0:0] mux_272_nl;
  wire[0:0] and_996_nl;
  wire[0:0] and_987_nl;
  wire[0:0] or_735_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] nor_436_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] nor_435_nl;
  wire[0:0] mux_276_nl;
  wire[0:0] nor_434_nl;
  wire[0:0] mux_277_nl;
  wire[0:0] nor_433_nl;
  wire[0:0] mux_278_nl;
  wire[0:0] nor_432_nl;
  wire[0:0] mux_279_nl;
  wire[0:0] nor_430_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] nor_431_nl;
  wire[0:0] nor_427_nl;
  wire[0:0] mux_282_nl;
  wire[0:0] nor_428_nl;
  wire[0:0] mux_283_nl;
  wire[0:0] nor_429_nl;
  wire[0:0] nor_423_nl;
  wire[0:0] nor_424_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] nor_425_nl;
  wire[0:0] mux_287_nl;
  wire[0:0] nor_426_nl;
  wire[0:0] nor_418_nl;
  wire[0:0] or_808_nl;
  wire[0:0] nor_419_nl;
  wire[0:0] nor_420_nl;
  wire[0:0] mux_291_nl;
  wire[0:0] nor_421_nl;
  wire[0:0] mux_292_nl;
  wire[0:0] nor_422_nl;
  wire[0:0] nor_409_nl;
  wire[0:0] or_823_nl;
  wire[0:0] nor_410_nl;
  wire[0:0] or_822_nl;
  wire[0:0] nor_411_nl;
  wire[0:0] or_821_nl;
  wire[0:0] nor_412_nl;
  wire[0:0] or_820_nl;
  wire[0:0] nor_413_nl;
  wire[0:0] or_819_nl;
  wire[0:0] nor_414_nl;
  wire[0:0] or_818_nl;
  wire[0:0] nor_415_nl;
  wire[0:0] or_817_nl;
  wire[0:0] nor_416_nl;
  wire[0:0] or_816_nl;
  wire[0:0] mux_301_nl;
  wire[0:0] nor_417_nl;
  wire[0:0] or_815_nl;
  wire[0:0] mux_302_nl;
  wire[0:0] nor_408_nl;
  wire[0:0] and_986_nl;
  wire[0:0] mux_304_nl;
  wire[0:0] nor_407_nl;
  wire[0:0] and_984_nl;
  wire[0:0] and_985_nl;
  wire[0:0] mux_307_nl;
  wire[0:0] nor_406_nl;
  wire[0:0] and_981_nl;
  wire[0:0] and_982_nl;
  wire[0:0] and_983_nl;
  wire[0:0] mux_311_nl;
  wire[0:0] nor_405_nl;
  wire[0:0] and_977_nl;
  wire[0:0] and_978_nl;
  wire[0:0] and_979_nl;
  wire[0:0] and_980_nl;
  wire[0:0] mux_316_nl;
  wire[0:0] nor_404_nl;
  wire[0:0] nor_402_nl;
  wire[0:0] and_973_nl;
  wire[0:0] and_974_nl;
  wire[0:0] and_975_nl;
  wire[0:0] and_976_nl;
  wire[0:0] mux_322_nl;
  wire[0:0] nor_403_nl;
  wire[0:0] nor_399_nl;
  wire[0:0] nor_400_nl;
  wire[0:0] and_969_nl;
  wire[0:0] and_970_nl;
  wire[0:0] and_971_nl;
  wire[0:0] and_972_nl;
  wire[0:0] mux_329_nl;
  wire[0:0] nor_401_nl;
  wire[0:0] nor_395_nl;
  wire[0:0] nor_396_nl;
  wire[0:0] nor_397_nl;
  wire[0:0] and_965_nl;
  wire[0:0] and_966_nl;
  wire[0:0] and_967_nl;
  wire[0:0] and_968_nl;
  wire[0:0] mux_337_nl;
  wire[0:0] nor_398_nl;
  wire[0:0] nor_390_nl;
  wire[0:0] or_919_nl;
  wire[0:0] nor_391_nl;
  wire[0:0] nor_392_nl;
  wire[0:0] nor_393_nl;
  wire[0:0] and_961_nl;
  wire[0:0] and_962_nl;
  wire[0:0] and_963_nl;
  wire[0:0] and_964_nl;
  wire[0:0] mux_346_nl;
  wire[0:0] nor_394_nl;
  wire[0:0] nor_380_nl;
  wire[0:0] or_938_nl;
  wire[0:0] nor_381_nl;
  wire[0:0] or_937_nl;
  wire[0:0] nor_382_nl;
  wire[0:0] or_936_nl;
  wire[0:0] nor_383_nl;
  wire[0:0] or_935_nl;
  wire[0:0] nor_384_nl;
  wire[0:0] or_934_nl;
  wire[0:0] nor_385_nl;
  wire[0:0] or_933_nl;
  wire[0:0] nor_386_nl;
  wire[0:0] or_932_nl;
  wire[0:0] nor_387_nl;
  wire[0:0] or_931_nl;
  wire[0:0] nor_388_nl;
  wire[0:0] or_930_nl;
  wire[0:0] nor_389_nl;
  wire[0:0] or_929_nl;
  wire[0:0] mux_357_nl;
  wire[0:0] nor_379_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] nor_378_nl;
  wire[0:0] mux_359_nl;
  wire[0:0] nor_377_nl;
  wire[0:0] mux_360_nl;
  wire[0:0] nor_376_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] nor_375_nl;
  wire[0:0] mux_362_nl;
  wire[0:0] nor_373_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] nor_374_nl;
  wire[0:0] nor_370_nl;
  wire[0:0] mux_365_nl;
  wire[0:0] nor_371_nl;
  wire[0:0] mux_366_nl;
  wire[0:0] nor_372_nl;
  wire[0:0] nor_366_nl;
  wire[0:0] nor_367_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] nor_368_nl;
  wire[0:0] mux_370_nl;
  wire[0:0] nor_369_nl;
  wire[0:0] nor_361_nl;
  wire[0:0] or_1012_nl;
  wire[0:0] nor_362_nl;
  wire[0:0] nor_363_nl;
  wire[0:0] mux_374_nl;
  wire[0:0] nor_364_nl;
  wire[0:0] mux_375_nl;
  wire[0:0] nor_365_nl;
  wire[0:0] nor_352_nl;
  wire[0:0] or_1027_nl;
  wire[0:0] nor_353_nl;
  wire[0:0] or_1026_nl;
  wire[0:0] nor_354_nl;
  wire[0:0] or_1025_nl;
  wire[0:0] nor_355_nl;
  wire[0:0] or_1024_nl;
  wire[0:0] nor_356_nl;
  wire[0:0] or_1023_nl;
  wire[0:0] nor_357_nl;
  wire[0:0] or_1022_nl;
  wire[0:0] nor_358_nl;
  wire[0:0] or_1021_nl;
  wire[0:0] nor_359_nl;
  wire[0:0] or_1020_nl;
  wire[0:0] mux_384_nl;
  wire[0:0] nor_360_nl;
  wire[0:0] or_1019_nl;
  wire[0:0] mux_385_nl;
  wire[0:0] nor_351_nl;
  wire[0:0] and_960_nl;
  wire[0:0] mux_387_nl;
  wire[0:0] nor_350_nl;
  wire[0:0] and_958_nl;
  wire[0:0] and_959_nl;
  wire[0:0] mux_390_nl;
  wire[0:0] nor_349_nl;
  wire[0:0] and_955_nl;
  wire[0:0] and_956_nl;
  wire[0:0] and_957_nl;
  wire[0:0] mux_394_nl;
  wire[0:0] nor_348_nl;
  wire[0:0] and_951_nl;
  wire[0:0] and_952_nl;
  wire[0:0] and_953_nl;
  wire[0:0] and_954_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] nor_347_nl;
  wire[0:0] nor_345_nl;
  wire[0:0] and_947_nl;
  wire[0:0] and_948_nl;
  wire[0:0] and_949_nl;
  wire[0:0] and_950_nl;
  wire[0:0] mux_405_nl;
  wire[0:0] nor_346_nl;
  wire[0:0] nor_342_nl;
  wire[0:0] nor_343_nl;
  wire[0:0] and_943_nl;
  wire[0:0] and_944_nl;
  wire[0:0] and_945_nl;
  wire[0:0] and_946_nl;
  wire[0:0] mux_412_nl;
  wire[0:0] nor_344_nl;
  wire[0:0] nor_338_nl;
  wire[0:0] nor_339_nl;
  wire[0:0] nor_340_nl;
  wire[0:0] and_939_nl;
  wire[0:0] and_940_nl;
  wire[0:0] and_941_nl;
  wire[0:0] and_942_nl;
  wire[0:0] mux_420_nl;
  wire[0:0] nor_341_nl;
  wire[0:0] nor_333_nl;
  wire[0:0] nand_12_nl;
  wire[0:0] nor_334_nl;
  wire[0:0] nor_335_nl;
  wire[0:0] nor_336_nl;
  wire[0:0] and_935_nl;
  wire[0:0] and_936_nl;
  wire[0:0] and_937_nl;
  wire[0:0] and_938_nl;
  wire[0:0] mux_429_nl;
  wire[0:0] nor_337_nl;
  wire[0:0] nor_324_nl;
  wire[0:0] nand_1_nl;
  wire[0:0] nor_325_nl;
  wire[0:0] nand_2_nl;
  wire[0:0] nor_326_nl;
  wire[0:0] nand_3_nl;
  wire[0:0] nor_327_nl;
  wire[0:0] nand_4_nl;
  wire[0:0] nor_328_nl;
  wire[0:0] nand_5_nl;
  wire[0:0] nor_329_nl;
  wire[0:0] nand_6_nl;
  wire[0:0] nor_330_nl;
  wire[0:0] nand_7_nl;
  wire[0:0] nor_331_nl;
  wire[0:0] nand_8_nl;
  wire[0:0] nor_332_nl;
  wire[0:0] nand_9_nl;
  wire[0:0] and_934_nl;
  wire[0:0] nand_11_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [64:0] nl_rem_13_cmp_a;
  assign nl_rem_13_cmp_a = {{1{rem_13_cmp_a_63_0[63]}}, rem_13_cmp_a_63_0};
  wire [64:0] nl_rem_13_cmp_b;
  assign nl_rem_13_cmp_b = {1'b0 , rem_13_cmp_b_63_0};
  wire [64:0] nl_rem_13_cmp_1_a;
  assign nl_rem_13_cmp_1_a = {{1{rem_13_cmp_1_a_63_0[63]}}, rem_13_cmp_1_a_63_0};
  wire [64:0] nl_rem_13_cmp_1_b;
  assign nl_rem_13_cmp_1_b = {1'b0 , rem_13_cmp_1_b_63_0};
  wire [64:0] nl_rem_13_cmp_2_a;
  assign nl_rem_13_cmp_2_a = {{1{rem_13_cmp_2_a_63_0[63]}}, rem_13_cmp_2_a_63_0};
  wire [64:0] nl_rem_13_cmp_2_b;
  assign nl_rem_13_cmp_2_b = {1'b0 , rem_13_cmp_2_b_63_0};
  wire [64:0] nl_rem_13_cmp_3_a;
  assign nl_rem_13_cmp_3_a = {{1{rem_13_cmp_3_a_63_0[63]}}, rem_13_cmp_3_a_63_0};
  wire [64:0] nl_rem_13_cmp_3_b;
  assign nl_rem_13_cmp_3_b = {1'b0 , rem_13_cmp_3_b_63_0};
  wire [64:0] nl_rem_13_cmp_4_a;
  assign nl_rem_13_cmp_4_a = {{1{rem_13_cmp_4_a_63_0[63]}}, rem_13_cmp_4_a_63_0};
  wire [64:0] nl_rem_13_cmp_4_b;
  assign nl_rem_13_cmp_4_b = {1'b0 , rem_13_cmp_4_b_63_0};
  wire [64:0] nl_rem_13_cmp_5_a;
  assign nl_rem_13_cmp_5_a = {{1{rem_13_cmp_5_a_63_0[63]}}, rem_13_cmp_5_a_63_0};
  wire [64:0] nl_rem_13_cmp_5_b;
  assign nl_rem_13_cmp_5_b = {1'b0 , rem_13_cmp_5_b_63_0};
  wire [64:0] nl_rem_13_cmp_6_a;
  assign nl_rem_13_cmp_6_a = {{1{rem_13_cmp_6_a_63_0[63]}}, rem_13_cmp_6_a_63_0};
  wire [64:0] nl_rem_13_cmp_6_b;
  assign nl_rem_13_cmp_6_b = {1'b0 , rem_13_cmp_6_b_63_0};
  wire [64:0] nl_rem_13_cmp_7_a;
  assign nl_rem_13_cmp_7_a = {{1{rem_13_cmp_7_a_63_0[63]}}, rem_13_cmp_7_a_63_0};
  wire [64:0] nl_rem_13_cmp_7_b;
  assign nl_rem_13_cmp_7_b = {1'b0 , rem_13_cmp_7_b_63_0};
  wire [64:0] nl_rem_13_cmp_8_a;
  assign nl_rem_13_cmp_8_a = {{1{rem_13_cmp_8_a_63_0[63]}}, rem_13_cmp_8_a_63_0};
  wire [64:0] nl_rem_13_cmp_8_b;
  assign nl_rem_13_cmp_8_b = {1'b0 , rem_13_cmp_8_b_63_0};
  wire [64:0] nl_rem_13_cmp_9_a;
  assign nl_rem_13_cmp_9_a = {{1{rem_13_cmp_9_a_63_0[63]}}, rem_13_cmp_9_a_63_0};
  wire [64:0] nl_rem_13_cmp_9_b;
  assign nl_rem_13_cmp_9_b = {1'b0 , rem_13_cmp_9_b_63_0};
  wire [64:0] nl_rem_13_cmp_10_a;
  assign nl_rem_13_cmp_10_a = {{1{rem_13_cmp_10_a_63_0[63]}}, rem_13_cmp_10_a_63_0};
  wire [64:0] nl_rem_13_cmp_10_b;
  assign nl_rem_13_cmp_10_b = {1'b0 , rem_13_cmp_10_b_63_0};
  wire [64:0] nl_rem_13_cmp_11_a;
  assign nl_rem_13_cmp_11_a = {{1{rem_13_cmp_11_a_63_0[63]}}, rem_13_cmp_11_a_63_0};
  wire [64:0] nl_rem_13_cmp_11_b;
  assign nl_rem_13_cmp_11_b = {1'b0 , rem_13_cmp_11_b_63_0};
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd64)) base_rsci (
      .dat(base_rsc_dat),
      .idat(base_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd3),
  .width(32'sd64)) return_rsci (
      .d(return_rsci_d),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd7),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp (
      .a(nl_rem_13_cmp_a[64:0]),
      .b(nl_rem_13_cmp_b[64:0]),
      .z(rem_13_cmp_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_1 (
      .a(nl_rem_13_cmp_1_a[64:0]),
      .b(nl_rem_13_cmp_1_b[64:0]),
      .z(rem_13_cmp_1_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_2 (
      .a(nl_rem_13_cmp_2_a[64:0]),
      .b(nl_rem_13_cmp_2_b[64:0]),
      .z(rem_13_cmp_2_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_3 (
      .a(nl_rem_13_cmp_3_a[64:0]),
      .b(nl_rem_13_cmp_3_b[64:0]),
      .z(rem_13_cmp_3_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_4 (
      .a(nl_rem_13_cmp_4_a[64:0]),
      .b(nl_rem_13_cmp_4_b[64:0]),
      .z(rem_13_cmp_4_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_5 (
      .a(nl_rem_13_cmp_5_a[64:0]),
      .b(nl_rem_13_cmp_5_b[64:0]),
      .z(rem_13_cmp_5_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_6 (
      .a(nl_rem_13_cmp_6_a[64:0]),
      .b(nl_rem_13_cmp_6_b[64:0]),
      .z(rem_13_cmp_6_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_7 (
      .a(nl_rem_13_cmp_7_a[64:0]),
      .b(nl_rem_13_cmp_7_b[64:0]),
      .z(rem_13_cmp_7_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_8 (
      .a(nl_rem_13_cmp_8_a[64:0]),
      .b(nl_rem_13_cmp_8_b[64:0]),
      .z(rem_13_cmp_8_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_9 (
      .a(nl_rem_13_cmp_9_a[64:0]),
      .b(nl_rem_13_cmp_9_b[64:0]),
      .z(rem_13_cmp_9_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_10 (
      .a(nl_rem_13_cmp_10_a[64:0]),
      .b(nl_rem_13_cmp_10_b[64:0]),
      .z(rem_13_cmp_10_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_13_cmp_11 (
      .a(nl_rem_13_cmp_11_a[64:0]),
      .b(nl_rem_13_cmp_11_b[64:0]),
      .z(rem_13_cmp_11_z)
    );
  assign and_1203_cse = ccs_ccore_en & main_stage_0_12 & asn_itm_11;
  assign and_1173_cse = ccs_ccore_en & (and_dcpl_294 | and_dcpl_300 | and_dcpl_306
      | and_dcpl_312 | and_dcpl_318 | and_dcpl_324 | and_dcpl_330 | and_dcpl_336
      | and_dcpl_342 | and_dcpl_348 | and_tmp_35);
  assign and_1175_cse = ccs_ccore_en & (and_dcpl_356 | and_dcpl_360 | and_dcpl_364
      | and_dcpl_368 | and_dcpl_372 | and_dcpl_376 | and_dcpl_379 | and_dcpl_382
      | and_dcpl_385 | and_dcpl_388 | mux_tmp_76);
  assign and_1177_cse = ccs_ccore_en & (and_dcpl_394 | and_dcpl_397 | and_dcpl_400
      | and_dcpl_403 | and_dcpl_406 | and_dcpl_409 | and_dcpl_413 | and_dcpl_417
      | and_dcpl_421 | and_dcpl_425 | and_tmp_80);
  assign and_1179_cse = ccs_ccore_en & (and_dcpl_431 | and_dcpl_433 | and_dcpl_435
      | and_dcpl_437 | and_dcpl_439 | and_dcpl_442 | and_dcpl_445 | and_dcpl_448
      | and_dcpl_451 | and_dcpl_454 | mux_tmp_141);
  assign and_1181_cse = ccs_ccore_en & (and_dcpl_461 | and_dcpl_465 | and_dcpl_469
      | and_dcpl_473 | and_dcpl_477 | and_dcpl_480 | and_dcpl_483 | and_dcpl_486
      | and_dcpl_489 | and_dcpl_492 | and_tmp_125);
  assign and_1183_cse = ccs_ccore_en & (and_dcpl_498 | and_dcpl_500 | and_dcpl_502
      | and_dcpl_504 | and_dcpl_506 | and_dcpl_508 | and_dcpl_510 | and_dcpl_512
      | and_dcpl_514 | and_dcpl_516 | mux_tmp_206);
  assign and_1185_cse = ccs_ccore_en & (and_dcpl_520 | and_dcpl_523 | and_dcpl_526
      | and_dcpl_529 | and_dcpl_532 | and_dcpl_534 | and_dcpl_536 | and_dcpl_538
      | and_dcpl_540 | and_dcpl_542 | and_tmp_170);
  assign and_1187_cse = ccs_ccore_en & (and_dcpl_546 | and_dcpl_548 | and_dcpl_550
      | and_dcpl_552 | and_dcpl_554 | and_dcpl_556 | and_dcpl_558 | and_dcpl_560
      | and_dcpl_562 | and_dcpl_564 | mux_tmp_271);
  assign and_1189_cse = ccs_ccore_en & (and_dcpl_569 | and_dcpl_573 | and_dcpl_577
      | and_dcpl_581 | and_dcpl_585 | and_dcpl_589 | and_dcpl_593 | and_dcpl_597
      | and_dcpl_601 | and_dcpl_605 | and_tmp_206);
  assign and_1191_cse = ccs_ccore_en & (and_dcpl_610 | and_dcpl_612 | and_dcpl_614
      | and_dcpl_616 | and_dcpl_618 | and_dcpl_622 | and_dcpl_625 | and_dcpl_628
      | and_dcpl_631 | and_dcpl_634 | mux_tmp_354);
  assign and_1193_cse = ccs_ccore_en & (and_dcpl_638 | and_dcpl_641 | and_dcpl_644
      | and_dcpl_647 | and_dcpl_650 | and_dcpl_653 | and_dcpl_657 | and_dcpl_661
      | and_dcpl_665 | and_dcpl_669 | and_tmp_233);
  assign and_1195_cse = ccs_ccore_en & (and_dcpl_673 | and_dcpl_675 | and_dcpl_677
      | and_dcpl_679 | and_dcpl_681 | and_dcpl_684 | and_dcpl_687 | and_dcpl_690
      | and_dcpl_693 | and_dcpl_696 | mux_tmp_437);
  assign and_1205_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_2;
  assign and_1207_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_6;
  assign and_1209_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_9;
  assign and_1211_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_11;
  assign and_1213_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_2;
  assign and_1215_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_6;
  assign and_1217_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_9;
  assign and_1219_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_11;
  assign and_1221_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_18 & (~ (rem_12cyc_st_10_1_0[0]));
  assign and_1223_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_18 & (rem_12cyc_st_10_1_0[0]);
  assign and_1225_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_23 & (~ (rem_12cyc_st_10_1_0[0]));
  assign and_1227_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_23 & (rem_12cyc_st_10_1_0[0]);
  assign and_1229_cse = ccs_ccore_en & and_dcpl_3;
  assign and_1231_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_29;
  assign and_1233_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_33;
  assign and_1235_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_36;
  assign and_1237_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_38;
  assign and_1239_cse = ccs_ccore_en & and_dcpl_40 & and_dcpl_29;
  assign and_1241_cse = ccs_ccore_en & and_dcpl_40 & and_dcpl_33;
  assign and_1243_cse = ccs_ccore_en & and_dcpl_40 & and_dcpl_36;
  assign and_1245_cse = ccs_ccore_en & and_dcpl_40 & and_dcpl_38;
  assign and_1247_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_45 & (~ (rem_12cyc_st_9_1_0[0]));
  assign and_1249_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_45 & (rem_12cyc_st_9_1_0[0]);
  assign and_1251_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_50 & (~ (rem_12cyc_st_9_1_0[0]));
  assign and_1253_cse = ccs_ccore_en & and_dcpl_31 & and_dcpl_50 & (rem_12cyc_st_9_1_0[0]);
  assign and_1255_cse = ccs_ccore_en & and_dcpl_30;
  assign and_1257_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_56;
  assign and_1259_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_60;
  assign and_1261_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_63;
  assign and_1263_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_65;
  assign and_1265_cse = ccs_ccore_en & and_dcpl_67 & and_dcpl_56;
  assign and_1267_cse = ccs_ccore_en & and_dcpl_67 & and_dcpl_60;
  assign and_1269_cse = ccs_ccore_en & and_dcpl_67 & and_dcpl_63;
  assign and_1271_cse = ccs_ccore_en & and_dcpl_67 & and_dcpl_65;
  assign and_1273_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_72 & (~ (rem_12cyc_st_8_1_0[0]));
  assign and_1275_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_72 & (rem_12cyc_st_8_1_0[0]);
  assign and_1277_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_77 & (~ (rem_12cyc_st_8_1_0[0]));
  assign and_1279_cse = ccs_ccore_en & and_dcpl_58 & and_dcpl_77 & (rem_12cyc_st_8_1_0[0]);
  assign and_1281_cse = ccs_ccore_en & and_dcpl_57;
  assign and_1283_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_83;
  assign and_1285_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_87;
  assign and_1287_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_90;
  assign and_1289_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_92;
  assign and_1291_cse = ccs_ccore_en & and_dcpl_94 & and_dcpl_83;
  assign and_1293_cse = ccs_ccore_en & and_dcpl_94 & and_dcpl_87;
  assign and_1295_cse = ccs_ccore_en & and_dcpl_94 & and_dcpl_90;
  assign and_1297_cse = ccs_ccore_en & and_dcpl_94 & and_dcpl_92;
  assign and_1299_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_99 & (~ (rem_12cyc_st_7_1_0[0]));
  assign and_1301_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_99 & (rem_12cyc_st_7_1_0[0]);
  assign and_1303_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_104 & (~ (rem_12cyc_st_7_1_0[0]));
  assign and_1305_cse = ccs_ccore_en & and_dcpl_85 & and_dcpl_104 & (rem_12cyc_st_7_1_0[0]);
  assign and_1307_cse = ccs_ccore_en & and_dcpl_84;
  assign and_1309_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_110;
  assign and_1311_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_115;
  assign and_1313_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_117;
  assign and_1315_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_119;
  assign and_1317_cse = ccs_ccore_en & and_dcpl_121 & and_dcpl_110;
  assign and_1319_cse = ccs_ccore_en & and_dcpl_121 & and_dcpl_115;
  assign and_1321_cse = ccs_ccore_en & and_dcpl_121 & and_dcpl_117;
  assign and_1323_cse = ccs_ccore_en & and_dcpl_121 & and_dcpl_119;
  assign and_1325_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_126 & (~ (rem_12cyc_st_6_1_0[1]));
  assign and_1327_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_129 & (~ (rem_12cyc_st_6_1_0[1]));
  assign and_1329_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_126 & (rem_12cyc_st_6_1_0[1]);
  assign and_1331_cse = ccs_ccore_en & and_dcpl_112 & and_dcpl_129 & (rem_12cyc_st_6_1_0[1]);
  assign and_1333_cse = ccs_ccore_en & and_dcpl_111;
  assign and_1335_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_137;
  assign and_1337_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_141;
  assign and_1339_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_144;
  assign and_1341_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_146;
  assign and_1343_cse = ccs_ccore_en & and_dcpl_148 & and_dcpl_137;
  assign and_1345_cse = ccs_ccore_en & and_dcpl_148 & and_dcpl_141;
  assign and_1347_cse = ccs_ccore_en & and_dcpl_148 & and_dcpl_144;
  assign and_1349_cse = ccs_ccore_en & and_dcpl_148 & and_dcpl_146;
  assign and_1351_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_153 & (~ (rem_12cyc_st_5_1_0[0]));
  assign and_1353_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_153 & (rem_12cyc_st_5_1_0[0]);
  assign and_1355_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_158 & (~ (rem_12cyc_st_5_1_0[0]));
  assign and_1357_cse = ccs_ccore_en & and_dcpl_139 & and_dcpl_158 & (rem_12cyc_st_5_1_0[0]);
  assign and_1359_cse = ccs_ccore_en & and_dcpl_138;
  assign and_1361_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_164;
  assign and_1363_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_168;
  assign and_1365_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_171;
  assign and_1367_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_173;
  assign and_1369_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_175 & (~ (rem_12cyc_st_4_1_0[0]));
  assign and_1371_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_175 & (rem_12cyc_st_4_1_0[0]);
  assign and_1373_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_180 & (~ (rem_12cyc_st_4_1_0[0]));
  assign and_1375_cse = ccs_ccore_en & and_dcpl_166 & and_dcpl_180 & (rem_12cyc_st_4_1_0[0]);
  assign and_1377_cse = ccs_ccore_en & and_dcpl_185 & and_dcpl_164;
  assign and_1379_cse = ccs_ccore_en & and_dcpl_185 & and_dcpl_168;
  assign and_1381_cse = ccs_ccore_en & and_dcpl_185 & and_dcpl_171;
  assign and_1383_cse = ccs_ccore_en & and_dcpl_185 & and_dcpl_173;
  assign and_1385_cse = ccs_ccore_en & and_dcpl_165;
  assign and_1387_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_191;
  assign and_1389_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_195;
  assign and_1391_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_198;
  assign and_1393_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_200;
  assign and_1395_cse = ccs_ccore_en & and_dcpl_202 & and_dcpl_191;
  assign and_1397_cse = ccs_ccore_en & and_dcpl_202 & and_dcpl_195;
  assign and_1399_cse = ccs_ccore_en & and_dcpl_202 & and_dcpl_198;
  assign and_1401_cse = ccs_ccore_en & and_dcpl_202 & and_dcpl_200;
  assign and_1403_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_207 & (~ (rem_12cyc_st_3_1_0[0]));
  assign and_1405_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_207 & (rem_12cyc_st_3_1_0[0]);
  assign and_1407_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_212 & (~ (rem_12cyc_st_3_1_0[0]));
  assign and_1409_cse = ccs_ccore_en & and_dcpl_193 & and_dcpl_212 & (rem_12cyc_st_3_1_0[0]);
  assign and_1411_cse = ccs_ccore_en & and_dcpl_192;
  assign and_1413_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_218;
  assign and_1415_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_222;
  assign and_1417_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_225;
  assign and_1419_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_227;
  assign and_1421_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_229 & (~ (rem_12cyc_st_2_1_0[0]));
  assign and_1423_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_229 & (rem_12cyc_st_2_1_0[0]);
  assign and_1425_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_234 & (~ (rem_12cyc_st_2_1_0[0]));
  assign and_1427_cse = ccs_ccore_en & and_dcpl_220 & and_dcpl_234 & (rem_12cyc_st_2_1_0[0]);
  assign and_1429_cse = ccs_ccore_en & and_dcpl_239 & and_dcpl_218;
  assign and_1431_cse = ccs_ccore_en & and_dcpl_239 & and_dcpl_222;
  assign and_1433_cse = ccs_ccore_en & and_dcpl_239 & and_dcpl_225;
  assign and_1435_cse = ccs_ccore_en & and_dcpl_239 & and_dcpl_227;
  assign and_1437_cse = ccs_ccore_en & and_dcpl_219;
  assign and_1439_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_245;
  assign and_1441_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_249;
  assign and_1443_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_252;
  assign and_1445_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_254;
  assign and_1447_cse = ccs_ccore_en & and_dcpl_256 & and_dcpl_245;
  assign and_1449_cse = ccs_ccore_en & and_dcpl_256 & and_dcpl_249;
  assign and_1451_cse = ccs_ccore_en & and_dcpl_256 & and_dcpl_252;
  assign and_1453_cse = ccs_ccore_en & and_dcpl_256 & and_dcpl_254;
  assign and_1455_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_261 & (~ (rem_12cyc_1_0[0]));
  assign and_1457_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_261 & (rem_12cyc_1_0[0]);
  assign and_1459_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_266 & (~ (rem_12cyc_1_0[0]));
  assign and_1461_cse = ccs_ccore_en & and_dcpl_247 & and_dcpl_266 & (rem_12cyc_1_0[0]);
  assign and_1463_cse = ccs_ccore_en & and_dcpl_246;
  assign and_1197_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  assign and_273_nl = and_dcpl_272 & and_dcpl_271;
  assign and_275_nl = and_dcpl_272 & and_dcpl_274;
  assign and_277_nl = and_dcpl_272 & and_dcpl_276;
  assign and_279_nl = and_dcpl_272 & and_dcpl_278;
  assign and_281_nl = and_dcpl_280 & and_dcpl_271;
  assign and_282_nl = and_dcpl_280 & and_dcpl_274;
  assign and_283_nl = and_dcpl_280 & and_dcpl_276;
  assign and_284_nl = and_dcpl_280 & and_dcpl_278;
  assign and_286_nl = and_dcpl_285 & and_dcpl_271;
  assign and_287_nl = and_dcpl_285 & and_dcpl_274;
  assign and_288_nl = and_dcpl_285 & and_dcpl_276;
  assign and_289_nl = and_dcpl_285 & and_dcpl_278;
  assign and_290_nl = (rem_12cyc_st_12_3_2==2'b11);
  assign result_sva_duc_mx0 = MUX1HOT_v_64_13_2((rem_13_cmp_1_z[63:0]), (rem_13_cmp_2_z[63:0]),
      (rem_13_cmp_3_z[63:0]), (rem_13_cmp_4_z[63:0]), (rem_13_cmp_5_z[63:0]), (rem_13_cmp_6_z[63:0]),
      (rem_13_cmp_7_z[63:0]), (rem_13_cmp_8_z[63:0]), (rem_13_cmp_9_z[63:0]), (rem_13_cmp_10_z[63:0]),
      (rem_13_cmp_11_z[63:0]), (rem_13_cmp_z[63:0]), result_sva_duc, {and_273_nl
      , and_275_nl , and_277_nl , and_279_nl , and_281_nl , and_282_nl , and_283_nl
      , and_284_nl , and_286_nl , and_287_nl , and_288_nl , and_289_nl , and_290_nl});
  assign nl_acc_1_tmp = ({rem_12cyc_3_2 , rem_12cyc_1_0}) + 4'b0001;
  assign acc_1_tmp = nl_acc_1_tmp[3:0];
  assign xor_nl = (acc_1_tmp[2]) ^ (acc_1_tmp[3]);
  assign nor_nl = ~((acc_1_tmp[3:2]!=2'b10));
  assign nl_acc_tmp = conv_u2u_1_2(xor_nl) + conv_u2u_1_2(nor_nl);
  assign acc_tmp = nl_acc_tmp[1:0];
  assign and_dcpl_1 = ~((rem_12cyc_st_10_3_2[1]) | (rem_12cyc_st_10_1_0[1]));
  assign and_dcpl_2 = and_dcpl_1 & (~ (rem_12cyc_st_10_1_0[0]));
  assign and_dcpl_3 = main_stage_0_11 & asn_itm_10;
  assign and_dcpl_4 = and_dcpl_3 & (~ (rem_12cyc_st_10_3_2[0]));
  assign and_dcpl_6 = and_dcpl_1 & (rem_12cyc_st_10_1_0[0]);
  assign and_dcpl_8 = (~ (rem_12cyc_st_10_3_2[1])) & (rem_12cyc_st_10_1_0[1]);
  assign and_dcpl_9 = and_dcpl_8 & (~ (rem_12cyc_st_10_1_0[0]));
  assign and_dcpl_11 = and_dcpl_8 & (rem_12cyc_st_10_1_0[0]);
  assign and_dcpl_13 = and_dcpl_3 & (rem_12cyc_st_10_3_2[0]);
  assign and_dcpl_18 = (rem_12cyc_st_10_3_2[1]) & (~ (rem_12cyc_st_10_1_0[1]));
  assign and_dcpl_23 = (rem_12cyc_st_10_3_2[1]) & (rem_12cyc_st_10_1_0[1]);
  assign and_dcpl_28 = ~((rem_12cyc_st_9_3_2[1]) | (rem_12cyc_st_9_1_0[1]));
  assign and_dcpl_29 = and_dcpl_28 & (~ (rem_12cyc_st_9_1_0[0]));
  assign and_dcpl_30 = main_stage_0_10 & asn_itm_9;
  assign and_dcpl_31 = and_dcpl_30 & (~ (rem_12cyc_st_9_3_2[0]));
  assign and_dcpl_33 = and_dcpl_28 & (rem_12cyc_st_9_1_0[0]);
  assign and_dcpl_35 = (~ (rem_12cyc_st_9_3_2[1])) & (rem_12cyc_st_9_1_0[1]);
  assign and_dcpl_36 = and_dcpl_35 & (~ (rem_12cyc_st_9_1_0[0]));
  assign and_dcpl_38 = and_dcpl_35 & (rem_12cyc_st_9_1_0[0]);
  assign and_dcpl_40 = and_dcpl_30 & (rem_12cyc_st_9_3_2[0]);
  assign and_dcpl_45 = (rem_12cyc_st_9_3_2[1]) & (~ (rem_12cyc_st_9_1_0[1]));
  assign and_dcpl_50 = (rem_12cyc_st_9_3_2[1]) & (rem_12cyc_st_9_1_0[1]);
  assign and_dcpl_55 = ~((rem_12cyc_st_8_3_2[1]) | (rem_12cyc_st_8_1_0[1]));
  assign and_dcpl_56 = and_dcpl_55 & (~ (rem_12cyc_st_8_1_0[0]));
  assign and_dcpl_57 = main_stage_0_9 & asn_itm_8;
  assign and_dcpl_58 = and_dcpl_57 & (~ (rem_12cyc_st_8_3_2[0]));
  assign and_dcpl_60 = and_dcpl_55 & (rem_12cyc_st_8_1_0[0]);
  assign and_dcpl_62 = (~ (rem_12cyc_st_8_3_2[1])) & (rem_12cyc_st_8_1_0[1]);
  assign and_dcpl_63 = and_dcpl_62 & (~ (rem_12cyc_st_8_1_0[0]));
  assign and_dcpl_65 = and_dcpl_62 & (rem_12cyc_st_8_1_0[0]);
  assign and_dcpl_67 = and_dcpl_57 & (rem_12cyc_st_8_3_2[0]);
  assign and_dcpl_72 = (rem_12cyc_st_8_3_2[1]) & (~ (rem_12cyc_st_8_1_0[1]));
  assign and_dcpl_77 = (rem_12cyc_st_8_3_2[1]) & (rem_12cyc_st_8_1_0[1]);
  assign and_dcpl_82 = ~((rem_12cyc_st_7_3_2[1]) | (rem_12cyc_st_7_1_0[1]));
  assign and_dcpl_83 = and_dcpl_82 & (~ (rem_12cyc_st_7_1_0[0]));
  assign and_dcpl_84 = main_stage_0_8 & asn_itm_7;
  assign and_dcpl_85 = and_dcpl_84 & (~ (rem_12cyc_st_7_3_2[0]));
  assign and_dcpl_87 = and_dcpl_82 & (rem_12cyc_st_7_1_0[0]);
  assign and_dcpl_89 = (~ (rem_12cyc_st_7_3_2[1])) & (rem_12cyc_st_7_1_0[1]);
  assign and_dcpl_90 = and_dcpl_89 & (~ (rem_12cyc_st_7_1_0[0]));
  assign and_dcpl_92 = and_dcpl_89 & (rem_12cyc_st_7_1_0[0]);
  assign and_dcpl_94 = and_dcpl_84 & (rem_12cyc_st_7_3_2[0]);
  assign and_dcpl_99 = (rem_12cyc_st_7_3_2[1]) & (~ (rem_12cyc_st_7_1_0[1]));
  assign and_dcpl_104 = (rem_12cyc_st_7_3_2[1]) & (rem_12cyc_st_7_1_0[1]);
  assign and_dcpl_109 = ~((rem_12cyc_st_6_3_2[1]) | (rem_12cyc_st_6_1_0[0]));
  assign and_dcpl_110 = and_dcpl_109 & (~ (rem_12cyc_st_6_1_0[1]));
  assign and_dcpl_111 = main_stage_0_7 & asn_itm_6;
  assign and_dcpl_112 = and_dcpl_111 & (~ (rem_12cyc_st_6_3_2[0]));
  assign and_dcpl_114 = (~ (rem_12cyc_st_6_3_2[1])) & (rem_12cyc_st_6_1_0[0]);
  assign and_dcpl_115 = and_dcpl_114 & (~ (rem_12cyc_st_6_1_0[1]));
  assign and_dcpl_117 = and_dcpl_109 & (rem_12cyc_st_6_1_0[1]);
  assign and_dcpl_119 = and_dcpl_114 & (rem_12cyc_st_6_1_0[1]);
  assign and_dcpl_121 = and_dcpl_111 & (rem_12cyc_st_6_3_2[0]);
  assign and_dcpl_126 = (rem_12cyc_st_6_3_2[1]) & (~ (rem_12cyc_st_6_1_0[0]));
  assign and_dcpl_129 = (rem_12cyc_st_6_3_2[1]) & (rem_12cyc_st_6_1_0[0]);
  assign and_dcpl_136 = ~((rem_12cyc_st_5_3_2[1]) | (rem_12cyc_st_5_1_0[1]));
  assign and_dcpl_137 = and_dcpl_136 & (~ (rem_12cyc_st_5_1_0[0]));
  assign and_dcpl_138 = main_stage_0_6 & asn_itm_5;
  assign and_dcpl_139 = and_dcpl_138 & (~ (rem_12cyc_st_5_3_2[0]));
  assign and_dcpl_141 = and_dcpl_136 & (rem_12cyc_st_5_1_0[0]);
  assign and_dcpl_143 = (~ (rem_12cyc_st_5_3_2[1])) & (rem_12cyc_st_5_1_0[1]);
  assign and_dcpl_144 = and_dcpl_143 & (~ (rem_12cyc_st_5_1_0[0]));
  assign and_dcpl_146 = and_dcpl_143 & (rem_12cyc_st_5_1_0[0]);
  assign and_dcpl_148 = and_dcpl_138 & (rem_12cyc_st_5_3_2[0]);
  assign and_dcpl_153 = (rem_12cyc_st_5_3_2[1]) & (~ (rem_12cyc_st_5_1_0[1]));
  assign and_dcpl_158 = (rem_12cyc_st_5_3_2[1]) & (rem_12cyc_st_5_1_0[1]);
  assign and_dcpl_163 = ~((rem_12cyc_st_4_3_2[0]) | (rem_12cyc_st_4_1_0[1]));
  assign and_dcpl_164 = and_dcpl_163 & (~ (rem_12cyc_st_4_1_0[0]));
  assign and_dcpl_165 = main_stage_0_5 & asn_itm_4;
  assign and_dcpl_166 = and_dcpl_165 & (~ (rem_12cyc_st_4_3_2[1]));
  assign and_dcpl_168 = and_dcpl_163 & (rem_12cyc_st_4_1_0[0]);
  assign and_dcpl_170 = (~ (rem_12cyc_st_4_3_2[0])) & (rem_12cyc_st_4_1_0[1]);
  assign and_dcpl_171 = and_dcpl_170 & (~ (rem_12cyc_st_4_1_0[0]));
  assign and_dcpl_173 = and_dcpl_170 & (rem_12cyc_st_4_1_0[0]);
  assign and_dcpl_175 = (rem_12cyc_st_4_3_2[0]) & (~ (rem_12cyc_st_4_1_0[1]));
  assign and_dcpl_180 = (rem_12cyc_st_4_3_2[0]) & (rem_12cyc_st_4_1_0[1]);
  assign and_dcpl_185 = and_dcpl_165 & (rem_12cyc_st_4_3_2[1]);
  assign and_dcpl_190 = ~((rem_12cyc_st_3_3_2[1]) | (rem_12cyc_st_3_1_0[1]));
  assign and_dcpl_191 = and_dcpl_190 & (~ (rem_12cyc_st_3_1_0[0]));
  assign and_dcpl_192 = main_stage_0_4 & asn_itm_3;
  assign and_dcpl_193 = and_dcpl_192 & (~ (rem_12cyc_st_3_3_2[0]));
  assign and_dcpl_195 = and_dcpl_190 & (rem_12cyc_st_3_1_0[0]);
  assign and_dcpl_197 = (~ (rem_12cyc_st_3_3_2[1])) & (rem_12cyc_st_3_1_0[1]);
  assign and_dcpl_198 = and_dcpl_197 & (~ (rem_12cyc_st_3_1_0[0]));
  assign and_dcpl_200 = and_dcpl_197 & (rem_12cyc_st_3_1_0[0]);
  assign and_dcpl_202 = and_dcpl_192 & (rem_12cyc_st_3_3_2[0]);
  assign and_dcpl_207 = (rem_12cyc_st_3_3_2[1]) & (~ (rem_12cyc_st_3_1_0[1]));
  assign and_dcpl_212 = (rem_12cyc_st_3_3_2[1]) & (rem_12cyc_st_3_1_0[1]);
  assign and_dcpl_217 = ~((rem_12cyc_st_2_3_2[0]) | (rem_12cyc_st_2_1_0[1]));
  assign and_dcpl_218 = and_dcpl_217 & (~ (rem_12cyc_st_2_1_0[0]));
  assign and_dcpl_219 = main_stage_0_3 & asn_itm_2;
  assign and_dcpl_220 = and_dcpl_219 & (~ (rem_12cyc_st_2_3_2[1]));
  assign and_dcpl_222 = and_dcpl_217 & (rem_12cyc_st_2_1_0[0]);
  assign and_dcpl_224 = (~ (rem_12cyc_st_2_3_2[0])) & (rem_12cyc_st_2_1_0[1]);
  assign and_dcpl_225 = and_dcpl_224 & (~ (rem_12cyc_st_2_1_0[0]));
  assign and_dcpl_227 = and_dcpl_224 & (rem_12cyc_st_2_1_0[0]);
  assign and_dcpl_229 = (rem_12cyc_st_2_3_2[0]) & (~ (rem_12cyc_st_2_1_0[1]));
  assign and_dcpl_234 = (rem_12cyc_st_2_3_2[0]) & (rem_12cyc_st_2_1_0[1]);
  assign and_dcpl_239 = and_dcpl_219 & (rem_12cyc_st_2_3_2[1]);
  assign and_dcpl_244 = ~((rem_12cyc_3_2[1]) | (rem_12cyc_1_0[1]));
  assign and_dcpl_245 = and_dcpl_244 & (~ (rem_12cyc_1_0[0]));
  assign and_dcpl_246 = main_stage_0_2 & asn_itm_1;
  assign and_dcpl_247 = and_dcpl_246 & (~ (rem_12cyc_3_2[0]));
  assign and_dcpl_249 = and_dcpl_244 & (rem_12cyc_1_0[0]);
  assign and_dcpl_251 = (~ (rem_12cyc_3_2[1])) & (rem_12cyc_1_0[1]);
  assign and_dcpl_252 = and_dcpl_251 & (~ (rem_12cyc_1_0[0]));
  assign and_dcpl_254 = and_dcpl_251 & (rem_12cyc_1_0[0]);
  assign and_dcpl_256 = and_dcpl_246 & (rem_12cyc_3_2[0]);
  assign and_dcpl_261 = (rem_12cyc_3_2[1]) & (~ (rem_12cyc_1_0[1]));
  assign and_dcpl_266 = (rem_12cyc_3_2[1]) & (rem_12cyc_1_0[1]);
  assign and_dcpl_271 = ~((rem_12cyc_st_12_1_0!=2'b00));
  assign and_dcpl_272 = ~((rem_12cyc_st_12_3_2!=2'b00));
  assign and_dcpl_274 = (rem_12cyc_st_12_1_0==2'b01);
  assign and_dcpl_276 = (rem_12cyc_st_12_1_0==2'b10);
  assign and_dcpl_278 = (rem_12cyc_st_12_1_0==2'b11);
  assign and_dcpl_280 = (rem_12cyc_st_12_3_2==2'b01);
  assign and_dcpl_285 = (rem_12cyc_st_12_3_2==2'b10);
  assign and_dcpl_291 = ~((acc_1_tmp[1:0]!=2'b00));
  assign and_dcpl_292 = ccs_ccore_start_rsci_idat & (~ (acc_tmp[0]));
  assign and_dcpl_293 = and_dcpl_292 & (~ (acc_tmp[1]));
  assign and_dcpl_294 = and_dcpl_293 & and_dcpl_291;
  assign and_dcpl_295 = ~((rem_12cyc_st_2_3_2!=2'b00));
  assign and_dcpl_296 = and_dcpl_295 & (~ (rem_12cyc_st_2_1_0[1]));
  assign and_dcpl_298 = (~ (rem_12cyc_st_2_1_0[0])) & main_stage_0_3 & asn_itm_2;
  assign not_tmp_54 = ~(asn_itm_1 & main_stage_0_2);
  assign or_tmp_2 = (rem_12cyc_1_0!=2'b00) | (rem_12cyc_3_2!=2'b00) | not_tmp_54;
  assign or_1_cse = (acc_1_tmp[1:0]!=2'b00) | (acc_tmp!=2'b00);
  assign nor_518_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_2));
  assign mux_14_nl = MUX_s_1_2_2(nor_518_nl, or_tmp_2, or_1_cse);
  assign and_dcpl_300 = mux_14_nl & and_dcpl_298 & and_dcpl_296;
  assign and_dcpl_301 = ~((rem_12cyc_st_3_3_2!=2'b00));
  assign and_dcpl_302 = and_dcpl_301 & (~ (rem_12cyc_st_3_1_0[1]));
  assign and_dcpl_304 = (~ (rem_12cyc_st_3_1_0[0])) & main_stage_0_4 & asn_itm_3;
  assign or_6_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2!=2'b00) | (~ asn_itm_2)
      | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp = or_6_cse & or_tmp_2;
  assign nor_517_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp));
  assign mux_15_nl = MUX_s_1_2_2(nor_517_nl, and_tmp, or_1_cse);
  assign and_dcpl_306 = mux_15_nl & and_dcpl_304 & and_dcpl_302;
  assign and_dcpl_307 = ~((rem_12cyc_st_4_3_2!=2'b00));
  assign and_dcpl_308 = and_dcpl_307 & (~ (rem_12cyc_st_4_1_0[1]));
  assign and_dcpl_310 = (~ (rem_12cyc_st_4_1_0[0])) & main_stage_0_5 & asn_itm_4;
  assign or_10_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2!=2'b00) | (~ asn_itm_3)
      | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_2 = or_6_cse & or_10_cse & or_tmp_2;
  assign nor_516_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_2));
  assign mux_16_nl = MUX_s_1_2_2(nor_516_nl, and_tmp_2, or_1_cse);
  assign and_dcpl_312 = mux_16_nl & and_dcpl_310 & and_dcpl_308;
  assign and_dcpl_313 = ~((rem_12cyc_st_5_3_2!=2'b00));
  assign and_dcpl_314 = and_dcpl_313 & (~ (rem_12cyc_st_5_1_0[1]));
  assign and_dcpl_316 = (~ (rem_12cyc_st_5_1_0[0])) & main_stage_0_6 & asn_itm_5;
  assign or_15_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2!=2'b00) | (~ asn_itm_4)
      | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_5 = or_6_cse & or_10_cse & or_15_cse & or_tmp_2;
  assign nor_515_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_5));
  assign mux_17_nl = MUX_s_1_2_2(nor_515_nl, and_tmp_5, or_1_cse);
  assign and_dcpl_318 = mux_17_nl & and_dcpl_316 & and_dcpl_314;
  assign or_21_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2!=2'b00) | (~ asn_itm_5)
      | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_9 = or_6_cse & or_10_cse & or_15_cse & or_21_cse & or_tmp_2;
  assign nor_514_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_9));
  assign mux_18_nl = MUX_s_1_2_2(nor_514_nl, and_tmp_9, or_1_cse);
  assign and_dcpl_324 = mux_18_nl & and_dcpl_112 & and_dcpl_110;
  assign or_28_cse = (rem_12cyc_st_6_1_0!=2'b00) | (rem_12cyc_st_6_3_2!=2'b00);
  assign nor_512_nl = ~(and_dcpl_111 | (~ or_tmp_2));
  assign mux_19_nl = MUX_s_1_2_2(nor_512_nl, or_tmp_2, or_28_cse);
  assign and_tmp_13 = or_6_cse & or_10_cse & or_15_cse & or_21_cse & mux_19_nl;
  assign nor_513_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_13));
  assign mux_20_nl = MUX_s_1_2_2(nor_513_nl, and_tmp_13, or_1_cse);
  assign and_dcpl_330 = mux_20_nl & and_dcpl_85 & and_dcpl_83;
  assign or_37_cse = (rem_12cyc_st_7_1_0!=2'b00) | (rem_12cyc_st_7_3_2!=2'b00);
  assign nor_509_nl = ~(and_dcpl_84 | (~ or_tmp_2));
  assign mux_tmp_19 = MUX_s_1_2_2(nor_509_nl, or_tmp_2, or_37_cse);
  assign nor_510_nl = ~(and_dcpl_111 | (~ mux_tmp_19));
  assign mux_22_nl = MUX_s_1_2_2(nor_510_nl, mux_tmp_19, or_28_cse);
  assign and_tmp_17 = or_6_cse & or_10_cse & or_15_cse & or_21_cse & mux_22_nl;
  assign nor_511_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_17));
  assign mux_23_nl = MUX_s_1_2_2(nor_511_nl, and_tmp_17, or_1_cse);
  assign and_dcpl_336 = mux_23_nl & and_dcpl_58 & and_dcpl_56;
  assign or_48_cse = (rem_12cyc_st_8_1_0!=2'b00) | (rem_12cyc_st_8_3_2!=2'b00);
  assign nor_505_nl = ~(and_dcpl_57 | (~ or_tmp_2));
  assign mux_tmp_22 = MUX_s_1_2_2(nor_505_nl, or_tmp_2, or_48_cse);
  assign nor_506_nl = ~(and_dcpl_84 | (~ mux_tmp_22));
  assign mux_tmp_23 = MUX_s_1_2_2(nor_506_nl, mux_tmp_22, or_37_cse);
  assign nor_507_nl = ~(and_dcpl_111 | (~ mux_tmp_23));
  assign mux_26_nl = MUX_s_1_2_2(nor_507_nl, mux_tmp_23, or_28_cse);
  assign and_tmp_21 = or_6_cse & or_10_cse & or_15_cse & or_21_cse & mux_26_nl;
  assign nor_508_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_21));
  assign mux_27_nl = MUX_s_1_2_2(nor_508_nl, and_tmp_21, or_1_cse);
  assign and_dcpl_342 = mux_27_nl & and_dcpl_31 & and_dcpl_29;
  assign nor_500_nl = ~(and_dcpl_30 | (~ or_tmp_2));
  assign or_61_nl = (rem_12cyc_st_9_1_0!=2'b00) | (rem_12cyc_st_9_3_2!=2'b00);
  assign mux_tmp_26 = MUX_s_1_2_2(nor_500_nl, or_tmp_2, or_61_nl);
  assign nor_501_nl = ~(and_dcpl_57 | (~ mux_tmp_26));
  assign mux_tmp_27 = MUX_s_1_2_2(nor_501_nl, mux_tmp_26, or_48_cse);
  assign nor_502_nl = ~(and_dcpl_84 | (~ mux_tmp_27));
  assign mux_tmp_28 = MUX_s_1_2_2(nor_502_nl, mux_tmp_27, or_37_cse);
  assign nor_503_nl = ~(and_dcpl_111 | (~ mux_tmp_28));
  assign mux_31_nl = MUX_s_1_2_2(nor_503_nl, mux_tmp_28, or_28_cse);
  assign and_tmp_25 = or_6_cse & or_10_cse & or_15_cse & or_21_cse & mux_31_nl;
  assign nor_504_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_25));
  assign mux_32_nl = MUX_s_1_2_2(nor_504_nl, and_tmp_25, or_1_cse);
  assign and_dcpl_348 = mux_32_nl & and_dcpl_4 & and_dcpl_2;
  assign and_tmp_35 = ((~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b00)
      | (rem_12cyc_1_0!=2'b00)) & ((~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b00)
      | (rem_12cyc_st_7_3_2!=2'b00)) & ((~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b00)
      | (rem_12cyc_st_8_3_2!=2'b00)) & ((~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b00)
      | (rem_12cyc_st_9_3_2!=2'b00)) & or_6_cse & or_10_cse & or_15_cse & or_21_cse
      & ((~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b00) | (rem_12cyc_st_6_3_2!=2'b00))
      & ((~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b00) | (rem_12cyc_st_10_3_2!=2'b00))
      & ((acc_tmp!=2'b00) | (acc_1_tmp[1:0]!=2'b00) | (~ ccs_ccore_start_rsci_idat));
  assign and_dcpl_355 = (acc_1_tmp[1:0]==2'b01);
  assign and_dcpl_356 = and_dcpl_293 & and_dcpl_355;
  assign and_dcpl_358 = (rem_12cyc_st_2_1_0[0]) & main_stage_0_3 & asn_itm_2;
  assign or_tmp_80 = (rem_12cyc_1_0!=2'b01) | (rem_12cyc_3_2!=2'b00) | not_tmp_54;
  assign or_83_cse = (acc_1_tmp[1:0]!=2'b01) | (acc_tmp!=2'b00);
  assign nor_499_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_80));
  assign mux_33_nl = MUX_s_1_2_2(nor_499_nl, or_tmp_80, or_83_cse);
  assign and_dcpl_360 = mux_33_nl & and_dcpl_358 & and_dcpl_296;
  assign and_dcpl_362 = (rem_12cyc_st_3_1_0[0]) & main_stage_0_4 & asn_itm_3;
  assign nand_276_cse = ~(asn_itm_2 & main_stage_0_3 & (rem_12cyc_st_2_1_0[0]));
  assign or_88_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2!=2'b00);
  assign and_1168_nl = nand_276_cse & or_tmp_80;
  assign mux_tmp_32 = MUX_s_1_2_2(and_1168_nl, or_tmp_80, or_88_cse);
  assign nor_498_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_32));
  assign mux_35_nl = MUX_s_1_2_2(nor_498_nl, mux_tmp_32, or_83_cse);
  assign and_dcpl_364 = mux_35_nl & and_dcpl_362 & and_dcpl_302;
  assign and_dcpl_366 = (rem_12cyc_st_4_1_0[0]) & main_stage_0_5 & asn_itm_4;
  assign nand_274_cse = ~(asn_itm_3 & main_stage_0_4 & (rem_12cyc_st_3_1_0[0]));
  assign or_93_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2!=2'b00);
  assign and_1166_nl = nand_274_cse & or_tmp_80;
  assign mux_tmp_34 = MUX_s_1_2_2(and_1166_nl, or_tmp_80, or_93_cse);
  assign and_1167_nl = nand_276_cse & mux_tmp_34;
  assign mux_tmp_35 = MUX_s_1_2_2(and_1167_nl, mux_tmp_34, or_88_cse);
  assign nor_497_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_35));
  assign mux_38_nl = MUX_s_1_2_2(nor_497_nl, mux_tmp_35, or_83_cse);
  assign and_dcpl_368 = mux_38_nl & and_dcpl_366 & and_dcpl_308;
  assign and_dcpl_370 = (rem_12cyc_st_5_1_0[0]) & main_stage_0_6 & asn_itm_5;
  assign nand_271_cse = ~(asn_itm_4 & main_stage_0_5 & (rem_12cyc_st_4_1_0[0]));
  assign or_100_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2!=2'b00);
  assign and_1163_nl = nand_271_cse & or_tmp_80;
  assign mux_tmp_37 = MUX_s_1_2_2(and_1163_nl, or_tmp_80, or_100_cse);
  assign and_1164_nl = nand_274_cse & mux_tmp_37;
  assign mux_tmp_38 = MUX_s_1_2_2(and_1164_nl, mux_tmp_37, or_93_cse);
  assign and_1165_nl = nand_276_cse & mux_tmp_38;
  assign mux_tmp_39 = MUX_s_1_2_2(and_1165_nl, mux_tmp_38, or_88_cse);
  assign nor_496_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_39));
  assign mux_42_nl = MUX_s_1_2_2(nor_496_nl, mux_tmp_39, or_83_cse);
  assign and_dcpl_372 = mux_42_nl & and_dcpl_370 & and_dcpl_314;
  assign nand_267_cse = ~(asn_itm_5 & main_stage_0_6 & (rem_12cyc_st_5_1_0[0]));
  assign or_109_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2!=2'b00);
  assign and_1159_nl = nand_267_cse & or_tmp_80;
  assign mux_tmp_41 = MUX_s_1_2_2(and_1159_nl, or_tmp_80, or_109_cse);
  assign and_1160_nl = nand_271_cse & mux_tmp_41;
  assign mux_tmp_42 = MUX_s_1_2_2(and_1160_nl, mux_tmp_41, or_100_cse);
  assign and_1161_nl = nand_274_cse & mux_tmp_42;
  assign mux_tmp_43 = MUX_s_1_2_2(and_1161_nl, mux_tmp_42, or_93_cse);
  assign and_1162_nl = nand_276_cse & mux_tmp_43;
  assign mux_tmp_44 = MUX_s_1_2_2(and_1162_nl, mux_tmp_43, or_88_cse);
  assign nor_495_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_44));
  assign mux_47_nl = MUX_s_1_2_2(nor_495_nl, mux_tmp_44, or_83_cse);
  assign and_dcpl_376 = mux_47_nl & and_dcpl_112 & and_dcpl_115;
  assign or_120_cse = (rem_12cyc_st_6_1_0!=2'b01) | (rem_12cyc_st_6_3_2!=2'b00);
  assign nor_493_nl = ~(and_dcpl_111 | (~ or_tmp_80));
  assign mux_tmp_46 = MUX_s_1_2_2(nor_493_nl, or_tmp_80, or_120_cse);
  assign and_1155_nl = nand_267_cse & mux_tmp_46;
  assign mux_tmp_47 = MUX_s_1_2_2(and_1155_nl, mux_tmp_46, or_109_cse);
  assign and_1156_nl = nand_271_cse & mux_tmp_47;
  assign mux_tmp_48 = MUX_s_1_2_2(and_1156_nl, mux_tmp_47, or_100_cse);
  assign and_1157_nl = nand_274_cse & mux_tmp_48;
  assign mux_tmp_49 = MUX_s_1_2_2(and_1157_nl, mux_tmp_48, or_93_cse);
  assign and_1158_nl = nand_276_cse & mux_tmp_49;
  assign mux_tmp_50 = MUX_s_1_2_2(and_1158_nl, mux_tmp_49, or_88_cse);
  assign nor_494_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_50));
  assign mux_53_nl = MUX_s_1_2_2(nor_494_nl, mux_tmp_50, or_83_cse);
  assign and_dcpl_379 = mux_53_nl & and_dcpl_85 & and_dcpl_87;
  assign or_133_cse = (rem_12cyc_st_7_1_0!=2'b01) | (rem_12cyc_st_7_3_2!=2'b00);
  assign nor_490_nl = ~(and_dcpl_84 | (~ or_tmp_80));
  assign mux_tmp_52 = MUX_s_1_2_2(nor_490_nl, or_tmp_80, or_133_cse);
  assign nor_491_nl = ~(and_dcpl_111 | (~ mux_tmp_52));
  assign mux_tmp_53 = MUX_s_1_2_2(nor_491_nl, mux_tmp_52, or_120_cse);
  assign and_1151_nl = nand_267_cse & mux_tmp_53;
  assign mux_tmp_54 = MUX_s_1_2_2(and_1151_nl, mux_tmp_53, or_109_cse);
  assign and_1152_nl = nand_271_cse & mux_tmp_54;
  assign mux_tmp_55 = MUX_s_1_2_2(and_1152_nl, mux_tmp_54, or_100_cse);
  assign and_1153_nl = nand_274_cse & mux_tmp_55;
  assign mux_tmp_56 = MUX_s_1_2_2(and_1153_nl, mux_tmp_55, or_93_cse);
  assign and_1154_nl = nand_276_cse & mux_tmp_56;
  assign mux_tmp_57 = MUX_s_1_2_2(and_1154_nl, mux_tmp_56, or_88_cse);
  assign nor_492_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_57));
  assign mux_60_nl = MUX_s_1_2_2(nor_492_nl, mux_tmp_57, or_83_cse);
  assign and_dcpl_382 = mux_60_nl & and_dcpl_58 & and_dcpl_60;
  assign or_148_cse = (rem_12cyc_st_8_1_0!=2'b01) | (rem_12cyc_st_8_3_2!=2'b00);
  assign nor_486_nl = ~(and_dcpl_57 | (~ or_tmp_80));
  assign mux_tmp_59 = MUX_s_1_2_2(nor_486_nl, or_tmp_80, or_148_cse);
  assign nor_487_nl = ~(and_dcpl_84 | (~ mux_tmp_59));
  assign mux_tmp_60 = MUX_s_1_2_2(nor_487_nl, mux_tmp_59, or_133_cse);
  assign nor_488_nl = ~(and_dcpl_111 | (~ mux_tmp_60));
  assign mux_tmp_61 = MUX_s_1_2_2(nor_488_nl, mux_tmp_60, or_120_cse);
  assign and_1147_nl = nand_267_cse & mux_tmp_61;
  assign mux_tmp_62 = MUX_s_1_2_2(and_1147_nl, mux_tmp_61, or_109_cse);
  assign and_1148_nl = nand_271_cse & mux_tmp_62;
  assign mux_tmp_63 = MUX_s_1_2_2(and_1148_nl, mux_tmp_62, or_100_cse);
  assign and_1149_nl = nand_274_cse & mux_tmp_63;
  assign mux_tmp_64 = MUX_s_1_2_2(and_1149_nl, mux_tmp_63, or_93_cse);
  assign and_1150_nl = nand_276_cse & mux_tmp_64;
  assign mux_tmp_65 = MUX_s_1_2_2(and_1150_nl, mux_tmp_64, or_88_cse);
  assign nor_489_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_65));
  assign mux_68_nl = MUX_s_1_2_2(nor_489_nl, mux_tmp_65, or_83_cse);
  assign and_dcpl_385 = mux_68_nl & and_dcpl_31 & and_dcpl_33;
  assign nor_481_nl = ~(and_dcpl_30 | (~ or_tmp_80));
  assign or_165_nl = (rem_12cyc_st_9_1_0!=2'b01) | (rem_12cyc_st_9_3_2!=2'b00);
  assign mux_tmp_67 = MUX_s_1_2_2(nor_481_nl, or_tmp_80, or_165_nl);
  assign nor_482_nl = ~(and_dcpl_57 | (~ mux_tmp_67));
  assign mux_tmp_68 = MUX_s_1_2_2(nor_482_nl, mux_tmp_67, or_148_cse);
  assign nor_483_nl = ~(and_dcpl_84 | (~ mux_tmp_68));
  assign mux_tmp_69 = MUX_s_1_2_2(nor_483_nl, mux_tmp_68, or_133_cse);
  assign nor_484_nl = ~(and_dcpl_111 | (~ mux_tmp_69));
  assign mux_tmp_70 = MUX_s_1_2_2(nor_484_nl, mux_tmp_69, or_120_cse);
  assign and_1143_nl = nand_267_cse & mux_tmp_70;
  assign mux_tmp_71 = MUX_s_1_2_2(and_1143_nl, mux_tmp_70, or_109_cse);
  assign and_1144_nl = nand_271_cse & mux_tmp_71;
  assign mux_tmp_72 = MUX_s_1_2_2(and_1144_nl, mux_tmp_71, or_100_cse);
  assign and_1145_nl = nand_274_cse & mux_tmp_72;
  assign mux_tmp_73 = MUX_s_1_2_2(and_1145_nl, mux_tmp_72, or_93_cse);
  assign and_1146_nl = nand_276_cse & mux_tmp_73;
  assign mux_tmp_74 = MUX_s_1_2_2(and_1146_nl, mux_tmp_73, or_88_cse);
  assign nor_485_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_74));
  assign mux_77_nl = MUX_s_1_2_2(nor_485_nl, mux_tmp_74, or_83_cse);
  assign and_dcpl_388 = mux_77_nl & and_dcpl_4 & and_dcpl_6;
  assign nand_250_cse = ~((acc_1_tmp[0]) & ccs_ccore_start_rsci_idat);
  assign and_tmp_44 = ((~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b01)
      | (rem_12cyc_st_7_3_2!=2'b00)) & ((~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b01)
      | (rem_12cyc_st_8_3_2!=2'b00)) & ((~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b01)
      | (rem_12cyc_st_9_3_2!=2'b00)) & ((~ main_stage_0_3) | (~ asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b01)
      | (rem_12cyc_st_2_3_2!=2'b00)) & ((~ main_stage_0_4) | (~ asn_itm_3) | (rem_12cyc_st_3_1_0!=2'b01)
      | (rem_12cyc_st_3_3_2!=2'b00)) & ((~ main_stage_0_5) | (~ asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b01)
      | (rem_12cyc_st_4_3_2!=2'b00)) & ((~ main_stage_0_6) | (~ asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b01)
      | (rem_12cyc_st_5_3_2!=2'b00)) & ((~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b01)
      | (rem_12cyc_st_6_3_2!=2'b00)) & ((~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b01)
      | (rem_12cyc_st_10_3_2!=2'b00)) & ((acc_tmp!=2'b00) | (acc_1_tmp[1]) | nand_250_cse);
  assign nor_480_nl = ~((rem_12cyc_1_0[0]) | (~ and_tmp_44));
  assign or_175_nl = (~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b00)
      | (rem_12cyc_1_0[1]);
  assign mux_tmp_76 = MUX_s_1_2_2(nor_480_nl, and_tmp_44, or_175_nl);
  assign and_dcpl_393 = (acc_1_tmp[1:0]==2'b10);
  assign and_dcpl_394 = and_dcpl_293 & and_dcpl_393;
  assign and_dcpl_395 = and_dcpl_295 & (rem_12cyc_st_2_1_0[1]);
  assign or_tmp_185 = (rem_12cyc_1_0!=2'b10) | (rem_12cyc_3_2!=2'b00) | not_tmp_54;
  assign or_190_cse = (acc_1_tmp[1:0]!=2'b10) | (acc_tmp!=2'b00);
  assign nor_479_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_185));
  assign mux_79_nl = MUX_s_1_2_2(nor_479_nl, or_tmp_185, or_190_cse);
  assign and_dcpl_397 = mux_79_nl & and_dcpl_298 & and_dcpl_395;
  assign and_dcpl_398 = and_dcpl_301 & (rem_12cyc_st_3_1_0[1]);
  assign or_195_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2!=2'b00) |
      (~ asn_itm_2) | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp_45 = or_195_cse & or_tmp_185;
  assign nor_478_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_45));
  assign mux_80_nl = MUX_s_1_2_2(nor_478_nl, and_tmp_45, or_190_cse);
  assign and_dcpl_400 = mux_80_nl & and_dcpl_304 & and_dcpl_398;
  assign and_dcpl_401 = and_dcpl_307 & (rem_12cyc_st_4_1_0[1]);
  assign or_199_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2!=2'b00) |
      (~ asn_itm_3) | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_47 = or_195_cse & or_199_cse & or_tmp_185;
  assign nor_477_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_47));
  assign mux_81_nl = MUX_s_1_2_2(nor_477_nl, and_tmp_47, or_190_cse);
  assign and_dcpl_403 = mux_81_nl & and_dcpl_310 & and_dcpl_401;
  assign and_dcpl_404 = and_dcpl_313 & (rem_12cyc_st_5_1_0[1]);
  assign or_204_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2!=2'b00) |
      (~ asn_itm_4) | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_50 = or_195_cse & or_199_cse & or_204_cse & or_tmp_185;
  assign nor_476_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_50));
  assign mux_82_nl = MUX_s_1_2_2(nor_476_nl, and_tmp_50, or_190_cse);
  assign and_dcpl_406 = mux_82_nl & and_dcpl_316 & and_dcpl_404;
  assign or_210_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2!=2'b00) |
      (~ asn_itm_5) | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_54 = or_195_cse & or_199_cse & or_204_cse & or_210_cse & or_tmp_185;
  assign nor_475_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_54));
  assign mux_83_nl = MUX_s_1_2_2(nor_475_nl, and_tmp_54, or_190_cse);
  assign and_dcpl_409 = mux_83_nl & and_dcpl_112 & and_dcpl_117;
  assign or_217_cse = (rem_12cyc_st_6_1_0!=2'b10) | (rem_12cyc_st_6_3_2!=2'b00);
  assign nor_473_nl = ~(and_dcpl_111 | (~ or_tmp_185));
  assign mux_84_nl = MUX_s_1_2_2(nor_473_nl, or_tmp_185, or_217_cse);
  assign and_tmp_58 = or_195_cse & or_199_cse & or_204_cse & or_210_cse & mux_84_nl;
  assign nor_474_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_58));
  assign mux_85_nl = MUX_s_1_2_2(nor_474_nl, and_tmp_58, or_190_cse);
  assign and_dcpl_413 = mux_85_nl & and_dcpl_85 & and_dcpl_90;
  assign or_226_cse = (rem_12cyc_st_7_1_0!=2'b10) | (rem_12cyc_st_7_3_2!=2'b00);
  assign nor_470_nl = ~(and_dcpl_84 | (~ or_tmp_185));
  assign mux_tmp_84 = MUX_s_1_2_2(nor_470_nl, or_tmp_185, or_226_cse);
  assign nor_471_nl = ~(and_dcpl_111 | (~ mux_tmp_84));
  assign mux_87_nl = MUX_s_1_2_2(nor_471_nl, mux_tmp_84, or_217_cse);
  assign and_tmp_62 = or_195_cse & or_199_cse & or_204_cse & or_210_cse & mux_87_nl;
  assign nor_472_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_62));
  assign mux_88_nl = MUX_s_1_2_2(nor_472_nl, and_tmp_62, or_190_cse);
  assign and_dcpl_417 = mux_88_nl & and_dcpl_58 & and_dcpl_63;
  assign or_237_cse = (rem_12cyc_st_8_1_0!=2'b10) | (rem_12cyc_st_8_3_2!=2'b00);
  assign nor_466_nl = ~(and_dcpl_57 | (~ or_tmp_185));
  assign mux_tmp_87 = MUX_s_1_2_2(nor_466_nl, or_tmp_185, or_237_cse);
  assign nor_467_nl = ~(and_dcpl_84 | (~ mux_tmp_87));
  assign mux_tmp_88 = MUX_s_1_2_2(nor_467_nl, mux_tmp_87, or_226_cse);
  assign nor_468_nl = ~(and_dcpl_111 | (~ mux_tmp_88));
  assign mux_91_nl = MUX_s_1_2_2(nor_468_nl, mux_tmp_88, or_217_cse);
  assign and_tmp_66 = or_195_cse & or_199_cse & or_204_cse & or_210_cse & mux_91_nl;
  assign nor_469_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_66));
  assign mux_92_nl = MUX_s_1_2_2(nor_469_nl, and_tmp_66, or_190_cse);
  assign and_dcpl_421 = mux_92_nl & and_dcpl_31 & and_dcpl_36;
  assign nor_461_nl = ~(and_dcpl_30 | (~ or_tmp_185));
  assign or_250_nl = (rem_12cyc_st_9_1_0!=2'b10) | (rem_12cyc_st_9_3_2!=2'b00);
  assign mux_tmp_91 = MUX_s_1_2_2(nor_461_nl, or_tmp_185, or_250_nl);
  assign nor_462_nl = ~(and_dcpl_57 | (~ mux_tmp_91));
  assign mux_tmp_92 = MUX_s_1_2_2(nor_462_nl, mux_tmp_91, or_237_cse);
  assign nor_463_nl = ~(and_dcpl_84 | (~ mux_tmp_92));
  assign mux_tmp_93 = MUX_s_1_2_2(nor_463_nl, mux_tmp_92, or_226_cse);
  assign nor_464_nl = ~(and_dcpl_111 | (~ mux_tmp_93));
  assign mux_96_nl = MUX_s_1_2_2(nor_464_nl, mux_tmp_93, or_217_cse);
  assign and_tmp_70 = or_195_cse & or_199_cse & or_204_cse & or_210_cse & mux_96_nl;
  assign nor_465_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_70));
  assign mux_97_nl = MUX_s_1_2_2(nor_465_nl, and_tmp_70, or_190_cse);
  assign and_dcpl_425 = mux_97_nl & and_dcpl_4 & and_dcpl_9;
  assign and_tmp_80 = ((~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b00)
      | (rem_12cyc_1_0!=2'b10)) & ((~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b10)
      | (rem_12cyc_st_7_3_2!=2'b00)) & ((~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b10)
      | (rem_12cyc_st_8_3_2!=2'b00)) & ((~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b10)
      | (rem_12cyc_st_9_3_2!=2'b00)) & or_195_cse & or_199_cse & or_204_cse & or_210_cse
      & ((~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b10) | (rem_12cyc_st_6_3_2!=2'b00))
      & ((~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b10) | (rem_12cyc_st_10_3_2!=2'b00))
      & ((acc_tmp!=2'b00) | (acc_1_tmp[1:0]!=2'b10) | (~ ccs_ccore_start_rsci_idat));
  assign and_dcpl_430 = (acc_1_tmp[1:0]==2'b11);
  assign and_dcpl_431 = and_dcpl_293 & and_dcpl_430;
  assign or_tmp_263 = (rem_12cyc_1_0!=2'b11) | (rem_12cyc_3_2!=2'b00) | not_tmp_54;
  assign or_270_cse = (acc_1_tmp[1:0]!=2'b11) | (acc_tmp!=2'b00);
  assign nor_460_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_263));
  assign mux_98_nl = MUX_s_1_2_2(nor_460_nl, or_tmp_263, or_270_cse);
  assign and_dcpl_433 = mux_98_nl & and_dcpl_358 & and_dcpl_395;
  assign or_275_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2!=2'b00);
  assign and_1142_nl = nand_276_cse & or_tmp_263;
  assign mux_tmp_97 = MUX_s_1_2_2(and_1142_nl, or_tmp_263, or_275_cse);
  assign nor_459_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_97));
  assign mux_100_nl = MUX_s_1_2_2(nor_459_nl, mux_tmp_97, or_270_cse);
  assign and_dcpl_435 = mux_100_nl & and_dcpl_362 & and_dcpl_398;
  assign or_280_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2!=2'b00);
  assign and_1140_nl = nand_274_cse & or_tmp_263;
  assign mux_tmp_99 = MUX_s_1_2_2(and_1140_nl, or_tmp_263, or_280_cse);
  assign and_1141_nl = nand_276_cse & mux_tmp_99;
  assign mux_tmp_100 = MUX_s_1_2_2(and_1141_nl, mux_tmp_99, or_275_cse);
  assign nor_458_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_100));
  assign mux_103_nl = MUX_s_1_2_2(nor_458_nl, mux_tmp_100, or_270_cse);
  assign and_dcpl_437 = mux_103_nl & and_dcpl_366 & and_dcpl_401;
  assign or_287_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2!=2'b00);
  assign and_1137_nl = nand_271_cse & or_tmp_263;
  assign mux_tmp_102 = MUX_s_1_2_2(and_1137_nl, or_tmp_263, or_287_cse);
  assign and_1138_nl = nand_274_cse & mux_tmp_102;
  assign mux_tmp_103 = MUX_s_1_2_2(and_1138_nl, mux_tmp_102, or_280_cse);
  assign and_1139_nl = nand_276_cse & mux_tmp_103;
  assign mux_tmp_104 = MUX_s_1_2_2(and_1139_nl, mux_tmp_103, or_275_cse);
  assign nor_457_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_104));
  assign mux_107_nl = MUX_s_1_2_2(nor_457_nl, mux_tmp_104, or_270_cse);
  assign and_dcpl_439 = mux_107_nl & and_dcpl_370 & and_dcpl_404;
  assign or_296_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2!=2'b00);
  assign and_1133_nl = nand_267_cse & or_tmp_263;
  assign mux_tmp_106 = MUX_s_1_2_2(and_1133_nl, or_tmp_263, or_296_cse);
  assign and_1134_nl = nand_271_cse & mux_tmp_106;
  assign mux_tmp_107 = MUX_s_1_2_2(and_1134_nl, mux_tmp_106, or_287_cse);
  assign and_1135_nl = nand_274_cse & mux_tmp_107;
  assign mux_tmp_108 = MUX_s_1_2_2(and_1135_nl, mux_tmp_107, or_280_cse);
  assign and_1136_nl = nand_276_cse & mux_tmp_108;
  assign mux_tmp_109 = MUX_s_1_2_2(and_1136_nl, mux_tmp_108, or_275_cse);
  assign nor_456_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_109));
  assign mux_112_nl = MUX_s_1_2_2(nor_456_nl, mux_tmp_109, or_270_cse);
  assign and_dcpl_442 = mux_112_nl & and_dcpl_112 & and_dcpl_119;
  assign or_307_cse = (rem_12cyc_st_6_1_0!=2'b11) | (rem_12cyc_st_6_3_2!=2'b00);
  assign nor_454_nl = ~(and_dcpl_111 | (~ or_tmp_263));
  assign mux_tmp_111 = MUX_s_1_2_2(nor_454_nl, or_tmp_263, or_307_cse);
  assign and_1129_nl = nand_267_cse & mux_tmp_111;
  assign mux_tmp_112 = MUX_s_1_2_2(and_1129_nl, mux_tmp_111, or_296_cse);
  assign and_1130_nl = nand_271_cse & mux_tmp_112;
  assign mux_tmp_113 = MUX_s_1_2_2(and_1130_nl, mux_tmp_112, or_287_cse);
  assign and_1131_nl = nand_274_cse & mux_tmp_113;
  assign mux_tmp_114 = MUX_s_1_2_2(and_1131_nl, mux_tmp_113, or_280_cse);
  assign and_1132_nl = nand_276_cse & mux_tmp_114;
  assign mux_tmp_115 = MUX_s_1_2_2(and_1132_nl, mux_tmp_114, or_275_cse);
  assign nor_455_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_115));
  assign mux_118_nl = MUX_s_1_2_2(nor_455_nl, mux_tmp_115, or_270_cse);
  assign and_dcpl_445 = mux_118_nl & and_dcpl_85 & and_dcpl_92;
  assign or_320_cse = (rem_12cyc_st_7_1_0!=2'b11) | (rem_12cyc_st_7_3_2!=2'b00);
  assign nor_451_nl = ~(and_dcpl_84 | (~ or_tmp_263));
  assign mux_tmp_117 = MUX_s_1_2_2(nor_451_nl, or_tmp_263, or_320_cse);
  assign nor_452_nl = ~(and_dcpl_111 | (~ mux_tmp_117));
  assign mux_tmp_118 = MUX_s_1_2_2(nor_452_nl, mux_tmp_117, or_307_cse);
  assign and_1125_nl = nand_267_cse & mux_tmp_118;
  assign mux_tmp_119 = MUX_s_1_2_2(and_1125_nl, mux_tmp_118, or_296_cse);
  assign and_1126_nl = nand_271_cse & mux_tmp_119;
  assign mux_tmp_120 = MUX_s_1_2_2(and_1126_nl, mux_tmp_119, or_287_cse);
  assign and_1127_nl = nand_274_cse & mux_tmp_120;
  assign mux_tmp_121 = MUX_s_1_2_2(and_1127_nl, mux_tmp_120, or_280_cse);
  assign and_1128_nl = nand_276_cse & mux_tmp_121;
  assign mux_tmp_122 = MUX_s_1_2_2(and_1128_nl, mux_tmp_121, or_275_cse);
  assign nor_453_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_122));
  assign mux_125_nl = MUX_s_1_2_2(nor_453_nl, mux_tmp_122, or_270_cse);
  assign and_dcpl_448 = mux_125_nl & and_dcpl_58 & and_dcpl_65;
  assign or_335_cse = (rem_12cyc_st_8_1_0!=2'b11) | (rem_12cyc_st_8_3_2!=2'b00);
  assign nor_447_nl = ~(and_dcpl_57 | (~ or_tmp_263));
  assign mux_tmp_124 = MUX_s_1_2_2(nor_447_nl, or_tmp_263, or_335_cse);
  assign nor_448_nl = ~(and_dcpl_84 | (~ mux_tmp_124));
  assign mux_tmp_125 = MUX_s_1_2_2(nor_448_nl, mux_tmp_124, or_320_cse);
  assign nor_449_nl = ~(and_dcpl_111 | (~ mux_tmp_125));
  assign mux_tmp_126 = MUX_s_1_2_2(nor_449_nl, mux_tmp_125, or_307_cse);
  assign and_1121_nl = nand_267_cse & mux_tmp_126;
  assign mux_tmp_127 = MUX_s_1_2_2(and_1121_nl, mux_tmp_126, or_296_cse);
  assign and_1122_nl = nand_271_cse & mux_tmp_127;
  assign mux_tmp_128 = MUX_s_1_2_2(and_1122_nl, mux_tmp_127, or_287_cse);
  assign and_1123_nl = nand_274_cse & mux_tmp_128;
  assign mux_tmp_129 = MUX_s_1_2_2(and_1123_nl, mux_tmp_128, or_280_cse);
  assign and_1124_nl = nand_276_cse & mux_tmp_129;
  assign mux_tmp_130 = MUX_s_1_2_2(and_1124_nl, mux_tmp_129, or_275_cse);
  assign nor_450_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_130));
  assign mux_133_nl = MUX_s_1_2_2(nor_450_nl, mux_tmp_130, or_270_cse);
  assign and_dcpl_451 = mux_133_nl & and_dcpl_31 & and_dcpl_38;
  assign nor_442_nl = ~(and_dcpl_30 | (~ or_tmp_263));
  assign or_352_nl = (rem_12cyc_st_9_1_0!=2'b11) | (rem_12cyc_st_9_3_2!=2'b00);
  assign mux_tmp_132 = MUX_s_1_2_2(nor_442_nl, or_tmp_263, or_352_nl);
  assign nor_443_nl = ~(and_dcpl_57 | (~ mux_tmp_132));
  assign mux_tmp_133 = MUX_s_1_2_2(nor_443_nl, mux_tmp_132, or_335_cse);
  assign nor_444_nl = ~(and_dcpl_84 | (~ mux_tmp_133));
  assign mux_tmp_134 = MUX_s_1_2_2(nor_444_nl, mux_tmp_133, or_320_cse);
  assign nor_445_nl = ~(and_dcpl_111 | (~ mux_tmp_134));
  assign mux_tmp_135 = MUX_s_1_2_2(nor_445_nl, mux_tmp_134, or_307_cse);
  assign and_1117_nl = nand_267_cse & mux_tmp_135;
  assign mux_tmp_136 = MUX_s_1_2_2(and_1117_nl, mux_tmp_135, or_296_cse);
  assign and_1118_nl = nand_271_cse & mux_tmp_136;
  assign mux_tmp_137 = MUX_s_1_2_2(and_1118_nl, mux_tmp_136, or_287_cse);
  assign and_1119_nl = nand_274_cse & mux_tmp_137;
  assign mux_tmp_138 = MUX_s_1_2_2(and_1119_nl, mux_tmp_137, or_280_cse);
  assign and_1120_nl = nand_276_cse & mux_tmp_138;
  assign mux_tmp_139 = MUX_s_1_2_2(and_1120_nl, mux_tmp_138, or_275_cse);
  assign nor_446_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_139));
  assign mux_142_nl = MUX_s_1_2_2(nor_446_nl, mux_tmp_139, or_270_cse);
  assign and_dcpl_454 = mux_142_nl & and_dcpl_4 & and_dcpl_11;
  assign nand_222_cse = ~((acc_1_tmp[1:0]==2'b11) & ccs_ccore_start_rsci_idat);
  assign and_tmp_89 = ((~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b11)
      | (rem_12cyc_st_7_3_2!=2'b00)) & ((~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b11)
      | (rem_12cyc_st_8_3_2!=2'b00)) & ((~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b11)
      | (rem_12cyc_st_9_3_2!=2'b00)) & ((~ main_stage_0_3) | (~ asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b11)
      | (rem_12cyc_st_2_3_2!=2'b00)) & ((~ main_stage_0_4) | (~ asn_itm_3) | (rem_12cyc_st_3_1_0!=2'b11)
      | (rem_12cyc_st_3_3_2!=2'b00)) & ((~ main_stage_0_5) | (~ asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b11)
      | (rem_12cyc_st_4_3_2!=2'b00)) & ((~ main_stage_0_6) | (~ asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b11)
      | (rem_12cyc_st_5_3_2!=2'b00)) & ((~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b11)
      | (rem_12cyc_st_6_3_2!=2'b00)) & ((~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b11)
      | (rem_12cyc_st_10_3_2!=2'b00)) & ((acc_tmp!=2'b00) | nand_222_cse);
  assign nand_223_cse = ~((rem_12cyc_1_0==2'b11));
  assign and_1116_nl = nand_223_cse & and_tmp_89;
  assign or_362_nl = (~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b00);
  assign mux_tmp_141 = MUX_s_1_2_2(and_1116_nl, and_tmp_89, or_362_nl);
  assign and_dcpl_460 = ccs_ccore_start_rsci_idat & (acc_tmp==2'b01);
  assign and_dcpl_461 = and_dcpl_460 & and_dcpl_291;
  assign and_dcpl_462 = (rem_12cyc_st_2_3_2==2'b01);
  assign and_dcpl_463 = and_dcpl_462 & (~ (rem_12cyc_st_2_1_0[1]));
  assign not_tmp_332 = ~((rem_12cyc_3_2[0]) & asn_itm_1 & main_stage_0_2);
  assign or_tmp_368 = (rem_12cyc_1_0!=2'b00) | (rem_12cyc_3_2[1]) | not_tmp_332;
  assign nand_281_cse = ~((acc_tmp[0]) & ccs_ccore_start_rsci_idat);
  assign or_377_cse = (acc_1_tmp[1:0]!=2'b00) | (acc_tmp[1]);
  assign and_1172_nl = nand_281_cse & or_tmp_368;
  assign mux_144_nl = MUX_s_1_2_2(and_1172_nl, or_tmp_368, or_377_cse);
  assign and_dcpl_465 = mux_144_nl & and_dcpl_298 & and_dcpl_463;
  assign and_dcpl_466 = (rem_12cyc_st_3_3_2==2'b01);
  assign and_dcpl_467 = and_dcpl_466 & (~ (rem_12cyc_st_3_1_0[1]));
  assign or_382_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2!=2'b01) | (~
      asn_itm_2) | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp_90 = or_382_cse & or_tmp_368;
  assign and_1114_nl = nand_281_cse & and_tmp_90;
  assign mux_145_nl = MUX_s_1_2_2(and_1114_nl, and_tmp_90, or_377_cse);
  assign and_dcpl_469 = mux_145_nl & and_dcpl_304 & and_dcpl_467;
  assign and_dcpl_470 = (rem_12cyc_st_4_3_2==2'b01);
  assign and_dcpl_471 = and_dcpl_470 & (~ (rem_12cyc_st_4_1_0[1]));
  assign or_386_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2!=2'b01) | (~
      asn_itm_3) | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_92 = or_382_cse & or_386_cse & or_tmp_368;
  assign and_1113_nl = nand_281_cse & and_tmp_92;
  assign mux_146_nl = MUX_s_1_2_2(and_1113_nl, and_tmp_92, or_377_cse);
  assign and_dcpl_473 = mux_146_nl & and_dcpl_310 & and_dcpl_471;
  assign and_dcpl_474 = (rem_12cyc_st_5_3_2==2'b01);
  assign and_dcpl_475 = and_dcpl_474 & (~ (rem_12cyc_st_5_1_0[1]));
  assign or_391_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2!=2'b01) | (~
      asn_itm_4) | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_95 = or_382_cse & or_386_cse & or_391_cse & or_tmp_368;
  assign and_1112_nl = nand_281_cse & and_tmp_95;
  assign mux_147_nl = MUX_s_1_2_2(and_1112_nl, and_tmp_95, or_377_cse);
  assign and_dcpl_477 = mux_147_nl & and_dcpl_316 & and_dcpl_475;
  assign or_397_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2!=2'b01) | (~
      asn_itm_5) | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_99 = or_382_cse & or_386_cse & or_391_cse & or_397_cse & or_tmp_368;
  assign and_1111_nl = nand_281_cse & and_tmp_99;
  assign mux_148_nl = MUX_s_1_2_2(and_1111_nl, and_tmp_99, or_377_cse);
  assign and_dcpl_480 = mux_148_nl & and_dcpl_121 & and_dcpl_110;
  assign nand_215_cse = ~((rem_12cyc_st_6_3_2[0]) & asn_itm_6 & main_stage_0_7);
  assign or_404_cse = (rem_12cyc_st_6_1_0!=2'b00) | (rem_12cyc_st_6_3_2[1]);
  assign and_1109_nl = nand_215_cse & or_tmp_368;
  assign mux_149_nl = MUX_s_1_2_2(and_1109_nl, or_tmp_368, or_404_cse);
  assign and_tmp_103 = or_382_cse & or_386_cse & or_391_cse & or_397_cse & mux_149_nl;
  assign and_1110_nl = nand_281_cse & and_tmp_103;
  assign mux_150_nl = MUX_s_1_2_2(and_1110_nl, and_tmp_103, or_377_cse);
  assign and_dcpl_483 = mux_150_nl & and_dcpl_94 & and_dcpl_83;
  assign nand_212_cse = ~((rem_12cyc_st_7_3_2[0]) & asn_itm_7 & main_stage_0_8);
  assign or_413_cse = (rem_12cyc_st_7_1_0!=2'b00) | (rem_12cyc_st_7_3_2[1]);
  assign and_1106_nl = nand_212_cse & or_tmp_368;
  assign mux_tmp_149 = MUX_s_1_2_2(and_1106_nl, or_tmp_368, or_413_cse);
  assign and_1107_nl = nand_215_cse & mux_tmp_149;
  assign mux_152_nl = MUX_s_1_2_2(and_1107_nl, mux_tmp_149, or_404_cse);
  assign and_tmp_107 = or_382_cse & or_386_cse & or_391_cse & or_397_cse & mux_152_nl;
  assign and_1108_nl = nand_281_cse & and_tmp_107;
  assign mux_153_nl = MUX_s_1_2_2(and_1108_nl, and_tmp_107, or_377_cse);
  assign and_dcpl_486 = mux_153_nl & and_dcpl_67 & and_dcpl_56;
  assign nand_208_cse = ~((rem_12cyc_st_8_3_2[0]) & asn_itm_8 & main_stage_0_9);
  assign or_424_cse = (rem_12cyc_st_8_1_0!=2'b00) | (rem_12cyc_st_8_3_2[1]);
  assign and_1102_nl = nand_208_cse & or_tmp_368;
  assign mux_tmp_152 = MUX_s_1_2_2(and_1102_nl, or_tmp_368, or_424_cse);
  assign and_1103_nl = nand_212_cse & mux_tmp_152;
  assign mux_tmp_153 = MUX_s_1_2_2(and_1103_nl, mux_tmp_152, or_413_cse);
  assign and_1104_nl = nand_215_cse & mux_tmp_153;
  assign mux_156_nl = MUX_s_1_2_2(and_1104_nl, mux_tmp_153, or_404_cse);
  assign and_tmp_111 = or_382_cse & or_386_cse & or_391_cse & or_397_cse & mux_156_nl;
  assign and_1105_nl = nand_281_cse & and_tmp_111;
  assign mux_157_nl = MUX_s_1_2_2(and_1105_nl, and_tmp_111, or_377_cse);
  assign and_dcpl_489 = mux_157_nl & and_dcpl_40 & and_dcpl_29;
  assign nand_203_cse = ~((rem_12cyc_st_9_3_2[0]) & asn_itm_9 & main_stage_0_10);
  assign and_1097_nl = nand_203_cse & or_tmp_368;
  assign or_437_nl = (rem_12cyc_st_9_1_0!=2'b00) | (rem_12cyc_st_9_3_2[1]);
  assign mux_tmp_156 = MUX_s_1_2_2(and_1097_nl, or_tmp_368, or_437_nl);
  assign and_1098_nl = nand_208_cse & mux_tmp_156;
  assign mux_tmp_157 = MUX_s_1_2_2(and_1098_nl, mux_tmp_156, or_424_cse);
  assign and_1099_nl = nand_212_cse & mux_tmp_157;
  assign mux_tmp_158 = MUX_s_1_2_2(and_1099_nl, mux_tmp_157, or_413_cse);
  assign and_1100_nl = nand_215_cse & mux_tmp_158;
  assign mux_161_nl = MUX_s_1_2_2(and_1100_nl, mux_tmp_158, or_404_cse);
  assign and_tmp_115 = or_382_cse & or_386_cse & or_391_cse & or_397_cse & mux_161_nl;
  assign and_1101_nl = nand_281_cse & and_tmp_115;
  assign mux_162_nl = MUX_s_1_2_2(and_1101_nl, and_tmp_115, or_377_cse);
  assign and_dcpl_492 = mux_162_nl & and_dcpl_13 & and_dcpl_2;
  assign and_tmp_125 = ((~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b01)
      | (rem_12cyc_1_0!=2'b00)) & ((~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b00)
      | (rem_12cyc_st_7_3_2!=2'b01)) & ((~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b00)
      | (rem_12cyc_st_8_3_2!=2'b01)) & ((~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b00)
      | (rem_12cyc_st_9_3_2!=2'b01)) & or_382_cse & or_386_cse & or_391_cse & or_397_cse
      & ((~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b00) | (rem_12cyc_st_6_3_2!=2'b01))
      & ((~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b00) | (rem_12cyc_st_10_3_2!=2'b01))
      & ((acc_tmp!=2'b01) | (acc_1_tmp[1:0]!=2'b00) | (~ ccs_ccore_start_rsci_idat));
  assign and_dcpl_498 = and_dcpl_460 & and_dcpl_355;
  assign or_tmp_446 = (rem_12cyc_1_0!=2'b01) | (rem_12cyc_3_2[1]) | not_tmp_332;
  assign or_458_cse = (acc_1_tmp[1:0]!=2'b01) | (acc_tmp[1]);
  assign and_1171_nl = nand_281_cse & or_tmp_446;
  assign mux_163_nl = MUX_s_1_2_2(and_1171_nl, or_tmp_446, or_458_cse);
  assign and_dcpl_500 = mux_163_nl & and_dcpl_358 & and_dcpl_463;
  assign or_463_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2!=2'b01);
  assign and_1094_nl = nand_276_cse & or_tmp_446;
  assign mux_tmp_162 = MUX_s_1_2_2(and_1094_nl, or_tmp_446, or_463_cse);
  assign and_1095_nl = nand_281_cse & mux_tmp_162;
  assign mux_165_nl = MUX_s_1_2_2(and_1095_nl, mux_tmp_162, or_458_cse);
  assign and_dcpl_502 = mux_165_nl & and_dcpl_362 & and_dcpl_467;
  assign nand_198_cse = ~((rem_12cyc_st_3_3_2[0]) & asn_itm_3 & main_stage_0_4 &
      (rem_12cyc_st_3_1_0[0]));
  assign or_468_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2[1]);
  assign and_1091_nl = nand_198_cse & or_tmp_446;
  assign mux_tmp_164 = MUX_s_1_2_2(and_1091_nl, or_tmp_446, or_468_cse);
  assign and_1092_nl = nand_276_cse & mux_tmp_164;
  assign mux_tmp_165 = MUX_s_1_2_2(and_1092_nl, mux_tmp_164, or_463_cse);
  assign and_1093_nl = nand_281_cse & mux_tmp_165;
  assign mux_168_nl = MUX_s_1_2_2(and_1093_nl, mux_tmp_165, or_458_cse);
  assign and_dcpl_504 = mux_168_nl & and_dcpl_366 & and_dcpl_471;
  assign or_475_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2!=2'b01);
  assign and_1087_nl = nand_271_cse & or_tmp_446;
  assign mux_tmp_167 = MUX_s_1_2_2(and_1087_nl, or_tmp_446, or_475_cse);
  assign and_1088_nl = nand_198_cse & mux_tmp_167;
  assign mux_tmp_168 = MUX_s_1_2_2(and_1088_nl, mux_tmp_167, or_468_cse);
  assign and_1089_nl = nand_276_cse & mux_tmp_168;
  assign mux_tmp_169 = MUX_s_1_2_2(and_1089_nl, mux_tmp_168, or_463_cse);
  assign and_1090_nl = nand_281_cse & mux_tmp_169;
  assign mux_172_nl = MUX_s_1_2_2(and_1090_nl, mux_tmp_169, or_458_cse);
  assign and_dcpl_506 = mux_172_nl & and_dcpl_370 & and_dcpl_475;
  assign nand_189_cse = ~((rem_12cyc_st_5_3_2[0]) & asn_itm_5 & main_stage_0_6 &
      (rem_12cyc_st_5_1_0[0]));
  assign or_484_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2[1]);
  assign and_1082_nl = nand_189_cse & or_tmp_446;
  assign mux_tmp_171 = MUX_s_1_2_2(and_1082_nl, or_tmp_446, or_484_cse);
  assign and_1083_nl = nand_271_cse & mux_tmp_171;
  assign mux_tmp_172 = MUX_s_1_2_2(and_1083_nl, mux_tmp_171, or_475_cse);
  assign and_1084_nl = nand_198_cse & mux_tmp_172;
  assign mux_tmp_173 = MUX_s_1_2_2(and_1084_nl, mux_tmp_172, or_468_cse);
  assign and_1085_nl = nand_276_cse & mux_tmp_173;
  assign mux_tmp_174 = MUX_s_1_2_2(and_1085_nl, mux_tmp_173, or_463_cse);
  assign and_1086_nl = nand_281_cse & mux_tmp_174;
  assign mux_177_nl = MUX_s_1_2_2(and_1086_nl, mux_tmp_174, or_458_cse);
  assign and_dcpl_508 = mux_177_nl & and_dcpl_121 & and_dcpl_115;
  assign or_495_cse = (rem_12cyc_st_6_1_0!=2'b01) | (rem_12cyc_st_6_3_2[1]);
  assign and_1076_nl = nand_215_cse & or_tmp_446;
  assign mux_tmp_176 = MUX_s_1_2_2(and_1076_nl, or_tmp_446, or_495_cse);
  assign and_1077_nl = nand_189_cse & mux_tmp_176;
  assign mux_tmp_177 = MUX_s_1_2_2(and_1077_nl, mux_tmp_176, or_484_cse);
  assign and_1078_nl = nand_271_cse & mux_tmp_177;
  assign mux_tmp_178 = MUX_s_1_2_2(and_1078_nl, mux_tmp_177, or_475_cse);
  assign and_1079_nl = nand_198_cse & mux_tmp_178;
  assign mux_tmp_179 = MUX_s_1_2_2(and_1079_nl, mux_tmp_178, or_468_cse);
  assign and_1080_nl = nand_276_cse & mux_tmp_179;
  assign mux_tmp_180 = MUX_s_1_2_2(and_1080_nl, mux_tmp_179, or_463_cse);
  assign and_1081_nl = nand_281_cse & mux_tmp_180;
  assign mux_183_nl = MUX_s_1_2_2(and_1081_nl, mux_tmp_180, or_458_cse);
  assign and_dcpl_510 = mux_183_nl & and_dcpl_94 & and_dcpl_87;
  assign or_508_cse = (rem_12cyc_st_7_1_0!=2'b01) | (rem_12cyc_st_7_3_2[1]);
  assign and_1069_nl = nand_212_cse & or_tmp_446;
  assign mux_tmp_182 = MUX_s_1_2_2(and_1069_nl, or_tmp_446, or_508_cse);
  assign and_1070_nl = nand_215_cse & mux_tmp_182;
  assign mux_tmp_183 = MUX_s_1_2_2(and_1070_nl, mux_tmp_182, or_495_cse);
  assign and_1071_nl = nand_189_cse & mux_tmp_183;
  assign mux_tmp_184 = MUX_s_1_2_2(and_1071_nl, mux_tmp_183, or_484_cse);
  assign and_1072_nl = nand_271_cse & mux_tmp_184;
  assign mux_tmp_185 = MUX_s_1_2_2(and_1072_nl, mux_tmp_184, or_475_cse);
  assign and_1073_nl = nand_198_cse & mux_tmp_185;
  assign mux_tmp_186 = MUX_s_1_2_2(and_1073_nl, mux_tmp_185, or_468_cse);
  assign and_1074_nl = nand_276_cse & mux_tmp_186;
  assign mux_tmp_187 = MUX_s_1_2_2(and_1074_nl, mux_tmp_186, or_463_cse);
  assign and_1075_nl = nand_281_cse & mux_tmp_187;
  assign mux_190_nl = MUX_s_1_2_2(and_1075_nl, mux_tmp_187, or_458_cse);
  assign and_dcpl_512 = mux_190_nl & and_dcpl_67 & and_dcpl_60;
  assign or_523_cse = (rem_12cyc_st_8_1_0!=2'b01) | (rem_12cyc_st_8_3_2[1]);
  assign and_1061_nl = nand_208_cse & or_tmp_446;
  assign mux_tmp_189 = MUX_s_1_2_2(and_1061_nl, or_tmp_446, or_523_cse);
  assign and_1062_nl = nand_212_cse & mux_tmp_189;
  assign mux_tmp_190 = MUX_s_1_2_2(and_1062_nl, mux_tmp_189, or_508_cse);
  assign and_1063_nl = nand_215_cse & mux_tmp_190;
  assign mux_tmp_191 = MUX_s_1_2_2(and_1063_nl, mux_tmp_190, or_495_cse);
  assign and_1064_nl = nand_189_cse & mux_tmp_191;
  assign mux_tmp_192 = MUX_s_1_2_2(and_1064_nl, mux_tmp_191, or_484_cse);
  assign and_1065_nl = nand_271_cse & mux_tmp_192;
  assign mux_tmp_193 = MUX_s_1_2_2(and_1065_nl, mux_tmp_192, or_475_cse);
  assign and_1066_nl = nand_198_cse & mux_tmp_193;
  assign mux_tmp_194 = MUX_s_1_2_2(and_1066_nl, mux_tmp_193, or_468_cse);
  assign and_1067_nl = nand_276_cse & mux_tmp_194;
  assign mux_tmp_195 = MUX_s_1_2_2(and_1067_nl, mux_tmp_194, or_463_cse);
  assign and_1068_nl = nand_281_cse & mux_tmp_195;
  assign mux_198_nl = MUX_s_1_2_2(and_1068_nl, mux_tmp_195, or_458_cse);
  assign and_dcpl_514 = mux_198_nl & and_dcpl_40 & and_dcpl_33;
  assign and_1052_nl = nand_203_cse & or_tmp_446;
  assign or_540_nl = (rem_12cyc_st_9_1_0!=2'b01) | (rem_12cyc_st_9_3_2[1]);
  assign mux_tmp_197 = MUX_s_1_2_2(and_1052_nl, or_tmp_446, or_540_nl);
  assign and_1053_nl = nand_208_cse & mux_tmp_197;
  assign mux_tmp_198 = MUX_s_1_2_2(and_1053_nl, mux_tmp_197, or_523_cse);
  assign and_1054_nl = nand_212_cse & mux_tmp_198;
  assign mux_tmp_199 = MUX_s_1_2_2(and_1054_nl, mux_tmp_198, or_508_cse);
  assign and_1055_nl = nand_215_cse & mux_tmp_199;
  assign mux_tmp_200 = MUX_s_1_2_2(and_1055_nl, mux_tmp_199, or_495_cse);
  assign and_1056_nl = nand_189_cse & mux_tmp_200;
  assign mux_tmp_201 = MUX_s_1_2_2(and_1056_nl, mux_tmp_200, or_484_cse);
  assign and_1057_nl = nand_271_cse & mux_tmp_201;
  assign mux_tmp_202 = MUX_s_1_2_2(and_1057_nl, mux_tmp_201, or_475_cse);
  assign and_1058_nl = nand_198_cse & mux_tmp_202;
  assign mux_tmp_203 = MUX_s_1_2_2(and_1058_nl, mux_tmp_202, or_468_cse);
  assign and_1059_nl = nand_276_cse & mux_tmp_203;
  assign mux_tmp_204 = MUX_s_1_2_2(and_1059_nl, mux_tmp_203, or_463_cse);
  assign and_1060_nl = nand_281_cse & mux_tmp_204;
  assign mux_207_nl = MUX_s_1_2_2(and_1060_nl, mux_tmp_204, or_458_cse);
  assign and_dcpl_516 = mux_207_nl & and_dcpl_13 & and_dcpl_6;
  assign and_tmp_134 = ((~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b01)
      | (rem_12cyc_st_7_3_2!=2'b01)) & ((~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b01)
      | (rem_12cyc_st_8_3_2!=2'b01)) & ((~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b01)
      | (rem_12cyc_st_9_3_2!=2'b01)) & ((~ main_stage_0_3) | (~ asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b01)
      | (rem_12cyc_st_2_3_2!=2'b01)) & ((~ main_stage_0_4) | (~ asn_itm_3) | (rem_12cyc_st_3_1_0!=2'b01)
      | (rem_12cyc_st_3_3_2!=2'b01)) & ((~ main_stage_0_5) | (~ asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b01)
      | (rem_12cyc_st_4_3_2!=2'b01)) & ((~ main_stage_0_6) | (~ asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b01)
      | (rem_12cyc_st_5_3_2!=2'b01)) & ((~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b01)
      | (rem_12cyc_st_6_3_2!=2'b01)) & ((~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b01)
      | (rem_12cyc_st_10_3_2!=2'b01)) & ((acc_tmp!=2'b01) | (acc_1_tmp[1]) | nand_250_cse);
  assign nor_439_nl = ~((rem_12cyc_1_0[0]) | (~ and_tmp_134));
  assign or_550_nl = (~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b01)
      | (rem_12cyc_1_0[1]);
  assign mux_tmp_206 = MUX_s_1_2_2(nor_439_nl, and_tmp_134, or_550_nl);
  assign and_dcpl_520 = and_dcpl_460 & and_dcpl_393;
  assign and_dcpl_521 = and_dcpl_462 & (rem_12cyc_st_2_1_0[1]);
  assign or_tmp_551 = (rem_12cyc_1_0!=2'b10) | (rem_12cyc_3_2[1]) | not_tmp_332;
  assign or_564_cse = (acc_1_tmp[1:0]!=2'b10) | (acc_tmp[1]);
  assign and_1170_nl = nand_281_cse & or_tmp_551;
  assign mux_209_nl = MUX_s_1_2_2(and_1170_nl, or_tmp_551, or_564_cse);
  assign and_dcpl_523 = mux_209_nl & and_dcpl_298 & and_dcpl_521;
  assign and_dcpl_524 = and_dcpl_466 & (rem_12cyc_st_3_1_0[1]);
  assign or_569_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2!=2'b01) |
      (~ asn_itm_2) | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp_135 = or_569_cse & or_tmp_551;
  assign and_1050_nl = nand_281_cse & and_tmp_135;
  assign mux_210_nl = MUX_s_1_2_2(and_1050_nl, and_tmp_135, or_564_cse);
  assign and_dcpl_526 = mux_210_nl & and_dcpl_304 & and_dcpl_524;
  assign and_dcpl_527 = and_dcpl_470 & (rem_12cyc_st_4_1_0[1]);
  assign or_573_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2!=2'b01) |
      (~ asn_itm_3) | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_137 = or_569_cse & or_573_cse & or_tmp_551;
  assign and_1049_nl = nand_281_cse & and_tmp_137;
  assign mux_211_nl = MUX_s_1_2_2(and_1049_nl, and_tmp_137, or_564_cse);
  assign and_dcpl_529 = mux_211_nl & and_dcpl_310 & and_dcpl_527;
  assign and_dcpl_530 = and_dcpl_474 & (rem_12cyc_st_5_1_0[1]);
  assign or_578_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2!=2'b01) |
      (~ asn_itm_4) | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_140 = or_569_cse & or_573_cse & or_578_cse & or_tmp_551;
  assign and_1048_nl = nand_281_cse & and_tmp_140;
  assign mux_212_nl = MUX_s_1_2_2(and_1048_nl, and_tmp_140, or_564_cse);
  assign and_dcpl_532 = mux_212_nl & and_dcpl_316 & and_dcpl_530;
  assign or_584_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2!=2'b01) |
      (~ asn_itm_5) | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_144 = or_569_cse & or_573_cse & or_578_cse & or_584_cse & or_tmp_551;
  assign and_1047_nl = nand_281_cse & and_tmp_144;
  assign mux_213_nl = MUX_s_1_2_2(and_1047_nl, and_tmp_144, or_564_cse);
  assign and_dcpl_534 = mux_213_nl & and_dcpl_121 & and_dcpl_117;
  assign or_591_cse = (rem_12cyc_st_6_1_0!=2'b10) | (rem_12cyc_st_6_3_2[1]);
  assign and_1045_nl = nand_215_cse & or_tmp_551;
  assign mux_214_nl = MUX_s_1_2_2(and_1045_nl, or_tmp_551, or_591_cse);
  assign and_tmp_148 = or_569_cse & or_573_cse & or_578_cse & or_584_cse & mux_214_nl;
  assign and_1046_nl = nand_281_cse & and_tmp_148;
  assign mux_215_nl = MUX_s_1_2_2(and_1046_nl, and_tmp_148, or_564_cse);
  assign and_dcpl_536 = mux_215_nl & and_dcpl_94 & and_dcpl_90;
  assign or_600_cse = (rem_12cyc_st_7_1_0!=2'b10) | (rem_12cyc_st_7_3_2[1]);
  assign and_1042_nl = nand_212_cse & or_tmp_551;
  assign mux_tmp_214 = MUX_s_1_2_2(and_1042_nl, or_tmp_551, or_600_cse);
  assign and_1043_nl = nand_215_cse & mux_tmp_214;
  assign mux_217_nl = MUX_s_1_2_2(and_1043_nl, mux_tmp_214, or_591_cse);
  assign and_tmp_152 = or_569_cse & or_573_cse & or_578_cse & or_584_cse & mux_217_nl;
  assign and_1044_nl = nand_281_cse & and_tmp_152;
  assign mux_218_nl = MUX_s_1_2_2(and_1044_nl, and_tmp_152, or_564_cse);
  assign and_dcpl_538 = mux_218_nl & and_dcpl_67 & and_dcpl_63;
  assign or_611_cse = (rem_12cyc_st_8_1_0!=2'b10) | (rem_12cyc_st_8_3_2[1]);
  assign and_1038_nl = nand_208_cse & or_tmp_551;
  assign mux_tmp_217 = MUX_s_1_2_2(and_1038_nl, or_tmp_551, or_611_cse);
  assign and_1039_nl = nand_212_cse & mux_tmp_217;
  assign mux_tmp_218 = MUX_s_1_2_2(and_1039_nl, mux_tmp_217, or_600_cse);
  assign and_1040_nl = nand_215_cse & mux_tmp_218;
  assign mux_221_nl = MUX_s_1_2_2(and_1040_nl, mux_tmp_218, or_591_cse);
  assign and_tmp_156 = or_569_cse & or_573_cse & or_578_cse & or_584_cse & mux_221_nl;
  assign and_1041_nl = nand_281_cse & and_tmp_156;
  assign mux_222_nl = MUX_s_1_2_2(and_1041_nl, and_tmp_156, or_564_cse);
  assign and_dcpl_540 = mux_222_nl & and_dcpl_40 & and_dcpl_36;
  assign and_1033_nl = nand_203_cse & or_tmp_551;
  assign or_624_nl = (rem_12cyc_st_9_1_0!=2'b10) | (rem_12cyc_st_9_3_2[1]);
  assign mux_tmp_221 = MUX_s_1_2_2(and_1033_nl, or_tmp_551, or_624_nl);
  assign and_1034_nl = nand_208_cse & mux_tmp_221;
  assign mux_tmp_222 = MUX_s_1_2_2(and_1034_nl, mux_tmp_221, or_611_cse);
  assign and_1035_nl = nand_212_cse & mux_tmp_222;
  assign mux_tmp_223 = MUX_s_1_2_2(and_1035_nl, mux_tmp_222, or_600_cse);
  assign and_1036_nl = nand_215_cse & mux_tmp_223;
  assign mux_226_nl = MUX_s_1_2_2(and_1036_nl, mux_tmp_223, or_591_cse);
  assign and_tmp_160 = or_569_cse & or_573_cse & or_578_cse & or_584_cse & mux_226_nl;
  assign and_1037_nl = nand_281_cse & and_tmp_160;
  assign mux_227_nl = MUX_s_1_2_2(and_1037_nl, and_tmp_160, or_564_cse);
  assign and_dcpl_542 = mux_227_nl & and_dcpl_13 & and_dcpl_9;
  assign and_tmp_170 = ((~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b01)
      | (rem_12cyc_1_0!=2'b10)) & ((~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b10)
      | (rem_12cyc_st_7_3_2!=2'b01)) & ((~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b10)
      | (rem_12cyc_st_8_3_2!=2'b01)) & ((~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b10)
      | (rem_12cyc_st_9_3_2!=2'b01)) & or_569_cse & or_573_cse & or_578_cse & or_584_cse
      & ((~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b10) | (rem_12cyc_st_6_3_2!=2'b01))
      & ((~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b10) | (rem_12cyc_st_10_3_2!=2'b01))
      & ((acc_tmp!=2'b01) | (acc_1_tmp[1:0]!=2'b10) | (~ ccs_ccore_start_rsci_idat));
  assign and_dcpl_546 = and_dcpl_460 & and_dcpl_430;
  assign or_tmp_629 = (rem_12cyc_1_0!=2'b11) | (rem_12cyc_3_2[1]) | not_tmp_332;
  assign or_643_cse = (acc_1_tmp[1:0]!=2'b11) | (acc_tmp[1]);
  assign and_1169_nl = nand_281_cse & or_tmp_629;
  assign mux_228_nl = MUX_s_1_2_2(and_1169_nl, or_tmp_629, or_643_cse);
  assign and_dcpl_548 = mux_228_nl & and_dcpl_358 & and_dcpl_521;
  assign or_648_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2!=2'b01);
  assign and_1030_nl = nand_276_cse & or_tmp_629;
  assign mux_tmp_227 = MUX_s_1_2_2(and_1030_nl, or_tmp_629, or_648_cse);
  assign and_1031_nl = nand_281_cse & mux_tmp_227;
  assign mux_230_nl = MUX_s_1_2_2(and_1031_nl, mux_tmp_227, or_643_cse);
  assign and_dcpl_550 = mux_230_nl & and_dcpl_362 & and_dcpl_524;
  assign or_653_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2[1]);
  assign and_1027_nl = nand_198_cse & or_tmp_629;
  assign mux_tmp_229 = MUX_s_1_2_2(and_1027_nl, or_tmp_629, or_653_cse);
  assign and_1028_nl = nand_276_cse & mux_tmp_229;
  assign mux_tmp_230 = MUX_s_1_2_2(and_1028_nl, mux_tmp_229, or_648_cse);
  assign and_1029_nl = nand_281_cse & mux_tmp_230;
  assign mux_233_nl = MUX_s_1_2_2(and_1029_nl, mux_tmp_230, or_643_cse);
  assign and_dcpl_552 = mux_233_nl & and_dcpl_366 & and_dcpl_527;
  assign or_660_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2!=2'b01);
  assign and_1023_nl = nand_271_cse & or_tmp_629;
  assign mux_tmp_232 = MUX_s_1_2_2(and_1023_nl, or_tmp_629, or_660_cse);
  assign and_1024_nl = nand_198_cse & mux_tmp_232;
  assign mux_tmp_233 = MUX_s_1_2_2(and_1024_nl, mux_tmp_232, or_653_cse);
  assign and_1025_nl = nand_276_cse & mux_tmp_233;
  assign mux_tmp_234 = MUX_s_1_2_2(and_1025_nl, mux_tmp_233, or_648_cse);
  assign and_1026_nl = nand_281_cse & mux_tmp_234;
  assign mux_237_nl = MUX_s_1_2_2(and_1026_nl, mux_tmp_234, or_643_cse);
  assign and_dcpl_554 = mux_237_nl & and_dcpl_370 & and_dcpl_530;
  assign or_669_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2[1]);
  assign and_1018_nl = nand_189_cse & or_tmp_629;
  assign mux_tmp_236 = MUX_s_1_2_2(and_1018_nl, or_tmp_629, or_669_cse);
  assign and_1019_nl = nand_271_cse & mux_tmp_236;
  assign mux_tmp_237 = MUX_s_1_2_2(and_1019_nl, mux_tmp_236, or_660_cse);
  assign and_1020_nl = nand_198_cse & mux_tmp_237;
  assign mux_tmp_238 = MUX_s_1_2_2(and_1020_nl, mux_tmp_237, or_653_cse);
  assign and_1021_nl = nand_276_cse & mux_tmp_238;
  assign mux_tmp_239 = MUX_s_1_2_2(and_1021_nl, mux_tmp_238, or_648_cse);
  assign and_1022_nl = nand_281_cse & mux_tmp_239;
  assign mux_242_nl = MUX_s_1_2_2(and_1022_nl, mux_tmp_239, or_643_cse);
  assign and_dcpl_556 = mux_242_nl & and_dcpl_121 & and_dcpl_119;
  assign or_680_cse = (rem_12cyc_st_6_1_0!=2'b11) | (rem_12cyc_st_6_3_2[1]);
  assign and_1012_nl = nand_215_cse & or_tmp_629;
  assign mux_tmp_241 = MUX_s_1_2_2(and_1012_nl, or_tmp_629, or_680_cse);
  assign and_1013_nl = nand_189_cse & mux_tmp_241;
  assign mux_tmp_242 = MUX_s_1_2_2(and_1013_nl, mux_tmp_241, or_669_cse);
  assign and_1014_nl = nand_271_cse & mux_tmp_242;
  assign mux_tmp_243 = MUX_s_1_2_2(and_1014_nl, mux_tmp_242, or_660_cse);
  assign and_1015_nl = nand_198_cse & mux_tmp_243;
  assign mux_tmp_244 = MUX_s_1_2_2(and_1015_nl, mux_tmp_243, or_653_cse);
  assign and_1016_nl = nand_276_cse & mux_tmp_244;
  assign mux_tmp_245 = MUX_s_1_2_2(and_1016_nl, mux_tmp_244, or_648_cse);
  assign and_1017_nl = nand_281_cse & mux_tmp_245;
  assign mux_248_nl = MUX_s_1_2_2(and_1017_nl, mux_tmp_245, or_643_cse);
  assign and_dcpl_558 = mux_248_nl & and_dcpl_94 & and_dcpl_92;
  assign or_693_cse = (rem_12cyc_st_7_1_0!=2'b11) | (rem_12cyc_st_7_3_2[1]);
  assign and_1005_nl = nand_212_cse & or_tmp_629;
  assign mux_tmp_247 = MUX_s_1_2_2(and_1005_nl, or_tmp_629, or_693_cse);
  assign and_1006_nl = nand_215_cse & mux_tmp_247;
  assign mux_tmp_248 = MUX_s_1_2_2(and_1006_nl, mux_tmp_247, or_680_cse);
  assign and_1007_nl = nand_189_cse & mux_tmp_248;
  assign mux_tmp_249 = MUX_s_1_2_2(and_1007_nl, mux_tmp_248, or_669_cse);
  assign and_1008_nl = nand_271_cse & mux_tmp_249;
  assign mux_tmp_250 = MUX_s_1_2_2(and_1008_nl, mux_tmp_249, or_660_cse);
  assign and_1009_nl = nand_198_cse & mux_tmp_250;
  assign mux_tmp_251 = MUX_s_1_2_2(and_1009_nl, mux_tmp_250, or_653_cse);
  assign and_1010_nl = nand_276_cse & mux_tmp_251;
  assign mux_tmp_252 = MUX_s_1_2_2(and_1010_nl, mux_tmp_251, or_648_cse);
  assign and_1011_nl = nand_281_cse & mux_tmp_252;
  assign mux_255_nl = MUX_s_1_2_2(and_1011_nl, mux_tmp_252, or_643_cse);
  assign and_dcpl_560 = mux_255_nl & and_dcpl_67 & and_dcpl_65;
  assign or_708_cse = (rem_12cyc_st_8_1_0!=2'b11) | (rem_12cyc_st_8_3_2[1]);
  assign and_997_nl = nand_208_cse & or_tmp_629;
  assign mux_tmp_254 = MUX_s_1_2_2(and_997_nl, or_tmp_629, or_708_cse);
  assign and_998_nl = nand_212_cse & mux_tmp_254;
  assign mux_tmp_255 = MUX_s_1_2_2(and_998_nl, mux_tmp_254, or_693_cse);
  assign and_999_nl = nand_215_cse & mux_tmp_255;
  assign mux_tmp_256 = MUX_s_1_2_2(and_999_nl, mux_tmp_255, or_680_cse);
  assign and_1000_nl = nand_189_cse & mux_tmp_256;
  assign mux_tmp_257 = MUX_s_1_2_2(and_1000_nl, mux_tmp_256, or_669_cse);
  assign and_1001_nl = nand_271_cse & mux_tmp_257;
  assign mux_tmp_258 = MUX_s_1_2_2(and_1001_nl, mux_tmp_257, or_660_cse);
  assign and_1002_nl = nand_198_cse & mux_tmp_258;
  assign mux_tmp_259 = MUX_s_1_2_2(and_1002_nl, mux_tmp_258, or_653_cse);
  assign and_1003_nl = nand_276_cse & mux_tmp_259;
  assign mux_tmp_260 = MUX_s_1_2_2(and_1003_nl, mux_tmp_259, or_648_cse);
  assign and_1004_nl = nand_281_cse & mux_tmp_260;
  assign mux_263_nl = MUX_s_1_2_2(and_1004_nl, mux_tmp_260, or_643_cse);
  assign and_dcpl_562 = mux_263_nl & and_dcpl_40 & and_dcpl_38;
  assign and_988_nl = nand_203_cse & or_tmp_629;
  assign or_725_nl = (rem_12cyc_st_9_1_0!=2'b11) | (rem_12cyc_st_9_3_2[1]);
  assign mux_tmp_262 = MUX_s_1_2_2(and_988_nl, or_tmp_629, or_725_nl);
  assign and_989_nl = nand_208_cse & mux_tmp_262;
  assign mux_tmp_263 = MUX_s_1_2_2(and_989_nl, mux_tmp_262, or_708_cse);
  assign and_990_nl = nand_212_cse & mux_tmp_263;
  assign mux_tmp_264 = MUX_s_1_2_2(and_990_nl, mux_tmp_263, or_693_cse);
  assign and_991_nl = nand_215_cse & mux_tmp_264;
  assign mux_tmp_265 = MUX_s_1_2_2(and_991_nl, mux_tmp_264, or_680_cse);
  assign and_992_nl = nand_189_cse & mux_tmp_265;
  assign mux_tmp_266 = MUX_s_1_2_2(and_992_nl, mux_tmp_265, or_669_cse);
  assign and_993_nl = nand_271_cse & mux_tmp_266;
  assign mux_tmp_267 = MUX_s_1_2_2(and_993_nl, mux_tmp_266, or_660_cse);
  assign and_994_nl = nand_198_cse & mux_tmp_267;
  assign mux_tmp_268 = MUX_s_1_2_2(and_994_nl, mux_tmp_267, or_653_cse);
  assign and_995_nl = nand_276_cse & mux_tmp_268;
  assign mux_tmp_269 = MUX_s_1_2_2(and_995_nl, mux_tmp_268, or_648_cse);
  assign and_996_nl = nand_281_cse & mux_tmp_269;
  assign mux_272_nl = MUX_s_1_2_2(and_996_nl, mux_tmp_269, or_643_cse);
  assign and_dcpl_564 = mux_272_nl & and_dcpl_13 & and_dcpl_11;
  assign and_tmp_179 = (~(main_stage_0_8 & asn_itm_7 & (rem_12cyc_st_7_1_0==2'b11)
      & (rem_12cyc_st_7_3_2==2'b01))) & (~(main_stage_0_9 & asn_itm_8 & (rem_12cyc_st_8_1_0==2'b11)
      & (rem_12cyc_st_8_3_2==2'b01))) & (~(main_stage_0_10 & asn_itm_9 & (rem_12cyc_st_9_1_0==2'b11)
      & (rem_12cyc_st_9_3_2==2'b01))) & (~(main_stage_0_3 & asn_itm_2 & (rem_12cyc_st_2_1_0==2'b11)
      & (rem_12cyc_st_2_3_2==2'b01))) & (~(main_stage_0_4 & asn_itm_3 & (rem_12cyc_st_3_1_0==2'b11)
      & (rem_12cyc_st_3_3_2==2'b01))) & (~(main_stage_0_5 & asn_itm_4 & (rem_12cyc_st_4_1_0==2'b11)
      & (rem_12cyc_st_4_3_2==2'b01))) & (~(main_stage_0_6 & asn_itm_5 & (rem_12cyc_st_5_1_0==2'b11)
      & (rem_12cyc_st_5_3_2==2'b01))) & (~(main_stage_0_7 & asn_itm_6 & (rem_12cyc_st_6_1_0==2'b11)
      & (rem_12cyc_st_6_3_2==2'b01))) & (~(main_stage_0_11 & asn_itm_10 & (rem_12cyc_st_10_1_0==2'b11)
      & (rem_12cyc_st_10_3_2==2'b01))) & ((acc_tmp[1]) | (~((acc_tmp[0]) & (acc_1_tmp[1:0]==2'b11)
      & ccs_ccore_start_rsci_idat)));
  assign and_987_nl = (~((rem_12cyc_3_2[0]) & (rem_12cyc_1_0==2'b11))) & and_tmp_179;
  assign or_735_nl = (~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2[1]);
  assign mux_tmp_271 = MUX_s_1_2_2(and_987_nl, and_tmp_179, or_735_nl);
  assign and_dcpl_568 = and_dcpl_292 & (acc_tmp[1]);
  assign and_dcpl_569 = and_dcpl_568 & and_dcpl_291;
  assign and_dcpl_570 = (rem_12cyc_st_2_3_2==2'b10);
  assign and_dcpl_571 = and_dcpl_570 & (~ (rem_12cyc_st_2_1_0[1]));
  assign or_tmp_733 = (rem_12cyc_1_0!=2'b00) | (rem_12cyc_3_2!=2'b10) | not_tmp_54;
  assign or_748_cse = (acc_1_tmp[1:0]!=2'b00) | (acc_tmp!=2'b10);
  assign nor_436_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_733));
  assign mux_274_nl = MUX_s_1_2_2(nor_436_nl, or_tmp_733, or_748_cse);
  assign and_dcpl_573 = mux_274_nl & and_dcpl_298 & and_dcpl_571;
  assign and_dcpl_574 = (rem_12cyc_st_3_3_2==2'b10);
  assign and_dcpl_575 = and_dcpl_574 & (~ (rem_12cyc_st_3_1_0[1]));
  assign or_753_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2!=2'b10) | (~
      asn_itm_2) | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp_180 = or_753_cse & or_tmp_733;
  assign nor_435_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_180));
  assign mux_275_nl = MUX_s_1_2_2(nor_435_nl, and_tmp_180, or_748_cse);
  assign and_dcpl_577 = mux_275_nl & and_dcpl_304 & and_dcpl_575;
  assign and_dcpl_578 = (rem_12cyc_st_4_3_2==2'b10);
  assign and_dcpl_579 = and_dcpl_578 & (~ (rem_12cyc_st_4_1_0[1]));
  assign or_757_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2!=2'b10) | (~
      asn_itm_3) | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_182 = or_753_cse & or_757_cse & or_tmp_733;
  assign nor_434_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_182));
  assign mux_276_nl = MUX_s_1_2_2(nor_434_nl, and_tmp_182, or_748_cse);
  assign and_dcpl_581 = mux_276_nl & and_dcpl_310 & and_dcpl_579;
  assign and_dcpl_582 = (rem_12cyc_st_5_3_2==2'b10);
  assign and_dcpl_583 = and_dcpl_582 & (~ (rem_12cyc_st_5_1_0[1]));
  assign or_762_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2!=2'b10) | (~
      asn_itm_4) | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_185 = or_753_cse & or_757_cse & or_762_cse & or_tmp_733;
  assign nor_433_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_185));
  assign mux_277_nl = MUX_s_1_2_2(nor_433_nl, and_tmp_185, or_748_cse);
  assign and_dcpl_585 = mux_277_nl & and_dcpl_316 & and_dcpl_583;
  assign or_768_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2!=2'b10) | (~
      asn_itm_5) | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_189 = or_753_cse & or_757_cse & or_762_cse & or_768_cse & or_tmp_733;
  assign nor_432_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_189));
  assign mux_278_nl = MUX_s_1_2_2(nor_432_nl, and_tmp_189, or_748_cse);
  assign and_dcpl_589 = mux_278_nl & and_dcpl_112 & and_dcpl_126 & (~ (rem_12cyc_st_6_1_0[1]));
  assign or_775_cse = (rem_12cyc_st_6_1_0!=2'b00) | (rem_12cyc_st_6_3_2!=2'b10);
  assign nor_430_nl = ~(and_dcpl_111 | (~ or_tmp_733));
  assign mux_279_nl = MUX_s_1_2_2(nor_430_nl, or_tmp_733, or_775_cse);
  assign and_tmp_193 = or_753_cse & or_757_cse & or_762_cse & or_768_cse & mux_279_nl;
  assign nor_431_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_193));
  assign mux_280_nl = MUX_s_1_2_2(nor_431_nl, and_tmp_193, or_748_cse);
  assign and_dcpl_593 = mux_280_nl & and_dcpl_85 & and_dcpl_99 & (~ (rem_12cyc_st_7_1_0[0]));
  assign or_784_cse = (rem_12cyc_st_7_1_0!=2'b00) | (rem_12cyc_st_7_3_2!=2'b10);
  assign nor_427_nl = ~(and_dcpl_84 | (~ or_tmp_733));
  assign mux_tmp_279 = MUX_s_1_2_2(nor_427_nl, or_tmp_733, or_784_cse);
  assign nor_428_nl = ~(and_dcpl_111 | (~ mux_tmp_279));
  assign mux_282_nl = MUX_s_1_2_2(nor_428_nl, mux_tmp_279, or_775_cse);
  assign and_tmp_197 = or_753_cse & or_757_cse & or_762_cse & or_768_cse & mux_282_nl;
  assign nor_429_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_197));
  assign mux_283_nl = MUX_s_1_2_2(nor_429_nl, and_tmp_197, or_748_cse);
  assign and_dcpl_597 = mux_283_nl & and_dcpl_58 & and_dcpl_72 & (~ (rem_12cyc_st_8_1_0[0]));
  assign or_795_cse = (rem_12cyc_st_8_1_0!=2'b00) | (rem_12cyc_st_8_3_2!=2'b10);
  assign nor_423_nl = ~(and_dcpl_57 | (~ or_tmp_733));
  assign mux_tmp_282 = MUX_s_1_2_2(nor_423_nl, or_tmp_733, or_795_cse);
  assign nor_424_nl = ~(and_dcpl_84 | (~ mux_tmp_282));
  assign mux_tmp_283 = MUX_s_1_2_2(nor_424_nl, mux_tmp_282, or_784_cse);
  assign nor_425_nl = ~(and_dcpl_111 | (~ mux_tmp_283));
  assign mux_286_nl = MUX_s_1_2_2(nor_425_nl, mux_tmp_283, or_775_cse);
  assign and_tmp_201 = or_753_cse & or_757_cse & or_762_cse & or_768_cse & mux_286_nl;
  assign nor_426_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_201));
  assign mux_287_nl = MUX_s_1_2_2(nor_426_nl, and_tmp_201, or_748_cse);
  assign and_dcpl_601 = mux_287_nl & and_dcpl_31 & and_dcpl_45 & (~ (rem_12cyc_st_9_1_0[0]));
  assign nor_418_nl = ~(and_dcpl_30 | (~ or_tmp_733));
  assign or_808_nl = (rem_12cyc_st_9_1_0!=2'b00) | (rem_12cyc_st_9_3_2!=2'b10);
  assign mux_tmp_286 = MUX_s_1_2_2(nor_418_nl, or_tmp_733, or_808_nl);
  assign nor_419_nl = ~(and_dcpl_57 | (~ mux_tmp_286));
  assign mux_tmp_287 = MUX_s_1_2_2(nor_419_nl, mux_tmp_286, or_795_cse);
  assign nor_420_nl = ~(and_dcpl_84 | (~ mux_tmp_287));
  assign mux_tmp_288 = MUX_s_1_2_2(nor_420_nl, mux_tmp_287, or_784_cse);
  assign nor_421_nl = ~(and_dcpl_111 | (~ mux_tmp_288));
  assign mux_291_nl = MUX_s_1_2_2(nor_421_nl, mux_tmp_288, or_775_cse);
  assign and_tmp_205 = or_753_cse & or_757_cse & or_762_cse & or_768_cse & mux_291_nl;
  assign nor_422_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_205));
  assign mux_292_nl = MUX_s_1_2_2(nor_422_nl, and_tmp_205, or_748_cse);
  assign and_dcpl_605 = mux_292_nl & and_dcpl_4 & and_dcpl_18 & (~ (rem_12cyc_st_10_1_0[0]));
  assign or_tmp_808 = (acc_tmp!=2'b10) | (acc_1_tmp[1:0]!=2'b00) | (~ ccs_ccore_start_rsci_idat);
  assign nor_409_nl = ~((rem_12cyc_st_10_3_2[1]) | (~ or_tmp_808));
  assign or_823_nl = (~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b00)
      | (rem_12cyc_st_10_3_2[0]);
  assign mux_tmp_291 = MUX_s_1_2_2(nor_409_nl, or_tmp_808, or_823_nl);
  assign nor_410_nl = ~((rem_12cyc_st_6_3_2[1]) | (~ mux_tmp_291));
  assign or_822_nl = (~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b00)
      | (rem_12cyc_st_6_3_2[0]);
  assign mux_tmp_292 = MUX_s_1_2_2(nor_410_nl, mux_tmp_291, or_822_nl);
  assign nor_411_nl = ~((rem_12cyc_st_5_3_2[1]) | (~ mux_tmp_292));
  assign or_821_nl = (~ main_stage_0_6) | (~ asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b00)
      | (rem_12cyc_st_5_3_2[0]);
  assign mux_tmp_293 = MUX_s_1_2_2(nor_411_nl, mux_tmp_292, or_821_nl);
  assign nor_412_nl = ~((rem_12cyc_st_4_3_2[1]) | (~ mux_tmp_293));
  assign or_820_nl = (~ main_stage_0_5) | (~ asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b00)
      | (rem_12cyc_st_4_3_2[0]);
  assign mux_tmp_294 = MUX_s_1_2_2(nor_412_nl, mux_tmp_293, or_820_nl);
  assign nor_413_nl = ~((rem_12cyc_st_3_3_2[1]) | (~ mux_tmp_294));
  assign or_819_nl = (~ main_stage_0_4) | (~ asn_itm_3) | (rem_12cyc_st_3_1_0!=2'b00)
      | (rem_12cyc_st_3_3_2[0]);
  assign mux_tmp_295 = MUX_s_1_2_2(nor_413_nl, mux_tmp_294, or_819_nl);
  assign nor_414_nl = ~((rem_12cyc_st_2_3_2[1]) | (~ mux_tmp_295));
  assign or_818_nl = (~ main_stage_0_3) | (~ asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b00)
      | (rem_12cyc_st_2_3_2[0]);
  assign mux_tmp_296 = MUX_s_1_2_2(nor_414_nl, mux_tmp_295, or_818_nl);
  assign nor_415_nl = ~((rem_12cyc_st_9_3_2[1]) | (~ mux_tmp_296));
  assign or_817_nl = (~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b00)
      | (rem_12cyc_st_9_3_2[0]);
  assign mux_tmp_297 = MUX_s_1_2_2(nor_415_nl, mux_tmp_296, or_817_nl);
  assign nor_416_nl = ~((rem_12cyc_st_8_3_2[1]) | (~ mux_tmp_297));
  assign or_816_nl = (~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b00)
      | (rem_12cyc_st_8_3_2[0]);
  assign mux_tmp_298 = MUX_s_1_2_2(nor_416_nl, mux_tmp_297, or_816_nl);
  assign nor_417_nl = ~((rem_12cyc_st_7_3_2[1]) | (~ mux_tmp_298));
  assign or_815_nl = (~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b00)
      | (rem_12cyc_st_7_3_2[0]);
  assign mux_301_nl = MUX_s_1_2_2(nor_417_nl, mux_tmp_298, or_815_nl);
  assign and_tmp_206 = ((~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b10)
      | (rem_12cyc_1_0!=2'b00)) & mux_301_nl;
  assign and_dcpl_610 = and_dcpl_568 & and_dcpl_355;
  assign or_tmp_820 = (rem_12cyc_1_0!=2'b01) | (rem_12cyc_3_2!=2'b10) | not_tmp_54;
  assign or_837_cse = (acc_1_tmp[1:0]!=2'b01) | (acc_tmp!=2'b10);
  assign nor_408_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_820));
  assign mux_302_nl = MUX_s_1_2_2(nor_408_nl, or_tmp_820, or_837_cse);
  assign and_dcpl_612 = mux_302_nl & and_dcpl_358 & and_dcpl_571;
  assign nand_84_cse = ~((rem_12cyc_st_2_3_2[1]) & asn_itm_2 & main_stage_0_3 & (rem_12cyc_st_2_1_0[0]));
  assign or_842_cse = (rem_12cyc_st_2_1_0[1]) | (rem_12cyc_st_2_3_2[0]);
  assign and_986_nl = nand_84_cse & or_tmp_820;
  assign mux_tmp_301 = MUX_s_1_2_2(and_986_nl, or_tmp_820, or_842_cse);
  assign nor_407_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_301));
  assign mux_304_nl = MUX_s_1_2_2(nor_407_nl, mux_tmp_301, or_837_cse);
  assign and_dcpl_614 = mux_304_nl & and_dcpl_362 & and_dcpl_575;
  assign or_847_cse = (rem_12cyc_st_3_1_0[1]) | (rem_12cyc_st_3_3_2!=2'b10);
  assign and_984_nl = nand_274_cse & or_tmp_820;
  assign mux_tmp_303 = MUX_s_1_2_2(and_984_nl, or_tmp_820, or_847_cse);
  assign and_985_nl = nand_84_cse & mux_tmp_303;
  assign mux_tmp_304 = MUX_s_1_2_2(and_985_nl, mux_tmp_303, or_842_cse);
  assign nor_406_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_304));
  assign mux_307_nl = MUX_s_1_2_2(nor_406_nl, mux_tmp_304, or_837_cse);
  assign and_dcpl_616 = mux_307_nl & and_dcpl_366 & and_dcpl_579;
  assign nand_79_cse = ~((rem_12cyc_st_4_3_2[1]) & asn_itm_4 & main_stage_0_5 & (rem_12cyc_st_4_1_0[0]));
  assign or_854_cse = (rem_12cyc_st_4_1_0[1]) | (rem_12cyc_st_4_3_2[0]);
  assign and_981_nl = nand_79_cse & or_tmp_820;
  assign mux_tmp_306 = MUX_s_1_2_2(and_981_nl, or_tmp_820, or_854_cse);
  assign and_982_nl = nand_274_cse & mux_tmp_306;
  assign mux_tmp_307 = MUX_s_1_2_2(and_982_nl, mux_tmp_306, or_847_cse);
  assign and_983_nl = nand_84_cse & mux_tmp_307;
  assign mux_tmp_308 = MUX_s_1_2_2(and_983_nl, mux_tmp_307, or_842_cse);
  assign nor_405_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_308));
  assign mux_311_nl = MUX_s_1_2_2(nor_405_nl, mux_tmp_308, or_837_cse);
  assign and_dcpl_618 = mux_311_nl & and_dcpl_370 & and_dcpl_583;
  assign or_863_cse = (rem_12cyc_st_5_1_0[1]) | (rem_12cyc_st_5_3_2!=2'b10);
  assign and_977_nl = nand_267_cse & or_tmp_820;
  assign mux_tmp_310 = MUX_s_1_2_2(and_977_nl, or_tmp_820, or_863_cse);
  assign and_978_nl = nand_79_cse & mux_tmp_310;
  assign mux_tmp_311 = MUX_s_1_2_2(and_978_nl, mux_tmp_310, or_854_cse);
  assign and_979_nl = nand_274_cse & mux_tmp_311;
  assign mux_tmp_312 = MUX_s_1_2_2(and_979_nl, mux_tmp_311, or_847_cse);
  assign and_980_nl = nand_84_cse & mux_tmp_312;
  assign mux_tmp_313 = MUX_s_1_2_2(and_980_nl, mux_tmp_312, or_842_cse);
  assign nor_404_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_313));
  assign mux_316_nl = MUX_s_1_2_2(nor_404_nl, mux_tmp_313, or_837_cse);
  assign and_dcpl_622 = mux_316_nl & and_dcpl_112 & and_dcpl_129 & (~ (rem_12cyc_st_6_1_0[1]));
  assign or_874_cse = (rem_12cyc_st_6_1_0!=2'b01) | (rem_12cyc_st_6_3_2!=2'b10);
  assign nor_402_nl = ~(and_dcpl_111 | (~ or_tmp_820));
  assign mux_tmp_315 = MUX_s_1_2_2(nor_402_nl, or_tmp_820, or_874_cse);
  assign and_973_nl = nand_267_cse & mux_tmp_315;
  assign mux_tmp_316 = MUX_s_1_2_2(and_973_nl, mux_tmp_315, or_863_cse);
  assign and_974_nl = nand_79_cse & mux_tmp_316;
  assign mux_tmp_317 = MUX_s_1_2_2(and_974_nl, mux_tmp_316, or_854_cse);
  assign and_975_nl = nand_274_cse & mux_tmp_317;
  assign mux_tmp_318 = MUX_s_1_2_2(and_975_nl, mux_tmp_317, or_847_cse);
  assign and_976_nl = nand_84_cse & mux_tmp_318;
  assign mux_tmp_319 = MUX_s_1_2_2(and_976_nl, mux_tmp_318, or_842_cse);
  assign nor_403_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_319));
  assign mux_322_nl = MUX_s_1_2_2(nor_403_nl, mux_tmp_319, or_837_cse);
  assign and_dcpl_625 = mux_322_nl & and_dcpl_85 & and_dcpl_99 & (rem_12cyc_st_7_1_0[0]);
  assign or_887_cse = (rem_12cyc_st_7_1_0!=2'b01) | (rem_12cyc_st_7_3_2!=2'b10);
  assign nor_399_nl = ~(and_dcpl_84 | (~ or_tmp_820));
  assign mux_tmp_321 = MUX_s_1_2_2(nor_399_nl, or_tmp_820, or_887_cse);
  assign nor_400_nl = ~(and_dcpl_111 | (~ mux_tmp_321));
  assign mux_tmp_322 = MUX_s_1_2_2(nor_400_nl, mux_tmp_321, or_874_cse);
  assign and_969_nl = nand_267_cse & mux_tmp_322;
  assign mux_tmp_323 = MUX_s_1_2_2(and_969_nl, mux_tmp_322, or_863_cse);
  assign and_970_nl = nand_79_cse & mux_tmp_323;
  assign mux_tmp_324 = MUX_s_1_2_2(and_970_nl, mux_tmp_323, or_854_cse);
  assign and_971_nl = nand_274_cse & mux_tmp_324;
  assign mux_tmp_325 = MUX_s_1_2_2(and_971_nl, mux_tmp_324, or_847_cse);
  assign and_972_nl = nand_84_cse & mux_tmp_325;
  assign mux_tmp_326 = MUX_s_1_2_2(and_972_nl, mux_tmp_325, or_842_cse);
  assign nor_401_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_326));
  assign mux_329_nl = MUX_s_1_2_2(nor_401_nl, mux_tmp_326, or_837_cse);
  assign and_dcpl_628 = mux_329_nl & and_dcpl_58 & and_dcpl_72 & (rem_12cyc_st_8_1_0[0]);
  assign or_902_cse = (rem_12cyc_st_8_1_0!=2'b01) | (rem_12cyc_st_8_3_2!=2'b10);
  assign nor_395_nl = ~(and_dcpl_57 | (~ or_tmp_820));
  assign mux_tmp_328 = MUX_s_1_2_2(nor_395_nl, or_tmp_820, or_902_cse);
  assign nor_396_nl = ~(and_dcpl_84 | (~ mux_tmp_328));
  assign mux_tmp_329 = MUX_s_1_2_2(nor_396_nl, mux_tmp_328, or_887_cse);
  assign nor_397_nl = ~(and_dcpl_111 | (~ mux_tmp_329));
  assign mux_tmp_330 = MUX_s_1_2_2(nor_397_nl, mux_tmp_329, or_874_cse);
  assign and_965_nl = nand_267_cse & mux_tmp_330;
  assign mux_tmp_331 = MUX_s_1_2_2(and_965_nl, mux_tmp_330, or_863_cse);
  assign and_966_nl = nand_79_cse & mux_tmp_331;
  assign mux_tmp_332 = MUX_s_1_2_2(and_966_nl, mux_tmp_331, or_854_cse);
  assign and_967_nl = nand_274_cse & mux_tmp_332;
  assign mux_tmp_333 = MUX_s_1_2_2(and_967_nl, mux_tmp_332, or_847_cse);
  assign and_968_nl = nand_84_cse & mux_tmp_333;
  assign mux_tmp_334 = MUX_s_1_2_2(and_968_nl, mux_tmp_333, or_842_cse);
  assign nor_398_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_334));
  assign mux_337_nl = MUX_s_1_2_2(nor_398_nl, mux_tmp_334, or_837_cse);
  assign and_dcpl_631 = mux_337_nl & and_dcpl_31 & and_dcpl_45 & (rem_12cyc_st_9_1_0[0]);
  assign nor_390_nl = ~(and_dcpl_30 | (~ or_tmp_820));
  assign or_919_nl = (rem_12cyc_st_9_1_0!=2'b01) | (rem_12cyc_st_9_3_2!=2'b10);
  assign mux_tmp_336 = MUX_s_1_2_2(nor_390_nl, or_tmp_820, or_919_nl);
  assign nor_391_nl = ~(and_dcpl_57 | (~ mux_tmp_336));
  assign mux_tmp_337 = MUX_s_1_2_2(nor_391_nl, mux_tmp_336, or_902_cse);
  assign nor_392_nl = ~(and_dcpl_84 | (~ mux_tmp_337));
  assign mux_tmp_338 = MUX_s_1_2_2(nor_392_nl, mux_tmp_337, or_887_cse);
  assign nor_393_nl = ~(and_dcpl_111 | (~ mux_tmp_338));
  assign mux_tmp_339 = MUX_s_1_2_2(nor_393_nl, mux_tmp_338, or_874_cse);
  assign and_961_nl = nand_267_cse & mux_tmp_339;
  assign mux_tmp_340 = MUX_s_1_2_2(and_961_nl, mux_tmp_339, or_863_cse);
  assign and_962_nl = nand_79_cse & mux_tmp_340;
  assign mux_tmp_341 = MUX_s_1_2_2(and_962_nl, mux_tmp_340, or_854_cse);
  assign and_963_nl = nand_274_cse & mux_tmp_341;
  assign mux_tmp_342 = MUX_s_1_2_2(and_963_nl, mux_tmp_341, or_847_cse);
  assign and_964_nl = nand_84_cse & mux_tmp_342;
  assign mux_tmp_343 = MUX_s_1_2_2(and_964_nl, mux_tmp_342, or_842_cse);
  assign nor_394_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_343));
  assign mux_346_nl = MUX_s_1_2_2(nor_394_nl, mux_tmp_343, or_837_cse);
  assign and_dcpl_634 = mux_346_nl & and_dcpl_4 & and_dcpl_18 & (rem_12cyc_st_10_1_0[0]);
  assign or_tmp_921 = (acc_tmp!=2'b10) | (acc_1_tmp[1]) | nand_250_cse;
  assign nor_380_nl = ~((rem_12cyc_st_10_3_2[1]) | (~ or_tmp_921));
  assign or_938_nl = (~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b01)
      | (rem_12cyc_st_10_3_2[0]);
  assign mux_tmp_345 = MUX_s_1_2_2(nor_380_nl, or_tmp_921, or_938_nl);
  assign nor_381_nl = ~((rem_12cyc_st_6_3_2[1]) | (~ mux_tmp_345));
  assign or_937_nl = (~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b01)
      | (rem_12cyc_st_6_3_2[0]);
  assign mux_tmp_346 = MUX_s_1_2_2(nor_381_nl, mux_tmp_345, or_937_nl);
  assign nor_382_nl = ~((rem_12cyc_st_5_3_2[1]) | (~ mux_tmp_346));
  assign or_936_nl = (~ main_stage_0_6) | (~ asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b01)
      | (rem_12cyc_st_5_3_2[0]);
  assign mux_tmp_347 = MUX_s_1_2_2(nor_382_nl, mux_tmp_346, or_936_nl);
  assign nor_383_nl = ~((rem_12cyc_st_4_3_2[1]) | (~ mux_tmp_347));
  assign or_935_nl = (~ main_stage_0_5) | (~ asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b01)
      | (rem_12cyc_st_4_3_2[0]);
  assign mux_tmp_348 = MUX_s_1_2_2(nor_383_nl, mux_tmp_347, or_935_nl);
  assign nor_384_nl = ~((rem_12cyc_st_3_3_2[1]) | (~ mux_tmp_348));
  assign or_934_nl = (~ main_stage_0_4) | (~ asn_itm_3) | (rem_12cyc_st_3_1_0!=2'b01)
      | (rem_12cyc_st_3_3_2[0]);
  assign mux_tmp_349 = MUX_s_1_2_2(nor_384_nl, mux_tmp_348, or_934_nl);
  assign nor_385_nl = ~((rem_12cyc_st_2_3_2[1]) | (~ mux_tmp_349));
  assign or_933_nl = (~ main_stage_0_3) | (~ asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b01)
      | (rem_12cyc_st_2_3_2[0]);
  assign mux_tmp_350 = MUX_s_1_2_2(nor_385_nl, mux_tmp_349, or_933_nl);
  assign nor_386_nl = ~((rem_12cyc_st_9_3_2[1]) | (~ mux_tmp_350));
  assign or_932_nl = (~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b01)
      | (rem_12cyc_st_9_3_2[0]);
  assign mux_tmp_351 = MUX_s_1_2_2(nor_386_nl, mux_tmp_350, or_932_nl);
  assign nor_387_nl = ~((rem_12cyc_st_8_3_2[1]) | (~ mux_tmp_351));
  assign or_931_nl = (~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b01)
      | (rem_12cyc_st_8_3_2[0]);
  assign mux_tmp_352 = MUX_s_1_2_2(nor_387_nl, mux_tmp_351, or_931_nl);
  assign nor_388_nl = ~((rem_12cyc_st_7_3_2[1]) | (~ mux_tmp_352));
  assign or_930_nl = (~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b01)
      | (rem_12cyc_st_7_3_2[0]);
  assign mux_tmp_353 = MUX_s_1_2_2(nor_388_nl, mux_tmp_352, or_930_nl);
  assign nor_389_nl = ~((rem_12cyc_1_0[0]) | (~ mux_tmp_353));
  assign or_929_nl = (~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b10)
      | (rem_12cyc_1_0[1]);
  assign mux_tmp_354 = MUX_s_1_2_2(nor_389_nl, mux_tmp_353, or_929_nl);
  assign and_dcpl_638 = and_dcpl_568 & and_dcpl_393;
  assign and_dcpl_639 = and_dcpl_570 & (rem_12cyc_st_2_1_0[1]);
  assign or_tmp_934 = (rem_12cyc_1_0!=2'b10) | (rem_12cyc_3_2!=2'b10) | not_tmp_54;
  assign or_952_cse = (acc_1_tmp[1:0]!=2'b10) | (acc_tmp!=2'b10);
  assign nor_379_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_934));
  assign mux_357_nl = MUX_s_1_2_2(nor_379_nl, or_tmp_934, or_952_cse);
  assign and_dcpl_641 = mux_357_nl & and_dcpl_298 & and_dcpl_639;
  assign and_dcpl_642 = and_dcpl_574 & (rem_12cyc_st_3_1_0[1]);
  assign or_957_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2!=2'b10) |
      (~ asn_itm_2) | (~ main_stage_0_3) | (rem_12cyc_st_2_1_0[0]);
  assign and_tmp_207 = or_957_cse & or_tmp_934;
  assign nor_378_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_207));
  assign mux_358_nl = MUX_s_1_2_2(nor_378_nl, and_tmp_207, or_952_cse);
  assign and_dcpl_644 = mux_358_nl & and_dcpl_304 & and_dcpl_642;
  assign and_dcpl_645 = and_dcpl_578 & (rem_12cyc_st_4_1_0[1]);
  assign or_961_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2!=2'b10) |
      (~ asn_itm_3) | (~ main_stage_0_4) | (rem_12cyc_st_3_1_0[0]);
  assign and_tmp_209 = or_957_cse & or_961_cse & or_tmp_934;
  assign nor_377_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_209));
  assign mux_359_nl = MUX_s_1_2_2(nor_377_nl, and_tmp_209, or_952_cse);
  assign and_dcpl_647 = mux_359_nl & and_dcpl_310 & and_dcpl_645;
  assign and_dcpl_648 = and_dcpl_582 & (rem_12cyc_st_5_1_0[1]);
  assign or_966_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2!=2'b10) |
      (~ asn_itm_4) | (~ main_stage_0_5) | (rem_12cyc_st_4_1_0[0]);
  assign and_tmp_212 = or_957_cse & or_961_cse & or_966_cse & or_tmp_934;
  assign nor_376_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_212));
  assign mux_360_nl = MUX_s_1_2_2(nor_376_nl, and_tmp_212, or_952_cse);
  assign and_dcpl_650 = mux_360_nl & and_dcpl_316 & and_dcpl_648;
  assign or_972_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2!=2'b10) |
      (~ asn_itm_5) | (~ main_stage_0_6) | (rem_12cyc_st_5_1_0[0]);
  assign and_tmp_216 = or_957_cse & or_961_cse & or_966_cse & or_972_cse & or_tmp_934;
  assign nor_375_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_216));
  assign mux_361_nl = MUX_s_1_2_2(nor_375_nl, and_tmp_216, or_952_cse);
  assign and_dcpl_653 = mux_361_nl & and_dcpl_112 & and_dcpl_126 & (rem_12cyc_st_6_1_0[1]);
  assign or_979_cse = (rem_12cyc_st_6_1_0!=2'b10) | (rem_12cyc_st_6_3_2!=2'b10);
  assign nor_373_nl = ~(and_dcpl_111 | (~ or_tmp_934));
  assign mux_362_nl = MUX_s_1_2_2(nor_373_nl, or_tmp_934, or_979_cse);
  assign and_tmp_220 = or_957_cse & or_961_cse & or_966_cse & or_972_cse & mux_362_nl;
  assign nor_374_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_220));
  assign mux_363_nl = MUX_s_1_2_2(nor_374_nl, and_tmp_220, or_952_cse);
  assign and_dcpl_657 = mux_363_nl & and_dcpl_85 & and_dcpl_104 & (~ (rem_12cyc_st_7_1_0[0]));
  assign or_988_cse = (rem_12cyc_st_7_1_0!=2'b10) | (rem_12cyc_st_7_3_2!=2'b10);
  assign nor_370_nl = ~(and_dcpl_84 | (~ or_tmp_934));
  assign mux_tmp_362 = MUX_s_1_2_2(nor_370_nl, or_tmp_934, or_988_cse);
  assign nor_371_nl = ~(and_dcpl_111 | (~ mux_tmp_362));
  assign mux_365_nl = MUX_s_1_2_2(nor_371_nl, mux_tmp_362, or_979_cse);
  assign and_tmp_224 = or_957_cse & or_961_cse & or_966_cse & or_972_cse & mux_365_nl;
  assign nor_372_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_224));
  assign mux_366_nl = MUX_s_1_2_2(nor_372_nl, and_tmp_224, or_952_cse);
  assign and_dcpl_661 = mux_366_nl & and_dcpl_58 & and_dcpl_77 & (~ (rem_12cyc_st_8_1_0[0]));
  assign or_999_cse = (rem_12cyc_st_8_1_0!=2'b10) | (rem_12cyc_st_8_3_2!=2'b10);
  assign nor_366_nl = ~(and_dcpl_57 | (~ or_tmp_934));
  assign mux_tmp_365 = MUX_s_1_2_2(nor_366_nl, or_tmp_934, or_999_cse);
  assign nor_367_nl = ~(and_dcpl_84 | (~ mux_tmp_365));
  assign mux_tmp_366 = MUX_s_1_2_2(nor_367_nl, mux_tmp_365, or_988_cse);
  assign nor_368_nl = ~(and_dcpl_111 | (~ mux_tmp_366));
  assign mux_369_nl = MUX_s_1_2_2(nor_368_nl, mux_tmp_366, or_979_cse);
  assign and_tmp_228 = or_957_cse & or_961_cse & or_966_cse & or_972_cse & mux_369_nl;
  assign nor_369_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_228));
  assign mux_370_nl = MUX_s_1_2_2(nor_369_nl, and_tmp_228, or_952_cse);
  assign and_dcpl_665 = mux_370_nl & and_dcpl_31 & and_dcpl_50 & (~ (rem_12cyc_st_9_1_0[0]));
  assign nor_361_nl = ~(and_dcpl_30 | (~ or_tmp_934));
  assign or_1012_nl = (rem_12cyc_st_9_1_0!=2'b10) | (rem_12cyc_st_9_3_2!=2'b10);
  assign mux_tmp_369 = MUX_s_1_2_2(nor_361_nl, or_tmp_934, or_1012_nl);
  assign nor_362_nl = ~(and_dcpl_57 | (~ mux_tmp_369));
  assign mux_tmp_370 = MUX_s_1_2_2(nor_362_nl, mux_tmp_369, or_999_cse);
  assign nor_363_nl = ~(and_dcpl_84 | (~ mux_tmp_370));
  assign mux_tmp_371 = MUX_s_1_2_2(nor_363_nl, mux_tmp_370, or_988_cse);
  assign nor_364_nl = ~(and_dcpl_111 | (~ mux_tmp_371));
  assign mux_374_nl = MUX_s_1_2_2(nor_364_nl, mux_tmp_371, or_979_cse);
  assign and_tmp_232 = or_957_cse & or_961_cse & or_966_cse & or_972_cse & mux_374_nl;
  assign nor_365_nl = ~(ccs_ccore_start_rsci_idat | (~ and_tmp_232));
  assign mux_375_nl = MUX_s_1_2_2(nor_365_nl, and_tmp_232, or_952_cse);
  assign and_dcpl_669 = mux_375_nl & and_dcpl_4 & and_dcpl_23 & (~ (rem_12cyc_st_10_1_0[0]));
  assign or_tmp_1009 = (acc_tmp!=2'b10) | (acc_1_tmp[1:0]!=2'b10) | (~ ccs_ccore_start_rsci_idat);
  assign nor_352_nl = ~((rem_12cyc_st_10_3_2[1]) | (~ or_tmp_1009));
  assign or_1027_nl = (~ main_stage_0_11) | (~ asn_itm_10) | (rem_12cyc_st_10_1_0!=2'b10)
      | (rem_12cyc_st_10_3_2[0]);
  assign mux_tmp_374 = MUX_s_1_2_2(nor_352_nl, or_tmp_1009, or_1027_nl);
  assign nor_353_nl = ~((rem_12cyc_st_6_3_2[1]) | (~ mux_tmp_374));
  assign or_1026_nl = (~ main_stage_0_7) | (~ asn_itm_6) | (rem_12cyc_st_6_1_0!=2'b10)
      | (rem_12cyc_st_6_3_2[0]);
  assign mux_tmp_375 = MUX_s_1_2_2(nor_353_nl, mux_tmp_374, or_1026_nl);
  assign nor_354_nl = ~((rem_12cyc_st_5_3_2[1]) | (~ mux_tmp_375));
  assign or_1025_nl = (~ main_stage_0_6) | (~ asn_itm_5) | (rem_12cyc_st_5_1_0!=2'b10)
      | (rem_12cyc_st_5_3_2[0]);
  assign mux_tmp_376 = MUX_s_1_2_2(nor_354_nl, mux_tmp_375, or_1025_nl);
  assign nor_355_nl = ~((rem_12cyc_st_4_3_2[1]) | (~ mux_tmp_376));
  assign or_1024_nl = (~ main_stage_0_5) | (~ asn_itm_4) | (rem_12cyc_st_4_1_0!=2'b10)
      | (rem_12cyc_st_4_3_2[0]);
  assign mux_tmp_377 = MUX_s_1_2_2(nor_355_nl, mux_tmp_376, or_1024_nl);
  assign nor_356_nl = ~((rem_12cyc_st_3_3_2[1]) | (~ mux_tmp_377));
  assign or_1023_nl = (~ main_stage_0_4) | (~ asn_itm_3) | (rem_12cyc_st_3_1_0!=2'b10)
      | (rem_12cyc_st_3_3_2[0]);
  assign mux_tmp_378 = MUX_s_1_2_2(nor_356_nl, mux_tmp_377, or_1023_nl);
  assign nor_357_nl = ~((rem_12cyc_st_2_3_2[1]) | (~ mux_tmp_378));
  assign or_1022_nl = (~ main_stage_0_3) | (~ asn_itm_2) | (rem_12cyc_st_2_1_0!=2'b10)
      | (rem_12cyc_st_2_3_2[0]);
  assign mux_tmp_379 = MUX_s_1_2_2(nor_357_nl, mux_tmp_378, or_1022_nl);
  assign nor_358_nl = ~((rem_12cyc_st_9_3_2[1]) | (~ mux_tmp_379));
  assign or_1021_nl = (~ main_stage_0_10) | (~ asn_itm_9) | (rem_12cyc_st_9_1_0!=2'b10)
      | (rem_12cyc_st_9_3_2[0]);
  assign mux_tmp_380 = MUX_s_1_2_2(nor_358_nl, mux_tmp_379, or_1021_nl);
  assign nor_359_nl = ~((rem_12cyc_st_8_3_2[1]) | (~ mux_tmp_380));
  assign or_1020_nl = (~ main_stage_0_9) | (~ asn_itm_8) | (rem_12cyc_st_8_1_0!=2'b10)
      | (rem_12cyc_st_8_3_2[0]);
  assign mux_tmp_381 = MUX_s_1_2_2(nor_359_nl, mux_tmp_380, or_1020_nl);
  assign nor_360_nl = ~((rem_12cyc_st_7_3_2[1]) | (~ mux_tmp_381));
  assign or_1019_nl = (~ main_stage_0_8) | (~ asn_itm_7) | (rem_12cyc_st_7_1_0!=2'b10)
      | (rem_12cyc_st_7_3_2[0]);
  assign mux_384_nl = MUX_s_1_2_2(nor_360_nl, mux_tmp_381, or_1019_nl);
  assign and_tmp_233 = ((~ main_stage_0_2) | (~ asn_itm_1) | (rem_12cyc_3_2!=2'b10)
      | (rem_12cyc_1_0!=2'b10)) & mux_384_nl;
  assign and_dcpl_673 = and_dcpl_568 & and_dcpl_430;
  assign or_tmp_1021 = (~((rem_12cyc_1_0==2'b11) & (rem_12cyc_3_2==2'b10))) | not_tmp_54;
  assign nand_57_cse = ~((acc_1_tmp[1:0]==2'b11) & (acc_tmp==2'b10));
  assign nor_351_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_1021));
  assign mux_385_nl = MUX_s_1_2_2(nor_351_nl, or_tmp_1021, nand_57_cse);
  assign and_dcpl_675 = mux_385_nl & and_dcpl_358 & and_dcpl_639;
  assign or_1045_cse = (~ (rem_12cyc_st_2_1_0[1])) | (rem_12cyc_st_2_3_2[0]);
  assign and_960_nl = nand_84_cse & or_tmp_1021;
  assign mux_tmp_384 = MUX_s_1_2_2(and_960_nl, or_tmp_1021, or_1045_cse);
  assign nor_350_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_384));
  assign mux_387_nl = MUX_s_1_2_2(nor_350_nl, mux_tmp_384, nand_57_cse);
  assign and_dcpl_677 = mux_387_nl & and_dcpl_362 & and_dcpl_642;
  assign or_1050_cse = (~ (rem_12cyc_st_3_1_0[1])) | (rem_12cyc_st_3_3_2!=2'b10);
  assign and_958_nl = nand_274_cse & or_tmp_1021;
  assign mux_tmp_386 = MUX_s_1_2_2(and_958_nl, or_tmp_1021, or_1050_cse);
  assign and_959_nl = nand_84_cse & mux_tmp_386;
  assign mux_tmp_387 = MUX_s_1_2_2(and_959_nl, mux_tmp_386, or_1045_cse);
  assign nor_349_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_387));
  assign mux_390_nl = MUX_s_1_2_2(nor_349_nl, mux_tmp_387, nand_57_cse);
  assign and_dcpl_679 = mux_390_nl & and_dcpl_366 & and_dcpl_645;
  assign or_1057_cse = (~ (rem_12cyc_st_4_1_0[1])) | (rem_12cyc_st_4_3_2[0]);
  assign and_955_nl = nand_79_cse & or_tmp_1021;
  assign mux_tmp_389 = MUX_s_1_2_2(and_955_nl, or_tmp_1021, or_1057_cse);
  assign and_956_nl = nand_274_cse & mux_tmp_389;
  assign mux_tmp_390 = MUX_s_1_2_2(and_956_nl, mux_tmp_389, or_1050_cse);
  assign and_957_nl = nand_84_cse & mux_tmp_390;
  assign mux_tmp_391 = MUX_s_1_2_2(and_957_nl, mux_tmp_390, or_1045_cse);
  assign nor_348_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_391));
  assign mux_394_nl = MUX_s_1_2_2(nor_348_nl, mux_tmp_391, nand_57_cse);
  assign and_dcpl_681 = mux_394_nl & and_dcpl_370 & and_dcpl_648;
  assign or_1066_cse = (~ (rem_12cyc_st_5_1_0[1])) | (rem_12cyc_st_5_3_2!=2'b10);
  assign and_951_nl = nand_267_cse & or_tmp_1021;
  assign mux_tmp_393 = MUX_s_1_2_2(and_951_nl, or_tmp_1021, or_1066_cse);
  assign and_952_nl = nand_79_cse & mux_tmp_393;
  assign mux_tmp_394 = MUX_s_1_2_2(and_952_nl, mux_tmp_393, or_1057_cse);
  assign and_953_nl = nand_274_cse & mux_tmp_394;
  assign mux_tmp_395 = MUX_s_1_2_2(and_953_nl, mux_tmp_394, or_1050_cse);
  assign and_954_nl = nand_84_cse & mux_tmp_395;
  assign mux_tmp_396 = MUX_s_1_2_2(and_954_nl, mux_tmp_395, or_1045_cse);
  assign nor_347_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_396));
  assign mux_399_nl = MUX_s_1_2_2(nor_347_nl, mux_tmp_396, nand_57_cse);
  assign and_dcpl_684 = mux_399_nl & and_dcpl_112 & and_dcpl_129 & (rem_12cyc_st_6_1_0[1]);
  assign nand_36_cse = ~((rem_12cyc_st_6_1_0==2'b11) & (rem_12cyc_st_6_3_2==2'b10));
  assign nor_345_nl = ~(and_dcpl_111 | (~ or_tmp_1021));
  assign mux_tmp_398 = MUX_s_1_2_2(nor_345_nl, or_tmp_1021, nand_36_cse);
  assign and_947_nl = nand_267_cse & mux_tmp_398;
  assign mux_tmp_399 = MUX_s_1_2_2(and_947_nl, mux_tmp_398, or_1066_cse);
  assign and_948_nl = nand_79_cse & mux_tmp_399;
  assign mux_tmp_400 = MUX_s_1_2_2(and_948_nl, mux_tmp_399, or_1057_cse);
  assign and_949_nl = nand_274_cse & mux_tmp_400;
  assign mux_tmp_401 = MUX_s_1_2_2(and_949_nl, mux_tmp_400, or_1050_cse);
  assign and_950_nl = nand_84_cse & mux_tmp_401;
  assign mux_tmp_402 = MUX_s_1_2_2(and_950_nl, mux_tmp_401, or_1045_cse);
  assign nor_346_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_402));
  assign mux_405_nl = MUX_s_1_2_2(nor_346_nl, mux_tmp_402, nand_57_cse);
  assign and_dcpl_687 = mux_405_nl & and_dcpl_85 & and_dcpl_104 & (rem_12cyc_st_7_1_0[0]);
  assign nand_29_cse = ~((rem_12cyc_st_7_1_0==2'b11) & (rem_12cyc_st_7_3_2==2'b10));
  assign nor_342_nl = ~(and_dcpl_84 | (~ or_tmp_1021));
  assign mux_tmp_404 = MUX_s_1_2_2(nor_342_nl, or_tmp_1021, nand_29_cse);
  assign nor_343_nl = ~(and_dcpl_111 | (~ mux_tmp_404));
  assign mux_tmp_405 = MUX_s_1_2_2(nor_343_nl, mux_tmp_404, nand_36_cse);
  assign and_943_nl = nand_267_cse & mux_tmp_405;
  assign mux_tmp_406 = MUX_s_1_2_2(and_943_nl, mux_tmp_405, or_1066_cse);
  assign and_944_nl = nand_79_cse & mux_tmp_406;
  assign mux_tmp_407 = MUX_s_1_2_2(and_944_nl, mux_tmp_406, or_1057_cse);
  assign and_945_nl = nand_274_cse & mux_tmp_407;
  assign mux_tmp_408 = MUX_s_1_2_2(and_945_nl, mux_tmp_407, or_1050_cse);
  assign and_946_nl = nand_84_cse & mux_tmp_408;
  assign mux_tmp_409 = MUX_s_1_2_2(and_946_nl, mux_tmp_408, or_1045_cse);
  assign nor_344_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_409));
  assign mux_412_nl = MUX_s_1_2_2(nor_344_nl, mux_tmp_409, nand_57_cse);
  assign and_dcpl_690 = mux_412_nl & and_dcpl_58 & and_dcpl_77 & (rem_12cyc_st_8_1_0[0]);
  assign nand_21_cse = ~((rem_12cyc_st_8_1_0==2'b11) & (rem_12cyc_st_8_3_2==2'b10));
  assign nor_338_nl = ~(and_dcpl_57 | (~ or_tmp_1021));
  assign mux_tmp_411 = MUX_s_1_2_2(nor_338_nl, or_tmp_1021, nand_21_cse);
  assign nor_339_nl = ~(and_dcpl_84 | (~ mux_tmp_411));
  assign mux_tmp_412 = MUX_s_1_2_2(nor_339_nl, mux_tmp_411, nand_29_cse);
  assign nor_340_nl = ~(and_dcpl_111 | (~ mux_tmp_412));
  assign mux_tmp_413 = MUX_s_1_2_2(nor_340_nl, mux_tmp_412, nand_36_cse);
  assign and_939_nl = nand_267_cse & mux_tmp_413;
  assign mux_tmp_414 = MUX_s_1_2_2(and_939_nl, mux_tmp_413, or_1066_cse);
  assign and_940_nl = nand_79_cse & mux_tmp_414;
  assign mux_tmp_415 = MUX_s_1_2_2(and_940_nl, mux_tmp_414, or_1057_cse);
  assign and_941_nl = nand_274_cse & mux_tmp_415;
  assign mux_tmp_416 = MUX_s_1_2_2(and_941_nl, mux_tmp_415, or_1050_cse);
  assign and_942_nl = nand_84_cse & mux_tmp_416;
  assign mux_tmp_417 = MUX_s_1_2_2(and_942_nl, mux_tmp_416, or_1045_cse);
  assign nor_341_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_417));
  assign mux_420_nl = MUX_s_1_2_2(nor_341_nl, mux_tmp_417, nand_57_cse);
  assign and_dcpl_693 = mux_420_nl & and_dcpl_31 & and_dcpl_50 & (rem_12cyc_st_9_1_0[0]);
  assign nor_333_nl = ~(and_dcpl_30 | (~ or_tmp_1021));
  assign nand_12_nl = ~((rem_12cyc_st_9_1_0==2'b11) & (rem_12cyc_st_9_3_2==2'b10));
  assign mux_tmp_419 = MUX_s_1_2_2(nor_333_nl, or_tmp_1021, nand_12_nl);
  assign nor_334_nl = ~(and_dcpl_57 | (~ mux_tmp_419));
  assign mux_tmp_420 = MUX_s_1_2_2(nor_334_nl, mux_tmp_419, nand_21_cse);
  assign nor_335_nl = ~(and_dcpl_84 | (~ mux_tmp_420));
  assign mux_tmp_421 = MUX_s_1_2_2(nor_335_nl, mux_tmp_420, nand_29_cse);
  assign nor_336_nl = ~(and_dcpl_111 | (~ mux_tmp_421));
  assign mux_tmp_422 = MUX_s_1_2_2(nor_336_nl, mux_tmp_421, nand_36_cse);
  assign and_935_nl = nand_267_cse & mux_tmp_422;
  assign mux_tmp_423 = MUX_s_1_2_2(and_935_nl, mux_tmp_422, or_1066_cse);
  assign and_936_nl = nand_79_cse & mux_tmp_423;
  assign mux_tmp_424 = MUX_s_1_2_2(and_936_nl, mux_tmp_423, or_1057_cse);
  assign and_937_nl = nand_274_cse & mux_tmp_424;
  assign mux_tmp_425 = MUX_s_1_2_2(and_937_nl, mux_tmp_424, or_1050_cse);
  assign and_938_nl = nand_84_cse & mux_tmp_425;
  assign mux_tmp_426 = MUX_s_1_2_2(and_938_nl, mux_tmp_425, or_1045_cse);
  assign nor_337_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_426));
  assign mux_429_nl = MUX_s_1_2_2(nor_337_nl, mux_tmp_426, nand_57_cse);
  assign and_dcpl_696 = mux_429_nl & and_dcpl_4 & and_dcpl_23 & (rem_12cyc_st_10_1_0[0]);
  assign or_tmp_1122 = (acc_tmp!=2'b10) | nand_222_cse;
  assign nor_324_nl = ~((rem_12cyc_st_10_3_2[1]) | (~ or_tmp_1122));
  assign nand_1_nl = ~(main_stage_0_11 & asn_itm_10 & (rem_12cyc_st_10_1_0==2'b11)
      & (~ (rem_12cyc_st_10_3_2[0])));
  assign mux_tmp_428 = MUX_s_1_2_2(nor_324_nl, or_tmp_1122, nand_1_nl);
  assign nor_325_nl = ~((rem_12cyc_st_6_3_2[1]) | (~ mux_tmp_428));
  assign nand_2_nl = ~(main_stage_0_7 & asn_itm_6 & (rem_12cyc_st_6_1_0==2'b11) &
      (~ (rem_12cyc_st_6_3_2[0])));
  assign mux_tmp_429 = MUX_s_1_2_2(nor_325_nl, mux_tmp_428, nand_2_nl);
  assign nor_326_nl = ~((rem_12cyc_st_5_3_2[1]) | (~ mux_tmp_429));
  assign nand_3_nl = ~(main_stage_0_6 & asn_itm_5 & (rem_12cyc_st_5_1_0==2'b11) &
      (~ (rem_12cyc_st_5_3_2[0])));
  assign mux_tmp_430 = MUX_s_1_2_2(nor_326_nl, mux_tmp_429, nand_3_nl);
  assign nor_327_nl = ~((rem_12cyc_st_4_3_2[1]) | (~ mux_tmp_430));
  assign nand_4_nl = ~(main_stage_0_5 & asn_itm_4 & (rem_12cyc_st_4_1_0==2'b11) &
      (~ (rem_12cyc_st_4_3_2[0])));
  assign mux_tmp_431 = MUX_s_1_2_2(nor_327_nl, mux_tmp_430, nand_4_nl);
  assign nor_328_nl = ~((rem_12cyc_st_3_3_2[1]) | (~ mux_tmp_431));
  assign nand_5_nl = ~(main_stage_0_4 & asn_itm_3 & (rem_12cyc_st_3_1_0==2'b11) &
      (~ (rem_12cyc_st_3_3_2[0])));
  assign mux_tmp_432 = MUX_s_1_2_2(nor_328_nl, mux_tmp_431, nand_5_nl);
  assign nor_329_nl = ~((rem_12cyc_st_2_3_2[1]) | (~ mux_tmp_432));
  assign nand_6_nl = ~(main_stage_0_3 & asn_itm_2 & (rem_12cyc_st_2_1_0==2'b11) &
      (~ (rem_12cyc_st_2_3_2[0])));
  assign mux_tmp_433 = MUX_s_1_2_2(nor_329_nl, mux_tmp_432, nand_6_nl);
  assign nor_330_nl = ~((rem_12cyc_st_9_3_2[1]) | (~ mux_tmp_433));
  assign nand_7_nl = ~(main_stage_0_10 & asn_itm_9 & (rem_12cyc_st_9_1_0==2'b11)
      & (~ (rem_12cyc_st_9_3_2[0])));
  assign mux_tmp_434 = MUX_s_1_2_2(nor_330_nl, mux_tmp_433, nand_7_nl);
  assign nor_331_nl = ~((rem_12cyc_st_8_3_2[1]) | (~ mux_tmp_434));
  assign nand_8_nl = ~(main_stage_0_9 & asn_itm_8 & (rem_12cyc_st_8_1_0==2'b11) &
      (~ (rem_12cyc_st_8_3_2[0])));
  assign mux_tmp_435 = MUX_s_1_2_2(nor_331_nl, mux_tmp_434, nand_8_nl);
  assign nor_332_nl = ~((rem_12cyc_st_7_3_2[1]) | (~ mux_tmp_435));
  assign nand_9_nl = ~(main_stage_0_8 & asn_itm_7 & (rem_12cyc_st_7_1_0==2'b11) &
      (~ (rem_12cyc_st_7_3_2[0])));
  assign mux_tmp_436 = MUX_s_1_2_2(nor_332_nl, mux_tmp_435, nand_9_nl);
  assign and_934_nl = nand_223_cse & mux_tmp_436;
  assign nand_11_nl = ~(main_stage_0_2 & asn_itm_1 & (rem_12cyc_3_2==2'b10));
  assign mux_tmp_437 = MUX_s_1_2_2(and_934_nl, mux_tmp_436, nand_11_nl);
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_en ) begin
      return_rsci_d <= MUX_v_64_2_2(result_sva_duc_mx0, qelse_acc_nl, mux_13_nl);
      m_buf_sva_12 <= m_buf_sva_11;
      m_buf_sva_11 <= m_buf_sva_10;
      m_buf_sva_10 <= m_buf_sva_9;
      m_buf_sva_9 <= m_buf_sva_8;
      m_buf_sva_8 <= m_buf_sva_7;
      m_buf_sva_7 <= m_buf_sva_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      asn_itm_12 <= 1'b0;
      asn_itm_11 <= 1'b0;
      asn_itm_10 <= 1'b0;
      asn_itm_9 <= 1'b0;
      asn_itm_8 <= 1'b0;
      asn_itm_7 <= 1'b0;
      asn_itm_6 <= 1'b0;
      asn_itm_5 <= 1'b0;
      asn_itm_4 <= 1'b0;
      asn_itm_3 <= 1'b0;
      asn_itm_2 <= 1'b0;
      asn_itm_1 <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
      main_stage_0_5 <= 1'b0;
      main_stage_0_6 <= 1'b0;
      main_stage_0_7 <= 1'b0;
      main_stage_0_8 <= 1'b0;
      main_stage_0_9 <= 1'b0;
      main_stage_0_10 <= 1'b0;
      main_stage_0_11 <= 1'b0;
      main_stage_0_12 <= 1'b0;
      main_stage_0_13 <= 1'b0;
    end
    else if ( ccs_ccore_en ) begin
      asn_itm_12 <= asn_itm_11;
      asn_itm_11 <= asn_itm_10;
      asn_itm_10 <= asn_itm_9;
      asn_itm_9 <= asn_itm_8;
      asn_itm_8 <= asn_itm_7;
      asn_itm_7 <= asn_itm_6;
      asn_itm_6 <= asn_itm_5;
      asn_itm_5 <= asn_itm_4;
      asn_itm_4 <= asn_itm_3;
      asn_itm_3 <= asn_itm_2;
      asn_itm_2 <= asn_itm_1;
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
      main_stage_0_4 <= main_stage_0_3;
      main_stage_0_5 <= main_stage_0_4;
      main_stage_0_6 <= main_stage_0_5;
      main_stage_0_7 <= main_stage_0_6;
      main_stage_0_8 <= main_stage_0_7;
      main_stage_0_9 <= main_stage_0_8;
      main_stage_0_10 <= main_stage_0_9;
      main_stage_0_11 <= main_stage_0_10;
      main_stage_0_12 <= main_stage_0_11;
      main_stage_0_13 <= main_stage_0_12;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_sva_duc <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( asn_itm_12 & main_stage_0_13 & ccs_ccore_en & (~((rem_12cyc_st_12_3_2==2'b11)))
        ) begin
      result_sva_duc <= result_sva_duc_mx0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_12_3_2 <= 2'b00;
      rem_12cyc_st_12_1_0 <= 2'b00;
    end
    else if ( and_1203_cse ) begin
      rem_12cyc_st_12_3_2 <= rem_12cyc_st_11_3_2;
      rem_12cyc_st_12_1_0 <= rem_12cyc_st_11_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1173_cse ) begin
      rem_13_cmp_1_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_3_2_63_0, mut_3_3_63_0,
          mut_3_4_63_0, mut_3_5_63_0, mut_3_6_63_0, mut_3_7_63_0, mut_3_8_63_0, mut_3_9_63_0,
          mut_3_10_63_0, mut_3_11_63_0, {and_dcpl_294 , and_dcpl_300 , and_dcpl_306
          , and_dcpl_312 , and_dcpl_318 , and_dcpl_324 , and_dcpl_330 , and_dcpl_336
          , and_dcpl_342 , and_dcpl_348 , and_tmp_35});
      rem_13_cmp_1_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_2_2_63_0, mut_2_3_63_0,
          mut_2_4_63_0, mut_2_5_63_0, mut_2_6_63_0, mut_2_7_63_0, mut_2_8_63_0, mut_2_9_63_0,
          mut_2_10_63_0, mut_2_11_63_0, {and_dcpl_294 , and_dcpl_300 , and_dcpl_306
          , and_dcpl_312 , and_dcpl_318 , and_dcpl_324 , and_dcpl_330 , and_dcpl_336
          , and_dcpl_342 , and_dcpl_348 , and_tmp_35});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1175_cse ) begin
      rem_13_cmp_2_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_5_2_63_0, mut_5_3_63_0,
          mut_5_4_63_0, mut_5_5_63_0, mut_5_6_63_0, mut_5_7_63_0, mut_5_8_63_0, mut_5_9_63_0,
          mut_5_10_63_0, mut_5_11_63_0, {and_dcpl_356 , and_dcpl_360 , and_dcpl_364
          , and_dcpl_368 , and_dcpl_372 , and_dcpl_376 , and_dcpl_379 , and_dcpl_382
          , and_dcpl_385 , and_dcpl_388 , mux_tmp_76});
      rem_13_cmp_2_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_4_2_63_0, mut_4_3_63_0,
          mut_4_4_63_0, mut_4_5_63_0, mut_4_6_63_0, mut_4_7_63_0, mut_4_8_63_0, mut_4_9_63_0,
          mut_4_10_63_0, mut_4_11_63_0, {and_dcpl_356 , and_dcpl_360 , and_dcpl_364
          , and_dcpl_368 , and_dcpl_372 , and_dcpl_376 , and_dcpl_379 , and_dcpl_382
          , and_dcpl_385 , and_dcpl_388 , mux_tmp_76});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1177_cse ) begin
      rem_13_cmp_3_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_7_2_63_0, mut_7_3_63_0,
          mut_7_4_63_0, mut_7_5_63_0, mut_7_6_63_0, mut_7_7_63_0, mut_7_8_63_0, mut_7_9_63_0,
          mut_7_10_63_0, mut_7_11_63_0, {and_dcpl_394 , and_dcpl_397 , and_dcpl_400
          , and_dcpl_403 , and_dcpl_406 , and_dcpl_409 , and_dcpl_413 , and_dcpl_417
          , and_dcpl_421 , and_dcpl_425 , and_tmp_80});
      rem_13_cmp_3_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_6_2_63_0, mut_6_3_63_0,
          mut_6_4_63_0, mut_6_5_63_0, mut_6_6_63_0, mut_6_7_63_0, mut_6_8_63_0, mut_6_9_63_0,
          mut_6_10_63_0, mut_6_11_63_0, {and_dcpl_394 , and_dcpl_397 , and_dcpl_400
          , and_dcpl_403 , and_dcpl_406 , and_dcpl_409 , and_dcpl_413 , and_dcpl_417
          , and_dcpl_421 , and_dcpl_425 , and_tmp_80});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1179_cse ) begin
      rem_13_cmp_4_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_9_2_63_0, mut_9_3_63_0,
          mut_9_4_63_0, mut_9_5_63_0, mut_9_6_63_0, mut_9_7_63_0, mut_9_8_63_0, mut_9_9_63_0,
          mut_9_10_63_0, mut_9_11_63_0, {and_dcpl_431 , and_dcpl_433 , and_dcpl_435
          , and_dcpl_437 , and_dcpl_439 , and_dcpl_442 , and_dcpl_445 , and_dcpl_448
          , and_dcpl_451 , and_dcpl_454 , mux_tmp_141});
      rem_13_cmp_4_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_8_2_63_0, mut_8_3_63_0,
          mut_8_4_63_0, mut_8_5_63_0, mut_8_6_63_0, mut_8_7_63_0, mut_8_8_63_0, mut_8_9_63_0,
          mut_8_10_63_0, mut_8_11_63_0, {and_dcpl_431 , and_dcpl_433 , and_dcpl_435
          , and_dcpl_437 , and_dcpl_439 , and_dcpl_442 , and_dcpl_445 , and_dcpl_448
          , and_dcpl_451 , and_dcpl_454 , mux_tmp_141});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1181_cse ) begin
      rem_13_cmp_5_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_11_2_63_0, mut_11_3_63_0,
          mut_11_4_63_0, mut_11_5_63_0, mut_11_6_63_0, mut_11_7_63_0, mut_11_8_63_0,
          mut_11_9_63_0, mut_11_10_63_0, mut_11_11_63_0, {and_dcpl_461 , and_dcpl_465
          , and_dcpl_469 , and_dcpl_473 , and_dcpl_477 , and_dcpl_480 , and_dcpl_483
          , and_dcpl_486 , and_dcpl_489 , and_dcpl_492 , and_tmp_125});
      rem_13_cmp_5_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_10_2_63_0, mut_10_3_63_0,
          mut_10_4_63_0, mut_10_5_63_0, mut_10_6_63_0, mut_10_7_63_0, mut_10_8_63_0,
          mut_10_9_63_0, mut_10_10_63_0, mut_10_11_63_0, {and_dcpl_461 , and_dcpl_465
          , and_dcpl_469 , and_dcpl_473 , and_dcpl_477 , and_dcpl_480 , and_dcpl_483
          , and_dcpl_486 , and_dcpl_489 , and_dcpl_492 , and_tmp_125});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1183_cse ) begin
      rem_13_cmp_6_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_13_2_63_0, mut_13_3_63_0,
          mut_13_4_63_0, mut_13_5_63_0, mut_13_6_63_0, mut_13_7_63_0, mut_13_8_63_0,
          mut_13_9_63_0, mut_13_10_63_0, mut_13_11_63_0, {and_dcpl_498 , and_dcpl_500
          , and_dcpl_502 , and_dcpl_504 , and_dcpl_506 , and_dcpl_508 , and_dcpl_510
          , and_dcpl_512 , and_dcpl_514 , and_dcpl_516 , mux_tmp_206});
      rem_13_cmp_6_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_12_2_63_0, mut_12_3_63_0,
          mut_12_4_63_0, mut_12_5_63_0, mut_12_6_63_0, mut_12_7_63_0, mut_12_8_63_0,
          mut_12_9_63_0, mut_12_10_63_0, mut_12_11_63_0, {and_dcpl_498 , and_dcpl_500
          , and_dcpl_502 , and_dcpl_504 , and_dcpl_506 , and_dcpl_508 , and_dcpl_510
          , and_dcpl_512 , and_dcpl_514 , and_dcpl_516 , mux_tmp_206});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1185_cse ) begin
      rem_13_cmp_7_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_15_2_63_0, mut_15_3_63_0,
          mut_15_4_63_0, mut_15_5_63_0, mut_15_6_63_0, mut_15_7_63_0, mut_15_8_63_0,
          mut_15_9_63_0, mut_15_10_63_0, mut_15_11_63_0, {and_dcpl_520 , and_dcpl_523
          , and_dcpl_526 , and_dcpl_529 , and_dcpl_532 , and_dcpl_534 , and_dcpl_536
          , and_dcpl_538 , and_dcpl_540 , and_dcpl_542 , and_tmp_170});
      rem_13_cmp_7_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_14_2_63_0, mut_14_3_63_0,
          mut_14_4_63_0, mut_14_5_63_0, mut_14_6_63_0, mut_14_7_63_0, mut_14_8_63_0,
          mut_14_9_63_0, mut_14_10_63_0, mut_14_11_63_0, {and_dcpl_520 , and_dcpl_523
          , and_dcpl_526 , and_dcpl_529 , and_dcpl_532 , and_dcpl_534 , and_dcpl_536
          , and_dcpl_538 , and_dcpl_540 , and_dcpl_542 , and_tmp_170});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1187_cse ) begin
      rem_13_cmp_8_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_17_2_63_0, mut_17_3_63_0,
          mut_17_4_63_0, mut_17_5_63_0, mut_17_6_63_0, mut_17_7_63_0, mut_17_8_63_0,
          mut_17_9_63_0, mut_17_10_63_0, mut_17_11_63_0, {and_dcpl_546 , and_dcpl_548
          , and_dcpl_550 , and_dcpl_552 , and_dcpl_554 , and_dcpl_556 , and_dcpl_558
          , and_dcpl_560 , and_dcpl_562 , and_dcpl_564 , mux_tmp_271});
      rem_13_cmp_8_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_16_2_63_0, mut_16_3_63_0,
          mut_16_4_63_0, mut_16_5_63_0, mut_16_6_63_0, mut_16_7_63_0, mut_16_8_63_0,
          mut_16_9_63_0, mut_16_10_63_0, mut_16_11_63_0, {and_dcpl_546 , and_dcpl_548
          , and_dcpl_550 , and_dcpl_552 , and_dcpl_554 , and_dcpl_556 , and_dcpl_558
          , and_dcpl_560 , and_dcpl_562 , and_dcpl_564 , mux_tmp_271});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1189_cse ) begin
      rem_13_cmp_9_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_19_2_63_0, mut_19_3_63_0,
          mut_19_4_63_0, mut_19_5_63_0, mut_19_6_63_0, mut_19_7_63_0, mut_19_8_63_0,
          mut_19_9_63_0, mut_19_10_63_0, mut_19_11_63_0, {and_dcpl_569 , and_dcpl_573
          , and_dcpl_577 , and_dcpl_581 , and_dcpl_585 , and_dcpl_589 , and_dcpl_593
          , and_dcpl_597 , and_dcpl_601 , and_dcpl_605 , and_tmp_206});
      rem_13_cmp_9_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_18_2_63_0, mut_18_3_63_0,
          mut_18_4_63_0, mut_18_5_63_0, mut_18_6_63_0, mut_18_7_63_0, mut_18_8_63_0,
          mut_18_9_63_0, mut_18_10_63_0, mut_18_11_63_0, {and_dcpl_569 , and_dcpl_573
          , and_dcpl_577 , and_dcpl_581 , and_dcpl_585 , and_dcpl_589 , and_dcpl_593
          , and_dcpl_597 , and_dcpl_601 , and_dcpl_605 , and_tmp_206});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1191_cse ) begin
      rem_13_cmp_10_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_21_2_63_0, mut_21_3_63_0,
          mut_21_4_63_0, mut_21_5_63_0, mut_21_6_63_0, mut_21_7_63_0, mut_21_8_63_0,
          mut_21_9_63_0, mut_21_10_63_0, mut_21_11_63_0, {and_dcpl_610 , and_dcpl_612
          , and_dcpl_614 , and_dcpl_616 , and_dcpl_618 , and_dcpl_622 , and_dcpl_625
          , and_dcpl_628 , and_dcpl_631 , and_dcpl_634 , mux_tmp_354});
      rem_13_cmp_10_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_20_2_63_0, mut_20_3_63_0,
          mut_20_4_63_0, mut_20_5_63_0, mut_20_6_63_0, mut_20_7_63_0, mut_20_8_63_0,
          mut_20_9_63_0, mut_20_10_63_0, mut_20_11_63_0, {and_dcpl_610 , and_dcpl_612
          , and_dcpl_614 , and_dcpl_616 , and_dcpl_618 , and_dcpl_622 , and_dcpl_625
          , and_dcpl_628 , and_dcpl_631 , and_dcpl_634 , mux_tmp_354});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1193_cse ) begin
      rem_13_cmp_11_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_23_2_63_0, mut_23_3_63_0,
          mut_23_4_63_0, mut_23_5_63_0, mut_23_6_63_0, mut_23_7_63_0, mut_23_8_63_0,
          mut_23_9_63_0, mut_23_10_63_0, mut_23_11_63_0, {and_dcpl_638 , and_dcpl_641
          , and_dcpl_644 , and_dcpl_647 , and_dcpl_650 , and_dcpl_653 , and_dcpl_657
          , and_dcpl_661 , and_dcpl_665 , and_dcpl_669 , and_tmp_233});
      rem_13_cmp_11_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_22_2_63_0, mut_22_3_63_0,
          mut_22_4_63_0, mut_22_5_63_0, mut_22_6_63_0, mut_22_7_63_0, mut_22_8_63_0,
          mut_22_9_63_0, mut_22_10_63_0, mut_22_11_63_0, {and_dcpl_638 , and_dcpl_641
          , and_dcpl_644 , and_dcpl_647 , and_dcpl_650 , and_dcpl_653 , and_dcpl_657
          , and_dcpl_661 , and_dcpl_665 , and_dcpl_669 , and_tmp_233});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1195_cse ) begin
      rem_13_cmp_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_1_2_63_0, mut_1_3_63_0,
          mut_1_4_63_0, mut_1_5_63_0, mut_1_6_63_0, mut_1_7_63_0, mut_1_8_63_0, mut_1_9_63_0,
          mut_1_10_63_0, mut_1_11_63_0, {and_dcpl_673 , and_dcpl_675 , and_dcpl_677
          , and_dcpl_679 , and_dcpl_681 , and_dcpl_684 , and_dcpl_687 , and_dcpl_690
          , and_dcpl_693 , and_dcpl_696 , mux_tmp_437});
      rem_13_cmp_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_2_63_0, mut_3_63_0,
          mut_4_63_0, mut_5_63_0, mut_6_63_0, mut_7_63_0, mut_8_63_0, mut_9_63_0,
          mut_10_63_0, mut_11_63_0, {and_dcpl_673 , and_dcpl_675 , and_dcpl_677 ,
          and_dcpl_679 , and_dcpl_681 , and_dcpl_684 , and_dcpl_687 , and_dcpl_690
          , and_dcpl_693 , and_dcpl_696 , mux_tmp_437});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1205_cse ) begin
      mut_3_11_63_0 <= mut_3_10_63_0;
      mut_2_11_63_0 <= mut_2_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1207_cse ) begin
      mut_5_11_63_0 <= mut_5_10_63_0;
      mut_4_11_63_0 <= mut_4_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1209_cse ) begin
      mut_7_11_63_0 <= mut_7_10_63_0;
      mut_6_11_63_0 <= mut_6_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1211_cse ) begin
      mut_9_11_63_0 <= mut_9_10_63_0;
      mut_8_11_63_0 <= mut_8_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1213_cse ) begin
      mut_11_11_63_0 <= mut_11_10_63_0;
      mut_10_11_63_0 <= mut_10_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1215_cse ) begin
      mut_13_11_63_0 <= mut_13_10_63_0;
      mut_12_11_63_0 <= mut_12_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1217_cse ) begin
      mut_15_11_63_0 <= mut_15_10_63_0;
      mut_14_11_63_0 <= mut_14_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1219_cse ) begin
      mut_17_11_63_0 <= mut_17_10_63_0;
      mut_16_11_63_0 <= mut_16_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1221_cse ) begin
      mut_19_11_63_0 <= mut_19_10_63_0;
      mut_18_11_63_0 <= mut_18_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1223_cse ) begin
      mut_21_11_63_0 <= mut_21_10_63_0;
      mut_20_11_63_0 <= mut_20_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1225_cse ) begin
      mut_23_11_63_0 <= mut_23_10_63_0;
      mut_22_11_63_0 <= mut_22_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1227_cse ) begin
      mut_1_11_63_0 <= mut_1_10_63_0;
      mut_11_63_0 <= mut_10_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_11_3_2 <= 2'b00;
      rem_12cyc_st_11_1_0 <= 2'b00;
    end
    else if ( and_1229_cse ) begin
      rem_12cyc_st_11_3_2 <= rem_12cyc_st_10_3_2;
      rem_12cyc_st_11_1_0 <= rem_12cyc_st_10_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1231_cse ) begin
      mut_3_10_63_0 <= mut_3_9_63_0;
      mut_2_10_63_0 <= mut_2_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1233_cse ) begin
      mut_5_10_63_0 <= mut_5_9_63_0;
      mut_4_10_63_0 <= mut_4_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1235_cse ) begin
      mut_7_10_63_0 <= mut_7_9_63_0;
      mut_6_10_63_0 <= mut_6_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1237_cse ) begin
      mut_9_10_63_0 <= mut_9_9_63_0;
      mut_8_10_63_0 <= mut_8_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1239_cse ) begin
      mut_11_10_63_0 <= mut_11_9_63_0;
      mut_10_10_63_0 <= mut_10_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1241_cse ) begin
      mut_13_10_63_0 <= mut_13_9_63_0;
      mut_12_10_63_0 <= mut_12_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1243_cse ) begin
      mut_15_10_63_0 <= mut_15_9_63_0;
      mut_14_10_63_0 <= mut_14_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1245_cse ) begin
      mut_17_10_63_0 <= mut_17_9_63_0;
      mut_16_10_63_0 <= mut_16_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1247_cse ) begin
      mut_19_10_63_0 <= mut_19_9_63_0;
      mut_18_10_63_0 <= mut_18_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1249_cse ) begin
      mut_21_10_63_0 <= mut_21_9_63_0;
      mut_20_10_63_0 <= mut_20_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1251_cse ) begin
      mut_23_10_63_0 <= mut_23_9_63_0;
      mut_22_10_63_0 <= mut_22_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1253_cse ) begin
      mut_1_10_63_0 <= mut_1_9_63_0;
      mut_10_63_0 <= mut_9_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_10_3_2 <= 2'b00;
      rem_12cyc_st_10_1_0 <= 2'b00;
    end
    else if ( and_1255_cse ) begin
      rem_12cyc_st_10_3_2 <= rem_12cyc_st_9_3_2;
      rem_12cyc_st_10_1_0 <= rem_12cyc_st_9_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1257_cse ) begin
      mut_3_9_63_0 <= mut_3_8_63_0;
      mut_2_9_63_0 <= mut_2_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1259_cse ) begin
      mut_5_9_63_0 <= mut_5_8_63_0;
      mut_4_9_63_0 <= mut_4_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1261_cse ) begin
      mut_7_9_63_0 <= mut_7_8_63_0;
      mut_6_9_63_0 <= mut_6_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1263_cse ) begin
      mut_9_9_63_0 <= mut_9_8_63_0;
      mut_8_9_63_0 <= mut_8_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1265_cse ) begin
      mut_11_9_63_0 <= mut_11_8_63_0;
      mut_10_9_63_0 <= mut_10_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1267_cse ) begin
      mut_13_9_63_0 <= mut_13_8_63_0;
      mut_12_9_63_0 <= mut_12_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1269_cse ) begin
      mut_15_9_63_0 <= mut_15_8_63_0;
      mut_14_9_63_0 <= mut_14_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1271_cse ) begin
      mut_17_9_63_0 <= mut_17_8_63_0;
      mut_16_9_63_0 <= mut_16_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1273_cse ) begin
      mut_19_9_63_0 <= mut_19_8_63_0;
      mut_18_9_63_0 <= mut_18_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1275_cse ) begin
      mut_21_9_63_0 <= mut_21_8_63_0;
      mut_20_9_63_0 <= mut_20_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1277_cse ) begin
      mut_23_9_63_0 <= mut_23_8_63_0;
      mut_22_9_63_0 <= mut_22_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1279_cse ) begin
      mut_1_9_63_0 <= mut_1_8_63_0;
      mut_9_63_0 <= mut_8_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_9_3_2 <= 2'b00;
      rem_12cyc_st_9_1_0 <= 2'b00;
    end
    else if ( and_1281_cse ) begin
      rem_12cyc_st_9_3_2 <= rem_12cyc_st_8_3_2;
      rem_12cyc_st_9_1_0 <= rem_12cyc_st_8_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1283_cse ) begin
      mut_3_8_63_0 <= mut_3_7_63_0;
      mut_2_8_63_0 <= mut_2_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1285_cse ) begin
      mut_5_8_63_0 <= mut_5_7_63_0;
      mut_4_8_63_0 <= mut_4_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1287_cse ) begin
      mut_7_8_63_0 <= mut_7_7_63_0;
      mut_6_8_63_0 <= mut_6_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1289_cse ) begin
      mut_9_8_63_0 <= mut_9_7_63_0;
      mut_8_8_63_0 <= mut_8_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1291_cse ) begin
      mut_11_8_63_0 <= mut_11_7_63_0;
      mut_10_8_63_0 <= mut_10_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1293_cse ) begin
      mut_13_8_63_0 <= mut_13_7_63_0;
      mut_12_8_63_0 <= mut_12_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1295_cse ) begin
      mut_15_8_63_0 <= mut_15_7_63_0;
      mut_14_8_63_0 <= mut_14_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1297_cse ) begin
      mut_17_8_63_0 <= mut_17_7_63_0;
      mut_16_8_63_0 <= mut_16_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1299_cse ) begin
      mut_19_8_63_0 <= mut_19_7_63_0;
      mut_18_8_63_0 <= mut_18_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1301_cse ) begin
      mut_21_8_63_0 <= mut_21_7_63_0;
      mut_20_8_63_0 <= mut_20_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1303_cse ) begin
      mut_23_8_63_0 <= mut_23_7_63_0;
      mut_22_8_63_0 <= mut_22_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1305_cse ) begin
      mut_1_8_63_0 <= mut_1_7_63_0;
      mut_8_63_0 <= mut_7_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_8_3_2 <= 2'b00;
      rem_12cyc_st_8_1_0 <= 2'b00;
    end
    else if ( and_1307_cse ) begin
      rem_12cyc_st_8_3_2 <= rem_12cyc_st_7_3_2;
      rem_12cyc_st_8_1_0 <= rem_12cyc_st_7_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1309_cse ) begin
      mut_3_7_63_0 <= mut_3_6_63_0;
      mut_2_7_63_0 <= mut_2_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1311_cse ) begin
      mut_5_7_63_0 <= mut_5_6_63_0;
      mut_4_7_63_0 <= mut_4_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1313_cse ) begin
      mut_7_7_63_0 <= mut_7_6_63_0;
      mut_6_7_63_0 <= mut_6_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1315_cse ) begin
      mut_9_7_63_0 <= mut_9_6_63_0;
      mut_8_7_63_0 <= mut_8_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1317_cse ) begin
      mut_11_7_63_0 <= mut_11_6_63_0;
      mut_10_7_63_0 <= mut_10_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1319_cse ) begin
      mut_13_7_63_0 <= mut_13_6_63_0;
      mut_12_7_63_0 <= mut_12_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1321_cse ) begin
      mut_15_7_63_0 <= mut_15_6_63_0;
      mut_14_7_63_0 <= mut_14_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1323_cse ) begin
      mut_17_7_63_0 <= mut_17_6_63_0;
      mut_16_7_63_0 <= mut_16_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1325_cse ) begin
      mut_19_7_63_0 <= mut_19_6_63_0;
      mut_18_7_63_0 <= mut_18_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1327_cse ) begin
      mut_21_7_63_0 <= mut_21_6_63_0;
      mut_20_7_63_0 <= mut_20_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1329_cse ) begin
      mut_23_7_63_0 <= mut_23_6_63_0;
      mut_22_7_63_0 <= mut_22_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1331_cse ) begin
      mut_1_7_63_0 <= mut_1_6_63_0;
      mut_7_63_0 <= mut_6_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_7_3_2 <= 2'b00;
      rem_12cyc_st_7_1_0 <= 2'b00;
    end
    else if ( and_1333_cse ) begin
      rem_12cyc_st_7_3_2 <= rem_12cyc_st_6_3_2;
      rem_12cyc_st_7_1_0 <= rem_12cyc_st_6_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1335_cse ) begin
      mut_3_6_63_0 <= mut_3_5_63_0;
      mut_2_6_63_0 <= mut_2_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1337_cse ) begin
      mut_5_6_63_0 <= mut_5_5_63_0;
      mut_4_6_63_0 <= mut_4_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1339_cse ) begin
      mut_7_6_63_0 <= mut_7_5_63_0;
      mut_6_6_63_0 <= mut_6_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1341_cse ) begin
      mut_9_6_63_0 <= mut_9_5_63_0;
      mut_8_6_63_0 <= mut_8_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1343_cse ) begin
      mut_11_6_63_0 <= mut_11_5_63_0;
      mut_10_6_63_0 <= mut_10_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1345_cse ) begin
      mut_13_6_63_0 <= mut_13_5_63_0;
      mut_12_6_63_0 <= mut_12_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1347_cse ) begin
      mut_15_6_63_0 <= mut_15_5_63_0;
      mut_14_6_63_0 <= mut_14_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1349_cse ) begin
      mut_17_6_63_0 <= mut_17_5_63_0;
      mut_16_6_63_0 <= mut_16_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1351_cse ) begin
      mut_19_6_63_0 <= mut_19_5_63_0;
      mut_18_6_63_0 <= mut_18_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1353_cse ) begin
      mut_21_6_63_0 <= mut_21_5_63_0;
      mut_20_6_63_0 <= mut_20_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1355_cse ) begin
      mut_23_6_63_0 <= mut_23_5_63_0;
      mut_22_6_63_0 <= mut_22_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1357_cse ) begin
      mut_1_6_63_0 <= mut_1_5_63_0;
      mut_6_63_0 <= mut_5_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1359_cse ) begin
      m_buf_sva_6 <= m_buf_sva_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_6_3_2 <= 2'b00;
      rem_12cyc_st_6_1_0 <= 2'b00;
    end
    else if ( and_1359_cse ) begin
      rem_12cyc_st_6_3_2 <= rem_12cyc_st_5_3_2;
      rem_12cyc_st_6_1_0 <= rem_12cyc_st_5_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1361_cse ) begin
      mut_3_5_63_0 <= mut_3_4_63_0;
      mut_2_5_63_0 <= mut_2_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1363_cse ) begin
      mut_5_5_63_0 <= mut_5_4_63_0;
      mut_4_5_63_0 <= mut_4_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1365_cse ) begin
      mut_7_5_63_0 <= mut_7_4_63_0;
      mut_6_5_63_0 <= mut_6_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1367_cse ) begin
      mut_9_5_63_0 <= mut_9_4_63_0;
      mut_8_5_63_0 <= mut_8_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1369_cse ) begin
      mut_11_5_63_0 <= mut_11_4_63_0;
      mut_10_5_63_0 <= mut_10_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1371_cse ) begin
      mut_13_5_63_0 <= mut_13_4_63_0;
      mut_12_5_63_0 <= mut_12_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1373_cse ) begin
      mut_15_5_63_0 <= mut_15_4_63_0;
      mut_14_5_63_0 <= mut_14_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1375_cse ) begin
      mut_17_5_63_0 <= mut_17_4_63_0;
      mut_16_5_63_0 <= mut_16_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1377_cse ) begin
      mut_19_5_63_0 <= mut_19_4_63_0;
      mut_18_5_63_0 <= mut_18_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1379_cse ) begin
      mut_21_5_63_0 <= mut_21_4_63_0;
      mut_20_5_63_0 <= mut_20_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1381_cse ) begin
      mut_23_5_63_0 <= mut_23_4_63_0;
      mut_22_5_63_0 <= mut_22_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1383_cse ) begin
      mut_1_5_63_0 <= mut_1_4_63_0;
      mut_5_63_0 <= mut_4_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1385_cse ) begin
      m_buf_sva_5 <= m_buf_sva_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_5_3_2 <= 2'b00;
      rem_12cyc_st_5_1_0 <= 2'b00;
    end
    else if ( and_1385_cse ) begin
      rem_12cyc_st_5_3_2 <= rem_12cyc_st_4_3_2;
      rem_12cyc_st_5_1_0 <= rem_12cyc_st_4_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1387_cse ) begin
      mut_3_4_63_0 <= mut_3_3_63_0;
      mut_2_4_63_0 <= mut_2_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1389_cse ) begin
      mut_5_4_63_0 <= mut_5_3_63_0;
      mut_4_4_63_0 <= mut_4_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1391_cse ) begin
      mut_7_4_63_0 <= mut_7_3_63_0;
      mut_6_4_63_0 <= mut_6_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1393_cse ) begin
      mut_9_4_63_0 <= mut_9_3_63_0;
      mut_8_4_63_0 <= mut_8_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1395_cse ) begin
      mut_11_4_63_0 <= mut_11_3_63_0;
      mut_10_4_63_0 <= mut_10_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1397_cse ) begin
      mut_13_4_63_0 <= mut_13_3_63_0;
      mut_12_4_63_0 <= mut_12_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1399_cse ) begin
      mut_15_4_63_0 <= mut_15_3_63_0;
      mut_14_4_63_0 <= mut_14_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1401_cse ) begin
      mut_17_4_63_0 <= mut_17_3_63_0;
      mut_16_4_63_0 <= mut_16_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1403_cse ) begin
      mut_19_4_63_0 <= mut_19_3_63_0;
      mut_18_4_63_0 <= mut_18_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1405_cse ) begin
      mut_21_4_63_0 <= mut_21_3_63_0;
      mut_20_4_63_0 <= mut_20_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1407_cse ) begin
      mut_23_4_63_0 <= mut_23_3_63_0;
      mut_22_4_63_0 <= mut_22_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1409_cse ) begin
      mut_1_4_63_0 <= mut_1_3_63_0;
      mut_4_63_0 <= mut_3_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1411_cse ) begin
      m_buf_sva_4 <= m_buf_sva_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_4_3_2 <= 2'b00;
      rem_12cyc_st_4_1_0 <= 2'b00;
    end
    else if ( and_1411_cse ) begin
      rem_12cyc_st_4_3_2 <= rem_12cyc_st_3_3_2;
      rem_12cyc_st_4_1_0 <= rem_12cyc_st_3_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1413_cse ) begin
      mut_3_3_63_0 <= mut_3_2_63_0;
      mut_2_3_63_0 <= mut_2_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1415_cse ) begin
      mut_5_3_63_0 <= mut_5_2_63_0;
      mut_4_3_63_0 <= mut_4_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1417_cse ) begin
      mut_7_3_63_0 <= mut_7_2_63_0;
      mut_6_3_63_0 <= mut_6_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1419_cse ) begin
      mut_9_3_63_0 <= mut_9_2_63_0;
      mut_8_3_63_0 <= mut_8_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1421_cse ) begin
      mut_11_3_63_0 <= mut_11_2_63_0;
      mut_10_3_63_0 <= mut_10_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1423_cse ) begin
      mut_13_3_63_0 <= mut_13_2_63_0;
      mut_12_3_63_0 <= mut_12_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1425_cse ) begin
      mut_15_3_63_0 <= mut_15_2_63_0;
      mut_14_3_63_0 <= mut_14_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1427_cse ) begin
      mut_17_3_63_0 <= mut_17_2_63_0;
      mut_16_3_63_0 <= mut_16_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1429_cse ) begin
      mut_19_3_63_0 <= mut_19_2_63_0;
      mut_18_3_63_0 <= mut_18_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1431_cse ) begin
      mut_21_3_63_0 <= mut_21_2_63_0;
      mut_20_3_63_0 <= mut_20_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1433_cse ) begin
      mut_23_3_63_0 <= mut_23_2_63_0;
      mut_22_3_63_0 <= mut_22_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1435_cse ) begin
      mut_1_3_63_0 <= mut_1_2_63_0;
      mut_3_63_0 <= mut_2_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1437_cse ) begin
      m_buf_sva_3 <= m_buf_sva_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_3_3_2 <= 2'b00;
      rem_12cyc_st_3_1_0 <= 2'b00;
    end
    else if ( and_1437_cse ) begin
      rem_12cyc_st_3_3_2 <= rem_12cyc_st_2_3_2;
      rem_12cyc_st_3_1_0 <= rem_12cyc_st_2_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1439_cse ) begin
      mut_3_2_63_0 <= rem_13_cmp_1_b_63_0;
      mut_2_2_63_0 <= rem_13_cmp_1_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1441_cse ) begin
      mut_5_2_63_0 <= rem_13_cmp_2_b_63_0;
      mut_4_2_63_0 <= rem_13_cmp_2_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1443_cse ) begin
      mut_7_2_63_0 <= rem_13_cmp_3_b_63_0;
      mut_6_2_63_0 <= rem_13_cmp_3_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1445_cse ) begin
      mut_9_2_63_0 <= rem_13_cmp_4_b_63_0;
      mut_8_2_63_0 <= rem_13_cmp_4_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1447_cse ) begin
      mut_11_2_63_0 <= rem_13_cmp_5_b_63_0;
      mut_10_2_63_0 <= rem_13_cmp_5_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1449_cse ) begin
      mut_13_2_63_0 <= rem_13_cmp_6_b_63_0;
      mut_12_2_63_0 <= rem_13_cmp_6_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1451_cse ) begin
      mut_15_2_63_0 <= rem_13_cmp_7_b_63_0;
      mut_14_2_63_0 <= rem_13_cmp_7_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1453_cse ) begin
      mut_17_2_63_0 <= rem_13_cmp_8_b_63_0;
      mut_16_2_63_0 <= rem_13_cmp_8_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1455_cse ) begin
      mut_19_2_63_0 <= rem_13_cmp_9_b_63_0;
      mut_18_2_63_0 <= rem_13_cmp_9_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1457_cse ) begin
      mut_21_2_63_0 <= rem_13_cmp_10_b_63_0;
      mut_20_2_63_0 <= rem_13_cmp_10_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1459_cse ) begin
      mut_23_2_63_0 <= rem_13_cmp_11_b_63_0;
      mut_22_2_63_0 <= rem_13_cmp_11_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1461_cse ) begin
      mut_1_2_63_0 <= rem_13_cmp_b_63_0;
      mut_2_63_0 <= rem_13_cmp_a_63_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1463_cse ) begin
      m_buf_sva_2 <= m_buf_sva_1;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_st_2_3_2 <= 2'b00;
      rem_12cyc_st_2_1_0 <= 2'b00;
    end
    else if ( and_1463_cse ) begin
      rem_12cyc_st_2_3_2 <= rem_12cyc_3_2;
      rem_12cyc_st_2_1_0 <= rem_12cyc_1_0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( and_1197_cse ) begin
      m_buf_sva_1 <= m_rsci_idat;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_12cyc_3_2 <= 2'b00;
      rem_12cyc_1_0 <= 2'b00;
    end
    else if ( and_1197_cse ) begin
      rem_12cyc_3_2 <= acc_tmp;
      rem_12cyc_1_0 <= acc_1_tmp[1:0];
    end
  end
  assign nl_qelse_acc_nl = result_sva_duc_mx0 + m_buf_sva_12;
  assign qelse_acc_nl = nl_qelse_acc_nl[63:0];
  assign mux_10_nl = MUX_s_1_2_2((rem_13_cmp_1_z[63]), (rem_13_cmp_3_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_9_nl = MUX_s_1_2_2((rem_13_cmp_2_z[63]), (rem_13_cmp_4_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_11_nl = MUX_s_1_2_2(mux_10_nl, mux_9_nl, rem_12cyc_st_12_1_0[0]);
  assign mux_7_nl = MUX_s_1_2_2((rem_13_cmp_9_z[63]), (rem_13_cmp_11_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_6_nl = MUX_s_1_2_2((rem_13_cmp_10_z[63]), (rem_13_cmp_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_8_nl = MUX_s_1_2_2(mux_7_nl, mux_6_nl, rem_12cyc_st_12_1_0[0]);
  assign mux_12_nl = MUX_s_1_2_2(mux_11_nl, mux_8_nl, rem_12cyc_st_12_3_2[1]);
  assign mux_3_nl = MUX_s_1_2_2((rem_13_cmp_5_z[63]), (rem_13_cmp_7_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_2_nl = MUX_s_1_2_2((rem_13_cmp_6_z[63]), (rem_13_cmp_8_z[63]), rem_12cyc_st_12_1_0[1]);
  assign mux_4_nl = MUX_s_1_2_2(mux_3_nl, mux_2_nl, rem_12cyc_st_12_1_0[0]);
  assign mux_5_nl = MUX_s_1_2_2(mux_4_nl, (result_sva_duc[63]), rem_12cyc_st_12_3_2[1]);
  assign mux_13_nl = MUX_s_1_2_2(mux_12_nl, mux_5_nl, rem_12cyc_st_12_3_2[0]);

  function automatic [63:0] MUX1HOT_v_64_11_2;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [10:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    MUX1HOT_v_64_11_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_13_2;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [12:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    MUX1HOT_v_64_13_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    modulo_dev
// ------------------------------------------------------------------


module modulo_dev (
  base_rsc_dat, m_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [63:0] base_rsc_dat;
  input [63:0] m_rsc_dat;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  modulo_dev_core modulo_dev_core_inst (
      .base_rsc_dat(base_rsc_dat),
      .m_rsc_dat(m_rsc_dat),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.v 
module mgc_div(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_a-1:0] z;  
   reg  [width_a-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  div_s(a,b,z);
	else
          div_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Thu Aug  5 01:56:25 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_6_64_64_64_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_6_64_64_64_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [5:0] radr;
  output we;
  output [63:0] d;
  output [5:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [5:0] radr_d;
  input [5:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core_core_fsm (
  clk, rst, fsm_output, STAGE_LOOP_C_3_tr0, modExp_dev_while_C_14_tr0, COMP_LOOP_C_1_tr0,
      COMP_LOOP_1_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_32_tr0, COMP_LOOP_2_modExp_dev_1_while_C_14_tr0,
      COMP_LOOP_C_64_tr0, COMP_LOOP_3_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_96_tr0,
      COMP_LOOP_4_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_128_tr0, COMP_LOOP_5_modExp_dev_1_while_C_14_tr0,
      COMP_LOOP_C_160_tr0, COMP_LOOP_6_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_192_tr0,
      COMP_LOOP_7_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_224_tr0, COMP_LOOP_8_modExp_dev_1_while_C_14_tr0,
      COMP_LOOP_C_256_tr0, COMP_LOOP_9_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_288_tr0,
      COMP_LOOP_10_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_320_tr0, COMP_LOOP_11_modExp_dev_1_while_C_14_tr0,
      COMP_LOOP_C_352_tr0, COMP_LOOP_12_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_384_tr0,
      COMP_LOOP_13_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_416_tr0, COMP_LOOP_14_modExp_dev_1_while_C_14_tr0,
      COMP_LOOP_C_448_tr0, COMP_LOOP_15_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_480_tr0,
      COMP_LOOP_16_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_512_tr0, VEC_LOOP_C_0_tr0,
      STAGE_LOOP_C_4_tr0
);
  input clk;
  input rst;
  output [9:0] fsm_output;
  reg [9:0] fsm_output;
  input STAGE_LOOP_C_3_tr0;
  input modExp_dev_while_C_14_tr0;
  input COMP_LOOP_C_1_tr0;
  input COMP_LOOP_1_modExp_dev_1_while_C_14_tr0;
  input COMP_LOOP_C_32_tr0;
  input COMP_LOOP_2_modExp_dev_1_while_C_14_tr0;
  input COMP_LOOP_C_64_tr0;
  input COMP_LOOP_3_modExp_dev_1_while_C_14_tr0;
  input COMP_LOOP_C_96_tr0;
  input COMP_LOOP_4_modExp_dev_1_while_C_14_tr0;
  input COMP_LOOP_C_128_tr0;
  input COMP_LOOP_5_modExp_dev_1_while_C_14_tr0;
  input COMP_LOOP_C_160_tr0;
  input COMP_LOOP_6_modExp_dev_1_while_C_14_tr0;
  input COMP_LOOP_C_192_tr0;
  input COMP_LOOP_7_modExp_dev_1_while_C_14_tr0;
  input COMP_LOOP_C_224_tr0;
  input COMP_LOOP_8_modExp_dev_1_while_C_14_tr0;
  input COMP_LOOP_C_256_tr0;
  input COMP_LOOP_9_modExp_dev_1_while_C_14_tr0;
  input COMP_LOOP_C_288_tr0;
  input COMP_LOOP_10_modExp_dev_1_while_C_14_tr0;
  input COMP_LOOP_C_320_tr0;
  input COMP_LOOP_11_modExp_dev_1_while_C_14_tr0;
  input COMP_LOOP_C_352_tr0;
  input COMP_LOOP_12_modExp_dev_1_while_C_14_tr0;
  input COMP_LOOP_C_384_tr0;
  input COMP_LOOP_13_modExp_dev_1_while_C_14_tr0;
  input COMP_LOOP_C_416_tr0;
  input COMP_LOOP_14_modExp_dev_1_while_C_14_tr0;
  input COMP_LOOP_C_448_tr0;
  input COMP_LOOP_15_modExp_dev_1_while_C_14_tr0;
  input COMP_LOOP_C_480_tr0;
  input COMP_LOOP_16_modExp_dev_1_while_C_14_tr0;
  input COMP_LOOP_C_512_tr0;
  input VEC_LOOP_C_0_tr0;
  input STAGE_LOOP_C_4_tr0;


  // FSM State Type Declaration for inPlaceNTT_DIT_core_core_fsm_1
  parameter
    main_C_0 = 10'd0,
    STAGE_LOOP_C_0 = 10'd1,
    STAGE_LOOP_C_1 = 10'd2,
    STAGE_LOOP_C_2 = 10'd3,
    STAGE_LOOP_C_3 = 10'd4,
    modExp_dev_while_C_0 = 10'd5,
    modExp_dev_while_C_1 = 10'd6,
    modExp_dev_while_C_2 = 10'd7,
    modExp_dev_while_C_3 = 10'd8,
    modExp_dev_while_C_4 = 10'd9,
    modExp_dev_while_C_5 = 10'd10,
    modExp_dev_while_C_6 = 10'd11,
    modExp_dev_while_C_7 = 10'd12,
    modExp_dev_while_C_8 = 10'd13,
    modExp_dev_while_C_9 = 10'd14,
    modExp_dev_while_C_10 = 10'd15,
    modExp_dev_while_C_11 = 10'd16,
    modExp_dev_while_C_12 = 10'd17,
    modExp_dev_while_C_13 = 10'd18,
    modExp_dev_while_C_14 = 10'd19,
    COMP_LOOP_C_0 = 10'd20,
    COMP_LOOP_C_1 = 10'd21,
    COMP_LOOP_1_modExp_dev_1_while_C_0 = 10'd22,
    COMP_LOOP_1_modExp_dev_1_while_C_1 = 10'd23,
    COMP_LOOP_1_modExp_dev_1_while_C_2 = 10'd24,
    COMP_LOOP_1_modExp_dev_1_while_C_3 = 10'd25,
    COMP_LOOP_1_modExp_dev_1_while_C_4 = 10'd26,
    COMP_LOOP_1_modExp_dev_1_while_C_5 = 10'd27,
    COMP_LOOP_1_modExp_dev_1_while_C_6 = 10'd28,
    COMP_LOOP_1_modExp_dev_1_while_C_7 = 10'd29,
    COMP_LOOP_1_modExp_dev_1_while_C_8 = 10'd30,
    COMP_LOOP_1_modExp_dev_1_while_C_9 = 10'd31,
    COMP_LOOP_1_modExp_dev_1_while_C_10 = 10'd32,
    COMP_LOOP_1_modExp_dev_1_while_C_11 = 10'd33,
    COMP_LOOP_1_modExp_dev_1_while_C_12 = 10'd34,
    COMP_LOOP_1_modExp_dev_1_while_C_13 = 10'd35,
    COMP_LOOP_1_modExp_dev_1_while_C_14 = 10'd36,
    COMP_LOOP_C_2 = 10'd37,
    COMP_LOOP_C_3 = 10'd38,
    COMP_LOOP_C_4 = 10'd39,
    COMP_LOOP_C_5 = 10'd40,
    COMP_LOOP_C_6 = 10'd41,
    COMP_LOOP_C_7 = 10'd42,
    COMP_LOOP_C_8 = 10'd43,
    COMP_LOOP_C_9 = 10'd44,
    COMP_LOOP_C_10 = 10'd45,
    COMP_LOOP_C_11 = 10'd46,
    COMP_LOOP_C_12 = 10'd47,
    COMP_LOOP_C_13 = 10'd48,
    COMP_LOOP_C_14 = 10'd49,
    COMP_LOOP_C_15 = 10'd50,
    COMP_LOOP_C_16 = 10'd51,
    COMP_LOOP_C_17 = 10'd52,
    COMP_LOOP_C_18 = 10'd53,
    COMP_LOOP_C_19 = 10'd54,
    COMP_LOOP_C_20 = 10'd55,
    COMP_LOOP_C_21 = 10'd56,
    COMP_LOOP_C_22 = 10'd57,
    COMP_LOOP_C_23 = 10'd58,
    COMP_LOOP_C_24 = 10'd59,
    COMP_LOOP_C_25 = 10'd60,
    COMP_LOOP_C_26 = 10'd61,
    COMP_LOOP_C_27 = 10'd62,
    COMP_LOOP_C_28 = 10'd63,
    COMP_LOOP_C_29 = 10'd64,
    COMP_LOOP_C_30 = 10'd65,
    COMP_LOOP_C_31 = 10'd66,
    COMP_LOOP_C_32 = 10'd67,
    COMP_LOOP_C_33 = 10'd68,
    COMP_LOOP_2_modExp_dev_1_while_C_0 = 10'd69,
    COMP_LOOP_2_modExp_dev_1_while_C_1 = 10'd70,
    COMP_LOOP_2_modExp_dev_1_while_C_2 = 10'd71,
    COMP_LOOP_2_modExp_dev_1_while_C_3 = 10'd72,
    COMP_LOOP_2_modExp_dev_1_while_C_4 = 10'd73,
    COMP_LOOP_2_modExp_dev_1_while_C_5 = 10'd74,
    COMP_LOOP_2_modExp_dev_1_while_C_6 = 10'd75,
    COMP_LOOP_2_modExp_dev_1_while_C_7 = 10'd76,
    COMP_LOOP_2_modExp_dev_1_while_C_8 = 10'd77,
    COMP_LOOP_2_modExp_dev_1_while_C_9 = 10'd78,
    COMP_LOOP_2_modExp_dev_1_while_C_10 = 10'd79,
    COMP_LOOP_2_modExp_dev_1_while_C_11 = 10'd80,
    COMP_LOOP_2_modExp_dev_1_while_C_12 = 10'd81,
    COMP_LOOP_2_modExp_dev_1_while_C_13 = 10'd82,
    COMP_LOOP_2_modExp_dev_1_while_C_14 = 10'd83,
    COMP_LOOP_C_34 = 10'd84,
    COMP_LOOP_C_35 = 10'd85,
    COMP_LOOP_C_36 = 10'd86,
    COMP_LOOP_C_37 = 10'd87,
    COMP_LOOP_C_38 = 10'd88,
    COMP_LOOP_C_39 = 10'd89,
    COMP_LOOP_C_40 = 10'd90,
    COMP_LOOP_C_41 = 10'd91,
    COMP_LOOP_C_42 = 10'd92,
    COMP_LOOP_C_43 = 10'd93,
    COMP_LOOP_C_44 = 10'd94,
    COMP_LOOP_C_45 = 10'd95,
    COMP_LOOP_C_46 = 10'd96,
    COMP_LOOP_C_47 = 10'd97,
    COMP_LOOP_C_48 = 10'd98,
    COMP_LOOP_C_49 = 10'd99,
    COMP_LOOP_C_50 = 10'd100,
    COMP_LOOP_C_51 = 10'd101,
    COMP_LOOP_C_52 = 10'd102,
    COMP_LOOP_C_53 = 10'd103,
    COMP_LOOP_C_54 = 10'd104,
    COMP_LOOP_C_55 = 10'd105,
    COMP_LOOP_C_56 = 10'd106,
    COMP_LOOP_C_57 = 10'd107,
    COMP_LOOP_C_58 = 10'd108,
    COMP_LOOP_C_59 = 10'd109,
    COMP_LOOP_C_60 = 10'd110,
    COMP_LOOP_C_61 = 10'd111,
    COMP_LOOP_C_62 = 10'd112,
    COMP_LOOP_C_63 = 10'd113,
    COMP_LOOP_C_64 = 10'd114,
    COMP_LOOP_C_65 = 10'd115,
    COMP_LOOP_3_modExp_dev_1_while_C_0 = 10'd116,
    COMP_LOOP_3_modExp_dev_1_while_C_1 = 10'd117,
    COMP_LOOP_3_modExp_dev_1_while_C_2 = 10'd118,
    COMP_LOOP_3_modExp_dev_1_while_C_3 = 10'd119,
    COMP_LOOP_3_modExp_dev_1_while_C_4 = 10'd120,
    COMP_LOOP_3_modExp_dev_1_while_C_5 = 10'd121,
    COMP_LOOP_3_modExp_dev_1_while_C_6 = 10'd122,
    COMP_LOOP_3_modExp_dev_1_while_C_7 = 10'd123,
    COMP_LOOP_3_modExp_dev_1_while_C_8 = 10'd124,
    COMP_LOOP_3_modExp_dev_1_while_C_9 = 10'd125,
    COMP_LOOP_3_modExp_dev_1_while_C_10 = 10'd126,
    COMP_LOOP_3_modExp_dev_1_while_C_11 = 10'd127,
    COMP_LOOP_3_modExp_dev_1_while_C_12 = 10'd128,
    COMP_LOOP_3_modExp_dev_1_while_C_13 = 10'd129,
    COMP_LOOP_3_modExp_dev_1_while_C_14 = 10'd130,
    COMP_LOOP_C_66 = 10'd131,
    COMP_LOOP_C_67 = 10'd132,
    COMP_LOOP_C_68 = 10'd133,
    COMP_LOOP_C_69 = 10'd134,
    COMP_LOOP_C_70 = 10'd135,
    COMP_LOOP_C_71 = 10'd136,
    COMP_LOOP_C_72 = 10'd137,
    COMP_LOOP_C_73 = 10'd138,
    COMP_LOOP_C_74 = 10'd139,
    COMP_LOOP_C_75 = 10'd140,
    COMP_LOOP_C_76 = 10'd141,
    COMP_LOOP_C_77 = 10'd142,
    COMP_LOOP_C_78 = 10'd143,
    COMP_LOOP_C_79 = 10'd144,
    COMP_LOOP_C_80 = 10'd145,
    COMP_LOOP_C_81 = 10'd146,
    COMP_LOOP_C_82 = 10'd147,
    COMP_LOOP_C_83 = 10'd148,
    COMP_LOOP_C_84 = 10'd149,
    COMP_LOOP_C_85 = 10'd150,
    COMP_LOOP_C_86 = 10'd151,
    COMP_LOOP_C_87 = 10'd152,
    COMP_LOOP_C_88 = 10'd153,
    COMP_LOOP_C_89 = 10'd154,
    COMP_LOOP_C_90 = 10'd155,
    COMP_LOOP_C_91 = 10'd156,
    COMP_LOOP_C_92 = 10'd157,
    COMP_LOOP_C_93 = 10'd158,
    COMP_LOOP_C_94 = 10'd159,
    COMP_LOOP_C_95 = 10'd160,
    COMP_LOOP_C_96 = 10'd161,
    COMP_LOOP_C_97 = 10'd162,
    COMP_LOOP_4_modExp_dev_1_while_C_0 = 10'd163,
    COMP_LOOP_4_modExp_dev_1_while_C_1 = 10'd164,
    COMP_LOOP_4_modExp_dev_1_while_C_2 = 10'd165,
    COMP_LOOP_4_modExp_dev_1_while_C_3 = 10'd166,
    COMP_LOOP_4_modExp_dev_1_while_C_4 = 10'd167,
    COMP_LOOP_4_modExp_dev_1_while_C_5 = 10'd168,
    COMP_LOOP_4_modExp_dev_1_while_C_6 = 10'd169,
    COMP_LOOP_4_modExp_dev_1_while_C_7 = 10'd170,
    COMP_LOOP_4_modExp_dev_1_while_C_8 = 10'd171,
    COMP_LOOP_4_modExp_dev_1_while_C_9 = 10'd172,
    COMP_LOOP_4_modExp_dev_1_while_C_10 = 10'd173,
    COMP_LOOP_4_modExp_dev_1_while_C_11 = 10'd174,
    COMP_LOOP_4_modExp_dev_1_while_C_12 = 10'd175,
    COMP_LOOP_4_modExp_dev_1_while_C_13 = 10'd176,
    COMP_LOOP_4_modExp_dev_1_while_C_14 = 10'd177,
    COMP_LOOP_C_98 = 10'd178,
    COMP_LOOP_C_99 = 10'd179,
    COMP_LOOP_C_100 = 10'd180,
    COMP_LOOP_C_101 = 10'd181,
    COMP_LOOP_C_102 = 10'd182,
    COMP_LOOP_C_103 = 10'd183,
    COMP_LOOP_C_104 = 10'd184,
    COMP_LOOP_C_105 = 10'd185,
    COMP_LOOP_C_106 = 10'd186,
    COMP_LOOP_C_107 = 10'd187,
    COMP_LOOP_C_108 = 10'd188,
    COMP_LOOP_C_109 = 10'd189,
    COMP_LOOP_C_110 = 10'd190,
    COMP_LOOP_C_111 = 10'd191,
    COMP_LOOP_C_112 = 10'd192,
    COMP_LOOP_C_113 = 10'd193,
    COMP_LOOP_C_114 = 10'd194,
    COMP_LOOP_C_115 = 10'd195,
    COMP_LOOP_C_116 = 10'd196,
    COMP_LOOP_C_117 = 10'd197,
    COMP_LOOP_C_118 = 10'd198,
    COMP_LOOP_C_119 = 10'd199,
    COMP_LOOP_C_120 = 10'd200,
    COMP_LOOP_C_121 = 10'd201,
    COMP_LOOP_C_122 = 10'd202,
    COMP_LOOP_C_123 = 10'd203,
    COMP_LOOP_C_124 = 10'd204,
    COMP_LOOP_C_125 = 10'd205,
    COMP_LOOP_C_126 = 10'd206,
    COMP_LOOP_C_127 = 10'd207,
    COMP_LOOP_C_128 = 10'd208,
    COMP_LOOP_C_129 = 10'd209,
    COMP_LOOP_5_modExp_dev_1_while_C_0 = 10'd210,
    COMP_LOOP_5_modExp_dev_1_while_C_1 = 10'd211,
    COMP_LOOP_5_modExp_dev_1_while_C_2 = 10'd212,
    COMP_LOOP_5_modExp_dev_1_while_C_3 = 10'd213,
    COMP_LOOP_5_modExp_dev_1_while_C_4 = 10'd214,
    COMP_LOOP_5_modExp_dev_1_while_C_5 = 10'd215,
    COMP_LOOP_5_modExp_dev_1_while_C_6 = 10'd216,
    COMP_LOOP_5_modExp_dev_1_while_C_7 = 10'd217,
    COMP_LOOP_5_modExp_dev_1_while_C_8 = 10'd218,
    COMP_LOOP_5_modExp_dev_1_while_C_9 = 10'd219,
    COMP_LOOP_5_modExp_dev_1_while_C_10 = 10'd220,
    COMP_LOOP_5_modExp_dev_1_while_C_11 = 10'd221,
    COMP_LOOP_5_modExp_dev_1_while_C_12 = 10'd222,
    COMP_LOOP_5_modExp_dev_1_while_C_13 = 10'd223,
    COMP_LOOP_5_modExp_dev_1_while_C_14 = 10'd224,
    COMP_LOOP_C_130 = 10'd225,
    COMP_LOOP_C_131 = 10'd226,
    COMP_LOOP_C_132 = 10'd227,
    COMP_LOOP_C_133 = 10'd228,
    COMP_LOOP_C_134 = 10'd229,
    COMP_LOOP_C_135 = 10'd230,
    COMP_LOOP_C_136 = 10'd231,
    COMP_LOOP_C_137 = 10'd232,
    COMP_LOOP_C_138 = 10'd233,
    COMP_LOOP_C_139 = 10'd234,
    COMP_LOOP_C_140 = 10'd235,
    COMP_LOOP_C_141 = 10'd236,
    COMP_LOOP_C_142 = 10'd237,
    COMP_LOOP_C_143 = 10'd238,
    COMP_LOOP_C_144 = 10'd239,
    COMP_LOOP_C_145 = 10'd240,
    COMP_LOOP_C_146 = 10'd241,
    COMP_LOOP_C_147 = 10'd242,
    COMP_LOOP_C_148 = 10'd243,
    COMP_LOOP_C_149 = 10'd244,
    COMP_LOOP_C_150 = 10'd245,
    COMP_LOOP_C_151 = 10'd246,
    COMP_LOOP_C_152 = 10'd247,
    COMP_LOOP_C_153 = 10'd248,
    COMP_LOOP_C_154 = 10'd249,
    COMP_LOOP_C_155 = 10'd250,
    COMP_LOOP_C_156 = 10'd251,
    COMP_LOOP_C_157 = 10'd252,
    COMP_LOOP_C_158 = 10'd253,
    COMP_LOOP_C_159 = 10'd254,
    COMP_LOOP_C_160 = 10'd255,
    COMP_LOOP_C_161 = 10'd256,
    COMP_LOOP_6_modExp_dev_1_while_C_0 = 10'd257,
    COMP_LOOP_6_modExp_dev_1_while_C_1 = 10'd258,
    COMP_LOOP_6_modExp_dev_1_while_C_2 = 10'd259,
    COMP_LOOP_6_modExp_dev_1_while_C_3 = 10'd260,
    COMP_LOOP_6_modExp_dev_1_while_C_4 = 10'd261,
    COMP_LOOP_6_modExp_dev_1_while_C_5 = 10'd262,
    COMP_LOOP_6_modExp_dev_1_while_C_6 = 10'd263,
    COMP_LOOP_6_modExp_dev_1_while_C_7 = 10'd264,
    COMP_LOOP_6_modExp_dev_1_while_C_8 = 10'd265,
    COMP_LOOP_6_modExp_dev_1_while_C_9 = 10'd266,
    COMP_LOOP_6_modExp_dev_1_while_C_10 = 10'd267,
    COMP_LOOP_6_modExp_dev_1_while_C_11 = 10'd268,
    COMP_LOOP_6_modExp_dev_1_while_C_12 = 10'd269,
    COMP_LOOP_6_modExp_dev_1_while_C_13 = 10'd270,
    COMP_LOOP_6_modExp_dev_1_while_C_14 = 10'd271,
    COMP_LOOP_C_162 = 10'd272,
    COMP_LOOP_C_163 = 10'd273,
    COMP_LOOP_C_164 = 10'd274,
    COMP_LOOP_C_165 = 10'd275,
    COMP_LOOP_C_166 = 10'd276,
    COMP_LOOP_C_167 = 10'd277,
    COMP_LOOP_C_168 = 10'd278,
    COMP_LOOP_C_169 = 10'd279,
    COMP_LOOP_C_170 = 10'd280,
    COMP_LOOP_C_171 = 10'd281,
    COMP_LOOP_C_172 = 10'd282,
    COMP_LOOP_C_173 = 10'd283,
    COMP_LOOP_C_174 = 10'd284,
    COMP_LOOP_C_175 = 10'd285,
    COMP_LOOP_C_176 = 10'd286,
    COMP_LOOP_C_177 = 10'd287,
    COMP_LOOP_C_178 = 10'd288,
    COMP_LOOP_C_179 = 10'd289,
    COMP_LOOP_C_180 = 10'd290,
    COMP_LOOP_C_181 = 10'd291,
    COMP_LOOP_C_182 = 10'd292,
    COMP_LOOP_C_183 = 10'd293,
    COMP_LOOP_C_184 = 10'd294,
    COMP_LOOP_C_185 = 10'd295,
    COMP_LOOP_C_186 = 10'd296,
    COMP_LOOP_C_187 = 10'd297,
    COMP_LOOP_C_188 = 10'd298,
    COMP_LOOP_C_189 = 10'd299,
    COMP_LOOP_C_190 = 10'd300,
    COMP_LOOP_C_191 = 10'd301,
    COMP_LOOP_C_192 = 10'd302,
    COMP_LOOP_C_193 = 10'd303,
    COMP_LOOP_7_modExp_dev_1_while_C_0 = 10'd304,
    COMP_LOOP_7_modExp_dev_1_while_C_1 = 10'd305,
    COMP_LOOP_7_modExp_dev_1_while_C_2 = 10'd306,
    COMP_LOOP_7_modExp_dev_1_while_C_3 = 10'd307,
    COMP_LOOP_7_modExp_dev_1_while_C_4 = 10'd308,
    COMP_LOOP_7_modExp_dev_1_while_C_5 = 10'd309,
    COMP_LOOP_7_modExp_dev_1_while_C_6 = 10'd310,
    COMP_LOOP_7_modExp_dev_1_while_C_7 = 10'd311,
    COMP_LOOP_7_modExp_dev_1_while_C_8 = 10'd312,
    COMP_LOOP_7_modExp_dev_1_while_C_9 = 10'd313,
    COMP_LOOP_7_modExp_dev_1_while_C_10 = 10'd314,
    COMP_LOOP_7_modExp_dev_1_while_C_11 = 10'd315,
    COMP_LOOP_7_modExp_dev_1_while_C_12 = 10'd316,
    COMP_LOOP_7_modExp_dev_1_while_C_13 = 10'd317,
    COMP_LOOP_7_modExp_dev_1_while_C_14 = 10'd318,
    COMP_LOOP_C_194 = 10'd319,
    COMP_LOOP_C_195 = 10'd320,
    COMP_LOOP_C_196 = 10'd321,
    COMP_LOOP_C_197 = 10'd322,
    COMP_LOOP_C_198 = 10'd323,
    COMP_LOOP_C_199 = 10'd324,
    COMP_LOOP_C_200 = 10'd325,
    COMP_LOOP_C_201 = 10'd326,
    COMP_LOOP_C_202 = 10'd327,
    COMP_LOOP_C_203 = 10'd328,
    COMP_LOOP_C_204 = 10'd329,
    COMP_LOOP_C_205 = 10'd330,
    COMP_LOOP_C_206 = 10'd331,
    COMP_LOOP_C_207 = 10'd332,
    COMP_LOOP_C_208 = 10'd333,
    COMP_LOOP_C_209 = 10'd334,
    COMP_LOOP_C_210 = 10'd335,
    COMP_LOOP_C_211 = 10'd336,
    COMP_LOOP_C_212 = 10'd337,
    COMP_LOOP_C_213 = 10'd338,
    COMP_LOOP_C_214 = 10'd339,
    COMP_LOOP_C_215 = 10'd340,
    COMP_LOOP_C_216 = 10'd341,
    COMP_LOOP_C_217 = 10'd342,
    COMP_LOOP_C_218 = 10'd343,
    COMP_LOOP_C_219 = 10'd344,
    COMP_LOOP_C_220 = 10'd345,
    COMP_LOOP_C_221 = 10'd346,
    COMP_LOOP_C_222 = 10'd347,
    COMP_LOOP_C_223 = 10'd348,
    COMP_LOOP_C_224 = 10'd349,
    COMP_LOOP_C_225 = 10'd350,
    COMP_LOOP_8_modExp_dev_1_while_C_0 = 10'd351,
    COMP_LOOP_8_modExp_dev_1_while_C_1 = 10'd352,
    COMP_LOOP_8_modExp_dev_1_while_C_2 = 10'd353,
    COMP_LOOP_8_modExp_dev_1_while_C_3 = 10'd354,
    COMP_LOOP_8_modExp_dev_1_while_C_4 = 10'd355,
    COMP_LOOP_8_modExp_dev_1_while_C_5 = 10'd356,
    COMP_LOOP_8_modExp_dev_1_while_C_6 = 10'd357,
    COMP_LOOP_8_modExp_dev_1_while_C_7 = 10'd358,
    COMP_LOOP_8_modExp_dev_1_while_C_8 = 10'd359,
    COMP_LOOP_8_modExp_dev_1_while_C_9 = 10'd360,
    COMP_LOOP_8_modExp_dev_1_while_C_10 = 10'd361,
    COMP_LOOP_8_modExp_dev_1_while_C_11 = 10'd362,
    COMP_LOOP_8_modExp_dev_1_while_C_12 = 10'd363,
    COMP_LOOP_8_modExp_dev_1_while_C_13 = 10'd364,
    COMP_LOOP_8_modExp_dev_1_while_C_14 = 10'd365,
    COMP_LOOP_C_226 = 10'd366,
    COMP_LOOP_C_227 = 10'd367,
    COMP_LOOP_C_228 = 10'd368,
    COMP_LOOP_C_229 = 10'd369,
    COMP_LOOP_C_230 = 10'd370,
    COMP_LOOP_C_231 = 10'd371,
    COMP_LOOP_C_232 = 10'd372,
    COMP_LOOP_C_233 = 10'd373,
    COMP_LOOP_C_234 = 10'd374,
    COMP_LOOP_C_235 = 10'd375,
    COMP_LOOP_C_236 = 10'd376,
    COMP_LOOP_C_237 = 10'd377,
    COMP_LOOP_C_238 = 10'd378,
    COMP_LOOP_C_239 = 10'd379,
    COMP_LOOP_C_240 = 10'd380,
    COMP_LOOP_C_241 = 10'd381,
    COMP_LOOP_C_242 = 10'd382,
    COMP_LOOP_C_243 = 10'd383,
    COMP_LOOP_C_244 = 10'd384,
    COMP_LOOP_C_245 = 10'd385,
    COMP_LOOP_C_246 = 10'd386,
    COMP_LOOP_C_247 = 10'd387,
    COMP_LOOP_C_248 = 10'd388,
    COMP_LOOP_C_249 = 10'd389,
    COMP_LOOP_C_250 = 10'd390,
    COMP_LOOP_C_251 = 10'd391,
    COMP_LOOP_C_252 = 10'd392,
    COMP_LOOP_C_253 = 10'd393,
    COMP_LOOP_C_254 = 10'd394,
    COMP_LOOP_C_255 = 10'd395,
    COMP_LOOP_C_256 = 10'd396,
    COMP_LOOP_C_257 = 10'd397,
    COMP_LOOP_9_modExp_dev_1_while_C_0 = 10'd398,
    COMP_LOOP_9_modExp_dev_1_while_C_1 = 10'd399,
    COMP_LOOP_9_modExp_dev_1_while_C_2 = 10'd400,
    COMP_LOOP_9_modExp_dev_1_while_C_3 = 10'd401,
    COMP_LOOP_9_modExp_dev_1_while_C_4 = 10'd402,
    COMP_LOOP_9_modExp_dev_1_while_C_5 = 10'd403,
    COMP_LOOP_9_modExp_dev_1_while_C_6 = 10'd404,
    COMP_LOOP_9_modExp_dev_1_while_C_7 = 10'd405,
    COMP_LOOP_9_modExp_dev_1_while_C_8 = 10'd406,
    COMP_LOOP_9_modExp_dev_1_while_C_9 = 10'd407,
    COMP_LOOP_9_modExp_dev_1_while_C_10 = 10'd408,
    COMP_LOOP_9_modExp_dev_1_while_C_11 = 10'd409,
    COMP_LOOP_9_modExp_dev_1_while_C_12 = 10'd410,
    COMP_LOOP_9_modExp_dev_1_while_C_13 = 10'd411,
    COMP_LOOP_9_modExp_dev_1_while_C_14 = 10'd412,
    COMP_LOOP_C_258 = 10'd413,
    COMP_LOOP_C_259 = 10'd414,
    COMP_LOOP_C_260 = 10'd415,
    COMP_LOOP_C_261 = 10'd416,
    COMP_LOOP_C_262 = 10'd417,
    COMP_LOOP_C_263 = 10'd418,
    COMP_LOOP_C_264 = 10'd419,
    COMP_LOOP_C_265 = 10'd420,
    COMP_LOOP_C_266 = 10'd421,
    COMP_LOOP_C_267 = 10'd422,
    COMP_LOOP_C_268 = 10'd423,
    COMP_LOOP_C_269 = 10'd424,
    COMP_LOOP_C_270 = 10'd425,
    COMP_LOOP_C_271 = 10'd426,
    COMP_LOOP_C_272 = 10'd427,
    COMP_LOOP_C_273 = 10'd428,
    COMP_LOOP_C_274 = 10'd429,
    COMP_LOOP_C_275 = 10'd430,
    COMP_LOOP_C_276 = 10'd431,
    COMP_LOOP_C_277 = 10'd432,
    COMP_LOOP_C_278 = 10'd433,
    COMP_LOOP_C_279 = 10'd434,
    COMP_LOOP_C_280 = 10'd435,
    COMP_LOOP_C_281 = 10'd436,
    COMP_LOOP_C_282 = 10'd437,
    COMP_LOOP_C_283 = 10'd438,
    COMP_LOOP_C_284 = 10'd439,
    COMP_LOOP_C_285 = 10'd440,
    COMP_LOOP_C_286 = 10'd441,
    COMP_LOOP_C_287 = 10'd442,
    COMP_LOOP_C_288 = 10'd443,
    COMP_LOOP_C_289 = 10'd444,
    COMP_LOOP_10_modExp_dev_1_while_C_0 = 10'd445,
    COMP_LOOP_10_modExp_dev_1_while_C_1 = 10'd446,
    COMP_LOOP_10_modExp_dev_1_while_C_2 = 10'd447,
    COMP_LOOP_10_modExp_dev_1_while_C_3 = 10'd448,
    COMP_LOOP_10_modExp_dev_1_while_C_4 = 10'd449,
    COMP_LOOP_10_modExp_dev_1_while_C_5 = 10'd450,
    COMP_LOOP_10_modExp_dev_1_while_C_6 = 10'd451,
    COMP_LOOP_10_modExp_dev_1_while_C_7 = 10'd452,
    COMP_LOOP_10_modExp_dev_1_while_C_8 = 10'd453,
    COMP_LOOP_10_modExp_dev_1_while_C_9 = 10'd454,
    COMP_LOOP_10_modExp_dev_1_while_C_10 = 10'd455,
    COMP_LOOP_10_modExp_dev_1_while_C_11 = 10'd456,
    COMP_LOOP_10_modExp_dev_1_while_C_12 = 10'd457,
    COMP_LOOP_10_modExp_dev_1_while_C_13 = 10'd458,
    COMP_LOOP_10_modExp_dev_1_while_C_14 = 10'd459,
    COMP_LOOP_C_290 = 10'd460,
    COMP_LOOP_C_291 = 10'd461,
    COMP_LOOP_C_292 = 10'd462,
    COMP_LOOP_C_293 = 10'd463,
    COMP_LOOP_C_294 = 10'd464,
    COMP_LOOP_C_295 = 10'd465,
    COMP_LOOP_C_296 = 10'd466,
    COMP_LOOP_C_297 = 10'd467,
    COMP_LOOP_C_298 = 10'd468,
    COMP_LOOP_C_299 = 10'd469,
    COMP_LOOP_C_300 = 10'd470,
    COMP_LOOP_C_301 = 10'd471,
    COMP_LOOP_C_302 = 10'd472,
    COMP_LOOP_C_303 = 10'd473,
    COMP_LOOP_C_304 = 10'd474,
    COMP_LOOP_C_305 = 10'd475,
    COMP_LOOP_C_306 = 10'd476,
    COMP_LOOP_C_307 = 10'd477,
    COMP_LOOP_C_308 = 10'd478,
    COMP_LOOP_C_309 = 10'd479,
    COMP_LOOP_C_310 = 10'd480,
    COMP_LOOP_C_311 = 10'd481,
    COMP_LOOP_C_312 = 10'd482,
    COMP_LOOP_C_313 = 10'd483,
    COMP_LOOP_C_314 = 10'd484,
    COMP_LOOP_C_315 = 10'd485,
    COMP_LOOP_C_316 = 10'd486,
    COMP_LOOP_C_317 = 10'd487,
    COMP_LOOP_C_318 = 10'd488,
    COMP_LOOP_C_319 = 10'd489,
    COMP_LOOP_C_320 = 10'd490,
    COMP_LOOP_C_321 = 10'd491,
    COMP_LOOP_11_modExp_dev_1_while_C_0 = 10'd492,
    COMP_LOOP_11_modExp_dev_1_while_C_1 = 10'd493,
    COMP_LOOP_11_modExp_dev_1_while_C_2 = 10'd494,
    COMP_LOOP_11_modExp_dev_1_while_C_3 = 10'd495,
    COMP_LOOP_11_modExp_dev_1_while_C_4 = 10'd496,
    COMP_LOOP_11_modExp_dev_1_while_C_5 = 10'd497,
    COMP_LOOP_11_modExp_dev_1_while_C_6 = 10'd498,
    COMP_LOOP_11_modExp_dev_1_while_C_7 = 10'd499,
    COMP_LOOP_11_modExp_dev_1_while_C_8 = 10'd500,
    COMP_LOOP_11_modExp_dev_1_while_C_9 = 10'd501,
    COMP_LOOP_11_modExp_dev_1_while_C_10 = 10'd502,
    COMP_LOOP_11_modExp_dev_1_while_C_11 = 10'd503,
    COMP_LOOP_11_modExp_dev_1_while_C_12 = 10'd504,
    COMP_LOOP_11_modExp_dev_1_while_C_13 = 10'd505,
    COMP_LOOP_11_modExp_dev_1_while_C_14 = 10'd506,
    COMP_LOOP_C_322 = 10'd507,
    COMP_LOOP_C_323 = 10'd508,
    COMP_LOOP_C_324 = 10'd509,
    COMP_LOOP_C_325 = 10'd510,
    COMP_LOOP_C_326 = 10'd511,
    COMP_LOOP_C_327 = 10'd512,
    COMP_LOOP_C_328 = 10'd513,
    COMP_LOOP_C_329 = 10'd514,
    COMP_LOOP_C_330 = 10'd515,
    COMP_LOOP_C_331 = 10'd516,
    COMP_LOOP_C_332 = 10'd517,
    COMP_LOOP_C_333 = 10'd518,
    COMP_LOOP_C_334 = 10'd519,
    COMP_LOOP_C_335 = 10'd520,
    COMP_LOOP_C_336 = 10'd521,
    COMP_LOOP_C_337 = 10'd522,
    COMP_LOOP_C_338 = 10'd523,
    COMP_LOOP_C_339 = 10'd524,
    COMP_LOOP_C_340 = 10'd525,
    COMP_LOOP_C_341 = 10'd526,
    COMP_LOOP_C_342 = 10'd527,
    COMP_LOOP_C_343 = 10'd528,
    COMP_LOOP_C_344 = 10'd529,
    COMP_LOOP_C_345 = 10'd530,
    COMP_LOOP_C_346 = 10'd531,
    COMP_LOOP_C_347 = 10'd532,
    COMP_LOOP_C_348 = 10'd533,
    COMP_LOOP_C_349 = 10'd534,
    COMP_LOOP_C_350 = 10'd535,
    COMP_LOOP_C_351 = 10'd536,
    COMP_LOOP_C_352 = 10'd537,
    COMP_LOOP_C_353 = 10'd538,
    COMP_LOOP_12_modExp_dev_1_while_C_0 = 10'd539,
    COMP_LOOP_12_modExp_dev_1_while_C_1 = 10'd540,
    COMP_LOOP_12_modExp_dev_1_while_C_2 = 10'd541,
    COMP_LOOP_12_modExp_dev_1_while_C_3 = 10'd542,
    COMP_LOOP_12_modExp_dev_1_while_C_4 = 10'd543,
    COMP_LOOP_12_modExp_dev_1_while_C_5 = 10'd544,
    COMP_LOOP_12_modExp_dev_1_while_C_6 = 10'd545,
    COMP_LOOP_12_modExp_dev_1_while_C_7 = 10'd546,
    COMP_LOOP_12_modExp_dev_1_while_C_8 = 10'd547,
    COMP_LOOP_12_modExp_dev_1_while_C_9 = 10'd548,
    COMP_LOOP_12_modExp_dev_1_while_C_10 = 10'd549,
    COMP_LOOP_12_modExp_dev_1_while_C_11 = 10'd550,
    COMP_LOOP_12_modExp_dev_1_while_C_12 = 10'd551,
    COMP_LOOP_12_modExp_dev_1_while_C_13 = 10'd552,
    COMP_LOOP_12_modExp_dev_1_while_C_14 = 10'd553,
    COMP_LOOP_C_354 = 10'd554,
    COMP_LOOP_C_355 = 10'd555,
    COMP_LOOP_C_356 = 10'd556,
    COMP_LOOP_C_357 = 10'd557,
    COMP_LOOP_C_358 = 10'd558,
    COMP_LOOP_C_359 = 10'd559,
    COMP_LOOP_C_360 = 10'd560,
    COMP_LOOP_C_361 = 10'd561,
    COMP_LOOP_C_362 = 10'd562,
    COMP_LOOP_C_363 = 10'd563,
    COMP_LOOP_C_364 = 10'd564,
    COMP_LOOP_C_365 = 10'd565,
    COMP_LOOP_C_366 = 10'd566,
    COMP_LOOP_C_367 = 10'd567,
    COMP_LOOP_C_368 = 10'd568,
    COMP_LOOP_C_369 = 10'd569,
    COMP_LOOP_C_370 = 10'd570,
    COMP_LOOP_C_371 = 10'd571,
    COMP_LOOP_C_372 = 10'd572,
    COMP_LOOP_C_373 = 10'd573,
    COMP_LOOP_C_374 = 10'd574,
    COMP_LOOP_C_375 = 10'd575,
    COMP_LOOP_C_376 = 10'd576,
    COMP_LOOP_C_377 = 10'd577,
    COMP_LOOP_C_378 = 10'd578,
    COMP_LOOP_C_379 = 10'd579,
    COMP_LOOP_C_380 = 10'd580,
    COMP_LOOP_C_381 = 10'd581,
    COMP_LOOP_C_382 = 10'd582,
    COMP_LOOP_C_383 = 10'd583,
    COMP_LOOP_C_384 = 10'd584,
    COMP_LOOP_C_385 = 10'd585,
    COMP_LOOP_13_modExp_dev_1_while_C_0 = 10'd586,
    COMP_LOOP_13_modExp_dev_1_while_C_1 = 10'd587,
    COMP_LOOP_13_modExp_dev_1_while_C_2 = 10'd588,
    COMP_LOOP_13_modExp_dev_1_while_C_3 = 10'd589,
    COMP_LOOP_13_modExp_dev_1_while_C_4 = 10'd590,
    COMP_LOOP_13_modExp_dev_1_while_C_5 = 10'd591,
    COMP_LOOP_13_modExp_dev_1_while_C_6 = 10'd592,
    COMP_LOOP_13_modExp_dev_1_while_C_7 = 10'd593,
    COMP_LOOP_13_modExp_dev_1_while_C_8 = 10'd594,
    COMP_LOOP_13_modExp_dev_1_while_C_9 = 10'd595,
    COMP_LOOP_13_modExp_dev_1_while_C_10 = 10'd596,
    COMP_LOOP_13_modExp_dev_1_while_C_11 = 10'd597,
    COMP_LOOP_13_modExp_dev_1_while_C_12 = 10'd598,
    COMP_LOOP_13_modExp_dev_1_while_C_13 = 10'd599,
    COMP_LOOP_13_modExp_dev_1_while_C_14 = 10'd600,
    COMP_LOOP_C_386 = 10'd601,
    COMP_LOOP_C_387 = 10'd602,
    COMP_LOOP_C_388 = 10'd603,
    COMP_LOOP_C_389 = 10'd604,
    COMP_LOOP_C_390 = 10'd605,
    COMP_LOOP_C_391 = 10'd606,
    COMP_LOOP_C_392 = 10'd607,
    COMP_LOOP_C_393 = 10'd608,
    COMP_LOOP_C_394 = 10'd609,
    COMP_LOOP_C_395 = 10'd610,
    COMP_LOOP_C_396 = 10'd611,
    COMP_LOOP_C_397 = 10'd612,
    COMP_LOOP_C_398 = 10'd613,
    COMP_LOOP_C_399 = 10'd614,
    COMP_LOOP_C_400 = 10'd615,
    COMP_LOOP_C_401 = 10'd616,
    COMP_LOOP_C_402 = 10'd617,
    COMP_LOOP_C_403 = 10'd618,
    COMP_LOOP_C_404 = 10'd619,
    COMP_LOOP_C_405 = 10'd620,
    COMP_LOOP_C_406 = 10'd621,
    COMP_LOOP_C_407 = 10'd622,
    COMP_LOOP_C_408 = 10'd623,
    COMP_LOOP_C_409 = 10'd624,
    COMP_LOOP_C_410 = 10'd625,
    COMP_LOOP_C_411 = 10'd626,
    COMP_LOOP_C_412 = 10'd627,
    COMP_LOOP_C_413 = 10'd628,
    COMP_LOOP_C_414 = 10'd629,
    COMP_LOOP_C_415 = 10'd630,
    COMP_LOOP_C_416 = 10'd631,
    COMP_LOOP_C_417 = 10'd632,
    COMP_LOOP_14_modExp_dev_1_while_C_0 = 10'd633,
    COMP_LOOP_14_modExp_dev_1_while_C_1 = 10'd634,
    COMP_LOOP_14_modExp_dev_1_while_C_2 = 10'd635,
    COMP_LOOP_14_modExp_dev_1_while_C_3 = 10'd636,
    COMP_LOOP_14_modExp_dev_1_while_C_4 = 10'd637,
    COMP_LOOP_14_modExp_dev_1_while_C_5 = 10'd638,
    COMP_LOOP_14_modExp_dev_1_while_C_6 = 10'd639,
    COMP_LOOP_14_modExp_dev_1_while_C_7 = 10'd640,
    COMP_LOOP_14_modExp_dev_1_while_C_8 = 10'd641,
    COMP_LOOP_14_modExp_dev_1_while_C_9 = 10'd642,
    COMP_LOOP_14_modExp_dev_1_while_C_10 = 10'd643,
    COMP_LOOP_14_modExp_dev_1_while_C_11 = 10'd644,
    COMP_LOOP_14_modExp_dev_1_while_C_12 = 10'd645,
    COMP_LOOP_14_modExp_dev_1_while_C_13 = 10'd646,
    COMP_LOOP_14_modExp_dev_1_while_C_14 = 10'd647,
    COMP_LOOP_C_418 = 10'd648,
    COMP_LOOP_C_419 = 10'd649,
    COMP_LOOP_C_420 = 10'd650,
    COMP_LOOP_C_421 = 10'd651,
    COMP_LOOP_C_422 = 10'd652,
    COMP_LOOP_C_423 = 10'd653,
    COMP_LOOP_C_424 = 10'd654,
    COMP_LOOP_C_425 = 10'd655,
    COMP_LOOP_C_426 = 10'd656,
    COMP_LOOP_C_427 = 10'd657,
    COMP_LOOP_C_428 = 10'd658,
    COMP_LOOP_C_429 = 10'd659,
    COMP_LOOP_C_430 = 10'd660,
    COMP_LOOP_C_431 = 10'd661,
    COMP_LOOP_C_432 = 10'd662,
    COMP_LOOP_C_433 = 10'd663,
    COMP_LOOP_C_434 = 10'd664,
    COMP_LOOP_C_435 = 10'd665,
    COMP_LOOP_C_436 = 10'd666,
    COMP_LOOP_C_437 = 10'd667,
    COMP_LOOP_C_438 = 10'd668,
    COMP_LOOP_C_439 = 10'd669,
    COMP_LOOP_C_440 = 10'd670,
    COMP_LOOP_C_441 = 10'd671,
    COMP_LOOP_C_442 = 10'd672,
    COMP_LOOP_C_443 = 10'd673,
    COMP_LOOP_C_444 = 10'd674,
    COMP_LOOP_C_445 = 10'd675,
    COMP_LOOP_C_446 = 10'd676,
    COMP_LOOP_C_447 = 10'd677,
    COMP_LOOP_C_448 = 10'd678,
    COMP_LOOP_C_449 = 10'd679,
    COMP_LOOP_15_modExp_dev_1_while_C_0 = 10'd680,
    COMP_LOOP_15_modExp_dev_1_while_C_1 = 10'd681,
    COMP_LOOP_15_modExp_dev_1_while_C_2 = 10'd682,
    COMP_LOOP_15_modExp_dev_1_while_C_3 = 10'd683,
    COMP_LOOP_15_modExp_dev_1_while_C_4 = 10'd684,
    COMP_LOOP_15_modExp_dev_1_while_C_5 = 10'd685,
    COMP_LOOP_15_modExp_dev_1_while_C_6 = 10'd686,
    COMP_LOOP_15_modExp_dev_1_while_C_7 = 10'd687,
    COMP_LOOP_15_modExp_dev_1_while_C_8 = 10'd688,
    COMP_LOOP_15_modExp_dev_1_while_C_9 = 10'd689,
    COMP_LOOP_15_modExp_dev_1_while_C_10 = 10'd690,
    COMP_LOOP_15_modExp_dev_1_while_C_11 = 10'd691,
    COMP_LOOP_15_modExp_dev_1_while_C_12 = 10'd692,
    COMP_LOOP_15_modExp_dev_1_while_C_13 = 10'd693,
    COMP_LOOP_15_modExp_dev_1_while_C_14 = 10'd694,
    COMP_LOOP_C_450 = 10'd695,
    COMP_LOOP_C_451 = 10'd696,
    COMP_LOOP_C_452 = 10'd697,
    COMP_LOOP_C_453 = 10'd698,
    COMP_LOOP_C_454 = 10'd699,
    COMP_LOOP_C_455 = 10'd700,
    COMP_LOOP_C_456 = 10'd701,
    COMP_LOOP_C_457 = 10'd702,
    COMP_LOOP_C_458 = 10'd703,
    COMP_LOOP_C_459 = 10'd704,
    COMP_LOOP_C_460 = 10'd705,
    COMP_LOOP_C_461 = 10'd706,
    COMP_LOOP_C_462 = 10'd707,
    COMP_LOOP_C_463 = 10'd708,
    COMP_LOOP_C_464 = 10'd709,
    COMP_LOOP_C_465 = 10'd710,
    COMP_LOOP_C_466 = 10'd711,
    COMP_LOOP_C_467 = 10'd712,
    COMP_LOOP_C_468 = 10'd713,
    COMP_LOOP_C_469 = 10'd714,
    COMP_LOOP_C_470 = 10'd715,
    COMP_LOOP_C_471 = 10'd716,
    COMP_LOOP_C_472 = 10'd717,
    COMP_LOOP_C_473 = 10'd718,
    COMP_LOOP_C_474 = 10'd719,
    COMP_LOOP_C_475 = 10'd720,
    COMP_LOOP_C_476 = 10'd721,
    COMP_LOOP_C_477 = 10'd722,
    COMP_LOOP_C_478 = 10'd723,
    COMP_LOOP_C_479 = 10'd724,
    COMP_LOOP_C_480 = 10'd725,
    COMP_LOOP_C_481 = 10'd726,
    COMP_LOOP_16_modExp_dev_1_while_C_0 = 10'd727,
    COMP_LOOP_16_modExp_dev_1_while_C_1 = 10'd728,
    COMP_LOOP_16_modExp_dev_1_while_C_2 = 10'd729,
    COMP_LOOP_16_modExp_dev_1_while_C_3 = 10'd730,
    COMP_LOOP_16_modExp_dev_1_while_C_4 = 10'd731,
    COMP_LOOP_16_modExp_dev_1_while_C_5 = 10'd732,
    COMP_LOOP_16_modExp_dev_1_while_C_6 = 10'd733,
    COMP_LOOP_16_modExp_dev_1_while_C_7 = 10'd734,
    COMP_LOOP_16_modExp_dev_1_while_C_8 = 10'd735,
    COMP_LOOP_16_modExp_dev_1_while_C_9 = 10'd736,
    COMP_LOOP_16_modExp_dev_1_while_C_10 = 10'd737,
    COMP_LOOP_16_modExp_dev_1_while_C_11 = 10'd738,
    COMP_LOOP_16_modExp_dev_1_while_C_12 = 10'd739,
    COMP_LOOP_16_modExp_dev_1_while_C_13 = 10'd740,
    COMP_LOOP_16_modExp_dev_1_while_C_14 = 10'd741,
    COMP_LOOP_C_482 = 10'd742,
    COMP_LOOP_C_483 = 10'd743,
    COMP_LOOP_C_484 = 10'd744,
    COMP_LOOP_C_485 = 10'd745,
    COMP_LOOP_C_486 = 10'd746,
    COMP_LOOP_C_487 = 10'd747,
    COMP_LOOP_C_488 = 10'd748,
    COMP_LOOP_C_489 = 10'd749,
    COMP_LOOP_C_490 = 10'd750,
    COMP_LOOP_C_491 = 10'd751,
    COMP_LOOP_C_492 = 10'd752,
    COMP_LOOP_C_493 = 10'd753,
    COMP_LOOP_C_494 = 10'd754,
    COMP_LOOP_C_495 = 10'd755,
    COMP_LOOP_C_496 = 10'd756,
    COMP_LOOP_C_497 = 10'd757,
    COMP_LOOP_C_498 = 10'd758,
    COMP_LOOP_C_499 = 10'd759,
    COMP_LOOP_C_500 = 10'd760,
    COMP_LOOP_C_501 = 10'd761,
    COMP_LOOP_C_502 = 10'd762,
    COMP_LOOP_C_503 = 10'd763,
    COMP_LOOP_C_504 = 10'd764,
    COMP_LOOP_C_505 = 10'd765,
    COMP_LOOP_C_506 = 10'd766,
    COMP_LOOP_C_507 = 10'd767,
    COMP_LOOP_C_508 = 10'd768,
    COMP_LOOP_C_509 = 10'd769,
    COMP_LOOP_C_510 = 10'd770,
    COMP_LOOP_C_511 = 10'd771,
    COMP_LOOP_C_512 = 10'd772,
    VEC_LOOP_C_0 = 10'd773,
    STAGE_LOOP_C_4 = 10'd774,
    main_C_1 = 10'd775;

  reg [9:0] state_var;
  reg [9:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : inPlaceNTT_DIT_core_core_fsm_1
    case (state_var)
      STAGE_LOOP_C_0 : begin
        fsm_output = 10'b0000000001;
        state_var_NS = STAGE_LOOP_C_1;
      end
      STAGE_LOOP_C_1 : begin
        fsm_output = 10'b0000000010;
        state_var_NS = STAGE_LOOP_C_2;
      end
      STAGE_LOOP_C_2 : begin
        fsm_output = 10'b0000000011;
        state_var_NS = STAGE_LOOP_C_3;
      end
      STAGE_LOOP_C_3 : begin
        fsm_output = 10'b0000000100;
        if ( STAGE_LOOP_C_3_tr0 ) begin
          state_var_NS = COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_dev_while_C_0;
        end
      end
      modExp_dev_while_C_0 : begin
        fsm_output = 10'b0000000101;
        state_var_NS = modExp_dev_while_C_1;
      end
      modExp_dev_while_C_1 : begin
        fsm_output = 10'b0000000110;
        state_var_NS = modExp_dev_while_C_2;
      end
      modExp_dev_while_C_2 : begin
        fsm_output = 10'b0000000111;
        state_var_NS = modExp_dev_while_C_3;
      end
      modExp_dev_while_C_3 : begin
        fsm_output = 10'b0000001000;
        state_var_NS = modExp_dev_while_C_4;
      end
      modExp_dev_while_C_4 : begin
        fsm_output = 10'b0000001001;
        state_var_NS = modExp_dev_while_C_5;
      end
      modExp_dev_while_C_5 : begin
        fsm_output = 10'b0000001010;
        state_var_NS = modExp_dev_while_C_6;
      end
      modExp_dev_while_C_6 : begin
        fsm_output = 10'b0000001011;
        state_var_NS = modExp_dev_while_C_7;
      end
      modExp_dev_while_C_7 : begin
        fsm_output = 10'b0000001100;
        state_var_NS = modExp_dev_while_C_8;
      end
      modExp_dev_while_C_8 : begin
        fsm_output = 10'b0000001101;
        state_var_NS = modExp_dev_while_C_9;
      end
      modExp_dev_while_C_9 : begin
        fsm_output = 10'b0000001110;
        state_var_NS = modExp_dev_while_C_10;
      end
      modExp_dev_while_C_10 : begin
        fsm_output = 10'b0000001111;
        state_var_NS = modExp_dev_while_C_11;
      end
      modExp_dev_while_C_11 : begin
        fsm_output = 10'b0000010000;
        state_var_NS = modExp_dev_while_C_12;
      end
      modExp_dev_while_C_12 : begin
        fsm_output = 10'b0000010001;
        state_var_NS = modExp_dev_while_C_13;
      end
      modExp_dev_while_C_13 : begin
        fsm_output = 10'b0000010010;
        state_var_NS = modExp_dev_while_C_14;
      end
      modExp_dev_while_C_14 : begin
        fsm_output = 10'b0000010011;
        if ( modExp_dev_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_dev_while_C_0;
        end
      end
      COMP_LOOP_C_0 : begin
        fsm_output = 10'b0000010100;
        state_var_NS = COMP_LOOP_C_1;
      end
      COMP_LOOP_C_1 : begin
        fsm_output = 10'b0000010101;
        if ( COMP_LOOP_C_1_tr0 ) begin
          state_var_NS = COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_1_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0000010110;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0000010111;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0000011000;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0000011001;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0000011010;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0000011011;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0000011100;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0000011101;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0000011110;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0000011111;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0000100000;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0000100001;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_12;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_12 : begin
        fsm_output = 10'b0000100010;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_13;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_13 : begin
        fsm_output = 10'b0000100011;
        state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_14;
      end
      COMP_LOOP_1_modExp_dev_1_while_C_14 : begin
        fsm_output = 10'b0000100100;
        if ( COMP_LOOP_1_modExp_dev_1_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = COMP_LOOP_1_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_2 : begin
        fsm_output = 10'b0000100101;
        state_var_NS = COMP_LOOP_C_3;
      end
      COMP_LOOP_C_3 : begin
        fsm_output = 10'b0000100110;
        state_var_NS = COMP_LOOP_C_4;
      end
      COMP_LOOP_C_4 : begin
        fsm_output = 10'b0000100111;
        state_var_NS = COMP_LOOP_C_5;
      end
      COMP_LOOP_C_5 : begin
        fsm_output = 10'b0000101000;
        state_var_NS = COMP_LOOP_C_6;
      end
      COMP_LOOP_C_6 : begin
        fsm_output = 10'b0000101001;
        state_var_NS = COMP_LOOP_C_7;
      end
      COMP_LOOP_C_7 : begin
        fsm_output = 10'b0000101010;
        state_var_NS = COMP_LOOP_C_8;
      end
      COMP_LOOP_C_8 : begin
        fsm_output = 10'b0000101011;
        state_var_NS = COMP_LOOP_C_9;
      end
      COMP_LOOP_C_9 : begin
        fsm_output = 10'b0000101100;
        state_var_NS = COMP_LOOP_C_10;
      end
      COMP_LOOP_C_10 : begin
        fsm_output = 10'b0000101101;
        state_var_NS = COMP_LOOP_C_11;
      end
      COMP_LOOP_C_11 : begin
        fsm_output = 10'b0000101110;
        state_var_NS = COMP_LOOP_C_12;
      end
      COMP_LOOP_C_12 : begin
        fsm_output = 10'b0000101111;
        state_var_NS = COMP_LOOP_C_13;
      end
      COMP_LOOP_C_13 : begin
        fsm_output = 10'b0000110000;
        state_var_NS = COMP_LOOP_C_14;
      end
      COMP_LOOP_C_14 : begin
        fsm_output = 10'b0000110001;
        state_var_NS = COMP_LOOP_C_15;
      end
      COMP_LOOP_C_15 : begin
        fsm_output = 10'b0000110010;
        state_var_NS = COMP_LOOP_C_16;
      end
      COMP_LOOP_C_16 : begin
        fsm_output = 10'b0000110011;
        state_var_NS = COMP_LOOP_C_17;
      end
      COMP_LOOP_C_17 : begin
        fsm_output = 10'b0000110100;
        state_var_NS = COMP_LOOP_C_18;
      end
      COMP_LOOP_C_18 : begin
        fsm_output = 10'b0000110101;
        state_var_NS = COMP_LOOP_C_19;
      end
      COMP_LOOP_C_19 : begin
        fsm_output = 10'b0000110110;
        state_var_NS = COMP_LOOP_C_20;
      end
      COMP_LOOP_C_20 : begin
        fsm_output = 10'b0000110111;
        state_var_NS = COMP_LOOP_C_21;
      end
      COMP_LOOP_C_21 : begin
        fsm_output = 10'b0000111000;
        state_var_NS = COMP_LOOP_C_22;
      end
      COMP_LOOP_C_22 : begin
        fsm_output = 10'b0000111001;
        state_var_NS = COMP_LOOP_C_23;
      end
      COMP_LOOP_C_23 : begin
        fsm_output = 10'b0000111010;
        state_var_NS = COMP_LOOP_C_24;
      end
      COMP_LOOP_C_24 : begin
        fsm_output = 10'b0000111011;
        state_var_NS = COMP_LOOP_C_25;
      end
      COMP_LOOP_C_25 : begin
        fsm_output = 10'b0000111100;
        state_var_NS = COMP_LOOP_C_26;
      end
      COMP_LOOP_C_26 : begin
        fsm_output = 10'b0000111101;
        state_var_NS = COMP_LOOP_C_27;
      end
      COMP_LOOP_C_27 : begin
        fsm_output = 10'b0000111110;
        state_var_NS = COMP_LOOP_C_28;
      end
      COMP_LOOP_C_28 : begin
        fsm_output = 10'b0000111111;
        state_var_NS = COMP_LOOP_C_29;
      end
      COMP_LOOP_C_29 : begin
        fsm_output = 10'b0001000000;
        state_var_NS = COMP_LOOP_C_30;
      end
      COMP_LOOP_C_30 : begin
        fsm_output = 10'b0001000001;
        state_var_NS = COMP_LOOP_C_31;
      end
      COMP_LOOP_C_31 : begin
        fsm_output = 10'b0001000010;
        state_var_NS = COMP_LOOP_C_32;
      end
      COMP_LOOP_C_32 : begin
        fsm_output = 10'b0001000011;
        if ( COMP_LOOP_C_32_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_33;
        end
      end
      COMP_LOOP_C_33 : begin
        fsm_output = 10'b0001000100;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0001000101;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0001000110;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0001000111;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0001001000;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0001001001;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0001001010;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0001001011;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0001001100;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0001001101;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0001001110;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0001001111;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0001010000;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_12;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_12 : begin
        fsm_output = 10'b0001010001;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_13;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_13 : begin
        fsm_output = 10'b0001010010;
        state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_14;
      end
      COMP_LOOP_2_modExp_dev_1_while_C_14 : begin
        fsm_output = 10'b0001010011;
        if ( COMP_LOOP_2_modExp_dev_1_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_34;
        end
        else begin
          state_var_NS = COMP_LOOP_2_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_34 : begin
        fsm_output = 10'b0001010100;
        state_var_NS = COMP_LOOP_C_35;
      end
      COMP_LOOP_C_35 : begin
        fsm_output = 10'b0001010101;
        state_var_NS = COMP_LOOP_C_36;
      end
      COMP_LOOP_C_36 : begin
        fsm_output = 10'b0001010110;
        state_var_NS = COMP_LOOP_C_37;
      end
      COMP_LOOP_C_37 : begin
        fsm_output = 10'b0001010111;
        state_var_NS = COMP_LOOP_C_38;
      end
      COMP_LOOP_C_38 : begin
        fsm_output = 10'b0001011000;
        state_var_NS = COMP_LOOP_C_39;
      end
      COMP_LOOP_C_39 : begin
        fsm_output = 10'b0001011001;
        state_var_NS = COMP_LOOP_C_40;
      end
      COMP_LOOP_C_40 : begin
        fsm_output = 10'b0001011010;
        state_var_NS = COMP_LOOP_C_41;
      end
      COMP_LOOP_C_41 : begin
        fsm_output = 10'b0001011011;
        state_var_NS = COMP_LOOP_C_42;
      end
      COMP_LOOP_C_42 : begin
        fsm_output = 10'b0001011100;
        state_var_NS = COMP_LOOP_C_43;
      end
      COMP_LOOP_C_43 : begin
        fsm_output = 10'b0001011101;
        state_var_NS = COMP_LOOP_C_44;
      end
      COMP_LOOP_C_44 : begin
        fsm_output = 10'b0001011110;
        state_var_NS = COMP_LOOP_C_45;
      end
      COMP_LOOP_C_45 : begin
        fsm_output = 10'b0001011111;
        state_var_NS = COMP_LOOP_C_46;
      end
      COMP_LOOP_C_46 : begin
        fsm_output = 10'b0001100000;
        state_var_NS = COMP_LOOP_C_47;
      end
      COMP_LOOP_C_47 : begin
        fsm_output = 10'b0001100001;
        state_var_NS = COMP_LOOP_C_48;
      end
      COMP_LOOP_C_48 : begin
        fsm_output = 10'b0001100010;
        state_var_NS = COMP_LOOP_C_49;
      end
      COMP_LOOP_C_49 : begin
        fsm_output = 10'b0001100011;
        state_var_NS = COMP_LOOP_C_50;
      end
      COMP_LOOP_C_50 : begin
        fsm_output = 10'b0001100100;
        state_var_NS = COMP_LOOP_C_51;
      end
      COMP_LOOP_C_51 : begin
        fsm_output = 10'b0001100101;
        state_var_NS = COMP_LOOP_C_52;
      end
      COMP_LOOP_C_52 : begin
        fsm_output = 10'b0001100110;
        state_var_NS = COMP_LOOP_C_53;
      end
      COMP_LOOP_C_53 : begin
        fsm_output = 10'b0001100111;
        state_var_NS = COMP_LOOP_C_54;
      end
      COMP_LOOP_C_54 : begin
        fsm_output = 10'b0001101000;
        state_var_NS = COMP_LOOP_C_55;
      end
      COMP_LOOP_C_55 : begin
        fsm_output = 10'b0001101001;
        state_var_NS = COMP_LOOP_C_56;
      end
      COMP_LOOP_C_56 : begin
        fsm_output = 10'b0001101010;
        state_var_NS = COMP_LOOP_C_57;
      end
      COMP_LOOP_C_57 : begin
        fsm_output = 10'b0001101011;
        state_var_NS = COMP_LOOP_C_58;
      end
      COMP_LOOP_C_58 : begin
        fsm_output = 10'b0001101100;
        state_var_NS = COMP_LOOP_C_59;
      end
      COMP_LOOP_C_59 : begin
        fsm_output = 10'b0001101101;
        state_var_NS = COMP_LOOP_C_60;
      end
      COMP_LOOP_C_60 : begin
        fsm_output = 10'b0001101110;
        state_var_NS = COMP_LOOP_C_61;
      end
      COMP_LOOP_C_61 : begin
        fsm_output = 10'b0001101111;
        state_var_NS = COMP_LOOP_C_62;
      end
      COMP_LOOP_C_62 : begin
        fsm_output = 10'b0001110000;
        state_var_NS = COMP_LOOP_C_63;
      end
      COMP_LOOP_C_63 : begin
        fsm_output = 10'b0001110001;
        state_var_NS = COMP_LOOP_C_64;
      end
      COMP_LOOP_C_64 : begin
        fsm_output = 10'b0001110010;
        if ( COMP_LOOP_C_64_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_65;
        end
      end
      COMP_LOOP_C_65 : begin
        fsm_output = 10'b0001110011;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0001110100;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0001110101;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0001110110;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0001110111;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0001111000;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0001111001;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0001111010;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0001111011;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0001111100;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0001111101;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0001111110;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0001111111;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_12;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_12 : begin
        fsm_output = 10'b0010000000;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_13;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_13 : begin
        fsm_output = 10'b0010000001;
        state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_14;
      end
      COMP_LOOP_3_modExp_dev_1_while_C_14 : begin
        fsm_output = 10'b0010000010;
        if ( COMP_LOOP_3_modExp_dev_1_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_66;
        end
        else begin
          state_var_NS = COMP_LOOP_3_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_66 : begin
        fsm_output = 10'b0010000011;
        state_var_NS = COMP_LOOP_C_67;
      end
      COMP_LOOP_C_67 : begin
        fsm_output = 10'b0010000100;
        state_var_NS = COMP_LOOP_C_68;
      end
      COMP_LOOP_C_68 : begin
        fsm_output = 10'b0010000101;
        state_var_NS = COMP_LOOP_C_69;
      end
      COMP_LOOP_C_69 : begin
        fsm_output = 10'b0010000110;
        state_var_NS = COMP_LOOP_C_70;
      end
      COMP_LOOP_C_70 : begin
        fsm_output = 10'b0010000111;
        state_var_NS = COMP_LOOP_C_71;
      end
      COMP_LOOP_C_71 : begin
        fsm_output = 10'b0010001000;
        state_var_NS = COMP_LOOP_C_72;
      end
      COMP_LOOP_C_72 : begin
        fsm_output = 10'b0010001001;
        state_var_NS = COMP_LOOP_C_73;
      end
      COMP_LOOP_C_73 : begin
        fsm_output = 10'b0010001010;
        state_var_NS = COMP_LOOP_C_74;
      end
      COMP_LOOP_C_74 : begin
        fsm_output = 10'b0010001011;
        state_var_NS = COMP_LOOP_C_75;
      end
      COMP_LOOP_C_75 : begin
        fsm_output = 10'b0010001100;
        state_var_NS = COMP_LOOP_C_76;
      end
      COMP_LOOP_C_76 : begin
        fsm_output = 10'b0010001101;
        state_var_NS = COMP_LOOP_C_77;
      end
      COMP_LOOP_C_77 : begin
        fsm_output = 10'b0010001110;
        state_var_NS = COMP_LOOP_C_78;
      end
      COMP_LOOP_C_78 : begin
        fsm_output = 10'b0010001111;
        state_var_NS = COMP_LOOP_C_79;
      end
      COMP_LOOP_C_79 : begin
        fsm_output = 10'b0010010000;
        state_var_NS = COMP_LOOP_C_80;
      end
      COMP_LOOP_C_80 : begin
        fsm_output = 10'b0010010001;
        state_var_NS = COMP_LOOP_C_81;
      end
      COMP_LOOP_C_81 : begin
        fsm_output = 10'b0010010010;
        state_var_NS = COMP_LOOP_C_82;
      end
      COMP_LOOP_C_82 : begin
        fsm_output = 10'b0010010011;
        state_var_NS = COMP_LOOP_C_83;
      end
      COMP_LOOP_C_83 : begin
        fsm_output = 10'b0010010100;
        state_var_NS = COMP_LOOP_C_84;
      end
      COMP_LOOP_C_84 : begin
        fsm_output = 10'b0010010101;
        state_var_NS = COMP_LOOP_C_85;
      end
      COMP_LOOP_C_85 : begin
        fsm_output = 10'b0010010110;
        state_var_NS = COMP_LOOP_C_86;
      end
      COMP_LOOP_C_86 : begin
        fsm_output = 10'b0010010111;
        state_var_NS = COMP_LOOP_C_87;
      end
      COMP_LOOP_C_87 : begin
        fsm_output = 10'b0010011000;
        state_var_NS = COMP_LOOP_C_88;
      end
      COMP_LOOP_C_88 : begin
        fsm_output = 10'b0010011001;
        state_var_NS = COMP_LOOP_C_89;
      end
      COMP_LOOP_C_89 : begin
        fsm_output = 10'b0010011010;
        state_var_NS = COMP_LOOP_C_90;
      end
      COMP_LOOP_C_90 : begin
        fsm_output = 10'b0010011011;
        state_var_NS = COMP_LOOP_C_91;
      end
      COMP_LOOP_C_91 : begin
        fsm_output = 10'b0010011100;
        state_var_NS = COMP_LOOP_C_92;
      end
      COMP_LOOP_C_92 : begin
        fsm_output = 10'b0010011101;
        state_var_NS = COMP_LOOP_C_93;
      end
      COMP_LOOP_C_93 : begin
        fsm_output = 10'b0010011110;
        state_var_NS = COMP_LOOP_C_94;
      end
      COMP_LOOP_C_94 : begin
        fsm_output = 10'b0010011111;
        state_var_NS = COMP_LOOP_C_95;
      end
      COMP_LOOP_C_95 : begin
        fsm_output = 10'b0010100000;
        state_var_NS = COMP_LOOP_C_96;
      end
      COMP_LOOP_C_96 : begin
        fsm_output = 10'b0010100001;
        if ( COMP_LOOP_C_96_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_97;
        end
      end
      COMP_LOOP_C_97 : begin
        fsm_output = 10'b0010100010;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0010100011;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0010100100;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0010100101;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0010100110;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0010100111;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0010101000;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0010101001;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0010101010;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0010101011;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0010101100;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0010101101;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0010101110;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_12;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_12 : begin
        fsm_output = 10'b0010101111;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_13;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_13 : begin
        fsm_output = 10'b0010110000;
        state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_14;
      end
      COMP_LOOP_4_modExp_dev_1_while_C_14 : begin
        fsm_output = 10'b0010110001;
        if ( COMP_LOOP_4_modExp_dev_1_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_98;
        end
        else begin
          state_var_NS = COMP_LOOP_4_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_98 : begin
        fsm_output = 10'b0010110010;
        state_var_NS = COMP_LOOP_C_99;
      end
      COMP_LOOP_C_99 : begin
        fsm_output = 10'b0010110011;
        state_var_NS = COMP_LOOP_C_100;
      end
      COMP_LOOP_C_100 : begin
        fsm_output = 10'b0010110100;
        state_var_NS = COMP_LOOP_C_101;
      end
      COMP_LOOP_C_101 : begin
        fsm_output = 10'b0010110101;
        state_var_NS = COMP_LOOP_C_102;
      end
      COMP_LOOP_C_102 : begin
        fsm_output = 10'b0010110110;
        state_var_NS = COMP_LOOP_C_103;
      end
      COMP_LOOP_C_103 : begin
        fsm_output = 10'b0010110111;
        state_var_NS = COMP_LOOP_C_104;
      end
      COMP_LOOP_C_104 : begin
        fsm_output = 10'b0010111000;
        state_var_NS = COMP_LOOP_C_105;
      end
      COMP_LOOP_C_105 : begin
        fsm_output = 10'b0010111001;
        state_var_NS = COMP_LOOP_C_106;
      end
      COMP_LOOP_C_106 : begin
        fsm_output = 10'b0010111010;
        state_var_NS = COMP_LOOP_C_107;
      end
      COMP_LOOP_C_107 : begin
        fsm_output = 10'b0010111011;
        state_var_NS = COMP_LOOP_C_108;
      end
      COMP_LOOP_C_108 : begin
        fsm_output = 10'b0010111100;
        state_var_NS = COMP_LOOP_C_109;
      end
      COMP_LOOP_C_109 : begin
        fsm_output = 10'b0010111101;
        state_var_NS = COMP_LOOP_C_110;
      end
      COMP_LOOP_C_110 : begin
        fsm_output = 10'b0010111110;
        state_var_NS = COMP_LOOP_C_111;
      end
      COMP_LOOP_C_111 : begin
        fsm_output = 10'b0010111111;
        state_var_NS = COMP_LOOP_C_112;
      end
      COMP_LOOP_C_112 : begin
        fsm_output = 10'b0011000000;
        state_var_NS = COMP_LOOP_C_113;
      end
      COMP_LOOP_C_113 : begin
        fsm_output = 10'b0011000001;
        state_var_NS = COMP_LOOP_C_114;
      end
      COMP_LOOP_C_114 : begin
        fsm_output = 10'b0011000010;
        state_var_NS = COMP_LOOP_C_115;
      end
      COMP_LOOP_C_115 : begin
        fsm_output = 10'b0011000011;
        state_var_NS = COMP_LOOP_C_116;
      end
      COMP_LOOP_C_116 : begin
        fsm_output = 10'b0011000100;
        state_var_NS = COMP_LOOP_C_117;
      end
      COMP_LOOP_C_117 : begin
        fsm_output = 10'b0011000101;
        state_var_NS = COMP_LOOP_C_118;
      end
      COMP_LOOP_C_118 : begin
        fsm_output = 10'b0011000110;
        state_var_NS = COMP_LOOP_C_119;
      end
      COMP_LOOP_C_119 : begin
        fsm_output = 10'b0011000111;
        state_var_NS = COMP_LOOP_C_120;
      end
      COMP_LOOP_C_120 : begin
        fsm_output = 10'b0011001000;
        state_var_NS = COMP_LOOP_C_121;
      end
      COMP_LOOP_C_121 : begin
        fsm_output = 10'b0011001001;
        state_var_NS = COMP_LOOP_C_122;
      end
      COMP_LOOP_C_122 : begin
        fsm_output = 10'b0011001010;
        state_var_NS = COMP_LOOP_C_123;
      end
      COMP_LOOP_C_123 : begin
        fsm_output = 10'b0011001011;
        state_var_NS = COMP_LOOP_C_124;
      end
      COMP_LOOP_C_124 : begin
        fsm_output = 10'b0011001100;
        state_var_NS = COMP_LOOP_C_125;
      end
      COMP_LOOP_C_125 : begin
        fsm_output = 10'b0011001101;
        state_var_NS = COMP_LOOP_C_126;
      end
      COMP_LOOP_C_126 : begin
        fsm_output = 10'b0011001110;
        state_var_NS = COMP_LOOP_C_127;
      end
      COMP_LOOP_C_127 : begin
        fsm_output = 10'b0011001111;
        state_var_NS = COMP_LOOP_C_128;
      end
      COMP_LOOP_C_128 : begin
        fsm_output = 10'b0011010000;
        if ( COMP_LOOP_C_128_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_129;
        end
      end
      COMP_LOOP_C_129 : begin
        fsm_output = 10'b0011010001;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0011010010;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0011010011;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0011010100;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0011010101;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0011010110;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0011010111;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0011011000;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0011011001;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0011011010;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0011011011;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0011011100;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0011011101;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_12;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_12 : begin
        fsm_output = 10'b0011011110;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_13;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_13 : begin
        fsm_output = 10'b0011011111;
        state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_14;
      end
      COMP_LOOP_5_modExp_dev_1_while_C_14 : begin
        fsm_output = 10'b0011100000;
        if ( COMP_LOOP_5_modExp_dev_1_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_130;
        end
        else begin
          state_var_NS = COMP_LOOP_5_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_130 : begin
        fsm_output = 10'b0011100001;
        state_var_NS = COMP_LOOP_C_131;
      end
      COMP_LOOP_C_131 : begin
        fsm_output = 10'b0011100010;
        state_var_NS = COMP_LOOP_C_132;
      end
      COMP_LOOP_C_132 : begin
        fsm_output = 10'b0011100011;
        state_var_NS = COMP_LOOP_C_133;
      end
      COMP_LOOP_C_133 : begin
        fsm_output = 10'b0011100100;
        state_var_NS = COMP_LOOP_C_134;
      end
      COMP_LOOP_C_134 : begin
        fsm_output = 10'b0011100101;
        state_var_NS = COMP_LOOP_C_135;
      end
      COMP_LOOP_C_135 : begin
        fsm_output = 10'b0011100110;
        state_var_NS = COMP_LOOP_C_136;
      end
      COMP_LOOP_C_136 : begin
        fsm_output = 10'b0011100111;
        state_var_NS = COMP_LOOP_C_137;
      end
      COMP_LOOP_C_137 : begin
        fsm_output = 10'b0011101000;
        state_var_NS = COMP_LOOP_C_138;
      end
      COMP_LOOP_C_138 : begin
        fsm_output = 10'b0011101001;
        state_var_NS = COMP_LOOP_C_139;
      end
      COMP_LOOP_C_139 : begin
        fsm_output = 10'b0011101010;
        state_var_NS = COMP_LOOP_C_140;
      end
      COMP_LOOP_C_140 : begin
        fsm_output = 10'b0011101011;
        state_var_NS = COMP_LOOP_C_141;
      end
      COMP_LOOP_C_141 : begin
        fsm_output = 10'b0011101100;
        state_var_NS = COMP_LOOP_C_142;
      end
      COMP_LOOP_C_142 : begin
        fsm_output = 10'b0011101101;
        state_var_NS = COMP_LOOP_C_143;
      end
      COMP_LOOP_C_143 : begin
        fsm_output = 10'b0011101110;
        state_var_NS = COMP_LOOP_C_144;
      end
      COMP_LOOP_C_144 : begin
        fsm_output = 10'b0011101111;
        state_var_NS = COMP_LOOP_C_145;
      end
      COMP_LOOP_C_145 : begin
        fsm_output = 10'b0011110000;
        state_var_NS = COMP_LOOP_C_146;
      end
      COMP_LOOP_C_146 : begin
        fsm_output = 10'b0011110001;
        state_var_NS = COMP_LOOP_C_147;
      end
      COMP_LOOP_C_147 : begin
        fsm_output = 10'b0011110010;
        state_var_NS = COMP_LOOP_C_148;
      end
      COMP_LOOP_C_148 : begin
        fsm_output = 10'b0011110011;
        state_var_NS = COMP_LOOP_C_149;
      end
      COMP_LOOP_C_149 : begin
        fsm_output = 10'b0011110100;
        state_var_NS = COMP_LOOP_C_150;
      end
      COMP_LOOP_C_150 : begin
        fsm_output = 10'b0011110101;
        state_var_NS = COMP_LOOP_C_151;
      end
      COMP_LOOP_C_151 : begin
        fsm_output = 10'b0011110110;
        state_var_NS = COMP_LOOP_C_152;
      end
      COMP_LOOP_C_152 : begin
        fsm_output = 10'b0011110111;
        state_var_NS = COMP_LOOP_C_153;
      end
      COMP_LOOP_C_153 : begin
        fsm_output = 10'b0011111000;
        state_var_NS = COMP_LOOP_C_154;
      end
      COMP_LOOP_C_154 : begin
        fsm_output = 10'b0011111001;
        state_var_NS = COMP_LOOP_C_155;
      end
      COMP_LOOP_C_155 : begin
        fsm_output = 10'b0011111010;
        state_var_NS = COMP_LOOP_C_156;
      end
      COMP_LOOP_C_156 : begin
        fsm_output = 10'b0011111011;
        state_var_NS = COMP_LOOP_C_157;
      end
      COMP_LOOP_C_157 : begin
        fsm_output = 10'b0011111100;
        state_var_NS = COMP_LOOP_C_158;
      end
      COMP_LOOP_C_158 : begin
        fsm_output = 10'b0011111101;
        state_var_NS = COMP_LOOP_C_159;
      end
      COMP_LOOP_C_159 : begin
        fsm_output = 10'b0011111110;
        state_var_NS = COMP_LOOP_C_160;
      end
      COMP_LOOP_C_160 : begin
        fsm_output = 10'b0011111111;
        if ( COMP_LOOP_C_160_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_161;
        end
      end
      COMP_LOOP_C_161 : begin
        fsm_output = 10'b0100000000;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0100000001;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0100000010;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0100000011;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0100000100;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0100000101;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0100000110;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0100000111;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0100001000;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0100001001;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0100001010;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0100001011;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0100001100;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_12;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_12 : begin
        fsm_output = 10'b0100001101;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_13;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_13 : begin
        fsm_output = 10'b0100001110;
        state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_14;
      end
      COMP_LOOP_6_modExp_dev_1_while_C_14 : begin
        fsm_output = 10'b0100001111;
        if ( COMP_LOOP_6_modExp_dev_1_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_162;
        end
        else begin
          state_var_NS = COMP_LOOP_6_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_162 : begin
        fsm_output = 10'b0100010000;
        state_var_NS = COMP_LOOP_C_163;
      end
      COMP_LOOP_C_163 : begin
        fsm_output = 10'b0100010001;
        state_var_NS = COMP_LOOP_C_164;
      end
      COMP_LOOP_C_164 : begin
        fsm_output = 10'b0100010010;
        state_var_NS = COMP_LOOP_C_165;
      end
      COMP_LOOP_C_165 : begin
        fsm_output = 10'b0100010011;
        state_var_NS = COMP_LOOP_C_166;
      end
      COMP_LOOP_C_166 : begin
        fsm_output = 10'b0100010100;
        state_var_NS = COMP_LOOP_C_167;
      end
      COMP_LOOP_C_167 : begin
        fsm_output = 10'b0100010101;
        state_var_NS = COMP_LOOP_C_168;
      end
      COMP_LOOP_C_168 : begin
        fsm_output = 10'b0100010110;
        state_var_NS = COMP_LOOP_C_169;
      end
      COMP_LOOP_C_169 : begin
        fsm_output = 10'b0100010111;
        state_var_NS = COMP_LOOP_C_170;
      end
      COMP_LOOP_C_170 : begin
        fsm_output = 10'b0100011000;
        state_var_NS = COMP_LOOP_C_171;
      end
      COMP_LOOP_C_171 : begin
        fsm_output = 10'b0100011001;
        state_var_NS = COMP_LOOP_C_172;
      end
      COMP_LOOP_C_172 : begin
        fsm_output = 10'b0100011010;
        state_var_NS = COMP_LOOP_C_173;
      end
      COMP_LOOP_C_173 : begin
        fsm_output = 10'b0100011011;
        state_var_NS = COMP_LOOP_C_174;
      end
      COMP_LOOP_C_174 : begin
        fsm_output = 10'b0100011100;
        state_var_NS = COMP_LOOP_C_175;
      end
      COMP_LOOP_C_175 : begin
        fsm_output = 10'b0100011101;
        state_var_NS = COMP_LOOP_C_176;
      end
      COMP_LOOP_C_176 : begin
        fsm_output = 10'b0100011110;
        state_var_NS = COMP_LOOP_C_177;
      end
      COMP_LOOP_C_177 : begin
        fsm_output = 10'b0100011111;
        state_var_NS = COMP_LOOP_C_178;
      end
      COMP_LOOP_C_178 : begin
        fsm_output = 10'b0100100000;
        state_var_NS = COMP_LOOP_C_179;
      end
      COMP_LOOP_C_179 : begin
        fsm_output = 10'b0100100001;
        state_var_NS = COMP_LOOP_C_180;
      end
      COMP_LOOP_C_180 : begin
        fsm_output = 10'b0100100010;
        state_var_NS = COMP_LOOP_C_181;
      end
      COMP_LOOP_C_181 : begin
        fsm_output = 10'b0100100011;
        state_var_NS = COMP_LOOP_C_182;
      end
      COMP_LOOP_C_182 : begin
        fsm_output = 10'b0100100100;
        state_var_NS = COMP_LOOP_C_183;
      end
      COMP_LOOP_C_183 : begin
        fsm_output = 10'b0100100101;
        state_var_NS = COMP_LOOP_C_184;
      end
      COMP_LOOP_C_184 : begin
        fsm_output = 10'b0100100110;
        state_var_NS = COMP_LOOP_C_185;
      end
      COMP_LOOP_C_185 : begin
        fsm_output = 10'b0100100111;
        state_var_NS = COMP_LOOP_C_186;
      end
      COMP_LOOP_C_186 : begin
        fsm_output = 10'b0100101000;
        state_var_NS = COMP_LOOP_C_187;
      end
      COMP_LOOP_C_187 : begin
        fsm_output = 10'b0100101001;
        state_var_NS = COMP_LOOP_C_188;
      end
      COMP_LOOP_C_188 : begin
        fsm_output = 10'b0100101010;
        state_var_NS = COMP_LOOP_C_189;
      end
      COMP_LOOP_C_189 : begin
        fsm_output = 10'b0100101011;
        state_var_NS = COMP_LOOP_C_190;
      end
      COMP_LOOP_C_190 : begin
        fsm_output = 10'b0100101100;
        state_var_NS = COMP_LOOP_C_191;
      end
      COMP_LOOP_C_191 : begin
        fsm_output = 10'b0100101101;
        state_var_NS = COMP_LOOP_C_192;
      end
      COMP_LOOP_C_192 : begin
        fsm_output = 10'b0100101110;
        if ( COMP_LOOP_C_192_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_193;
        end
      end
      COMP_LOOP_C_193 : begin
        fsm_output = 10'b0100101111;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0100110000;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0100110001;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0100110010;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0100110011;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0100110100;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0100110101;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0100110110;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0100110111;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0100111000;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0100111001;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0100111010;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0100111011;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_12;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_12 : begin
        fsm_output = 10'b0100111100;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_13;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_13 : begin
        fsm_output = 10'b0100111101;
        state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_14;
      end
      COMP_LOOP_7_modExp_dev_1_while_C_14 : begin
        fsm_output = 10'b0100111110;
        if ( COMP_LOOP_7_modExp_dev_1_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_194;
        end
        else begin
          state_var_NS = COMP_LOOP_7_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_194 : begin
        fsm_output = 10'b0100111111;
        state_var_NS = COMP_LOOP_C_195;
      end
      COMP_LOOP_C_195 : begin
        fsm_output = 10'b0101000000;
        state_var_NS = COMP_LOOP_C_196;
      end
      COMP_LOOP_C_196 : begin
        fsm_output = 10'b0101000001;
        state_var_NS = COMP_LOOP_C_197;
      end
      COMP_LOOP_C_197 : begin
        fsm_output = 10'b0101000010;
        state_var_NS = COMP_LOOP_C_198;
      end
      COMP_LOOP_C_198 : begin
        fsm_output = 10'b0101000011;
        state_var_NS = COMP_LOOP_C_199;
      end
      COMP_LOOP_C_199 : begin
        fsm_output = 10'b0101000100;
        state_var_NS = COMP_LOOP_C_200;
      end
      COMP_LOOP_C_200 : begin
        fsm_output = 10'b0101000101;
        state_var_NS = COMP_LOOP_C_201;
      end
      COMP_LOOP_C_201 : begin
        fsm_output = 10'b0101000110;
        state_var_NS = COMP_LOOP_C_202;
      end
      COMP_LOOP_C_202 : begin
        fsm_output = 10'b0101000111;
        state_var_NS = COMP_LOOP_C_203;
      end
      COMP_LOOP_C_203 : begin
        fsm_output = 10'b0101001000;
        state_var_NS = COMP_LOOP_C_204;
      end
      COMP_LOOP_C_204 : begin
        fsm_output = 10'b0101001001;
        state_var_NS = COMP_LOOP_C_205;
      end
      COMP_LOOP_C_205 : begin
        fsm_output = 10'b0101001010;
        state_var_NS = COMP_LOOP_C_206;
      end
      COMP_LOOP_C_206 : begin
        fsm_output = 10'b0101001011;
        state_var_NS = COMP_LOOP_C_207;
      end
      COMP_LOOP_C_207 : begin
        fsm_output = 10'b0101001100;
        state_var_NS = COMP_LOOP_C_208;
      end
      COMP_LOOP_C_208 : begin
        fsm_output = 10'b0101001101;
        state_var_NS = COMP_LOOP_C_209;
      end
      COMP_LOOP_C_209 : begin
        fsm_output = 10'b0101001110;
        state_var_NS = COMP_LOOP_C_210;
      end
      COMP_LOOP_C_210 : begin
        fsm_output = 10'b0101001111;
        state_var_NS = COMP_LOOP_C_211;
      end
      COMP_LOOP_C_211 : begin
        fsm_output = 10'b0101010000;
        state_var_NS = COMP_LOOP_C_212;
      end
      COMP_LOOP_C_212 : begin
        fsm_output = 10'b0101010001;
        state_var_NS = COMP_LOOP_C_213;
      end
      COMP_LOOP_C_213 : begin
        fsm_output = 10'b0101010010;
        state_var_NS = COMP_LOOP_C_214;
      end
      COMP_LOOP_C_214 : begin
        fsm_output = 10'b0101010011;
        state_var_NS = COMP_LOOP_C_215;
      end
      COMP_LOOP_C_215 : begin
        fsm_output = 10'b0101010100;
        state_var_NS = COMP_LOOP_C_216;
      end
      COMP_LOOP_C_216 : begin
        fsm_output = 10'b0101010101;
        state_var_NS = COMP_LOOP_C_217;
      end
      COMP_LOOP_C_217 : begin
        fsm_output = 10'b0101010110;
        state_var_NS = COMP_LOOP_C_218;
      end
      COMP_LOOP_C_218 : begin
        fsm_output = 10'b0101010111;
        state_var_NS = COMP_LOOP_C_219;
      end
      COMP_LOOP_C_219 : begin
        fsm_output = 10'b0101011000;
        state_var_NS = COMP_LOOP_C_220;
      end
      COMP_LOOP_C_220 : begin
        fsm_output = 10'b0101011001;
        state_var_NS = COMP_LOOP_C_221;
      end
      COMP_LOOP_C_221 : begin
        fsm_output = 10'b0101011010;
        state_var_NS = COMP_LOOP_C_222;
      end
      COMP_LOOP_C_222 : begin
        fsm_output = 10'b0101011011;
        state_var_NS = COMP_LOOP_C_223;
      end
      COMP_LOOP_C_223 : begin
        fsm_output = 10'b0101011100;
        state_var_NS = COMP_LOOP_C_224;
      end
      COMP_LOOP_C_224 : begin
        fsm_output = 10'b0101011101;
        if ( COMP_LOOP_C_224_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_225;
        end
      end
      COMP_LOOP_C_225 : begin
        fsm_output = 10'b0101011110;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0101011111;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0101100000;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0101100001;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0101100010;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0101100011;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0101100100;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0101100101;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0101100110;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0101100111;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0101101000;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0101101001;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0101101010;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_12;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_12 : begin
        fsm_output = 10'b0101101011;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_13;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_13 : begin
        fsm_output = 10'b0101101100;
        state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_14;
      end
      COMP_LOOP_8_modExp_dev_1_while_C_14 : begin
        fsm_output = 10'b0101101101;
        if ( COMP_LOOP_8_modExp_dev_1_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_226;
        end
        else begin
          state_var_NS = COMP_LOOP_8_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_226 : begin
        fsm_output = 10'b0101101110;
        state_var_NS = COMP_LOOP_C_227;
      end
      COMP_LOOP_C_227 : begin
        fsm_output = 10'b0101101111;
        state_var_NS = COMP_LOOP_C_228;
      end
      COMP_LOOP_C_228 : begin
        fsm_output = 10'b0101110000;
        state_var_NS = COMP_LOOP_C_229;
      end
      COMP_LOOP_C_229 : begin
        fsm_output = 10'b0101110001;
        state_var_NS = COMP_LOOP_C_230;
      end
      COMP_LOOP_C_230 : begin
        fsm_output = 10'b0101110010;
        state_var_NS = COMP_LOOP_C_231;
      end
      COMP_LOOP_C_231 : begin
        fsm_output = 10'b0101110011;
        state_var_NS = COMP_LOOP_C_232;
      end
      COMP_LOOP_C_232 : begin
        fsm_output = 10'b0101110100;
        state_var_NS = COMP_LOOP_C_233;
      end
      COMP_LOOP_C_233 : begin
        fsm_output = 10'b0101110101;
        state_var_NS = COMP_LOOP_C_234;
      end
      COMP_LOOP_C_234 : begin
        fsm_output = 10'b0101110110;
        state_var_NS = COMP_LOOP_C_235;
      end
      COMP_LOOP_C_235 : begin
        fsm_output = 10'b0101110111;
        state_var_NS = COMP_LOOP_C_236;
      end
      COMP_LOOP_C_236 : begin
        fsm_output = 10'b0101111000;
        state_var_NS = COMP_LOOP_C_237;
      end
      COMP_LOOP_C_237 : begin
        fsm_output = 10'b0101111001;
        state_var_NS = COMP_LOOP_C_238;
      end
      COMP_LOOP_C_238 : begin
        fsm_output = 10'b0101111010;
        state_var_NS = COMP_LOOP_C_239;
      end
      COMP_LOOP_C_239 : begin
        fsm_output = 10'b0101111011;
        state_var_NS = COMP_LOOP_C_240;
      end
      COMP_LOOP_C_240 : begin
        fsm_output = 10'b0101111100;
        state_var_NS = COMP_LOOP_C_241;
      end
      COMP_LOOP_C_241 : begin
        fsm_output = 10'b0101111101;
        state_var_NS = COMP_LOOP_C_242;
      end
      COMP_LOOP_C_242 : begin
        fsm_output = 10'b0101111110;
        state_var_NS = COMP_LOOP_C_243;
      end
      COMP_LOOP_C_243 : begin
        fsm_output = 10'b0101111111;
        state_var_NS = COMP_LOOP_C_244;
      end
      COMP_LOOP_C_244 : begin
        fsm_output = 10'b0110000000;
        state_var_NS = COMP_LOOP_C_245;
      end
      COMP_LOOP_C_245 : begin
        fsm_output = 10'b0110000001;
        state_var_NS = COMP_LOOP_C_246;
      end
      COMP_LOOP_C_246 : begin
        fsm_output = 10'b0110000010;
        state_var_NS = COMP_LOOP_C_247;
      end
      COMP_LOOP_C_247 : begin
        fsm_output = 10'b0110000011;
        state_var_NS = COMP_LOOP_C_248;
      end
      COMP_LOOP_C_248 : begin
        fsm_output = 10'b0110000100;
        state_var_NS = COMP_LOOP_C_249;
      end
      COMP_LOOP_C_249 : begin
        fsm_output = 10'b0110000101;
        state_var_NS = COMP_LOOP_C_250;
      end
      COMP_LOOP_C_250 : begin
        fsm_output = 10'b0110000110;
        state_var_NS = COMP_LOOP_C_251;
      end
      COMP_LOOP_C_251 : begin
        fsm_output = 10'b0110000111;
        state_var_NS = COMP_LOOP_C_252;
      end
      COMP_LOOP_C_252 : begin
        fsm_output = 10'b0110001000;
        state_var_NS = COMP_LOOP_C_253;
      end
      COMP_LOOP_C_253 : begin
        fsm_output = 10'b0110001001;
        state_var_NS = COMP_LOOP_C_254;
      end
      COMP_LOOP_C_254 : begin
        fsm_output = 10'b0110001010;
        state_var_NS = COMP_LOOP_C_255;
      end
      COMP_LOOP_C_255 : begin
        fsm_output = 10'b0110001011;
        state_var_NS = COMP_LOOP_C_256;
      end
      COMP_LOOP_C_256 : begin
        fsm_output = 10'b0110001100;
        if ( COMP_LOOP_C_256_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_257;
        end
      end
      COMP_LOOP_C_257 : begin
        fsm_output = 10'b0110001101;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0110001110;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0110001111;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0110010000;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0110010001;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0110010010;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0110010011;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0110010100;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0110010101;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0110010110;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0110010111;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0110011000;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0110011001;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_12;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_12 : begin
        fsm_output = 10'b0110011010;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_13;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_13 : begin
        fsm_output = 10'b0110011011;
        state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_14;
      end
      COMP_LOOP_9_modExp_dev_1_while_C_14 : begin
        fsm_output = 10'b0110011100;
        if ( COMP_LOOP_9_modExp_dev_1_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_258;
        end
        else begin
          state_var_NS = COMP_LOOP_9_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_258 : begin
        fsm_output = 10'b0110011101;
        state_var_NS = COMP_LOOP_C_259;
      end
      COMP_LOOP_C_259 : begin
        fsm_output = 10'b0110011110;
        state_var_NS = COMP_LOOP_C_260;
      end
      COMP_LOOP_C_260 : begin
        fsm_output = 10'b0110011111;
        state_var_NS = COMP_LOOP_C_261;
      end
      COMP_LOOP_C_261 : begin
        fsm_output = 10'b0110100000;
        state_var_NS = COMP_LOOP_C_262;
      end
      COMP_LOOP_C_262 : begin
        fsm_output = 10'b0110100001;
        state_var_NS = COMP_LOOP_C_263;
      end
      COMP_LOOP_C_263 : begin
        fsm_output = 10'b0110100010;
        state_var_NS = COMP_LOOP_C_264;
      end
      COMP_LOOP_C_264 : begin
        fsm_output = 10'b0110100011;
        state_var_NS = COMP_LOOP_C_265;
      end
      COMP_LOOP_C_265 : begin
        fsm_output = 10'b0110100100;
        state_var_NS = COMP_LOOP_C_266;
      end
      COMP_LOOP_C_266 : begin
        fsm_output = 10'b0110100101;
        state_var_NS = COMP_LOOP_C_267;
      end
      COMP_LOOP_C_267 : begin
        fsm_output = 10'b0110100110;
        state_var_NS = COMP_LOOP_C_268;
      end
      COMP_LOOP_C_268 : begin
        fsm_output = 10'b0110100111;
        state_var_NS = COMP_LOOP_C_269;
      end
      COMP_LOOP_C_269 : begin
        fsm_output = 10'b0110101000;
        state_var_NS = COMP_LOOP_C_270;
      end
      COMP_LOOP_C_270 : begin
        fsm_output = 10'b0110101001;
        state_var_NS = COMP_LOOP_C_271;
      end
      COMP_LOOP_C_271 : begin
        fsm_output = 10'b0110101010;
        state_var_NS = COMP_LOOP_C_272;
      end
      COMP_LOOP_C_272 : begin
        fsm_output = 10'b0110101011;
        state_var_NS = COMP_LOOP_C_273;
      end
      COMP_LOOP_C_273 : begin
        fsm_output = 10'b0110101100;
        state_var_NS = COMP_LOOP_C_274;
      end
      COMP_LOOP_C_274 : begin
        fsm_output = 10'b0110101101;
        state_var_NS = COMP_LOOP_C_275;
      end
      COMP_LOOP_C_275 : begin
        fsm_output = 10'b0110101110;
        state_var_NS = COMP_LOOP_C_276;
      end
      COMP_LOOP_C_276 : begin
        fsm_output = 10'b0110101111;
        state_var_NS = COMP_LOOP_C_277;
      end
      COMP_LOOP_C_277 : begin
        fsm_output = 10'b0110110000;
        state_var_NS = COMP_LOOP_C_278;
      end
      COMP_LOOP_C_278 : begin
        fsm_output = 10'b0110110001;
        state_var_NS = COMP_LOOP_C_279;
      end
      COMP_LOOP_C_279 : begin
        fsm_output = 10'b0110110010;
        state_var_NS = COMP_LOOP_C_280;
      end
      COMP_LOOP_C_280 : begin
        fsm_output = 10'b0110110011;
        state_var_NS = COMP_LOOP_C_281;
      end
      COMP_LOOP_C_281 : begin
        fsm_output = 10'b0110110100;
        state_var_NS = COMP_LOOP_C_282;
      end
      COMP_LOOP_C_282 : begin
        fsm_output = 10'b0110110101;
        state_var_NS = COMP_LOOP_C_283;
      end
      COMP_LOOP_C_283 : begin
        fsm_output = 10'b0110110110;
        state_var_NS = COMP_LOOP_C_284;
      end
      COMP_LOOP_C_284 : begin
        fsm_output = 10'b0110110111;
        state_var_NS = COMP_LOOP_C_285;
      end
      COMP_LOOP_C_285 : begin
        fsm_output = 10'b0110111000;
        state_var_NS = COMP_LOOP_C_286;
      end
      COMP_LOOP_C_286 : begin
        fsm_output = 10'b0110111001;
        state_var_NS = COMP_LOOP_C_287;
      end
      COMP_LOOP_C_287 : begin
        fsm_output = 10'b0110111010;
        state_var_NS = COMP_LOOP_C_288;
      end
      COMP_LOOP_C_288 : begin
        fsm_output = 10'b0110111011;
        if ( COMP_LOOP_C_288_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_289;
        end
      end
      COMP_LOOP_C_289 : begin
        fsm_output = 10'b0110111100;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0110111101;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0110111110;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0110111111;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0111000000;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0111000001;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0111000010;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0111000011;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0111000100;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0111000101;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0111000110;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0111000111;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0111001000;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_12;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_12 : begin
        fsm_output = 10'b0111001001;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_13;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_13 : begin
        fsm_output = 10'b0111001010;
        state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_14;
      end
      COMP_LOOP_10_modExp_dev_1_while_C_14 : begin
        fsm_output = 10'b0111001011;
        if ( COMP_LOOP_10_modExp_dev_1_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_290;
        end
        else begin
          state_var_NS = COMP_LOOP_10_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_290 : begin
        fsm_output = 10'b0111001100;
        state_var_NS = COMP_LOOP_C_291;
      end
      COMP_LOOP_C_291 : begin
        fsm_output = 10'b0111001101;
        state_var_NS = COMP_LOOP_C_292;
      end
      COMP_LOOP_C_292 : begin
        fsm_output = 10'b0111001110;
        state_var_NS = COMP_LOOP_C_293;
      end
      COMP_LOOP_C_293 : begin
        fsm_output = 10'b0111001111;
        state_var_NS = COMP_LOOP_C_294;
      end
      COMP_LOOP_C_294 : begin
        fsm_output = 10'b0111010000;
        state_var_NS = COMP_LOOP_C_295;
      end
      COMP_LOOP_C_295 : begin
        fsm_output = 10'b0111010001;
        state_var_NS = COMP_LOOP_C_296;
      end
      COMP_LOOP_C_296 : begin
        fsm_output = 10'b0111010010;
        state_var_NS = COMP_LOOP_C_297;
      end
      COMP_LOOP_C_297 : begin
        fsm_output = 10'b0111010011;
        state_var_NS = COMP_LOOP_C_298;
      end
      COMP_LOOP_C_298 : begin
        fsm_output = 10'b0111010100;
        state_var_NS = COMP_LOOP_C_299;
      end
      COMP_LOOP_C_299 : begin
        fsm_output = 10'b0111010101;
        state_var_NS = COMP_LOOP_C_300;
      end
      COMP_LOOP_C_300 : begin
        fsm_output = 10'b0111010110;
        state_var_NS = COMP_LOOP_C_301;
      end
      COMP_LOOP_C_301 : begin
        fsm_output = 10'b0111010111;
        state_var_NS = COMP_LOOP_C_302;
      end
      COMP_LOOP_C_302 : begin
        fsm_output = 10'b0111011000;
        state_var_NS = COMP_LOOP_C_303;
      end
      COMP_LOOP_C_303 : begin
        fsm_output = 10'b0111011001;
        state_var_NS = COMP_LOOP_C_304;
      end
      COMP_LOOP_C_304 : begin
        fsm_output = 10'b0111011010;
        state_var_NS = COMP_LOOP_C_305;
      end
      COMP_LOOP_C_305 : begin
        fsm_output = 10'b0111011011;
        state_var_NS = COMP_LOOP_C_306;
      end
      COMP_LOOP_C_306 : begin
        fsm_output = 10'b0111011100;
        state_var_NS = COMP_LOOP_C_307;
      end
      COMP_LOOP_C_307 : begin
        fsm_output = 10'b0111011101;
        state_var_NS = COMP_LOOP_C_308;
      end
      COMP_LOOP_C_308 : begin
        fsm_output = 10'b0111011110;
        state_var_NS = COMP_LOOP_C_309;
      end
      COMP_LOOP_C_309 : begin
        fsm_output = 10'b0111011111;
        state_var_NS = COMP_LOOP_C_310;
      end
      COMP_LOOP_C_310 : begin
        fsm_output = 10'b0111100000;
        state_var_NS = COMP_LOOP_C_311;
      end
      COMP_LOOP_C_311 : begin
        fsm_output = 10'b0111100001;
        state_var_NS = COMP_LOOP_C_312;
      end
      COMP_LOOP_C_312 : begin
        fsm_output = 10'b0111100010;
        state_var_NS = COMP_LOOP_C_313;
      end
      COMP_LOOP_C_313 : begin
        fsm_output = 10'b0111100011;
        state_var_NS = COMP_LOOP_C_314;
      end
      COMP_LOOP_C_314 : begin
        fsm_output = 10'b0111100100;
        state_var_NS = COMP_LOOP_C_315;
      end
      COMP_LOOP_C_315 : begin
        fsm_output = 10'b0111100101;
        state_var_NS = COMP_LOOP_C_316;
      end
      COMP_LOOP_C_316 : begin
        fsm_output = 10'b0111100110;
        state_var_NS = COMP_LOOP_C_317;
      end
      COMP_LOOP_C_317 : begin
        fsm_output = 10'b0111100111;
        state_var_NS = COMP_LOOP_C_318;
      end
      COMP_LOOP_C_318 : begin
        fsm_output = 10'b0111101000;
        state_var_NS = COMP_LOOP_C_319;
      end
      COMP_LOOP_C_319 : begin
        fsm_output = 10'b0111101001;
        state_var_NS = COMP_LOOP_C_320;
      end
      COMP_LOOP_C_320 : begin
        fsm_output = 10'b0111101010;
        if ( COMP_LOOP_C_320_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_321;
        end
      end
      COMP_LOOP_C_321 : begin
        fsm_output = 10'b0111101011;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b0111101100;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b0111101101;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b0111101110;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b0111101111;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b0111110000;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b0111110001;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b0111110010;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b0111110011;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b0111110100;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b0111110101;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b0111110110;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b0111110111;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_12;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_12 : begin
        fsm_output = 10'b0111111000;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_13;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_13 : begin
        fsm_output = 10'b0111111001;
        state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_14;
      end
      COMP_LOOP_11_modExp_dev_1_while_C_14 : begin
        fsm_output = 10'b0111111010;
        if ( COMP_LOOP_11_modExp_dev_1_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_322;
        end
        else begin
          state_var_NS = COMP_LOOP_11_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_322 : begin
        fsm_output = 10'b0111111011;
        state_var_NS = COMP_LOOP_C_323;
      end
      COMP_LOOP_C_323 : begin
        fsm_output = 10'b0111111100;
        state_var_NS = COMP_LOOP_C_324;
      end
      COMP_LOOP_C_324 : begin
        fsm_output = 10'b0111111101;
        state_var_NS = COMP_LOOP_C_325;
      end
      COMP_LOOP_C_325 : begin
        fsm_output = 10'b0111111110;
        state_var_NS = COMP_LOOP_C_326;
      end
      COMP_LOOP_C_326 : begin
        fsm_output = 10'b0111111111;
        state_var_NS = COMP_LOOP_C_327;
      end
      COMP_LOOP_C_327 : begin
        fsm_output = 10'b1000000000;
        state_var_NS = COMP_LOOP_C_328;
      end
      COMP_LOOP_C_328 : begin
        fsm_output = 10'b1000000001;
        state_var_NS = COMP_LOOP_C_329;
      end
      COMP_LOOP_C_329 : begin
        fsm_output = 10'b1000000010;
        state_var_NS = COMP_LOOP_C_330;
      end
      COMP_LOOP_C_330 : begin
        fsm_output = 10'b1000000011;
        state_var_NS = COMP_LOOP_C_331;
      end
      COMP_LOOP_C_331 : begin
        fsm_output = 10'b1000000100;
        state_var_NS = COMP_LOOP_C_332;
      end
      COMP_LOOP_C_332 : begin
        fsm_output = 10'b1000000101;
        state_var_NS = COMP_LOOP_C_333;
      end
      COMP_LOOP_C_333 : begin
        fsm_output = 10'b1000000110;
        state_var_NS = COMP_LOOP_C_334;
      end
      COMP_LOOP_C_334 : begin
        fsm_output = 10'b1000000111;
        state_var_NS = COMP_LOOP_C_335;
      end
      COMP_LOOP_C_335 : begin
        fsm_output = 10'b1000001000;
        state_var_NS = COMP_LOOP_C_336;
      end
      COMP_LOOP_C_336 : begin
        fsm_output = 10'b1000001001;
        state_var_NS = COMP_LOOP_C_337;
      end
      COMP_LOOP_C_337 : begin
        fsm_output = 10'b1000001010;
        state_var_NS = COMP_LOOP_C_338;
      end
      COMP_LOOP_C_338 : begin
        fsm_output = 10'b1000001011;
        state_var_NS = COMP_LOOP_C_339;
      end
      COMP_LOOP_C_339 : begin
        fsm_output = 10'b1000001100;
        state_var_NS = COMP_LOOP_C_340;
      end
      COMP_LOOP_C_340 : begin
        fsm_output = 10'b1000001101;
        state_var_NS = COMP_LOOP_C_341;
      end
      COMP_LOOP_C_341 : begin
        fsm_output = 10'b1000001110;
        state_var_NS = COMP_LOOP_C_342;
      end
      COMP_LOOP_C_342 : begin
        fsm_output = 10'b1000001111;
        state_var_NS = COMP_LOOP_C_343;
      end
      COMP_LOOP_C_343 : begin
        fsm_output = 10'b1000010000;
        state_var_NS = COMP_LOOP_C_344;
      end
      COMP_LOOP_C_344 : begin
        fsm_output = 10'b1000010001;
        state_var_NS = COMP_LOOP_C_345;
      end
      COMP_LOOP_C_345 : begin
        fsm_output = 10'b1000010010;
        state_var_NS = COMP_LOOP_C_346;
      end
      COMP_LOOP_C_346 : begin
        fsm_output = 10'b1000010011;
        state_var_NS = COMP_LOOP_C_347;
      end
      COMP_LOOP_C_347 : begin
        fsm_output = 10'b1000010100;
        state_var_NS = COMP_LOOP_C_348;
      end
      COMP_LOOP_C_348 : begin
        fsm_output = 10'b1000010101;
        state_var_NS = COMP_LOOP_C_349;
      end
      COMP_LOOP_C_349 : begin
        fsm_output = 10'b1000010110;
        state_var_NS = COMP_LOOP_C_350;
      end
      COMP_LOOP_C_350 : begin
        fsm_output = 10'b1000010111;
        state_var_NS = COMP_LOOP_C_351;
      end
      COMP_LOOP_C_351 : begin
        fsm_output = 10'b1000011000;
        state_var_NS = COMP_LOOP_C_352;
      end
      COMP_LOOP_C_352 : begin
        fsm_output = 10'b1000011001;
        if ( COMP_LOOP_C_352_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_353;
        end
      end
      COMP_LOOP_C_353 : begin
        fsm_output = 10'b1000011010;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b1000011011;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b1000011100;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b1000011101;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b1000011110;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b1000011111;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b1000100000;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b1000100001;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b1000100010;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b1000100011;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b1000100100;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b1000100101;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b1000100110;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_12;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_12 : begin
        fsm_output = 10'b1000100111;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_13;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_13 : begin
        fsm_output = 10'b1000101000;
        state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_14;
      end
      COMP_LOOP_12_modExp_dev_1_while_C_14 : begin
        fsm_output = 10'b1000101001;
        if ( COMP_LOOP_12_modExp_dev_1_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_354;
        end
        else begin
          state_var_NS = COMP_LOOP_12_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_354 : begin
        fsm_output = 10'b1000101010;
        state_var_NS = COMP_LOOP_C_355;
      end
      COMP_LOOP_C_355 : begin
        fsm_output = 10'b1000101011;
        state_var_NS = COMP_LOOP_C_356;
      end
      COMP_LOOP_C_356 : begin
        fsm_output = 10'b1000101100;
        state_var_NS = COMP_LOOP_C_357;
      end
      COMP_LOOP_C_357 : begin
        fsm_output = 10'b1000101101;
        state_var_NS = COMP_LOOP_C_358;
      end
      COMP_LOOP_C_358 : begin
        fsm_output = 10'b1000101110;
        state_var_NS = COMP_LOOP_C_359;
      end
      COMP_LOOP_C_359 : begin
        fsm_output = 10'b1000101111;
        state_var_NS = COMP_LOOP_C_360;
      end
      COMP_LOOP_C_360 : begin
        fsm_output = 10'b1000110000;
        state_var_NS = COMP_LOOP_C_361;
      end
      COMP_LOOP_C_361 : begin
        fsm_output = 10'b1000110001;
        state_var_NS = COMP_LOOP_C_362;
      end
      COMP_LOOP_C_362 : begin
        fsm_output = 10'b1000110010;
        state_var_NS = COMP_LOOP_C_363;
      end
      COMP_LOOP_C_363 : begin
        fsm_output = 10'b1000110011;
        state_var_NS = COMP_LOOP_C_364;
      end
      COMP_LOOP_C_364 : begin
        fsm_output = 10'b1000110100;
        state_var_NS = COMP_LOOP_C_365;
      end
      COMP_LOOP_C_365 : begin
        fsm_output = 10'b1000110101;
        state_var_NS = COMP_LOOP_C_366;
      end
      COMP_LOOP_C_366 : begin
        fsm_output = 10'b1000110110;
        state_var_NS = COMP_LOOP_C_367;
      end
      COMP_LOOP_C_367 : begin
        fsm_output = 10'b1000110111;
        state_var_NS = COMP_LOOP_C_368;
      end
      COMP_LOOP_C_368 : begin
        fsm_output = 10'b1000111000;
        state_var_NS = COMP_LOOP_C_369;
      end
      COMP_LOOP_C_369 : begin
        fsm_output = 10'b1000111001;
        state_var_NS = COMP_LOOP_C_370;
      end
      COMP_LOOP_C_370 : begin
        fsm_output = 10'b1000111010;
        state_var_NS = COMP_LOOP_C_371;
      end
      COMP_LOOP_C_371 : begin
        fsm_output = 10'b1000111011;
        state_var_NS = COMP_LOOP_C_372;
      end
      COMP_LOOP_C_372 : begin
        fsm_output = 10'b1000111100;
        state_var_NS = COMP_LOOP_C_373;
      end
      COMP_LOOP_C_373 : begin
        fsm_output = 10'b1000111101;
        state_var_NS = COMP_LOOP_C_374;
      end
      COMP_LOOP_C_374 : begin
        fsm_output = 10'b1000111110;
        state_var_NS = COMP_LOOP_C_375;
      end
      COMP_LOOP_C_375 : begin
        fsm_output = 10'b1000111111;
        state_var_NS = COMP_LOOP_C_376;
      end
      COMP_LOOP_C_376 : begin
        fsm_output = 10'b1001000000;
        state_var_NS = COMP_LOOP_C_377;
      end
      COMP_LOOP_C_377 : begin
        fsm_output = 10'b1001000001;
        state_var_NS = COMP_LOOP_C_378;
      end
      COMP_LOOP_C_378 : begin
        fsm_output = 10'b1001000010;
        state_var_NS = COMP_LOOP_C_379;
      end
      COMP_LOOP_C_379 : begin
        fsm_output = 10'b1001000011;
        state_var_NS = COMP_LOOP_C_380;
      end
      COMP_LOOP_C_380 : begin
        fsm_output = 10'b1001000100;
        state_var_NS = COMP_LOOP_C_381;
      end
      COMP_LOOP_C_381 : begin
        fsm_output = 10'b1001000101;
        state_var_NS = COMP_LOOP_C_382;
      end
      COMP_LOOP_C_382 : begin
        fsm_output = 10'b1001000110;
        state_var_NS = COMP_LOOP_C_383;
      end
      COMP_LOOP_C_383 : begin
        fsm_output = 10'b1001000111;
        state_var_NS = COMP_LOOP_C_384;
      end
      COMP_LOOP_C_384 : begin
        fsm_output = 10'b1001001000;
        if ( COMP_LOOP_C_384_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_385;
        end
      end
      COMP_LOOP_C_385 : begin
        fsm_output = 10'b1001001001;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b1001001010;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b1001001011;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b1001001100;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b1001001101;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b1001001110;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b1001001111;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b1001010000;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b1001010001;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b1001010010;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b1001010011;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b1001010100;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b1001010101;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_12;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_12 : begin
        fsm_output = 10'b1001010110;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_13;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_13 : begin
        fsm_output = 10'b1001010111;
        state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_14;
      end
      COMP_LOOP_13_modExp_dev_1_while_C_14 : begin
        fsm_output = 10'b1001011000;
        if ( COMP_LOOP_13_modExp_dev_1_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_386;
        end
        else begin
          state_var_NS = COMP_LOOP_13_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_386 : begin
        fsm_output = 10'b1001011001;
        state_var_NS = COMP_LOOP_C_387;
      end
      COMP_LOOP_C_387 : begin
        fsm_output = 10'b1001011010;
        state_var_NS = COMP_LOOP_C_388;
      end
      COMP_LOOP_C_388 : begin
        fsm_output = 10'b1001011011;
        state_var_NS = COMP_LOOP_C_389;
      end
      COMP_LOOP_C_389 : begin
        fsm_output = 10'b1001011100;
        state_var_NS = COMP_LOOP_C_390;
      end
      COMP_LOOP_C_390 : begin
        fsm_output = 10'b1001011101;
        state_var_NS = COMP_LOOP_C_391;
      end
      COMP_LOOP_C_391 : begin
        fsm_output = 10'b1001011110;
        state_var_NS = COMP_LOOP_C_392;
      end
      COMP_LOOP_C_392 : begin
        fsm_output = 10'b1001011111;
        state_var_NS = COMP_LOOP_C_393;
      end
      COMP_LOOP_C_393 : begin
        fsm_output = 10'b1001100000;
        state_var_NS = COMP_LOOP_C_394;
      end
      COMP_LOOP_C_394 : begin
        fsm_output = 10'b1001100001;
        state_var_NS = COMP_LOOP_C_395;
      end
      COMP_LOOP_C_395 : begin
        fsm_output = 10'b1001100010;
        state_var_NS = COMP_LOOP_C_396;
      end
      COMP_LOOP_C_396 : begin
        fsm_output = 10'b1001100011;
        state_var_NS = COMP_LOOP_C_397;
      end
      COMP_LOOP_C_397 : begin
        fsm_output = 10'b1001100100;
        state_var_NS = COMP_LOOP_C_398;
      end
      COMP_LOOP_C_398 : begin
        fsm_output = 10'b1001100101;
        state_var_NS = COMP_LOOP_C_399;
      end
      COMP_LOOP_C_399 : begin
        fsm_output = 10'b1001100110;
        state_var_NS = COMP_LOOP_C_400;
      end
      COMP_LOOP_C_400 : begin
        fsm_output = 10'b1001100111;
        state_var_NS = COMP_LOOP_C_401;
      end
      COMP_LOOP_C_401 : begin
        fsm_output = 10'b1001101000;
        state_var_NS = COMP_LOOP_C_402;
      end
      COMP_LOOP_C_402 : begin
        fsm_output = 10'b1001101001;
        state_var_NS = COMP_LOOP_C_403;
      end
      COMP_LOOP_C_403 : begin
        fsm_output = 10'b1001101010;
        state_var_NS = COMP_LOOP_C_404;
      end
      COMP_LOOP_C_404 : begin
        fsm_output = 10'b1001101011;
        state_var_NS = COMP_LOOP_C_405;
      end
      COMP_LOOP_C_405 : begin
        fsm_output = 10'b1001101100;
        state_var_NS = COMP_LOOP_C_406;
      end
      COMP_LOOP_C_406 : begin
        fsm_output = 10'b1001101101;
        state_var_NS = COMP_LOOP_C_407;
      end
      COMP_LOOP_C_407 : begin
        fsm_output = 10'b1001101110;
        state_var_NS = COMP_LOOP_C_408;
      end
      COMP_LOOP_C_408 : begin
        fsm_output = 10'b1001101111;
        state_var_NS = COMP_LOOP_C_409;
      end
      COMP_LOOP_C_409 : begin
        fsm_output = 10'b1001110000;
        state_var_NS = COMP_LOOP_C_410;
      end
      COMP_LOOP_C_410 : begin
        fsm_output = 10'b1001110001;
        state_var_NS = COMP_LOOP_C_411;
      end
      COMP_LOOP_C_411 : begin
        fsm_output = 10'b1001110010;
        state_var_NS = COMP_LOOP_C_412;
      end
      COMP_LOOP_C_412 : begin
        fsm_output = 10'b1001110011;
        state_var_NS = COMP_LOOP_C_413;
      end
      COMP_LOOP_C_413 : begin
        fsm_output = 10'b1001110100;
        state_var_NS = COMP_LOOP_C_414;
      end
      COMP_LOOP_C_414 : begin
        fsm_output = 10'b1001110101;
        state_var_NS = COMP_LOOP_C_415;
      end
      COMP_LOOP_C_415 : begin
        fsm_output = 10'b1001110110;
        state_var_NS = COMP_LOOP_C_416;
      end
      COMP_LOOP_C_416 : begin
        fsm_output = 10'b1001110111;
        if ( COMP_LOOP_C_416_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_417;
        end
      end
      COMP_LOOP_C_417 : begin
        fsm_output = 10'b1001111000;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b1001111001;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b1001111010;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b1001111011;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b1001111100;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b1001111101;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b1001111110;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b1001111111;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b1010000000;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b1010000001;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b1010000010;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b1010000011;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b1010000100;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_12;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_12 : begin
        fsm_output = 10'b1010000101;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_13;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_13 : begin
        fsm_output = 10'b1010000110;
        state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_14;
      end
      COMP_LOOP_14_modExp_dev_1_while_C_14 : begin
        fsm_output = 10'b1010000111;
        if ( COMP_LOOP_14_modExp_dev_1_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_418;
        end
        else begin
          state_var_NS = COMP_LOOP_14_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_418 : begin
        fsm_output = 10'b1010001000;
        state_var_NS = COMP_LOOP_C_419;
      end
      COMP_LOOP_C_419 : begin
        fsm_output = 10'b1010001001;
        state_var_NS = COMP_LOOP_C_420;
      end
      COMP_LOOP_C_420 : begin
        fsm_output = 10'b1010001010;
        state_var_NS = COMP_LOOP_C_421;
      end
      COMP_LOOP_C_421 : begin
        fsm_output = 10'b1010001011;
        state_var_NS = COMP_LOOP_C_422;
      end
      COMP_LOOP_C_422 : begin
        fsm_output = 10'b1010001100;
        state_var_NS = COMP_LOOP_C_423;
      end
      COMP_LOOP_C_423 : begin
        fsm_output = 10'b1010001101;
        state_var_NS = COMP_LOOP_C_424;
      end
      COMP_LOOP_C_424 : begin
        fsm_output = 10'b1010001110;
        state_var_NS = COMP_LOOP_C_425;
      end
      COMP_LOOP_C_425 : begin
        fsm_output = 10'b1010001111;
        state_var_NS = COMP_LOOP_C_426;
      end
      COMP_LOOP_C_426 : begin
        fsm_output = 10'b1010010000;
        state_var_NS = COMP_LOOP_C_427;
      end
      COMP_LOOP_C_427 : begin
        fsm_output = 10'b1010010001;
        state_var_NS = COMP_LOOP_C_428;
      end
      COMP_LOOP_C_428 : begin
        fsm_output = 10'b1010010010;
        state_var_NS = COMP_LOOP_C_429;
      end
      COMP_LOOP_C_429 : begin
        fsm_output = 10'b1010010011;
        state_var_NS = COMP_LOOP_C_430;
      end
      COMP_LOOP_C_430 : begin
        fsm_output = 10'b1010010100;
        state_var_NS = COMP_LOOP_C_431;
      end
      COMP_LOOP_C_431 : begin
        fsm_output = 10'b1010010101;
        state_var_NS = COMP_LOOP_C_432;
      end
      COMP_LOOP_C_432 : begin
        fsm_output = 10'b1010010110;
        state_var_NS = COMP_LOOP_C_433;
      end
      COMP_LOOP_C_433 : begin
        fsm_output = 10'b1010010111;
        state_var_NS = COMP_LOOP_C_434;
      end
      COMP_LOOP_C_434 : begin
        fsm_output = 10'b1010011000;
        state_var_NS = COMP_LOOP_C_435;
      end
      COMP_LOOP_C_435 : begin
        fsm_output = 10'b1010011001;
        state_var_NS = COMP_LOOP_C_436;
      end
      COMP_LOOP_C_436 : begin
        fsm_output = 10'b1010011010;
        state_var_NS = COMP_LOOP_C_437;
      end
      COMP_LOOP_C_437 : begin
        fsm_output = 10'b1010011011;
        state_var_NS = COMP_LOOP_C_438;
      end
      COMP_LOOP_C_438 : begin
        fsm_output = 10'b1010011100;
        state_var_NS = COMP_LOOP_C_439;
      end
      COMP_LOOP_C_439 : begin
        fsm_output = 10'b1010011101;
        state_var_NS = COMP_LOOP_C_440;
      end
      COMP_LOOP_C_440 : begin
        fsm_output = 10'b1010011110;
        state_var_NS = COMP_LOOP_C_441;
      end
      COMP_LOOP_C_441 : begin
        fsm_output = 10'b1010011111;
        state_var_NS = COMP_LOOP_C_442;
      end
      COMP_LOOP_C_442 : begin
        fsm_output = 10'b1010100000;
        state_var_NS = COMP_LOOP_C_443;
      end
      COMP_LOOP_C_443 : begin
        fsm_output = 10'b1010100001;
        state_var_NS = COMP_LOOP_C_444;
      end
      COMP_LOOP_C_444 : begin
        fsm_output = 10'b1010100010;
        state_var_NS = COMP_LOOP_C_445;
      end
      COMP_LOOP_C_445 : begin
        fsm_output = 10'b1010100011;
        state_var_NS = COMP_LOOP_C_446;
      end
      COMP_LOOP_C_446 : begin
        fsm_output = 10'b1010100100;
        state_var_NS = COMP_LOOP_C_447;
      end
      COMP_LOOP_C_447 : begin
        fsm_output = 10'b1010100101;
        state_var_NS = COMP_LOOP_C_448;
      end
      COMP_LOOP_C_448 : begin
        fsm_output = 10'b1010100110;
        if ( COMP_LOOP_C_448_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_449;
        end
      end
      COMP_LOOP_C_449 : begin
        fsm_output = 10'b1010100111;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b1010101000;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b1010101001;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b1010101010;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b1010101011;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b1010101100;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b1010101101;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b1010101110;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b1010101111;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b1010110000;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b1010110001;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b1010110010;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b1010110011;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_12;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_12 : begin
        fsm_output = 10'b1010110100;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_13;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_13 : begin
        fsm_output = 10'b1010110101;
        state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_14;
      end
      COMP_LOOP_15_modExp_dev_1_while_C_14 : begin
        fsm_output = 10'b1010110110;
        if ( COMP_LOOP_15_modExp_dev_1_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_450;
        end
        else begin
          state_var_NS = COMP_LOOP_15_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_450 : begin
        fsm_output = 10'b1010110111;
        state_var_NS = COMP_LOOP_C_451;
      end
      COMP_LOOP_C_451 : begin
        fsm_output = 10'b1010111000;
        state_var_NS = COMP_LOOP_C_452;
      end
      COMP_LOOP_C_452 : begin
        fsm_output = 10'b1010111001;
        state_var_NS = COMP_LOOP_C_453;
      end
      COMP_LOOP_C_453 : begin
        fsm_output = 10'b1010111010;
        state_var_NS = COMP_LOOP_C_454;
      end
      COMP_LOOP_C_454 : begin
        fsm_output = 10'b1010111011;
        state_var_NS = COMP_LOOP_C_455;
      end
      COMP_LOOP_C_455 : begin
        fsm_output = 10'b1010111100;
        state_var_NS = COMP_LOOP_C_456;
      end
      COMP_LOOP_C_456 : begin
        fsm_output = 10'b1010111101;
        state_var_NS = COMP_LOOP_C_457;
      end
      COMP_LOOP_C_457 : begin
        fsm_output = 10'b1010111110;
        state_var_NS = COMP_LOOP_C_458;
      end
      COMP_LOOP_C_458 : begin
        fsm_output = 10'b1010111111;
        state_var_NS = COMP_LOOP_C_459;
      end
      COMP_LOOP_C_459 : begin
        fsm_output = 10'b1011000000;
        state_var_NS = COMP_LOOP_C_460;
      end
      COMP_LOOP_C_460 : begin
        fsm_output = 10'b1011000001;
        state_var_NS = COMP_LOOP_C_461;
      end
      COMP_LOOP_C_461 : begin
        fsm_output = 10'b1011000010;
        state_var_NS = COMP_LOOP_C_462;
      end
      COMP_LOOP_C_462 : begin
        fsm_output = 10'b1011000011;
        state_var_NS = COMP_LOOP_C_463;
      end
      COMP_LOOP_C_463 : begin
        fsm_output = 10'b1011000100;
        state_var_NS = COMP_LOOP_C_464;
      end
      COMP_LOOP_C_464 : begin
        fsm_output = 10'b1011000101;
        state_var_NS = COMP_LOOP_C_465;
      end
      COMP_LOOP_C_465 : begin
        fsm_output = 10'b1011000110;
        state_var_NS = COMP_LOOP_C_466;
      end
      COMP_LOOP_C_466 : begin
        fsm_output = 10'b1011000111;
        state_var_NS = COMP_LOOP_C_467;
      end
      COMP_LOOP_C_467 : begin
        fsm_output = 10'b1011001000;
        state_var_NS = COMP_LOOP_C_468;
      end
      COMP_LOOP_C_468 : begin
        fsm_output = 10'b1011001001;
        state_var_NS = COMP_LOOP_C_469;
      end
      COMP_LOOP_C_469 : begin
        fsm_output = 10'b1011001010;
        state_var_NS = COMP_LOOP_C_470;
      end
      COMP_LOOP_C_470 : begin
        fsm_output = 10'b1011001011;
        state_var_NS = COMP_LOOP_C_471;
      end
      COMP_LOOP_C_471 : begin
        fsm_output = 10'b1011001100;
        state_var_NS = COMP_LOOP_C_472;
      end
      COMP_LOOP_C_472 : begin
        fsm_output = 10'b1011001101;
        state_var_NS = COMP_LOOP_C_473;
      end
      COMP_LOOP_C_473 : begin
        fsm_output = 10'b1011001110;
        state_var_NS = COMP_LOOP_C_474;
      end
      COMP_LOOP_C_474 : begin
        fsm_output = 10'b1011001111;
        state_var_NS = COMP_LOOP_C_475;
      end
      COMP_LOOP_C_475 : begin
        fsm_output = 10'b1011010000;
        state_var_NS = COMP_LOOP_C_476;
      end
      COMP_LOOP_C_476 : begin
        fsm_output = 10'b1011010001;
        state_var_NS = COMP_LOOP_C_477;
      end
      COMP_LOOP_C_477 : begin
        fsm_output = 10'b1011010010;
        state_var_NS = COMP_LOOP_C_478;
      end
      COMP_LOOP_C_478 : begin
        fsm_output = 10'b1011010011;
        state_var_NS = COMP_LOOP_C_479;
      end
      COMP_LOOP_C_479 : begin
        fsm_output = 10'b1011010100;
        state_var_NS = COMP_LOOP_C_480;
      end
      COMP_LOOP_C_480 : begin
        fsm_output = 10'b1011010101;
        if ( COMP_LOOP_C_480_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_481;
        end
      end
      COMP_LOOP_C_481 : begin
        fsm_output = 10'b1011010110;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_0;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_0 : begin
        fsm_output = 10'b1011010111;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_1;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_1 : begin
        fsm_output = 10'b1011011000;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_2;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_2 : begin
        fsm_output = 10'b1011011001;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_3;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_3 : begin
        fsm_output = 10'b1011011010;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_4;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_4 : begin
        fsm_output = 10'b1011011011;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_5;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_5 : begin
        fsm_output = 10'b1011011100;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_6;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_6 : begin
        fsm_output = 10'b1011011101;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_7;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_7 : begin
        fsm_output = 10'b1011011110;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_8;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_8 : begin
        fsm_output = 10'b1011011111;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_9;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_9 : begin
        fsm_output = 10'b1011100000;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_10;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_10 : begin
        fsm_output = 10'b1011100001;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_11;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_11 : begin
        fsm_output = 10'b1011100010;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_12;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_12 : begin
        fsm_output = 10'b1011100011;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_13;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_13 : begin
        fsm_output = 10'b1011100100;
        state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_14;
      end
      COMP_LOOP_16_modExp_dev_1_while_C_14 : begin
        fsm_output = 10'b1011100101;
        if ( COMP_LOOP_16_modExp_dev_1_while_C_14_tr0 ) begin
          state_var_NS = COMP_LOOP_C_482;
        end
        else begin
          state_var_NS = COMP_LOOP_16_modExp_dev_1_while_C_0;
        end
      end
      COMP_LOOP_C_482 : begin
        fsm_output = 10'b1011100110;
        state_var_NS = COMP_LOOP_C_483;
      end
      COMP_LOOP_C_483 : begin
        fsm_output = 10'b1011100111;
        state_var_NS = COMP_LOOP_C_484;
      end
      COMP_LOOP_C_484 : begin
        fsm_output = 10'b1011101000;
        state_var_NS = COMP_LOOP_C_485;
      end
      COMP_LOOP_C_485 : begin
        fsm_output = 10'b1011101001;
        state_var_NS = COMP_LOOP_C_486;
      end
      COMP_LOOP_C_486 : begin
        fsm_output = 10'b1011101010;
        state_var_NS = COMP_LOOP_C_487;
      end
      COMP_LOOP_C_487 : begin
        fsm_output = 10'b1011101011;
        state_var_NS = COMP_LOOP_C_488;
      end
      COMP_LOOP_C_488 : begin
        fsm_output = 10'b1011101100;
        state_var_NS = COMP_LOOP_C_489;
      end
      COMP_LOOP_C_489 : begin
        fsm_output = 10'b1011101101;
        state_var_NS = COMP_LOOP_C_490;
      end
      COMP_LOOP_C_490 : begin
        fsm_output = 10'b1011101110;
        state_var_NS = COMP_LOOP_C_491;
      end
      COMP_LOOP_C_491 : begin
        fsm_output = 10'b1011101111;
        state_var_NS = COMP_LOOP_C_492;
      end
      COMP_LOOP_C_492 : begin
        fsm_output = 10'b1011110000;
        state_var_NS = COMP_LOOP_C_493;
      end
      COMP_LOOP_C_493 : begin
        fsm_output = 10'b1011110001;
        state_var_NS = COMP_LOOP_C_494;
      end
      COMP_LOOP_C_494 : begin
        fsm_output = 10'b1011110010;
        state_var_NS = COMP_LOOP_C_495;
      end
      COMP_LOOP_C_495 : begin
        fsm_output = 10'b1011110011;
        state_var_NS = COMP_LOOP_C_496;
      end
      COMP_LOOP_C_496 : begin
        fsm_output = 10'b1011110100;
        state_var_NS = COMP_LOOP_C_497;
      end
      COMP_LOOP_C_497 : begin
        fsm_output = 10'b1011110101;
        state_var_NS = COMP_LOOP_C_498;
      end
      COMP_LOOP_C_498 : begin
        fsm_output = 10'b1011110110;
        state_var_NS = COMP_LOOP_C_499;
      end
      COMP_LOOP_C_499 : begin
        fsm_output = 10'b1011110111;
        state_var_NS = COMP_LOOP_C_500;
      end
      COMP_LOOP_C_500 : begin
        fsm_output = 10'b1011111000;
        state_var_NS = COMP_LOOP_C_501;
      end
      COMP_LOOP_C_501 : begin
        fsm_output = 10'b1011111001;
        state_var_NS = COMP_LOOP_C_502;
      end
      COMP_LOOP_C_502 : begin
        fsm_output = 10'b1011111010;
        state_var_NS = COMP_LOOP_C_503;
      end
      COMP_LOOP_C_503 : begin
        fsm_output = 10'b1011111011;
        state_var_NS = COMP_LOOP_C_504;
      end
      COMP_LOOP_C_504 : begin
        fsm_output = 10'b1011111100;
        state_var_NS = COMP_LOOP_C_505;
      end
      COMP_LOOP_C_505 : begin
        fsm_output = 10'b1011111101;
        state_var_NS = COMP_LOOP_C_506;
      end
      COMP_LOOP_C_506 : begin
        fsm_output = 10'b1011111110;
        state_var_NS = COMP_LOOP_C_507;
      end
      COMP_LOOP_C_507 : begin
        fsm_output = 10'b1011111111;
        state_var_NS = COMP_LOOP_C_508;
      end
      COMP_LOOP_C_508 : begin
        fsm_output = 10'b1100000000;
        state_var_NS = COMP_LOOP_C_509;
      end
      COMP_LOOP_C_509 : begin
        fsm_output = 10'b1100000001;
        state_var_NS = COMP_LOOP_C_510;
      end
      COMP_LOOP_C_510 : begin
        fsm_output = 10'b1100000010;
        state_var_NS = COMP_LOOP_C_511;
      end
      COMP_LOOP_C_511 : begin
        fsm_output = 10'b1100000011;
        state_var_NS = COMP_LOOP_C_512;
      end
      COMP_LOOP_C_512 : begin
        fsm_output = 10'b1100000100;
        if ( COMP_LOOP_C_512_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_C_0 : begin
        fsm_output = 10'b1100000101;
        if ( VEC_LOOP_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_4;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      STAGE_LOOP_C_4 : begin
        fsm_output = 10'b1100000110;
        if ( STAGE_LOOP_C_4_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = STAGE_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 10'b1100000111;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 10'b0000000000;
        state_var_NS = STAGE_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core_wait_dp
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core_wait_dp (
  ensig_cgo_iro, ensig_cgo, modulo_dev_cmp_ccs_ccore_en
);
  input ensig_cgo_iro;
  input ensig_cgo;
  output modulo_dev_cmp_ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  assign modulo_dev_cmp_ccs_ccore_en = ensig_cgo | ensig_cgo_iro;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core (
  clk, rst, vec_rsc_triosy_0_0_lz, vec_rsc_triosy_0_1_lz, vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz, vec_rsc_triosy_0_4_lz, vec_rsc_triosy_0_5_lz, vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz, vec_rsc_triosy_0_8_lz, vec_rsc_triosy_0_9_lz, vec_rsc_triosy_0_10_lz,
      vec_rsc_triosy_0_11_lz, vec_rsc_triosy_0_12_lz, vec_rsc_triosy_0_13_lz, vec_rsc_triosy_0_14_lz,
      vec_rsc_triosy_0_15_lz, p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz,
      vec_rsc_0_0_i_q_d, vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_1_i_q_d,
      vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_2_i_q_d, vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_q_d, vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_4_i_q_d,
      vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_5_i_q_d, vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_q_d, vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_7_i_q_d,
      vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_8_i_q_d, vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_9_i_q_d, vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_10_i_q_d,
      vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_11_i_q_d, vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_12_i_q_d, vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_13_i_q_d,
      vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_14_i_q_d, vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_15_i_q_d, vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_0_i_d_d_pff,
      vec_rsc_0_0_i_radr_d_pff, vec_rsc_0_0_i_wadr_d_pff, vec_rsc_0_0_i_we_d_pff,
      vec_rsc_0_1_i_we_d_pff, vec_rsc_0_2_i_we_d_pff, vec_rsc_0_3_i_we_d_pff, vec_rsc_0_4_i_we_d_pff,
      vec_rsc_0_5_i_we_d_pff, vec_rsc_0_6_i_we_d_pff, vec_rsc_0_7_i_we_d_pff, vec_rsc_0_8_i_we_d_pff,
      vec_rsc_0_9_i_we_d_pff, vec_rsc_0_10_i_we_d_pff, vec_rsc_0_11_i_we_d_pff, vec_rsc_0_12_i_we_d_pff,
      vec_rsc_0_13_i_we_d_pff, vec_rsc_0_14_i_we_d_pff, vec_rsc_0_15_i_we_d_pff
);
  input clk;
  input rst;
  output vec_rsc_triosy_0_0_lz;
  output vec_rsc_triosy_0_1_lz;
  output vec_rsc_triosy_0_2_lz;
  output vec_rsc_triosy_0_3_lz;
  output vec_rsc_triosy_0_4_lz;
  output vec_rsc_triosy_0_5_lz;
  output vec_rsc_triosy_0_6_lz;
  output vec_rsc_triosy_0_7_lz;
  output vec_rsc_triosy_0_8_lz;
  output vec_rsc_triosy_0_9_lz;
  output vec_rsc_triosy_0_10_lz;
  output vec_rsc_triosy_0_11_lz;
  output vec_rsc_triosy_0_12_lz;
  output vec_rsc_triosy_0_13_lz;
  output vec_rsc_triosy_0_14_lz;
  output vec_rsc_triosy_0_15_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  input [63:0] vec_rsc_0_0_i_q_d;
  output vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_1_i_q_d;
  output vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_2_i_q_d;
  output vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_3_i_q_d;
  output vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_4_i_q_d;
  output vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_5_i_q_d;
  output vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_6_i_q_d;
  output vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_7_i_q_d;
  output vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_8_i_q_d;
  output vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_9_i_q_d;
  output vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_10_i_q_d;
  output vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_11_i_q_d;
  output vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_12_i_q_d;
  output vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_13_i_q_d;
  output vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_14_i_q_d;
  output vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_15_i_q_d;
  output vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d;
  output [63:0] vec_rsc_0_0_i_d_d_pff;
  output [5:0] vec_rsc_0_0_i_radr_d_pff;
  output [5:0] vec_rsc_0_0_i_wadr_d_pff;
  output vec_rsc_0_0_i_we_d_pff;
  output vec_rsc_0_1_i_we_d_pff;
  output vec_rsc_0_2_i_we_d_pff;
  output vec_rsc_0_3_i_we_d_pff;
  output vec_rsc_0_4_i_we_d_pff;
  output vec_rsc_0_5_i_we_d_pff;
  output vec_rsc_0_6_i_we_d_pff;
  output vec_rsc_0_7_i_we_d_pff;
  output vec_rsc_0_8_i_we_d_pff;
  output vec_rsc_0_9_i_we_d_pff;
  output vec_rsc_0_10_i_we_d_pff;
  output vec_rsc_0_11_i_we_d_pff;
  output vec_rsc_0_12_i_we_d_pff;
  output vec_rsc_0_13_i_we_d_pff;
  output vec_rsc_0_14_i_we_d_pff;
  output vec_rsc_0_15_i_we_d_pff;


  // Interconnect Declarations
  wire [63:0] p_rsci_idat;
  wire [63:0] r_rsci_idat;
  wire [63:0] modulo_dev_cmp_return_rsc_z;
  wire modulo_dev_cmp_ccs_ccore_en;
  reg [64:0] operator_66_true_div_cmp_a;
  wire [64:0] operator_66_true_div_cmp_z;
  reg [9:0] operator_66_true_div_cmp_b_9_0;
  wire [9:0] fsm_output;
  wire nand_tmp;
  wire or_tmp_20;
  wire nor_tmp_14;
  wire or_tmp_74;
  wire nor_tmp_40;
  wire and_dcpl_13;
  wire and_dcpl_14;
  wire and_dcpl_15;
  wire and_dcpl_16;
  wire and_dcpl_17;
  wire and_dcpl_18;
  wire and_dcpl_19;
  wire and_dcpl_23;
  wire not_tmp_121;
  wire and_dcpl_26;
  wire and_dcpl_27;
  wire and_dcpl_28;
  wire and_dcpl_29;
  wire and_dcpl_30;
  wire and_dcpl_32;
  wire and_dcpl_33;
  wire and_dcpl_34;
  wire and_dcpl_35;
  wire and_dcpl_36;
  wire and_dcpl_37;
  wire and_dcpl_38;
  wire and_dcpl_39;
  wire and_dcpl_40;
  wire and_dcpl_42;
  wire and_dcpl_43;
  wire and_dcpl_44;
  wire and_dcpl_45;
  wire and_dcpl_47;
  wire and_dcpl_48;
  wire and_dcpl_49;
  wire and_dcpl_50;
  wire and_dcpl_51;
  wire and_dcpl_52;
  wire and_dcpl_54;
  wire and_dcpl_55;
  wire and_dcpl_57;
  wire and_dcpl_58;
  wire and_dcpl_59;
  wire and_dcpl_60;
  wire and_dcpl_61;
  wire and_dcpl_63;
  wire and_dcpl_64;
  wire and_dcpl_65;
  wire and_dcpl_66;
  wire and_dcpl_67;
  wire and_dcpl_68;
  wire and_dcpl_70;
  wire and_dcpl_71;
  wire and_dcpl_72;
  wire and_dcpl_73;
  wire and_dcpl_74;
  wire and_dcpl_75;
  wire and_dcpl_78;
  wire and_dcpl_79;
  wire and_dcpl_80;
  wire and_dcpl_81;
  wire and_dcpl_83;
  wire and_dcpl_84;
  wire and_dcpl_85;
  wire and_dcpl_86;
  wire and_dcpl_87;
  wire and_dcpl_89;
  wire and_dcpl_90;
  wire and_dcpl_91;
  wire and_dcpl_93;
  wire and_dcpl_94;
  wire and_dcpl_95;
  wire and_dcpl_97;
  wire and_dcpl_98;
  wire and_dcpl_99;
  wire and_dcpl_101;
  wire and_dcpl_102;
  wire and_dcpl_103;
  wire and_dcpl_106;
  wire and_dcpl_107;
  wire and_dcpl_108;
  wire and_dcpl_110;
  wire and_dcpl_111;
  wire and_dcpl_112;
  wire and_dcpl_115;
  wire and_dcpl_116;
  wire and_dcpl_117;
  wire and_dcpl_119;
  wire or_tmp_237;
  wire nand_tmp_6;
  wire or_tmp_239;
  wire or_tmp_241;
  wire nand_tmp_7;
  wire and_dcpl_122;
  wire and_dcpl_130;
  wire and_dcpl_132;
  wire and_dcpl_136;
  wire and_dcpl_138;
  wire or_tmp_252;
  wire or_tmp_253;
  wire or_tmp_258;
  wire or_tmp_259;
  wire not_tmp_133;
  wire not_tmp_134;
  wire or_tmp_346;
  wire or_tmp_352;
  wire or_tmp_353;
  wire or_tmp_362;
  wire or_tmp_438;
  wire or_tmp_439;
  wire or_tmp_444;
  wire or_tmp_445;
  wire or_tmp_531;
  wire or_tmp_532;
  wire or_tmp_537;
  wire or_tmp_538;
  wire or_tmp_624;
  wire or_tmp_625;
  wire or_tmp_630;
  wire or_tmp_631;
  wire or_tmp_718;
  wire or_tmp_724;
  wire or_tmp_725;
  wire or_tmp_734;
  wire or_tmp_810;
  wire or_tmp_811;
  wire or_tmp_816;
  wire or_tmp_817;
  wire or_tmp_903;
  wire or_tmp_904;
  wire or_tmp_909;
  wire or_tmp_910;
  wire or_tmp_997;
  wire or_tmp_999;
  wire or_tmp_1005;
  wire or_tmp_1007;
  wire or_tmp_1097;
  wire or_tmp_1104;
  wire or_tmp_1106;
  wire or_tmp_1116;
  wire or_tmp_1195;
  wire or_tmp_1197;
  wire or_tmp_1203;
  wire or_tmp_1205;
  wire or_tmp_1294;
  wire or_tmp_1296;
  wire or_tmp_1302;
  wire or_tmp_1304;
  wire not_tmp_289;
  wire or_tmp_1393;
  wire or_tmp_1395;
  wire or_tmp_1401;
  wire or_tmp_1403;
  wire not_tmp_304;
  wire or_tmp_1493;
  wire or_tmp_1500;
  wire or_tmp_1502;
  wire or_tmp_1512;
  wire or_tmp_1590;
  wire or_tmp_1592;
  wire or_tmp_1598;
  wire or_tmp_1600;
  wire not_tmp_335;
  wire or_tmp_1687;
  wire or_tmp_1689;
  wire not_tmp_336;
  wire or_tmp_1694;
  wire nor_tmp_186;
  wire mux_tmp_1470;
  wire mux_tmp_1471;
  wire mux_tmp_1472;
  wire mux_tmp_1473;
  wire mux_tmp_1476;
  wire nor_tmp_188;
  wire mux_tmp_1477;
  wire nor_tmp_190;
  wire mux_tmp_1482;
  wire mux_tmp_1483;
  wire mux_tmp_1484;
  wire mux_tmp_1485;
  wire mux_tmp_1488;
  wire mux_tmp_1489;
  wire mux_tmp_1496;
  wire mux_tmp_1498;
  wire mux_tmp_1501;
  wire mux_tmp_1503;
  wire mux_tmp_1514;
  wire or_tmp_1788;
  wire or_tmp_1793;
  wire or_tmp_1794;
  wire mux_tmp_1534;
  wire or_tmp_1796;
  wire mux_tmp_1537;
  wire or_tmp_1799;
  wire nand_tmp_106;
  wire not_tmp_370;
  wire or_tmp_1816;
  wire or_tmp_1818;
  wire mux_tmp_1562;
  wire mux_tmp_1563;
  wire or_tmp_1823;
  wire or_tmp_1824;
  wire mux_tmp_1566;
  wire or_tmp_1825;
  wire or_tmp_1827;
  wire or_tmp_1830;
  wire or_tmp_1831;
  wire mux_tmp_1573;
  wire or_tmp_1835;
  wire mux_tmp_1579;
  wire or_tmp_1838;
  wire or_tmp_1840;
  wire or_tmp_1841;
  wire and_dcpl_169;
  wire or_tmp_1845;
  wire and_tmp_12;
  wire mux_tmp_1610;
  wire mux_tmp_1612;
  wire or_tmp_1854;
  wire mux_tmp_1615;
  wire or_tmp_1855;
  wire mux_tmp_1618;
  wire mux_tmp_1621;
  wire mux_tmp_1623;
  wire mux_tmp_1625;
  wire mux_tmp_1626;
  wire mux_tmp_1629;
  wire mux_tmp_1688;
  wire or_tmp_1899;
  wire and_dcpl_183;
  wire not_tmp_402;
  wire nor_tmp_203;
  wire not_tmp_418;
  wire or_tmp_1989;
  wire or_tmp_1990;
  wire mux_tmp_1782;
  wire mux_tmp_1786;
  wire mux_tmp_1793;
  wire mux_tmp_1799;
  wire mux_tmp_1801;
  wire mux_tmp_1803;
  wire mux_tmp_1808;
  wire mux_tmp_1809;
  wire not_tmp_431;
  wire nor_tmp_215;
  wire not_tmp_439;
  wire mux_tmp_1839;
  wire and_dcpl_199;
  wire and_dcpl_200;
  wire and_dcpl_201;
  wire and_dcpl_202;
  wire and_dcpl_203;
  wire and_dcpl_204;
  wire and_dcpl_206;
  wire and_dcpl_207;
  wire and_dcpl_208;
  wire and_dcpl_210;
  wire and_dcpl_212;
  wire and_dcpl_214;
  wire and_dcpl_215;
  wire and_dcpl_217;
  wire and_dcpl_219;
  wire and_dcpl_220;
  wire and_dcpl_221;
  wire or_tmp_2035;
  wire mux_tmp_1861;
  wire or_tmp_2037;
  wire mux_tmp_1863;
  wire or_tmp_2040;
  wire or_tmp_2041;
  wire mux_tmp_1866;
  wire or_tmp_2043;
  wire or_tmp_2044;
  wire mux_tmp_1870;
  wire mux_tmp_1872;
  wire or_tmp_2047;
  wire mux_tmp_1874;
  wire mux_tmp_1875;
  wire nand_tmp_134;
  wire mux_tmp_1876;
  wire mux_tmp_1877;
  wire mux_tmp_1882;
  wire mux_tmp_1883;
  wire mux_tmp_1888;
  wire mux_tmp_1891;
  reg COMP_LOOP_COMP_LOOP_and_137_itm;
  reg COMP_LOOP_COMP_LOOP_and_10_itm;
  wire [10:0] VEC_LOOP_acc_1_psp_1;
  wire [11:0] nl_VEC_LOOP_acc_1_psp_1;
  reg COMP_LOOP_nor_11_itm;
  wire [7:0] COMP_LOOP_acc_13_psp_sva_1;
  wire [8:0] nl_COMP_LOOP_acc_13_psp_sva_1;
  reg [4:0] COMP_LOOP_k_9_4_sva_4_0;
  reg [9:0] VEC_LOOP_j_sva_9_0;
  reg COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  reg COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  reg [9:0] COMP_LOOP_acc_1_cse_6_sva;
  reg [7:0] COMP_LOOP_acc_13_psp_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_4_sva;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_4_sva;
  reg [8:0] COMP_LOOP_acc_11_psp_sva;
  wire [9:0] nl_COMP_LOOP_acc_11_psp_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_14_sva;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_14_sva;
  reg [7:0] COMP_LOOP_acc_19_psp_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_12_sva;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_12_sva;
  reg [8:0] COMP_LOOP_acc_17_psp_sva;
  wire [9:0] nl_COMP_LOOP_acc_17_psp_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_10_sva;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_10_sva;
  reg [6:0] COMP_LOOP_acc_16_psp_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_8_sva;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_8_sva;
  reg [8:0] COMP_LOOP_acc_14_psp_sva;
  wire [9:0] nl_COMP_LOOP_acc_14_psp_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_sva;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_sva;
  reg [8:0] COMP_LOOP_acc_20_psp_sva;
  wire [9:0] nl_COMP_LOOP_acc_20_psp_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_2_sva;
  wire [9:0] COMP_LOOP_acc_1_cse_2_sva_1;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_2_sva_1;
  wire nand_308_cse;
  wire nand_264_cse;
  reg reg_vec_rsc_triosy_0_15_obj_ld_cse;
  reg reg_ensig_cgo_cse;
  wire or_1973_cse;
  wire nor_256_cse;
  wire or_1916_cse;
  wire and_267_cse;
  wire or_2186_cse;
  wire and_418_cse;
  wire or_2040_cse;
  wire or_1982_cse;
  wire or_1967_cse;
  wire or_214_cse;
  wire nor_697_cse;
  wire or_279_cse;
  wire or_1977_cse;
  wire and_375_cse;
  wire mux_424_cse;
  wire or_212_cse;
  wire nand_321_cse;
  wire and_247_cse;
  wire or_2151_cse;
  wire and_376_cse;
  wire nor_728_cse;
  wire or_1820_cse;
  wire or_2012_cse;
  wire or_103_cse;
  wire nand_357_cse;
  wire mux_1802_cse;
  wire mux_1788_cse;
  wire mux_1797_cse;
  wire mux_461_cse;
  wire mux_460_cse;
  wire mux_1789_cse;
  wire mux_1583_cse;
  wire mux_1784_cse;
  wire or_1880_cse;
  wire nor_760_cse;
  wire mux_1602_cse;
  wire mux_1785_cse;
  wire and_259_cse;
  wire mux_1726_cse;
  wire mux_1909_cse;
  wire mux_1911_cse;
  reg [63:0] COMP_LOOP_1_mul_itm;
  wire signed [128:0] nl_COMP_LOOP_1_mul_itm;
  reg [63:0] tmp_10_lpi_4_dfm;
  reg [63:0] p_sva;
  reg [5:0] COMP_LOOP_acc_psp_sva;
  wire mux_1581_itm;
  wire mux_1832_itm;
  wire mux_1834_itm;
  wire mux_tmp_2006;
  wire and_dcpl_231;
  wire and_dcpl_232;
  wire and_dcpl_233;
  wire and_dcpl_234;
  wire and_dcpl_236;
  wire and_dcpl_237;
  wire and_dcpl_238;
  wire and_dcpl_242;
  wire and_dcpl_243;
  wire and_dcpl_244;
  wire and_dcpl_246;
  wire and_dcpl_248;
  wire and_dcpl_250;
  wire and_dcpl_251;
  wire and_dcpl_252;
  wire and_dcpl_255;
  wire and_dcpl_256;
  wire and_dcpl_260;
  wire and_dcpl_265;
  wire and_dcpl_267;
  wire and_dcpl_271;
  wire and_dcpl_272;
  wire and_dcpl_274;
  wire and_dcpl_277;
  wire and_dcpl_278;
  wire and_dcpl_279;
  wire and_dcpl_281;
  wire and_dcpl_284;
  wire [9:0] z_out_1;
  wire and_dcpl_293;
  wire and_dcpl_300;
  wire and_dcpl_308;
  wire [7:0] z_out_2;
  wire [5:0] z_out_3;
  wire [6:0] nl_z_out_3;
  wire and_dcpl_344;
  wire [5:0] z_out_4;
  wire and_dcpl_361;
  wire [6:0] z_out_5;
  wire and_dcpl_376;
  wire and_dcpl_382;
  wire and_dcpl_396;
  wire and_dcpl_398;
  wire and_dcpl_402;
  wire and_dcpl_403;
  wire and_dcpl_406;
  wire and_dcpl_407;
  wire and_dcpl_416;
  wire and_dcpl_417;
  wire and_dcpl_425;
  wire and_dcpl_444;
  wire [64:0] z_out_7;
  wire [65:0] nl_z_out_7;
  wire and_dcpl_460;
  wire and_dcpl_464;
  wire [64:0] z_out_9;
  wire [65:0] nl_z_out_9;
  reg [63:0] r_sva;
  reg [3:0] STAGE_LOOP_i_3_0_sva;
  reg [9:0] STAGE_LOOP_lshift_psp_sva;
  reg [63:0] modExp_dev_exp_sva;
  reg [63:0] modExp_dev_result_sva;
  reg COMP_LOOP_COMP_LOOP_nor_itm;
  reg COMP_LOOP_COMP_LOOP_and_2_itm;
  reg COMP_LOOP_COMP_LOOP_and_4_itm;
  reg COMP_LOOP_COMP_LOOP_and_5_itm;
  reg COMP_LOOP_COMP_LOOP_and_6_itm;
  reg COMP_LOOP_COMP_LOOP_and_8_itm;
  reg COMP_LOOP_COMP_LOOP_and_9_itm;
  reg COMP_LOOP_COMP_LOOP_and_11_itm;
  reg COMP_LOOP_COMP_LOOP_and_12_itm;
  reg COMP_LOOP_COMP_LOOP_and_13_itm;
  reg COMP_LOOP_COMP_LOOP_and_14_itm;
  reg COMP_LOOP_COMP_LOOP_nor_1_itm;
  reg COMP_LOOP_nor_12_itm;
  reg COMP_LOOP_COMP_LOOP_and_62_itm;
  reg COMP_LOOP_COMP_LOOP_and_64_itm;
  reg COMP_LOOP_COMP_LOOP_and_68_itm;
  reg COMP_LOOP_COMP_LOOP_and_139_itm;
  reg COMP_LOOP_COMP_LOOP_and_140_itm;
  reg COMP_LOOP_COMP_LOOP_and_141_itm;
  reg COMP_LOOP_COMP_LOOP_and_143_itm;
  reg COMP_LOOP_COMP_LOOP_and_144_itm;
  reg COMP_LOOP_COMP_LOOP_and_145_itm;
  reg COMP_LOOP_COMP_LOOP_and_146_itm;
  reg COMP_LOOP_COMP_LOOP_and_147_itm;
  reg COMP_LOOP_COMP_LOOP_and_148_itm;
  reg COMP_LOOP_COMP_LOOP_and_149_itm;
  reg COMP_LOOP_nor_134_itm;
  reg COMP_LOOP_nor_137_itm;
  reg COMP_LOOP_COMP_LOOP_and_244_itm;
  reg [54:0] modExp_dev_exp_1_sva_63_9;
  reg [3:0] modExp_dev_exp_1_sva_3_0;
  wire STAGE_LOOP_i_3_0_sva_mx0c1;
  wire [9:0] STAGE_LOOP_lshift_psp_sva_mx0w0;
  wire VEC_LOOP_j_sva_9_0_mx0c1;
  wire and_195_rgt;
  wire and_551_ssc;
  wire nand_270_cse_1;
  wire nand_260_cse_1;
  wire modExp_dev_while_or_2_cse;
  wire nor_678_cse;
  wire or_368_cse;
  wire or_369_cse;
  wire nor_650_cse;
  wire or_462_cse;
  wire nor_624_cse;
  wire or_554_cse;
  wire or_555_cse;
  wire nor_598_cse;
  wire or_648_cse;
  wire nor_572_cse;
  wire or_740_cse;
  wire or_741_cse;
  wire nor_544_cse;
  wire or_834_cse;
  wire nor_518_cse;
  wire or_926_cse;
  wire or_927_cse;
  wire nor_492_cse;
  wire nand_280_cse;
  wire nand_275_cse;
  wire nor_467_cse;
  wire or_1119_cse;
  wire nor_439_cse;
  wire or_1218_cse;
  wire nor_413_cse;
  wire or_1317_cse;
  wire nor_387_cse;
  wire nand_241_cse;
  wire nor_362_cse;
  wire or_1515_cse;
  wire nor_335_cse;
  wire nand_217_cse;
  wire nor_310_cse;
  wire nand_202_cse;
  wire nand_197_cse;
  wire and_291_cse;
  wire nand_161_cse;
  wire nand_160_cse;
  wire or_1995_cse;
  wire or_1976_cse;
  wire mux_1768_cse;
  wire mux_2066_cse;
  wire nand_tmp_139;
  wire or_tmp_2154;
  wire mux_tmp_2041;
  wire or_tmp_2156;
  wire mux_tmp_2043;
  wire mux_tmp_2046;
  wire or_tmp_2166;
  wire or_tmp_2168;
  wire mux_tmp_2052;
  wire or_tmp_2171;
  wire mux_tmp_2058;
  wire or_tmp_2183;
  wire mux_tmp_2072;
  wire not_tmp_571;
  wire or_tmp_2191;
  wire or_tmp_2193;
  wire mux_tmp_2081;
  wire mux_tmp_2083;
  wire [64:0] operator_64_false_operator_64_false_mux_rgt;
  wire mux_tmp_2108;
  wire or_tmp_2223;
  wire mux_tmp_2112;
  wire or_tmp_2227;
  wire mux_tmp_2119;
  wire mux_tmp_2124;
  wire mux_tmp_2128;
  wire or_tmp_2236;
  wire mux_tmp_2150;
  wire mux_tmp_2153;
  wire mux_tmp_2154;
  wire mux_tmp_2156;
  wire mux_tmp_2159;
  wire mux_tmp_2164;
  wire mux_tmp_2165;
  wire mux_tmp_2167;
  wire mux_tmp_2169;
  wire mux_tmp_2170;
  wire mux_tmp_2179;
  wire mux_tmp_2180;
  wire or_tmp_2243;
  wire or_tmp_2244;
  wire mux_tmp_2192;
  wire mux_tmp_2193;
  wire or_tmp_2245;
  wire mux_tmp_2196;
  wire mux_tmp_2199;
  wire mux_tmp_2204;
  wire [9:0] COMP_LOOP_mux1h_192_rgt;
  reg [4:0] COMP_LOOP_acc_10_cse_10_1_1_sva_9_5;
  reg [4:0] COMP_LOOP_acc_10_cse_10_1_1_sva_4_0;
  reg operator_64_false_acc_mut_64;
  reg [63:0] operator_64_false_acc_mut_63_0;
  wire or_2306_cse;
  wire or_2348_cse;
  wire or_2336_cse;
  wire nor_810_cse;
  wire or_2086_cse;
  wire or_2146_cse;
  wire and_357_cse;
  wire mux_1949_cse;
  wire mux_1920_cse;
  wire mux_1922_cse;
  wire mux_1938_cse;
  wire mux_2249_itm;
  wire [9:0] z_out_6_10_1;
  wire [62:0] z_out_8_64_2;
  wire nor_761_cse;

  wire[0:0] mux_1580_nl;
  wire[0:0] mux_1579_nl;
  wire[0:0] mux_1578_nl;
  wire[0:0] mux_1577_nl;
  wire[0:0] mux_1576_nl;
  wire[0:0] mux_1575_nl;
  wire[0:0] mux_1574_nl;
  wire[0:0] mux_1573_nl;
  wire[0:0] mux_1572_nl;
  wire[0:0] mux_1571_nl;
  wire[0:0] mux_1570_nl;
  wire[0:0] and_278_nl;
  wire[0:0] mux_1569_nl;
  wire[0:0] mux_1568_nl;
  wire[0:0] mux_1567_nl;
  wire[0:0] mux_1566_nl;
  wire[0:0] mux_1563_nl;
  wire[0:0] mux_1562_nl;
  wire[0:0] and_280_nl;
  wire[0:0] mux_1561_nl;
  wire[0:0] mux_1560_nl;
  wire[0:0] mux_1559_nl;
  wire[0:0] mux_1558_nl;
  wire[0:0] mux_1557_nl;
  wire[0:0] mux_1556_nl;
  wire[0:0] mux_1555_nl;
  wire[0:0] mux_1553_nl;
  wire[0:0] mux_1551_nl;
  wire[0:0] mux_1550_nl;
  wire[0:0] mux_1546_nl;
  wire[0:0] mux_1545_nl;
  wire[0:0] mux_1544_nl;
  wire[0:0] mux_1543_nl;
  wire[0:0] mux_1542_nl;
  wire[0:0] mux_1541_nl;
  wire[0:0] mux_1532_nl;
  wire[0:0] mux_1531_nl;
  wire[0:0] mux_1530_nl;
  wire[0:0] mux_1529_nl;
  wire[0:0] mux_1525_nl;
  wire[0:0] nor_271_nl;
  wire[0:0] or_1980_nl;
  wire[0:0] mux_1725_nl;
  wire[63:0] modExp_dev_while_mux1h_nl;
  wire[63:0] mul_nl;
  wire[127:0] nl_mul_nl;
  wire[63:0] modExp_dev_while_mux_2_nl;
  wire[63:0] modExp_dev_while_mux_3_nl;
  wire[63:0] COMP_LOOP_1_acc_8_nl;
  wire[64:0] nl_COMP_LOOP_1_acc_8_nl;
  wire[0:0] modExp_dev_while_or_1_nl;
  wire[0:0] mux_1792_nl;
  wire[0:0] mux_1791_nl;
  wire[0:0] mux_1790_nl;
  wire[0:0] and_258_nl;
  wire[0:0] nor_255_nl;
  wire[0:0] mux_1787_nl;
  wire[0:0] mux_1786_nl;
  wire[0:0] and_260_nl;
  wire[0:0] nor_257_nl;
  wire[0:0] mux_1783_nl;
  wire[0:0] mux_1698_nl;
  wire[0:0] mux_1697_nl;
  wire[0:0] mux_1696_nl;
  wire[0:0] mux_1695_nl;
  wire[0:0] mux_1694_nl;
  wire[0:0] or_1896_nl;
  wire[0:0] mux_1693_nl;
  wire[0:0] mux_1692_nl;
  wire[0:0] mux_1691_nl;
  wire[0:0] mux_1690_nl;
  wire[0:0] mux_1689_nl;
  wire[0:0] mux_1688_nl;
  wire[0:0] mux_1727_nl;
  wire[0:0] mux_1686_nl;
  wire[0:0] mux_1685_nl;
  wire[0:0] mux_1684_nl;
  wire[0:0] mux_1683_nl;
  wire[0:0] mux_1678_nl;
  wire[0:0] mux_1713_nl;
  wire[0:0] mux_1673_nl;
  wire[0:0] mux_1668_nl;
  wire[0:0] mux_1667_nl;
  wire[0:0] mux_1703_nl;
  wire[0:0] mux_1664_nl;
  wire[0:0] mux_2121_nl;
  wire[0:0] mux_2120_nl;
  wire[0:0] mux_2119_nl;
  wire[0:0] mux_2118_nl;
  wire[0:0] mux_2117_nl;
  wire[0:0] or_2287_nl;
  wire[0:0] mux_2116_nl;
  wire[0:0] or_2286_nl;
  wire[0:0] or_2284_nl;
  wire[0:0] mux_2115_nl;
  wire[0:0] mux_2114_nl;
  wire[0:0] mux_2113_nl;
  wire[0:0] or_2283_nl;
  wire[0:0] mux_2112_nl;
  wire[0:0] mux_2111_nl;
  wire[0:0] mux_2109_nl;
  wire[0:0] or_2280_nl;
  wire[0:0] mux_2108_nl;
  wire[0:0] mux_2107_nl;
  wire[0:0] mux_2106_nl;
  wire[0:0] mux_2105_nl;
  wire[0:0] nand_390_nl;
  wire[0:0] mux_2100_nl;
  wire[0:0] mux_2099_nl;
  wire[0:0] mux_2096_nl;
  wire[0:0] or_2265_nl;
  wire[0:0] mux_2094_nl;
  wire[0:0] mux_nl;
  wire[0:0] or_2258_nl;
  wire[0:0] mux_2153_nl;
  wire[0:0] mux_2152_nl;
  wire[0:0] mux_2151_nl;
  wire[0:0] mux_2150_nl;
  wire[0:0] mux_2149_nl;
  wire[0:0] or_2310_nl;
  wire[0:0] or_2309_nl;
  wire[0:0] mux_2148_nl;
  wire[0:0] mux_2147_nl;
  wire[0:0] mux_2146_nl;
  wire[0:0] or_2308_nl;
  wire[0:0] mux_2145_nl;
  wire[0:0] mux_2144_nl;
  wire[0:0] mux_2143_nl;
  wire[0:0] mux_2142_nl;
  wire[0:0] or_2305_nl;
  wire[0:0] mux_2141_nl;
  wire[0:0] nand_392_nl;
  wire[0:0] or_2304_nl;
  wire[0:0] mux_2140_nl;
  wire[0:0] mux_2139_nl;
  wire[0:0] mux_2138_nl;
  wire[0:0] mux_2137_nl;
  wire[0:0] mux_2136_nl;
  wire[0:0] or_2303_nl;
  wire[0:0] mux_2130_nl;
  wire[0:0] mux_2129_nl;
  wire[0:0] mux_2128_nl;
  wire[0:0] mux_2127_nl;
  wire[0:0] mux_2126_nl;
  wire[0:0] or_2367_nl;
  wire[0:0] or_2292_nl;
  wire[0:0] or_nl;
  wire[0:0] mux_1740_nl;
  wire[0:0] or_1923_nl;
  wire[0:0] or_1922_nl;
  wire[0:0] mux_2156_nl;
  wire[0:0] or_2365_nl;
  wire[0:0] mux_2155_nl;
  wire[0:0] or_2316_nl;
  wire[0:0] mux_2154_nl;
  wire[0:0] or_2315_nl;
  wire[0:0] or_2313_nl;
  wire[0:0] or_2366_nl;
  wire[0:0] mux_1749_nl;
  wire[0:0] nor_269_nl;
  wire[0:0] mux_1748_nl;
  wire[0:0] mux_1747_nl;
  wire[0:0] mux_1754_nl;
  wire[0:0] mux_1753_nl;
  wire[0:0] mux_1752_nl;
  wire[0:0] or_1936_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_17_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_10_nl;
  wire[9:0] COMP_LOOP_1_acc_nl;
  wire[10:0] nl_COMP_LOOP_1_acc_nl;
  wire[0:0] mux_1842_nl;
  wire[0:0] mux_1841_nl;
  wire[0:0] mux_1840_nl;
  wire[0:0] mux_1839_nl;
  wire[0:0] mux_1838_nl;
  wire[0:0] mux_1836_nl;
  wire[0:0] mux_1835_nl;
  wire[0:0] or_2033_nl;
  wire[0:0] nand_146_nl;
  wire[0:0] mux_1845_nl;
  wire[0:0] nand_338_nl;
  wire[0:0] mux_1848_nl;
  wire[0:0] mux_67_nl;
  wire[0:0] mux_66_nl;
  wire[0:0] or_23_nl;
  wire[0:0] nand_145_nl;
  wire[0:0] mux_1858_nl;
  wire[0:0] mux_1857_nl;
  wire[0:0] mux_1856_nl;
  wire[0:0] mux_1855_nl;
  wire[0:0] mux_1853_nl;
  wire[0:0] mux_1851_nl;
  wire[0:0] mux_1849_nl;
  wire[0:0] mux_1862_nl;
  wire[0:0] mux_1861_nl;
  wire[0:0] mux_1866_nl;
  wire[0:0] or_2041_nl;
  wire[0:0] mux_1865_nl;
  wire[0:0] mux_1864_nl;
  wire[0:0] mux_1863_nl;
  wire[0:0] mux_1869_nl;
  wire[0:0] mux_1868_nl;
  wire[0:0] mux_1867_nl;
  wire[0:0] or_2043_nl;
  wire[0:0] mux_1872_nl;
  wire[0:0] mux_1871_nl;
  wire[0:0] mux_1870_nl;
  wire[0:0] or_2175_nl;
  wire[0:0] mux_1874_nl;
  wire[0:0] mux_1873_nl;
  wire[0:0] and_248_nl;
  wire[0:0] mux_1875_nl;
  wire[0:0] and_213_nl;
  wire[0:0] mux_1877_nl;
  wire[0:0] or_2047_nl;
  wire[0:0] mux_1876_nl;
  wire[0:0] mux_1880_nl;
  wire[0:0] mux_1879_nl;
  wire[0:0] mux_1885_nl;
  wire[0:0] mux_1884_nl;
  wire[0:0] mux_1883_nl;
  wire[0:0] mux_1882_nl;
  wire[0:0] or_110_nl;
  wire[0:0] mux_1888_nl;
  wire[0:0] mux_1887_nl;
  wire[0:0] and_245_nl;
  wire[0:0] mux_459_nl;
  wire[0:0] mux_1896_nl;
  wire[0:0] mux_1895_nl;
  wire[0:0] mux_1894_nl;
  wire[0:0] mux_1893_nl;
  wire[0:0] mux_1892_nl;
  wire[0:0] mux_1891_nl;
  wire[0:0] nor_nl;
  wire[0:0] and_nl;
  wire[0:0] COMP_LOOP_nor_11_nl;
  wire[0:0] mux_1904_nl;
  wire[0:0] nor_758_nl;
  wire[0:0] and_256_nl;
  wire[0:0] mux_1910_nl;
  wire[0:0] mux_1907_nl;
  wire[0:0] and_445_nl;
  wire[0:0] mux_1800_nl;
  wire[0:0] mux_1905_nl;
  wire[0:0] and_446_nl;
  wire[0:0] mux_1901_nl;
  wire[0:0] mux_1794_nl;
  wire[0:0] COMP_LOOP_or_6_nl;
  wire[0:0] COMP_LOOP_or_7_nl;
  wire[0:0] COMP_LOOP_or_8_nl;
  wire[0:0] COMP_LOOP_or_9_nl;
  wire[0:0] COMP_LOOP_or_10_nl;
  wire[0:0] COMP_LOOP_or_11_nl;
  wire[0:0] COMP_LOOP_or_12_nl;
  wire[0:0] COMP_LOOP_or_13_nl;
  wire[0:0] COMP_LOOP_or_14_nl;
  wire[0:0] COMP_LOOP_or_15_nl;
  wire[0:0] COMP_LOOP_or_16_nl;
  wire[0:0] COMP_LOOP_or_17_nl;
  wire[0:0] COMP_LOOP_or_18_nl;
  wire[0:0] COMP_LOOP_or_19_nl;
  wire[0:0] COMP_LOOP_or_20_nl;
  wire[0:0] COMP_LOOP_or_21_nl;
  wire[3:0] COMP_LOOP_and_nl;
  wire[3:0] COMP_LOOP_mux1h_186_nl;
  wire[0:0] mux_1955_nl;
  wire[0:0] mux_1954_nl;
  wire[0:0] mux_1953_nl;
  wire[0:0] mux_1952_nl;
  wire[0:0] mux_1951_nl;
  wire[0:0] mux_1950_nl;
  wire[0:0] mux_1948_nl;
  wire[0:0] mux_1947_nl;
  wire[0:0] mux_1946_nl;
  wire[0:0] mux_1945_nl;
  wire[0:0] mux_1944_nl;
  wire[0:0] mux_1943_nl;
  wire[0:0] mux_1941_nl;
  wire[0:0] mux_1940_nl;
  wire[0:0] mux_1937_nl;
  wire[0:0] mux_1936_nl;
  wire[0:0] mux_1935_nl;
  wire[0:0] mux_1932_nl;
  wire[0:0] mux_1931_nl;
  wire[0:0] mux_1930_nl;
  wire[0:0] mux_1929_nl;
  wire[0:0] mux_1924_nl;
  wire[0:0] mux_1919_nl;
  wire[0:0] mux_1918_nl;
  wire[0:0] mux_1916_nl;
  wire[0:0] mux_1915_nl;
  wire[0:0] mux_1913_nl;
  wire[0:0] not_4628_nl;
  wire[0:0] not_nl;
  wire[0:0] mux_2196_nl;
  wire[0:0] mux_2195_nl;
  wire[0:0] mux_2194_nl;
  wire[0:0] mux_2193_nl;
  wire[0:0] mux_2192_nl;
  wire[0:0] mux_2191_nl;
  wire[0:0] mux_2190_nl;
  wire[0:0] mux_2189_nl;
  wire[0:0] mux_2187_nl;
  wire[0:0] mux_2186_nl;
  wire[0:0] mux_2185_nl;
  wire[0:0] mux_2184_nl;
  wire[0:0] mux_2183_nl;
  wire[0:0] mux_2182_nl;
  wire[0:0] mux_2181_nl;
  wire[0:0] mux_2177_nl;
  wire[0:0] mux_2174_nl;
  wire[0:0] mux_2173_nl;
  wire[0:0] mux_2172_nl;
  wire[0:0] mux_2165_nl;
  wire[0:0] mux_2161_nl;
  wire[0:0] mux_2157_nl;
  wire[4:0] COMP_LOOP_k_COMP_LOOP_k_mux_nl;
  wire[0:0] mux_2243_nl;
  wire[0:0] mux_2242_nl;
  wire[0:0] mux_2241_nl;
  wire[0:0] mux_2240_nl;
  wire[0:0] mux_2239_nl;
  wire[0:0] mux_2238_nl;
  wire[0:0] mux_2237_nl;
  wire[0:0] or_2347_nl;
  wire[0:0] mux_2236_nl;
  wire[0:0] mux_2235_nl;
  wire[0:0] mux_2234_nl;
  wire[0:0] mux_2233_nl;
  wire[0:0] mux_2230_nl;
  wire[0:0] mux_2228_nl;
  wire[0:0] mux_2227_nl;
  wire[0:0] mux_2226_nl;
  wire[0:0] mux_2225_nl;
  wire[0:0] mux_2224_nl;
  wire[0:0] mux_2223_nl;
  wire[0:0] mux_2218_nl;
  wire[0:0] mux_2213_nl;
  wire[0:0] mux_2212_nl;
  wire[0:0] mux_2210_nl;
  wire[0:0] mux_2209_nl;
  wire[0:0] mux_2207_nl;
  wire[0:0] mux_2204_nl;
  wire[0:0] mux_2203_nl;
  wire[0:0] mux_2201_nl;
  wire[0:0] mux_2200_nl;
  wire[0:0] mux_2198_nl;
  wire[0:0] mux_2262_nl;
  wire[0:0] nor_797_nl;
  wire[0:0] mux_2261_nl;
  wire[0:0] mux_2260_nl;
  wire[0:0] nand_396_nl;
  wire[0:0] mux_2259_nl;
  wire[0:0] or_2362_nl;
  wire[0:0] mux_2258_nl;
  wire[0:0] mux_2257_nl;
  wire[0:0] nand_397_nl;
  wire[0:0] mux_2255_nl;
  wire[0:0] and_700_nl;
  wire[0:0] mux_2254_nl;
  wire[0:0] nor_798_nl;
  wire[0:0] mux_2253_nl;
  wire[0:0] nor_799_nl;
  wire[0:0] nor_800_nl;
  wire[0:0] mux_2252_nl;
  wire[0:0] or_2356_nl;
  wire[0:0] mux_2250_nl;
  wire[0:0] nand_394_nl;
  wire[0:0] mux_2247_nl;
  wire[0:0] nand_398_nl;
  wire[0:0] mux_2246_nl;
  wire[63:0] COMP_LOOP_mux1h_209_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_930_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_932_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_934_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_936_nl;
  wire[0:0] COMP_LOOP_or_27_nl;
  wire[0:0] mux_51_nl;
  wire[0:0] nor_727_nl;
  wire[0:0] or_2152_nl;
  wire[0:0] nand_314_nl;
  wire[0:0] mux_514_nl;
  wire[0:0] or_265_nl;
  wire[0:0] mux_520_nl;
  wire[0:0] mux_1520_nl;
  wire[0:0] mux_1548_nl;
  wire[0:0] mux_1564_nl;
  wire[0:0] mux_1584_nl;
  wire[0:0] mux_1587_nl;
  wire[0:0] mux_1601_nl;
  wire[0:0] nor_275_nl;
  wire[0:0] mux_1611_nl;
  wire[0:0] and_272_nl;
  wire[0:0] mux_1610_nl;
  wire[0:0] nor_272_nl;
  wire[0:0] mux_1606_nl;
  wire[0:0] mux_1605_nl;
  wire[0:0] nor_273_nl;
  wire[0:0] and_273_nl;
  wire[0:0] mux_1603_nl;
  wire[0:0] nor_274_nl;
  wire[0:0] or_1849_nl;
  wire[0:0] or_1863_nl;
  wire[0:0] mux_1671_nl;
  wire[0:0] nand_111_nl;
  wire[0:0] mux_1670_nl;
  wire[0:0] nand_110_nl;
  wire[0:0] mux_1679_nl;
  wire[0:0] nand_151_nl;
  wire[0:0] nand_342_nl;
  wire[0:0] or_2000_nl;
  wire[0:0] mux_1779_nl;
  wire[0:0] and_261_nl;
  wire[0:0] mux_1804_nl;
  wire[0:0] mux_1803_nl;
  wire[0:0] or_1996_nl;
  wire[0:0] mux_1774_nl;
  wire[0:0] mux_1770_nl;
  wire[0:0] and_263_nl;
  wire[0:0] mux_1769_nl;
  wire[0:0] mux_1831_nl;
  wire[0:0] mux_1830_nl;
  wire[0:0] mux_1829_nl;
  wire[0:0] mux_1828_nl;
  wire[0:0] mux_1827_nl;
  wire[0:0] nor_248_nl;
  wire[0:0] mux_1843_nl;
  wire[0:0] nor_244_nl;
  wire[0:0] and_368_nl;
  wire[0:0] or_2091_nl;
  wire[0:0] and_42_nl;
  wire[0:0] and_52_nl;
  wire[0:0] and_57_nl;
  wire[0:0] and_67_nl;
  wire[0:0] and_73_nl;
  wire[0:0] and_80_nl;
  wire[0:0] and_87_nl;
  wire[0:0] and_93_nl;
  wire[0:0] and_99_nl;
  wire[0:0] and_103_nl;
  wire[0:0] and_107_nl;
  wire[0:0] and_111_nl;
  wire[0:0] and_116_nl;
  wire[0:0] and_120_nl;
  wire[0:0] and_124_nl;
  wire[0:0] and_129_nl;
  wire[0:0] and_131_nl;
  wire[0:0] mux_526_nl;
  wire[0:0] mux_525_nl;
  wire[0:0] or_280_nl;
  wire[0:0] mux_524_nl;
  wire[0:0] mux_523_nl;
  wire[0:0] mux_522_nl;
  wire[0:0] mux_521_nl;
  wire[0:0] or_275_nl;
  wire[0:0] mux_519_nl;
  wire[0:0] or_274_nl;
  wire[0:0] mux_518_nl;
  wire[0:0] mux_517_nl;
  wire[0:0] or_272_nl;
  wire[0:0] mux_516_nl;
  wire[0:0] or_271_nl;
  wire[0:0] or_269_nl;
  wire[0:0] mux_515_nl;
  wire[0:0] and_132_nl;
  wire[0:0] and_134_nl;
  wire[0:0] and_135_nl;
  wire[0:0] and_136_nl;
  wire[0:0] and_137_nl;
  wire[0:0] and_138_nl;
  wire[0:0] and_139_nl;
  wire[0:0] and_140_nl;
  wire[0:0] and_142_nl;
  wire[0:0] and_144_nl;
  wire[0:0] and_145_nl;
  wire[0:0] and_146_nl;
  wire[0:0] and_148_nl;
  wire[0:0] and_150_nl;
  wire[0:0] and_152_nl;
  wire[0:0] mux_556_nl;
  wire[0:0] mux_555_nl;
  wire[0:0] nor_689_nl;
  wire[0:0] mux_554_nl;
  wire[0:0] nand_10_nl;
  wire[0:0] mux_553_nl;
  wire[0:0] mux_552_nl;
  wire[0:0] or_319_nl;
  wire[0:0] mux_551_nl;
  wire[0:0] or_318_nl;
  wire[0:0] or_317_nl;
  wire[0:0] mux_550_nl;
  wire[0:0] nor_690_nl;
  wire[0:0] nor_691_nl;
  wire[0:0] mux_549_nl;
  wire[0:0] or_313_nl;
  wire[0:0] mux_548_nl;
  wire[0:0] and_344_nl;
  wire[0:0] mux_547_nl;
  wire[0:0] or_310_nl;
  wire[0:0] mux_546_nl;
  wire[0:0] mux_545_nl;
  wire[0:0] mux_544_nl;
  wire[0:0] or_308_nl;
  wire[0:0] mux_543_nl;
  wire[0:0] or_306_nl;
  wire[0:0] or_305_nl;
  wire[0:0] mux_542_nl;
  wire[0:0] or_304_nl;
  wire[0:0] nor_692_nl;
  wire[0:0] mux_541_nl;
  wire[0:0] nor_693_nl;
  wire[0:0] mux_540_nl;
  wire[0:0] mux_539_nl;
  wire[0:0] or_301_nl;
  wire[0:0] mux_538_nl;
  wire[0:0] mux_537_nl;
  wire[0:0] or_299_nl;
  wire[0:0] mux_536_nl;
  wire[0:0] or_297_nl;
  wire[0:0] mux_535_nl;
  wire[0:0] or_296_nl;
  wire[0:0] mux_534_nl;
  wire[0:0] or_295_nl;
  wire[0:0] nor_694_nl;
  wire[0:0] mux_533_nl;
  wire[0:0] nand_8_nl;
  wire[0:0] mux_532_nl;
  wire[0:0] or_292_nl;
  wire[0:0] mux_531_nl;
  wire[0:0] mux_530_nl;
  wire[0:0] or_290_nl;
  wire[0:0] mux_529_nl;
  wire[0:0] or_286_nl;
  wire[0:0] or_285_nl;
  wire[0:0] mux_528_nl;
  wire[0:0] or_284_nl;
  wire[0:0] mux_527_nl;
  wire[0:0] or_283_nl;
  wire[0:0] mux_587_nl;
  wire[0:0] mux_586_nl;
  wire[0:0] nor_669_nl;
  wire[0:0] mux_585_nl;
  wire[0:0] mux_584_nl;
  wire[0:0] or_372_nl;
  wire[0:0] mux_583_nl;
  wire[0:0] or_371_nl;
  wire[0:0] mux_582_nl;
  wire[0:0] mux_581_nl;
  wire[0:0] or_366_nl;
  wire[0:0] mux_580_nl;
  wire[0:0] or_365_nl;
  wire[0:0] or_363_nl;
  wire[0:0] mux_579_nl;
  wire[0:0] nor_670_nl;
  wire[0:0] mux_578_nl;
  wire[0:0] mux_577_nl;
  wire[0:0] or_361_nl;
  wire[0:0] or_359_nl;
  wire[0:0] or_358_nl;
  wire[0:0] nor_671_nl;
  wire[0:0] mux_576_nl;
  wire[0:0] mux_575_nl;
  wire[0:0] nor_672_nl;
  wire[0:0] and_342_nl;
  wire[0:0] mux_574_nl;
  wire[0:0] nor_673_nl;
  wire[0:0] mux_573_nl;
  wire[0:0] nor_674_nl;
  wire[0:0] nor_675_nl;
  wire[0:0] and_343_nl;
  wire[0:0] mux_572_nl;
  wire[0:0] mux_571_nl;
  wire[0:0] mux_570_nl;
  wire[0:0] nor_676_nl;
  wire[0:0] nor_677_nl;
  wire[0:0] mux_569_nl;
  wire[0:0] nor_679_nl;
  wire[0:0] mux_568_nl;
  wire[0:0] mux_567_nl;
  wire[0:0] nor_680_nl;
  wire[0:0] nor_681_nl;
  wire[0:0] nor_682_nl;
  wire[0:0] nor_683_nl;
  wire[0:0] mux_566_nl;
  wire[0:0] nand_11_nl;
  wire[0:0] mux_565_nl;
  wire[0:0] mux_564_nl;
  wire[0:0] mux_563_nl;
  wire[0:0] nor_685_nl;
  wire[0:0] mux_562_nl;
  wire[0:0] nor_686_nl;
  wire[0:0] nor_687_nl;
  wire[0:0] nor_688_nl;
  wire[0:0] or_329_nl;
  wire[0:0] mux_561_nl;
  wire[0:0] or_328_nl;
  wire[0:0] mux_560_nl;
  wire[0:0] mux_559_nl;
  wire[0:0] or_326_nl;
  wire[0:0] mux_558_nl;
  wire[0:0] or_322_nl;
  wire[0:0] mux_618_nl;
  wire[0:0] mux_617_nl;
  wire[0:0] mux_616_nl;
  wire[0:0] nor_661_nl;
  wire[0:0] mux_615_nl;
  wire[0:0] mux_614_nl;
  wire[0:0] or_413_nl;
  wire[0:0] mux_613_nl;
  wire[0:0] or_412_nl;
  wire[0:0] and_341_nl;
  wire[0:0] mux_612_nl;
  wire[0:0] or_410_nl;
  wire[0:0] mux_611_nl;
  wire[0:0] mux_610_nl;
  wire[0:0] or_409_nl;
  wire[0:0] mux_609_nl;
  wire[0:0] or_408_nl;
  wire[0:0] nor_662_nl;
  wire[0:0] mux_608_nl;
  wire[0:0] or_405_nl;
  wire[0:0] nor_663_nl;
  wire[0:0] mux_607_nl;
  wire[0:0] mux_606_nl;
  wire[0:0] or_402_nl;
  wire[0:0] or_401_nl;
  wire[0:0] nand_14_nl;
  wire[0:0] mux_605_nl;
  wire[0:0] or_400_nl;
  wire[0:0] mux_604_nl;
  wire[0:0] or_399_nl;
  wire[0:0] mux_603_nl;
  wire[0:0] mux_602_nl;
  wire[0:0] nor_664_nl;
  wire[0:0] mux_601_nl;
  wire[0:0] nor_665_nl;
  wire[0:0] nor_666_nl;
  wire[0:0] mux_600_nl;
  wire[0:0] or_394_nl;
  wire[0:0] mux_599_nl;
  wire[0:0] or_393_nl;
  wire[0:0] mux_598_nl;
  wire[0:0] nor_667_nl;
  wire[0:0] mux_597_nl;
  wire[0:0] or_389_nl;
  wire[0:0] mux_596_nl;
  wire[0:0] mux_595_nl;
  wire[0:0] or_388_nl;
  wire[0:0] mux_594_nl;
  wire[0:0] or_387_nl;
  wire[0:0] nor_668_nl;
  wire[0:0] mux_593_nl;
  wire[0:0] mux_592_nl;
  wire[0:0] mux_591_nl;
  wire[0:0] or_383_nl;
  wire[0:0] mux_590_nl;
  wire[0:0] or_380_nl;
  wire[0:0] or_378_nl;
  wire[0:0] mux_589_nl;
  wire[0:0] or_377_nl;
  wire[0:0] mux_649_nl;
  wire[0:0] mux_648_nl;
  wire[0:0] nor_641_nl;
  wire[0:0] mux_647_nl;
  wire[0:0] mux_646_nl;
  wire[0:0] or_465_nl;
  wire[0:0] mux_645_nl;
  wire[0:0] or_464_nl;
  wire[0:0] mux_644_nl;
  wire[0:0] mux_643_nl;
  wire[0:0] or_461_nl;
  wire[0:0] or_459_nl;
  wire[0:0] mux_642_nl;
  wire[0:0] or_458_nl;
  wire[0:0] or_456_nl;
  wire[0:0] mux_641_nl;
  wire[0:0] nor_642_nl;
  wire[0:0] mux_640_nl;
  wire[0:0] mux_639_nl;
  wire[0:0] or_454_nl;
  wire[0:0] or_452_nl;
  wire[0:0] or_451_nl;
  wire[0:0] nor_643_nl;
  wire[0:0] mux_638_nl;
  wire[0:0] mux_637_nl;
  wire[0:0] nor_644_nl;
  wire[0:0] and_339_nl;
  wire[0:0] mux_636_nl;
  wire[0:0] nor_645_nl;
  wire[0:0] mux_635_nl;
  wire[0:0] nor_646_nl;
  wire[0:0] nor_647_nl;
  wire[0:0] and_340_nl;
  wire[0:0] mux_634_nl;
  wire[0:0] mux_633_nl;
  wire[0:0] mux_632_nl;
  wire[0:0] nor_648_nl;
  wire[0:0] nor_649_nl;
  wire[0:0] mux_631_nl;
  wire[0:0] nor_651_nl;
  wire[0:0] mux_630_nl;
  wire[0:0] mux_629_nl;
  wire[0:0] nor_652_nl;
  wire[0:0] nor_653_nl;
  wire[0:0] nor_654_nl;
  wire[0:0] nor_655_nl;
  wire[0:0] mux_628_nl;
  wire[0:0] nand_17_nl;
  wire[0:0] mux_627_nl;
  wire[0:0] mux_626_nl;
  wire[0:0] mux_625_nl;
  wire[0:0] nor_657_nl;
  wire[0:0] mux_624_nl;
  wire[0:0] nor_658_nl;
  wire[0:0] nor_659_nl;
  wire[0:0] nor_660_nl;
  wire[0:0] or_422_nl;
  wire[0:0] mux_623_nl;
  wire[0:0] or_421_nl;
  wire[0:0] mux_622_nl;
  wire[0:0] mux_621_nl;
  wire[0:0] or_419_nl;
  wire[0:0] or_418_nl;
  wire[0:0] mux_620_nl;
  wire[0:0] or_415_nl;
  wire[0:0] mux_680_nl;
  wire[0:0] mux_679_nl;
  wire[0:0] nor_635_nl;
  wire[0:0] mux_678_nl;
  wire[0:0] nand_22_nl;
  wire[0:0] mux_677_nl;
  wire[0:0] mux_676_nl;
  wire[0:0] or_505_nl;
  wire[0:0] mux_675_nl;
  wire[0:0] or_504_nl;
  wire[0:0] or_503_nl;
  wire[0:0] mux_674_nl;
  wire[0:0] nor_636_nl;
  wire[0:0] nor_637_nl;
  wire[0:0] mux_673_nl;
  wire[0:0] or_499_nl;
  wire[0:0] mux_672_nl;
  wire[0:0] and_338_nl;
  wire[0:0] mux_671_nl;
  wire[0:0] or_496_nl;
  wire[0:0] mux_670_nl;
  wire[0:0] mux_669_nl;
  wire[0:0] mux_668_nl;
  wire[0:0] or_494_nl;
  wire[0:0] mux_667_nl;
  wire[0:0] or_492_nl;
  wire[0:0] or_491_nl;
  wire[0:0] mux_666_nl;
  wire[0:0] or_490_nl;
  wire[0:0] nor_638_nl;
  wire[0:0] mux_665_nl;
  wire[0:0] nor_639_nl;
  wire[0:0] mux_664_nl;
  wire[0:0] mux_663_nl;
  wire[0:0] or_487_nl;
  wire[0:0] mux_662_nl;
  wire[0:0] mux_661_nl;
  wire[0:0] or_485_nl;
  wire[0:0] mux_660_nl;
  wire[0:0] or_483_nl;
  wire[0:0] mux_659_nl;
  wire[0:0] or_482_nl;
  wire[0:0] mux_658_nl;
  wire[0:0] or_481_nl;
  wire[0:0] nor_640_nl;
  wire[0:0] mux_657_nl;
  wire[0:0] nand_20_nl;
  wire[0:0] mux_656_nl;
  wire[0:0] or_478_nl;
  wire[0:0] mux_655_nl;
  wire[0:0] mux_654_nl;
  wire[0:0] or_476_nl;
  wire[0:0] mux_653_nl;
  wire[0:0] or_472_nl;
  wire[0:0] or_471_nl;
  wire[0:0] mux_652_nl;
  wire[0:0] or_470_nl;
  wire[0:0] mux_651_nl;
  wire[0:0] or_469_nl;
  wire[0:0] mux_711_nl;
  wire[0:0] mux_710_nl;
  wire[0:0] nor_615_nl;
  wire[0:0] mux_709_nl;
  wire[0:0] mux_708_nl;
  wire[0:0] or_558_nl;
  wire[0:0] mux_707_nl;
  wire[0:0] or_557_nl;
  wire[0:0] mux_706_nl;
  wire[0:0] mux_705_nl;
  wire[0:0] or_552_nl;
  wire[0:0] mux_704_nl;
  wire[0:0] or_551_nl;
  wire[0:0] or_549_nl;
  wire[0:0] mux_703_nl;
  wire[0:0] nor_616_nl;
  wire[0:0] mux_702_nl;
  wire[0:0] mux_701_nl;
  wire[0:0] or_547_nl;
  wire[0:0] or_545_nl;
  wire[0:0] or_544_nl;
  wire[0:0] nor_617_nl;
  wire[0:0] mux_700_nl;
  wire[0:0] mux_699_nl;
  wire[0:0] nor_618_nl;
  wire[0:0] and_336_nl;
  wire[0:0] mux_698_nl;
  wire[0:0] nor_619_nl;
  wire[0:0] mux_697_nl;
  wire[0:0] nor_620_nl;
  wire[0:0] nor_621_nl;
  wire[0:0] and_337_nl;
  wire[0:0] mux_696_nl;
  wire[0:0] mux_695_nl;
  wire[0:0] mux_694_nl;
  wire[0:0] nor_622_nl;
  wire[0:0] nor_623_nl;
  wire[0:0] mux_693_nl;
  wire[0:0] nor_625_nl;
  wire[0:0] mux_692_nl;
  wire[0:0] mux_691_nl;
  wire[0:0] nor_626_nl;
  wire[0:0] nor_627_nl;
  wire[0:0] nor_628_nl;
  wire[0:0] nor_629_nl;
  wire[0:0] mux_690_nl;
  wire[0:0] nand_23_nl;
  wire[0:0] mux_689_nl;
  wire[0:0] mux_688_nl;
  wire[0:0] mux_687_nl;
  wire[0:0] nor_631_nl;
  wire[0:0] mux_686_nl;
  wire[0:0] nor_632_nl;
  wire[0:0] nor_633_nl;
  wire[0:0] nor_634_nl;
  wire[0:0] or_515_nl;
  wire[0:0] mux_685_nl;
  wire[0:0] or_514_nl;
  wire[0:0] mux_684_nl;
  wire[0:0] mux_683_nl;
  wire[0:0] or_512_nl;
  wire[0:0] mux_682_nl;
  wire[0:0] or_508_nl;
  wire[0:0] mux_742_nl;
  wire[0:0] mux_741_nl;
  wire[0:0] nor_609_nl;
  wire[0:0] mux_740_nl;
  wire[0:0] nand_28_nl;
  wire[0:0] mux_739_nl;
  wire[0:0] mux_738_nl;
  wire[0:0] or_598_nl;
  wire[0:0] mux_737_nl;
  wire[0:0] or_597_nl;
  wire[0:0] or_596_nl;
  wire[0:0] mux_736_nl;
  wire[0:0] and_439_nl;
  wire[0:0] nor_611_nl;
  wire[0:0] mux_735_nl;
  wire[0:0] or_592_nl;
  wire[0:0] mux_734_nl;
  wire[0:0] and_335_nl;
  wire[0:0] mux_733_nl;
  wire[0:0] or_589_nl;
  wire[0:0] mux_732_nl;
  wire[0:0] mux_731_nl;
  wire[0:0] mux_730_nl;
  wire[0:0] or_587_nl;
  wire[0:0] mux_729_nl;
  wire[0:0] or_585_nl;
  wire[0:0] or_584_nl;
  wire[0:0] mux_728_nl;
  wire[0:0] or_583_nl;
  wire[0:0] nor_612_nl;
  wire[0:0] mux_727_nl;
  wire[0:0] nor_613_nl;
  wire[0:0] mux_726_nl;
  wire[0:0] mux_725_nl;
  wire[0:0] or_580_nl;
  wire[0:0] mux_724_nl;
  wire[0:0] mux_723_nl;
  wire[0:0] or_578_nl;
  wire[0:0] mux_722_nl;
  wire[0:0] or_576_nl;
  wire[0:0] mux_721_nl;
  wire[0:0] or_575_nl;
  wire[0:0] mux_720_nl;
  wire[0:0] or_574_nl;
  wire[0:0] nor_614_nl;
  wire[0:0] mux_719_nl;
  wire[0:0] nand_26_nl;
  wire[0:0] mux_718_nl;
  wire[0:0] or_571_nl;
  wire[0:0] mux_717_nl;
  wire[0:0] mux_716_nl;
  wire[0:0] or_569_nl;
  wire[0:0] mux_715_nl;
  wire[0:0] or_565_nl;
  wire[0:0] or_564_nl;
  wire[0:0] mux_714_nl;
  wire[0:0] or_563_nl;
  wire[0:0] mux_713_nl;
  wire[0:0] or_562_nl;
  wire[0:0] mux_773_nl;
  wire[0:0] mux_772_nl;
  wire[0:0] nor_589_nl;
  wire[0:0] mux_771_nl;
  wire[0:0] mux_770_nl;
  wire[0:0] or_651_nl;
  wire[0:0] mux_769_nl;
  wire[0:0] or_650_nl;
  wire[0:0] mux_768_nl;
  wire[0:0] mux_767_nl;
  wire[0:0] or_647_nl;
  wire[0:0] or_645_nl;
  wire[0:0] mux_766_nl;
  wire[0:0] or_644_nl;
  wire[0:0] or_642_nl;
  wire[0:0] mux_765_nl;
  wire[0:0] nor_590_nl;
  wire[0:0] mux_764_nl;
  wire[0:0] mux_763_nl;
  wire[0:0] or_640_nl;
  wire[0:0] or_638_nl;
  wire[0:0] or_637_nl;
  wire[0:0] nor_591_nl;
  wire[0:0] mux_762_nl;
  wire[0:0] mux_761_nl;
  wire[0:0] nor_592_nl;
  wire[0:0] and_333_nl;
  wire[0:0] mux_760_nl;
  wire[0:0] nor_593_nl;
  wire[0:0] mux_759_nl;
  wire[0:0] nor_594_nl;
  wire[0:0] nor_595_nl;
  wire[0:0] and_334_nl;
  wire[0:0] mux_758_nl;
  wire[0:0] mux_757_nl;
  wire[0:0] mux_756_nl;
  wire[0:0] nor_596_nl;
  wire[0:0] nor_597_nl;
  wire[0:0] mux_755_nl;
  wire[0:0] nor_599_nl;
  wire[0:0] mux_754_nl;
  wire[0:0] mux_753_nl;
  wire[0:0] nor_600_nl;
  wire[0:0] nor_601_nl;
  wire[0:0] nor_602_nl;
  wire[0:0] nor_603_nl;
  wire[0:0] mux_752_nl;
  wire[0:0] nand_29_nl;
  wire[0:0] mux_751_nl;
  wire[0:0] mux_750_nl;
  wire[0:0] mux_749_nl;
  wire[0:0] nor_605_nl;
  wire[0:0] mux_748_nl;
  wire[0:0] nor_606_nl;
  wire[0:0] nor_607_nl;
  wire[0:0] nor_608_nl;
  wire[0:0] or_608_nl;
  wire[0:0] mux_747_nl;
  wire[0:0] or_607_nl;
  wire[0:0] mux_746_nl;
  wire[0:0] mux_745_nl;
  wire[0:0] or_605_nl;
  wire[0:0] or_604_nl;
  wire[0:0] mux_744_nl;
  wire[0:0] or_601_nl;
  wire[0:0] mux_804_nl;
  wire[0:0] mux_803_nl;
  wire[0:0] nor_583_nl;
  wire[0:0] mux_802_nl;
  wire[0:0] nand_34_nl;
  wire[0:0] mux_801_nl;
  wire[0:0] mux_800_nl;
  wire[0:0] or_691_nl;
  wire[0:0] mux_799_nl;
  wire[0:0] or_690_nl;
  wire[0:0] or_689_nl;
  wire[0:0] mux_798_nl;
  wire[0:0] nor_584_nl;
  wire[0:0] nor_585_nl;
  wire[0:0] mux_797_nl;
  wire[0:0] or_685_nl;
  wire[0:0] mux_796_nl;
  wire[0:0] and_332_nl;
  wire[0:0] mux_795_nl;
  wire[0:0] or_682_nl;
  wire[0:0] mux_794_nl;
  wire[0:0] mux_793_nl;
  wire[0:0] mux_792_nl;
  wire[0:0] or_680_nl;
  wire[0:0] mux_791_nl;
  wire[0:0] or_678_nl;
  wire[0:0] or_677_nl;
  wire[0:0] mux_790_nl;
  wire[0:0] or_676_nl;
  wire[0:0] nor_586_nl;
  wire[0:0] mux_789_nl;
  wire[0:0] nor_587_nl;
  wire[0:0] mux_788_nl;
  wire[0:0] mux_787_nl;
  wire[0:0] or_673_nl;
  wire[0:0] mux_786_nl;
  wire[0:0] mux_785_nl;
  wire[0:0] or_671_nl;
  wire[0:0] mux_784_nl;
  wire[0:0] or_669_nl;
  wire[0:0] mux_783_nl;
  wire[0:0] or_668_nl;
  wire[0:0] mux_782_nl;
  wire[0:0] or_667_nl;
  wire[0:0] nor_588_nl;
  wire[0:0] mux_781_nl;
  wire[0:0] nand_32_nl;
  wire[0:0] mux_780_nl;
  wire[0:0] or_664_nl;
  wire[0:0] mux_779_nl;
  wire[0:0] mux_778_nl;
  wire[0:0] or_662_nl;
  wire[0:0] mux_777_nl;
  wire[0:0] or_658_nl;
  wire[0:0] or_657_nl;
  wire[0:0] mux_776_nl;
  wire[0:0] or_656_nl;
  wire[0:0] mux_775_nl;
  wire[0:0] or_655_nl;
  wire[0:0] mux_835_nl;
  wire[0:0] mux_834_nl;
  wire[0:0] nor_563_nl;
  wire[0:0] mux_833_nl;
  wire[0:0] mux_832_nl;
  wire[0:0] or_744_nl;
  wire[0:0] mux_831_nl;
  wire[0:0] or_743_nl;
  wire[0:0] mux_830_nl;
  wire[0:0] mux_829_nl;
  wire[0:0] or_738_nl;
  wire[0:0] mux_828_nl;
  wire[0:0] or_737_nl;
  wire[0:0] or_735_nl;
  wire[0:0] mux_827_nl;
  wire[0:0] nor_564_nl;
  wire[0:0] mux_826_nl;
  wire[0:0] mux_825_nl;
  wire[0:0] or_733_nl;
  wire[0:0] or_731_nl;
  wire[0:0] or_730_nl;
  wire[0:0] nor_565_nl;
  wire[0:0] mux_824_nl;
  wire[0:0] mux_823_nl;
  wire[0:0] nor_566_nl;
  wire[0:0] and_330_nl;
  wire[0:0] mux_822_nl;
  wire[0:0] nor_567_nl;
  wire[0:0] mux_821_nl;
  wire[0:0] nor_568_nl;
  wire[0:0] nor_569_nl;
  wire[0:0] and_331_nl;
  wire[0:0] mux_820_nl;
  wire[0:0] mux_819_nl;
  wire[0:0] mux_818_nl;
  wire[0:0] nor_570_nl;
  wire[0:0] nor_571_nl;
  wire[0:0] mux_817_nl;
  wire[0:0] nor_573_nl;
  wire[0:0] mux_816_nl;
  wire[0:0] mux_815_nl;
  wire[0:0] nor_574_nl;
  wire[0:0] nor_575_nl;
  wire[0:0] nor_576_nl;
  wire[0:0] nor_577_nl;
  wire[0:0] mux_814_nl;
  wire[0:0] nand_35_nl;
  wire[0:0] mux_813_nl;
  wire[0:0] mux_812_nl;
  wire[0:0] mux_811_nl;
  wire[0:0] nor_579_nl;
  wire[0:0] mux_810_nl;
  wire[0:0] nor_580_nl;
  wire[0:0] nor_581_nl;
  wire[0:0] nor_582_nl;
  wire[0:0] or_701_nl;
  wire[0:0] mux_809_nl;
  wire[0:0] or_700_nl;
  wire[0:0] mux_808_nl;
  wire[0:0] mux_807_nl;
  wire[0:0] or_698_nl;
  wire[0:0] mux_806_nl;
  wire[0:0] or_694_nl;
  wire[0:0] mux_866_nl;
  wire[0:0] mux_865_nl;
  wire[0:0] mux_864_nl;
  wire[0:0] nor_555_nl;
  wire[0:0] mux_863_nl;
  wire[0:0] mux_862_nl;
  wire[0:0] or_785_nl;
  wire[0:0] mux_861_nl;
  wire[0:0] or_784_nl;
  wire[0:0] and_329_nl;
  wire[0:0] mux_860_nl;
  wire[0:0] or_782_nl;
  wire[0:0] mux_859_nl;
  wire[0:0] mux_858_nl;
  wire[0:0] or_781_nl;
  wire[0:0] mux_857_nl;
  wire[0:0] or_780_nl;
  wire[0:0] nor_556_nl;
  wire[0:0] mux_856_nl;
  wire[0:0] or_777_nl;
  wire[0:0] nor_557_nl;
  wire[0:0] mux_855_nl;
  wire[0:0] mux_854_nl;
  wire[0:0] or_774_nl;
  wire[0:0] or_773_nl;
  wire[0:0] nand_38_nl;
  wire[0:0] mux_853_nl;
  wire[0:0] or_772_nl;
  wire[0:0] mux_852_nl;
  wire[0:0] or_771_nl;
  wire[0:0] mux_851_nl;
  wire[0:0] mux_850_nl;
  wire[0:0] nor_558_nl;
  wire[0:0] mux_849_nl;
  wire[0:0] nor_559_nl;
  wire[0:0] nor_560_nl;
  wire[0:0] mux_848_nl;
  wire[0:0] or_766_nl;
  wire[0:0] mux_847_nl;
  wire[0:0] or_765_nl;
  wire[0:0] mux_846_nl;
  wire[0:0] nor_561_nl;
  wire[0:0] mux_845_nl;
  wire[0:0] or_761_nl;
  wire[0:0] mux_844_nl;
  wire[0:0] mux_843_nl;
  wire[0:0] or_760_nl;
  wire[0:0] mux_842_nl;
  wire[0:0] or_759_nl;
  wire[0:0] nor_562_nl;
  wire[0:0] mux_841_nl;
  wire[0:0] mux_840_nl;
  wire[0:0] mux_839_nl;
  wire[0:0] or_755_nl;
  wire[0:0] mux_838_nl;
  wire[0:0] or_752_nl;
  wire[0:0] or_750_nl;
  wire[0:0] mux_837_nl;
  wire[0:0] or_749_nl;
  wire[0:0] mux_897_nl;
  wire[0:0] mux_896_nl;
  wire[0:0] nor_535_nl;
  wire[0:0] mux_895_nl;
  wire[0:0] mux_894_nl;
  wire[0:0] or_837_nl;
  wire[0:0] mux_893_nl;
  wire[0:0] or_836_nl;
  wire[0:0] mux_892_nl;
  wire[0:0] mux_891_nl;
  wire[0:0] or_833_nl;
  wire[0:0] or_831_nl;
  wire[0:0] mux_890_nl;
  wire[0:0] or_830_nl;
  wire[0:0] or_828_nl;
  wire[0:0] mux_889_nl;
  wire[0:0] nor_536_nl;
  wire[0:0] mux_888_nl;
  wire[0:0] mux_887_nl;
  wire[0:0] or_826_nl;
  wire[0:0] or_824_nl;
  wire[0:0] or_823_nl;
  wire[0:0] nor_537_nl;
  wire[0:0] mux_886_nl;
  wire[0:0] mux_885_nl;
  wire[0:0] nor_538_nl;
  wire[0:0] and_327_nl;
  wire[0:0] mux_884_nl;
  wire[0:0] nor_539_nl;
  wire[0:0] mux_883_nl;
  wire[0:0] nor_540_nl;
  wire[0:0] nor_541_nl;
  wire[0:0] and_328_nl;
  wire[0:0] mux_882_nl;
  wire[0:0] mux_881_nl;
  wire[0:0] mux_880_nl;
  wire[0:0] nor_542_nl;
  wire[0:0] nor_543_nl;
  wire[0:0] mux_879_nl;
  wire[0:0] nor_545_nl;
  wire[0:0] mux_878_nl;
  wire[0:0] mux_877_nl;
  wire[0:0] nor_546_nl;
  wire[0:0] nor_547_nl;
  wire[0:0] nor_548_nl;
  wire[0:0] nor_549_nl;
  wire[0:0] mux_876_nl;
  wire[0:0] nand_41_nl;
  wire[0:0] mux_875_nl;
  wire[0:0] mux_874_nl;
  wire[0:0] mux_873_nl;
  wire[0:0] nor_551_nl;
  wire[0:0] mux_872_nl;
  wire[0:0] nor_552_nl;
  wire[0:0] nor_553_nl;
  wire[0:0] nor_554_nl;
  wire[0:0] or_794_nl;
  wire[0:0] mux_871_nl;
  wire[0:0] or_793_nl;
  wire[0:0] mux_870_nl;
  wire[0:0] mux_869_nl;
  wire[0:0] or_791_nl;
  wire[0:0] or_790_nl;
  wire[0:0] mux_868_nl;
  wire[0:0] or_787_nl;
  wire[0:0] mux_928_nl;
  wire[0:0] mux_927_nl;
  wire[0:0] nor_529_nl;
  wire[0:0] mux_926_nl;
  wire[0:0] nand_46_nl;
  wire[0:0] mux_925_nl;
  wire[0:0] mux_924_nl;
  wire[0:0] or_877_nl;
  wire[0:0] mux_923_nl;
  wire[0:0] or_876_nl;
  wire[0:0] or_875_nl;
  wire[0:0] mux_922_nl;
  wire[0:0] and_438_nl;
  wire[0:0] nor_531_nl;
  wire[0:0] mux_921_nl;
  wire[0:0] or_871_nl;
  wire[0:0] mux_920_nl;
  wire[0:0] and_326_nl;
  wire[0:0] mux_919_nl;
  wire[0:0] or_868_nl;
  wire[0:0] mux_918_nl;
  wire[0:0] mux_917_nl;
  wire[0:0] mux_916_nl;
  wire[0:0] or_866_nl;
  wire[0:0] mux_915_nl;
  wire[0:0] or_864_nl;
  wire[0:0] or_863_nl;
  wire[0:0] mux_914_nl;
  wire[0:0] or_862_nl;
  wire[0:0] nor_532_nl;
  wire[0:0] mux_913_nl;
  wire[0:0] nor_533_nl;
  wire[0:0] mux_912_nl;
  wire[0:0] mux_911_nl;
  wire[0:0] or_859_nl;
  wire[0:0] mux_910_nl;
  wire[0:0] mux_909_nl;
  wire[0:0] or_857_nl;
  wire[0:0] mux_908_nl;
  wire[0:0] or_855_nl;
  wire[0:0] mux_907_nl;
  wire[0:0] or_854_nl;
  wire[0:0] mux_906_nl;
  wire[0:0] or_853_nl;
  wire[0:0] nor_534_nl;
  wire[0:0] mux_905_nl;
  wire[0:0] nand_44_nl;
  wire[0:0] mux_904_nl;
  wire[0:0] or_850_nl;
  wire[0:0] mux_903_nl;
  wire[0:0] mux_902_nl;
  wire[0:0] or_848_nl;
  wire[0:0] mux_901_nl;
  wire[0:0] or_844_nl;
  wire[0:0] or_843_nl;
  wire[0:0] mux_900_nl;
  wire[0:0] or_842_nl;
  wire[0:0] mux_899_nl;
  wire[0:0] or_841_nl;
  wire[0:0] mux_959_nl;
  wire[0:0] mux_958_nl;
  wire[0:0] nor_509_nl;
  wire[0:0] mux_957_nl;
  wire[0:0] mux_956_nl;
  wire[0:0] or_930_nl;
  wire[0:0] mux_955_nl;
  wire[0:0] or_929_nl;
  wire[0:0] mux_954_nl;
  wire[0:0] mux_953_nl;
  wire[0:0] or_924_nl;
  wire[0:0] mux_952_nl;
  wire[0:0] or_923_nl;
  wire[0:0] or_921_nl;
  wire[0:0] mux_951_nl;
  wire[0:0] nor_510_nl;
  wire[0:0] mux_950_nl;
  wire[0:0] mux_949_nl;
  wire[0:0] or_919_nl;
  wire[0:0] or_917_nl;
  wire[0:0] or_916_nl;
  wire[0:0] nor_511_nl;
  wire[0:0] mux_948_nl;
  wire[0:0] mux_947_nl;
  wire[0:0] nor_512_nl;
  wire[0:0] and_324_nl;
  wire[0:0] mux_946_nl;
  wire[0:0] nor_513_nl;
  wire[0:0] mux_945_nl;
  wire[0:0] nor_514_nl;
  wire[0:0] nor_515_nl;
  wire[0:0] and_325_nl;
  wire[0:0] mux_944_nl;
  wire[0:0] mux_943_nl;
  wire[0:0] mux_942_nl;
  wire[0:0] nor_516_nl;
  wire[0:0] nor_517_nl;
  wire[0:0] mux_941_nl;
  wire[0:0] nor_519_nl;
  wire[0:0] mux_940_nl;
  wire[0:0] mux_939_nl;
  wire[0:0] nor_520_nl;
  wire[0:0] nor_521_nl;
  wire[0:0] nor_522_nl;
  wire[0:0] nor_523_nl;
  wire[0:0] mux_938_nl;
  wire[0:0] nand_47_nl;
  wire[0:0] mux_937_nl;
  wire[0:0] mux_936_nl;
  wire[0:0] mux_935_nl;
  wire[0:0] nor_525_nl;
  wire[0:0] mux_934_nl;
  wire[0:0] nor_526_nl;
  wire[0:0] nor_527_nl;
  wire[0:0] nor_528_nl;
  wire[0:0] or_887_nl;
  wire[0:0] mux_933_nl;
  wire[0:0] or_886_nl;
  wire[0:0] mux_932_nl;
  wire[0:0] mux_931_nl;
  wire[0:0] or_884_nl;
  wire[0:0] mux_930_nl;
  wire[0:0] or_880_nl;
  wire[0:0] mux_990_nl;
  wire[0:0] mux_989_nl;
  wire[0:0] nor_503_nl;
  wire[0:0] mux_988_nl;
  wire[0:0] nand_52_nl;
  wire[0:0] mux_987_nl;
  wire[0:0] mux_986_nl;
  wire[0:0] or_970_nl;
  wire[0:0] mux_985_nl;
  wire[0:0] or_969_nl;
  wire[0:0] or_968_nl;
  wire[0:0] mux_984_nl;
  wire[0:0] and_437_nl;
  wire[0:0] nor_505_nl;
  wire[0:0] mux_983_nl;
  wire[0:0] or_964_nl;
  wire[0:0] mux_982_nl;
  wire[0:0] and_323_nl;
  wire[0:0] mux_981_nl;
  wire[0:0] nand_376_nl;
  wire[0:0] mux_980_nl;
  wire[0:0] mux_979_nl;
  wire[0:0] mux_978_nl;
  wire[0:0] or_959_nl;
  wire[0:0] mux_977_nl;
  wire[0:0] or_957_nl;
  wire[0:0] or_956_nl;
  wire[0:0] mux_976_nl;
  wire[0:0] or_955_nl;
  wire[0:0] nor_506_nl;
  wire[0:0] mux_975_nl;
  wire[0:0] nor_507_nl;
  wire[0:0] mux_974_nl;
  wire[0:0] mux_973_nl;
  wire[0:0] nand_371_nl;
  wire[0:0] mux_972_nl;
  wire[0:0] mux_971_nl;
  wire[0:0] or_950_nl;
  wire[0:0] mux_970_nl;
  wire[0:0] or_948_nl;
  wire[0:0] mux_969_nl;
  wire[0:0] or_947_nl;
  wire[0:0] mux_968_nl;
  wire[0:0] or_946_nl;
  wire[0:0] nor_508_nl;
  wire[0:0] mux_967_nl;
  wire[0:0] nand_50_nl;
  wire[0:0] mux_966_nl;
  wire[0:0] nand_360_nl;
  wire[0:0] mux_965_nl;
  wire[0:0] mux_964_nl;
  wire[0:0] or_941_nl;
  wire[0:0] mux_963_nl;
  wire[0:0] or_937_nl;
  wire[0:0] or_936_nl;
  wire[0:0] mux_962_nl;
  wire[0:0] or_935_nl;
  wire[0:0] mux_961_nl;
  wire[0:0] or_934_nl;
  wire[0:0] mux_1021_nl;
  wire[0:0] mux_1020_nl;
  wire[0:0] nor_484_nl;
  wire[0:0] mux_1019_nl;
  wire[0:0] mux_1018_nl;
  wire[0:0] nand_274_nl;
  wire[0:0] mux_1017_nl;
  wire[0:0] or_1022_nl;
  wire[0:0] mux_1016_nl;
  wire[0:0] mux_1015_nl;
  wire[0:0] or_1019_nl;
  wire[0:0] or_1017_nl;
  wire[0:0] mux_1014_nl;
  wire[0:0] nand_370_nl;
  wire[0:0] or_1014_nl;
  wire[0:0] mux_1013_nl;
  wire[0:0] nor_485_nl;
  wire[0:0] mux_1012_nl;
  wire[0:0] mux_1011_nl;
  wire[0:0] or_1012_nl;
  wire[0:0] or_1010_nl;
  wire[0:0] or_1009_nl;
  wire[0:0] nor_486_nl;
  wire[0:0] mux_1010_nl;
  wire[0:0] mux_1009_nl;
  wire[0:0] nor_487_nl;
  wire[0:0] and_320_nl;
  wire[0:0] mux_1008_nl;
  wire[0:0] nor_488_nl;
  wire[0:0] mux_1007_nl;
  wire[0:0] and_321_nl;
  wire[0:0] nor_489_nl;
  wire[0:0] and_322_nl;
  wire[0:0] mux_1006_nl;
  wire[0:0] mux_1005_nl;
  wire[0:0] mux_1004_nl;
  wire[0:0] nor_490_nl;
  wire[0:0] nor_491_nl;
  wire[0:0] mux_1003_nl;
  wire[0:0] nor_493_nl;
  wire[0:0] mux_1002_nl;
  wire[0:0] mux_1001_nl;
  wire[0:0] nor_494_nl;
  wire[0:0] and_432_nl;
  wire[0:0] nor_496_nl;
  wire[0:0] nor_497_nl;
  wire[0:0] mux_1000_nl;
  wire[0:0] nand_53_nl;
  wire[0:0] mux_999_nl;
  wire[0:0] mux_998_nl;
  wire[0:0] mux_997_nl;
  wire[0:0] nor_499_nl;
  wire[0:0] mux_996_nl;
  wire[0:0] nor_500_nl;
  wire[0:0] nor_501_nl;
  wire[0:0] nor_502_nl;
  wire[0:0] or_980_nl;
  wire[0:0] mux_995_nl;
  wire[0:0] or_979_nl;
  wire[0:0] mux_994_nl;
  wire[0:0] mux_993_nl;
  wire[0:0] nand_282_nl;
  wire[0:0] or_976_nl;
  wire[0:0] mux_992_nl;
  wire[0:0] nand_354_nl;
  wire[0:0] mux_1052_nl;
  wire[0:0] mux_1051_nl;
  wire[0:0] nor_478_nl;
  wire[0:0] mux_1050_nl;
  wire[0:0] nand_58_nl;
  wire[0:0] mux_1049_nl;
  wire[0:0] mux_1048_nl;
  wire[0:0] or_1069_nl;
  wire[0:0] mux_1047_nl;
  wire[0:0] or_1068_nl;
  wire[0:0] or_1067_nl;
  wire[0:0] mux_1046_nl;
  wire[0:0] nor_479_nl;
  wire[0:0] nor_480_nl;
  wire[0:0] mux_1045_nl;
  wire[0:0] or_1062_nl;
  wire[0:0] mux_1044_nl;
  wire[0:0] and_319_nl;
  wire[0:0] mux_1043_nl;
  wire[0:0] or_1059_nl;
  wire[0:0] mux_1042_nl;
  wire[0:0] mux_1041_nl;
  wire[0:0] mux_1040_nl;
  wire[0:0] or_1057_nl;
  wire[0:0] mux_1039_nl;
  wire[0:0] or_1055_nl;
  wire[0:0] or_1054_nl;
  wire[0:0] mux_1038_nl;
  wire[0:0] or_1053_nl;
  wire[0:0] nor_481_nl;
  wire[0:0] mux_1037_nl;
  wire[0:0] nor_482_nl;
  wire[0:0] mux_1036_nl;
  wire[0:0] mux_1035_nl;
  wire[0:0] or_1049_nl;
  wire[0:0] mux_1034_nl;
  wire[0:0] mux_1033_nl;
  wire[0:0] or_1047_nl;
  wire[0:0] mux_1032_nl;
  wire[0:0] or_1045_nl;
  wire[0:0] mux_1031_nl;
  wire[0:0] or_1044_nl;
  wire[0:0] mux_1030_nl;
  wire[0:0] or_1043_nl;
  wire[0:0] nor_483_nl;
  wire[0:0] mux_1029_nl;
  wire[0:0] nand_56_nl;
  wire[0:0] mux_1028_nl;
  wire[0:0] or_1040_nl;
  wire[0:0] mux_1027_nl;
  wire[0:0] mux_1026_nl;
  wire[0:0] or_1038_nl;
  wire[0:0] mux_1025_nl;
  wire[0:0] or_1032_nl;
  wire[0:0] or_1031_nl;
  wire[0:0] mux_1024_nl;
  wire[0:0] or_1030_nl;
  wire[0:0] mux_1023_nl;
  wire[0:0] or_1029_nl;
  wire[0:0] mux_1083_nl;
  wire[0:0] mux_1082_nl;
  wire[0:0] nor_458_nl;
  wire[0:0] mux_1081_nl;
  wire[0:0] mux_1080_nl;
  wire[0:0] or_1122_nl;
  wire[0:0] mux_1079_nl;
  wire[0:0] or_1121_nl;
  wire[0:0] mux_1078_nl;
  wire[0:0] mux_1077_nl;
  wire[0:0] or_1118_nl;
  wire[0:0] or_1116_nl;
  wire[0:0] mux_1076_nl;
  wire[0:0] or_1115_nl;
  wire[0:0] or_1113_nl;
  wire[0:0] mux_1075_nl;
  wire[0:0] nor_459_nl;
  wire[0:0] mux_1074_nl;
  wire[0:0] mux_1073_nl;
  wire[0:0] or_1111_nl;
  wire[0:0] or_1109_nl;
  wire[0:0] or_1108_nl;
  wire[0:0] nor_460_nl;
  wire[0:0] mux_1072_nl;
  wire[0:0] mux_1071_nl;
  wire[0:0] nor_461_nl;
  wire[0:0] and_317_nl;
  wire[0:0] mux_1070_nl;
  wire[0:0] nor_462_nl;
  wire[0:0] mux_1069_nl;
  wire[0:0] nor_463_nl;
  wire[0:0] nor_464_nl;
  wire[0:0] and_318_nl;
  wire[0:0] mux_1068_nl;
  wire[0:0] mux_1067_nl;
  wire[0:0] mux_1066_nl;
  wire[0:0] nor_465_nl;
  wire[0:0] nor_466_nl;
  wire[0:0] mux_1065_nl;
  wire[0:0] nor_468_nl;
  wire[0:0] mux_1064_nl;
  wire[0:0] mux_1063_nl;
  wire[0:0] nor_469_nl;
  wire[0:0] nor_470_nl;
  wire[0:0] nor_471_nl;
  wire[0:0] nor_472_nl;
  wire[0:0] mux_1062_nl;
  wire[0:0] nand_59_nl;
  wire[0:0] mux_1061_nl;
  wire[0:0] mux_1060_nl;
  wire[0:0] mux_1059_nl;
  wire[0:0] nor_474_nl;
  wire[0:0] mux_1058_nl;
  wire[0:0] nor_475_nl;
  wire[0:0] nor_476_nl;
  wire[0:0] nor_477_nl;
  wire[0:0] or_1079_nl;
  wire[0:0] mux_1057_nl;
  wire[0:0] or_1078_nl;
  wire[0:0] mux_1056_nl;
  wire[0:0] mux_1055_nl;
  wire[0:0] or_1076_nl;
  wire[0:0] or_1075_nl;
  wire[0:0] mux_1054_nl;
  wire[0:0] or_1072_nl;
  wire[0:0] mux_1114_nl;
  wire[0:0] mux_1113_nl;
  wire[0:0] mux_1112_nl;
  wire[0:0] nor_450_nl;
  wire[0:0] mux_1111_nl;
  wire[0:0] mux_1110_nl;
  wire[0:0] or_1169_nl;
  wire[0:0] mux_1109_nl;
  wire[0:0] or_1168_nl;
  wire[0:0] and_316_nl;
  wire[0:0] mux_1108_nl;
  wire[0:0] or_1166_nl;
  wire[0:0] mux_1107_nl;
  wire[0:0] mux_1106_nl;
  wire[0:0] or_1165_nl;
  wire[0:0] mux_1105_nl;
  wire[0:0] or_1164_nl;
  wire[0:0] nor_451_nl;
  wire[0:0] mux_1104_nl;
  wire[0:0] or_1161_nl;
  wire[0:0] nor_452_nl;
  wire[0:0] mux_1103_nl;
  wire[0:0] mux_1102_nl;
  wire[0:0] or_1158_nl;
  wire[0:0] or_1156_nl;
  wire[0:0] nand_62_nl;
  wire[0:0] mux_1101_nl;
  wire[0:0] or_1155_nl;
  wire[0:0] mux_1100_nl;
  wire[0:0] or_1154_nl;
  wire[0:0] mux_1099_nl;
  wire[0:0] mux_1098_nl;
  wire[0:0] nor_453_nl;
  wire[0:0] mux_1097_nl;
  wire[0:0] nor_454_nl;
  wire[0:0] nor_455_nl;
  wire[0:0] mux_1096_nl;
  wire[0:0] or_1148_nl;
  wire[0:0] mux_1095_nl;
  wire[0:0] or_1147_nl;
  wire[0:0] mux_1094_nl;
  wire[0:0] nor_456_nl;
  wire[0:0] mux_1093_nl;
  wire[0:0] or_1142_nl;
  wire[0:0] mux_1092_nl;
  wire[0:0] mux_1091_nl;
  wire[0:0] or_1141_nl;
  wire[0:0] mux_1090_nl;
  wire[0:0] or_1140_nl;
  wire[0:0] nor_457_nl;
  wire[0:0] mux_1089_nl;
  wire[0:0] mux_1088_nl;
  wire[0:0] mux_1087_nl;
  wire[0:0] or_1136_nl;
  wire[0:0] mux_1086_nl;
  wire[0:0] or_1131_nl;
  wire[0:0] or_1129_nl;
  wire[0:0] mux_1085_nl;
  wire[0:0] or_1128_nl;
  wire[0:0] mux_1145_nl;
  wire[0:0] mux_1144_nl;
  wire[0:0] nor_430_nl;
  wire[0:0] mux_1143_nl;
  wire[0:0] mux_1142_nl;
  wire[0:0] or_1221_nl;
  wire[0:0] mux_1141_nl;
  wire[0:0] or_1220_nl;
  wire[0:0] mux_1140_nl;
  wire[0:0] mux_1139_nl;
  wire[0:0] or_1217_nl;
  wire[0:0] or_1215_nl;
  wire[0:0] mux_1138_nl;
  wire[0:0] or_1214_nl;
  wire[0:0] or_1212_nl;
  wire[0:0] mux_1137_nl;
  wire[0:0] nor_431_nl;
  wire[0:0] mux_1136_nl;
  wire[0:0] mux_1135_nl;
  wire[0:0] or_1210_nl;
  wire[0:0] or_1208_nl;
  wire[0:0] or_1207_nl;
  wire[0:0] nor_432_nl;
  wire[0:0] mux_1134_nl;
  wire[0:0] mux_1133_nl;
  wire[0:0] nor_433_nl;
  wire[0:0] and_314_nl;
  wire[0:0] mux_1132_nl;
  wire[0:0] nor_434_nl;
  wire[0:0] mux_1131_nl;
  wire[0:0] nor_435_nl;
  wire[0:0] nor_436_nl;
  wire[0:0] and_315_nl;
  wire[0:0] mux_1130_nl;
  wire[0:0] mux_1129_nl;
  wire[0:0] mux_1128_nl;
  wire[0:0] nor_437_nl;
  wire[0:0] nor_438_nl;
  wire[0:0] mux_1127_nl;
  wire[0:0] nor_440_nl;
  wire[0:0] mux_1126_nl;
  wire[0:0] mux_1125_nl;
  wire[0:0] nor_441_nl;
  wire[0:0] nor_442_nl;
  wire[0:0] nor_443_nl;
  wire[0:0] nor_444_nl;
  wire[0:0] mux_1124_nl;
  wire[0:0] nand_65_nl;
  wire[0:0] mux_1123_nl;
  wire[0:0] mux_1122_nl;
  wire[0:0] mux_1121_nl;
  wire[0:0] nor_446_nl;
  wire[0:0] mux_1120_nl;
  wire[0:0] nor_447_nl;
  wire[0:0] nor_448_nl;
  wire[0:0] nor_449_nl;
  wire[0:0] or_1178_nl;
  wire[0:0] mux_1119_nl;
  wire[0:0] or_1177_nl;
  wire[0:0] mux_1118_nl;
  wire[0:0] mux_1117_nl;
  wire[0:0] or_1175_nl;
  wire[0:0] or_1174_nl;
  wire[0:0] mux_1116_nl;
  wire[0:0] or_1171_nl;
  wire[0:0] mux_1176_nl;
  wire[0:0] mux_1175_nl;
  wire[0:0] nor_424_nl;
  wire[0:0] mux_1174_nl;
  wire[0:0] nand_70_nl;
  wire[0:0] mux_1173_nl;
  wire[0:0] mux_1172_nl;
  wire[0:0] or_1267_nl;
  wire[0:0] mux_1171_nl;
  wire[0:0] or_1266_nl;
  wire[0:0] or_1265_nl;
  wire[0:0] mux_1170_nl;
  wire[0:0] and_442_nl;
  wire[0:0] nor_426_nl;
  wire[0:0] mux_1169_nl;
  wire[0:0] or_1260_nl;
  wire[0:0] mux_1168_nl;
  wire[0:0] and_313_nl;
  wire[0:0] mux_1167_nl;
  wire[0:0] or_1257_nl;
  wire[0:0] mux_1166_nl;
  wire[0:0] mux_1165_nl;
  wire[0:0] mux_1164_nl;
  wire[0:0] or_1255_nl;
  wire[0:0] mux_1163_nl;
  wire[0:0] or_1253_nl;
  wire[0:0] or_1252_nl;
  wire[0:0] mux_1162_nl;
  wire[0:0] or_1251_nl;
  wire[0:0] nor_427_nl;
  wire[0:0] mux_1161_nl;
  wire[0:0] nor_428_nl;
  wire[0:0] mux_1160_nl;
  wire[0:0] mux_1159_nl;
  wire[0:0] or_1247_nl;
  wire[0:0] mux_1158_nl;
  wire[0:0] mux_1157_nl;
  wire[0:0] or_1245_nl;
  wire[0:0] mux_1156_nl;
  wire[0:0] or_1243_nl;
  wire[0:0] mux_1155_nl;
  wire[0:0] or_1242_nl;
  wire[0:0] mux_1154_nl;
  wire[0:0] or_1241_nl;
  wire[0:0] nor_429_nl;
  wire[0:0] mux_1153_nl;
  wire[0:0] nand_68_nl;
  wire[0:0] mux_1152_nl;
  wire[0:0] or_1238_nl;
  wire[0:0] mux_1151_nl;
  wire[0:0] mux_1150_nl;
  wire[0:0] or_1236_nl;
  wire[0:0] mux_1149_nl;
  wire[0:0] or_1230_nl;
  wire[0:0] or_1229_nl;
  wire[0:0] mux_1148_nl;
  wire[0:0] or_1228_nl;
  wire[0:0] mux_1147_nl;
  wire[0:0] or_1227_nl;
  wire[0:0] mux_1207_nl;
  wire[0:0] mux_1206_nl;
  wire[0:0] nor_404_nl;
  wire[0:0] mux_1205_nl;
  wire[0:0] mux_1204_nl;
  wire[0:0] or_1320_nl;
  wire[0:0] mux_1203_nl;
  wire[0:0] or_1319_nl;
  wire[0:0] mux_1202_nl;
  wire[0:0] mux_1201_nl;
  wire[0:0] or_1316_nl;
  wire[0:0] or_1314_nl;
  wire[0:0] mux_1200_nl;
  wire[0:0] or_1313_nl;
  wire[0:0] or_1311_nl;
  wire[0:0] mux_1199_nl;
  wire[0:0] nor_405_nl;
  wire[0:0] mux_1198_nl;
  wire[0:0] mux_1197_nl;
  wire[0:0] or_1309_nl;
  wire[0:0] or_1307_nl;
  wire[0:0] or_1306_nl;
  wire[0:0] nor_406_nl;
  wire[0:0] mux_1196_nl;
  wire[0:0] mux_1195_nl;
  wire[0:0] nor_407_nl;
  wire[0:0] and_311_nl;
  wire[0:0] mux_1194_nl;
  wire[0:0] nor_408_nl;
  wire[0:0] mux_1193_nl;
  wire[0:0] nor_409_nl;
  wire[0:0] nor_410_nl;
  wire[0:0] and_312_nl;
  wire[0:0] mux_1192_nl;
  wire[0:0] mux_1191_nl;
  wire[0:0] mux_1190_nl;
  wire[0:0] nor_411_nl;
  wire[0:0] nor_412_nl;
  wire[0:0] mux_1189_nl;
  wire[0:0] nor_414_nl;
  wire[0:0] mux_1188_nl;
  wire[0:0] mux_1187_nl;
  wire[0:0] nor_415_nl;
  wire[0:0] nor_416_nl;
  wire[0:0] nor_417_nl;
  wire[0:0] nor_418_nl;
  wire[0:0] mux_1186_nl;
  wire[0:0] nand_71_nl;
  wire[0:0] mux_1185_nl;
  wire[0:0] mux_1184_nl;
  wire[0:0] mux_1183_nl;
  wire[0:0] nor_420_nl;
  wire[0:0] mux_1182_nl;
  wire[0:0] nor_421_nl;
  wire[0:0] nor_422_nl;
  wire[0:0] nor_423_nl;
  wire[0:0] or_1277_nl;
  wire[0:0] mux_1181_nl;
  wire[0:0] or_1276_nl;
  wire[0:0] mux_1180_nl;
  wire[0:0] mux_1179_nl;
  wire[0:0] or_1274_nl;
  wire[0:0] or_1273_nl;
  wire[0:0] mux_1178_nl;
  wire[0:0] or_1270_nl;
  wire[0:0] mux_1238_nl;
  wire[0:0] mux_1237_nl;
  wire[0:0] nor_398_nl;
  wire[0:0] mux_1236_nl;
  wire[0:0] nand_76_nl;
  wire[0:0] mux_1235_nl;
  wire[0:0] mux_1234_nl;
  wire[0:0] or_1366_nl;
  wire[0:0] mux_1233_nl;
  wire[0:0] or_1365_nl;
  wire[0:0] or_1364_nl;
  wire[0:0] mux_1232_nl;
  wire[0:0] and_441_nl;
  wire[0:0] nor_400_nl;
  wire[0:0] mux_1231_nl;
  wire[0:0] or_1359_nl;
  wire[0:0] mux_1230_nl;
  wire[0:0] and_310_nl;
  wire[0:0] mux_1229_nl;
  wire[0:0] nand_378_nl;
  wire[0:0] mux_1228_nl;
  wire[0:0] mux_1227_nl;
  wire[0:0] mux_1226_nl;
  wire[0:0] or_1354_nl;
  wire[0:0] mux_1225_nl;
  wire[0:0] or_1352_nl;
  wire[0:0] or_1351_nl;
  wire[0:0] mux_1224_nl;
  wire[0:0] or_1350_nl;
  wire[0:0] nor_401_nl;
  wire[0:0] mux_1223_nl;
  wire[0:0] nor_402_nl;
  wire[0:0] mux_1222_nl;
  wire[0:0] mux_1221_nl;
  wire[0:0] nand_373_nl;
  wire[0:0] mux_1220_nl;
  wire[0:0] mux_1219_nl;
  wire[0:0] or_1344_nl;
  wire[0:0] mux_1218_nl;
  wire[0:0] or_1342_nl;
  wire[0:0] mux_1217_nl;
  wire[0:0] or_1341_nl;
  wire[0:0] mux_1216_nl;
  wire[0:0] or_1340_nl;
  wire[0:0] nor_403_nl;
  wire[0:0] mux_1215_nl;
  wire[0:0] nand_74_nl;
  wire[0:0] mux_1214_nl;
  wire[0:0] nand_363_nl;
  wire[0:0] mux_1213_nl;
  wire[0:0] mux_1212_nl;
  wire[0:0] or_1335_nl;
  wire[0:0] mux_1211_nl;
  wire[0:0] or_1329_nl;
  wire[0:0] or_1328_nl;
  wire[0:0] mux_1210_nl;
  wire[0:0] or_1327_nl;
  wire[0:0] mux_1209_nl;
  wire[0:0] or_1326_nl;
  wire[0:0] mux_1269_nl;
  wire[0:0] mux_1268_nl;
  wire[0:0] nor_379_nl;
  wire[0:0] mux_1267_nl;
  wire[0:0] mux_1266_nl;
  wire[0:0] nand_240_nl;
  wire[0:0] mux_1265_nl;
  wire[0:0] or_1418_nl;
  wire[0:0] mux_1264_nl;
  wire[0:0] mux_1263_nl;
  wire[0:0] or_1415_nl;
  wire[0:0] or_1413_nl;
  wire[0:0] mux_1262_nl;
  wire[0:0] nand_369_nl;
  wire[0:0] or_1410_nl;
  wire[0:0] mux_1261_nl;
  wire[0:0] nor_380_nl;
  wire[0:0] mux_1260_nl;
  wire[0:0] mux_1259_nl;
  wire[0:0] or_1408_nl;
  wire[0:0] or_1406_nl;
  wire[0:0] or_1405_nl;
  wire[0:0] nor_381_nl;
  wire[0:0] mux_1258_nl;
  wire[0:0] mux_1257_nl;
  wire[0:0] nor_382_nl;
  wire[0:0] and_307_nl;
  wire[0:0] mux_1256_nl;
  wire[0:0] nor_383_nl;
  wire[0:0] mux_1255_nl;
  wire[0:0] and_308_nl;
  wire[0:0] nor_384_nl;
  wire[0:0] and_309_nl;
  wire[0:0] mux_1254_nl;
  wire[0:0] mux_1253_nl;
  wire[0:0] mux_1252_nl;
  wire[0:0] nor_385_nl;
  wire[0:0] nor_386_nl;
  wire[0:0] mux_1251_nl;
  wire[0:0] nor_388_nl;
  wire[0:0] mux_1250_nl;
  wire[0:0] mux_1249_nl;
  wire[0:0] nor_389_nl;
  wire[0:0] and_431_nl;
  wire[0:0] nor_391_nl;
  wire[0:0] nor_392_nl;
  wire[0:0] mux_1248_nl;
  wire[0:0] nand_77_nl;
  wire[0:0] mux_1247_nl;
  wire[0:0] mux_1246_nl;
  wire[0:0] mux_1245_nl;
  wire[0:0] nor_394_nl;
  wire[0:0] mux_1244_nl;
  wire[0:0] nor_395_nl;
  wire[0:0] nor_396_nl;
  wire[0:0] nor_397_nl;
  wire[0:0] or_1376_nl;
  wire[0:0] mux_1243_nl;
  wire[0:0] or_1375_nl;
  wire[0:0] mux_1242_nl;
  wire[0:0] mux_1241_nl;
  wire[0:0] nand_248_nl;
  wire[0:0] or_1372_nl;
  wire[0:0] mux_1240_nl;
  wire[0:0] nand_352_nl;
  wire[0:0] mux_1300_nl;
  wire[0:0] mux_1299_nl;
  wire[0:0] nor_373_nl;
  wire[0:0] mux_1298_nl;
  wire[0:0] nand_82_nl;
  wire[0:0] mux_1297_nl;
  wire[0:0] mux_1296_nl;
  wire[0:0] or_1465_nl;
  wire[0:0] mux_1295_nl;
  wire[0:0] or_1464_nl;
  wire[0:0] or_1463_nl;
  wire[0:0] mux_1294_nl;
  wire[0:0] and_436_nl;
  wire[0:0] nor_375_nl;
  wire[0:0] mux_1293_nl;
  wire[0:0] or_1458_nl;
  wire[0:0] mux_1292_nl;
  wire[0:0] and_306_nl;
  wire[0:0] mux_1291_nl;
  wire[0:0] or_1455_nl;
  wire[0:0] mux_1290_nl;
  wire[0:0] mux_1289_nl;
  wire[0:0] mux_1288_nl;
  wire[0:0] or_1453_nl;
  wire[0:0] mux_1287_nl;
  wire[0:0] or_1451_nl;
  wire[0:0] or_1450_nl;
  wire[0:0] mux_1286_nl;
  wire[0:0] or_1449_nl;
  wire[0:0] nor_376_nl;
  wire[0:0] mux_1285_nl;
  wire[0:0] nor_377_nl;
  wire[0:0] mux_1284_nl;
  wire[0:0] mux_1283_nl;
  wire[0:0] or_1445_nl;
  wire[0:0] mux_1282_nl;
  wire[0:0] mux_1281_nl;
  wire[0:0] or_1443_nl;
  wire[0:0] mux_1280_nl;
  wire[0:0] or_1441_nl;
  wire[0:0] mux_1279_nl;
  wire[0:0] or_1440_nl;
  wire[0:0] mux_1278_nl;
  wire[0:0] or_1439_nl;
  wire[0:0] nor_378_nl;
  wire[0:0] mux_1277_nl;
  wire[0:0] nand_80_nl;
  wire[0:0] mux_1276_nl;
  wire[0:0] or_1436_nl;
  wire[0:0] mux_1275_nl;
  wire[0:0] mux_1274_nl;
  wire[0:0] or_1434_nl;
  wire[0:0] mux_1273_nl;
  wire[0:0] or_1428_nl;
  wire[0:0] or_1427_nl;
  wire[0:0] mux_1272_nl;
  wire[0:0] or_1426_nl;
  wire[0:0] mux_1271_nl;
  wire[0:0] or_1425_nl;
  wire[0:0] mux_1331_nl;
  wire[0:0] mux_1330_nl;
  wire[0:0] nor_353_nl;
  wire[0:0] mux_1329_nl;
  wire[0:0] mux_1328_nl;
  wire[0:0] or_1518_nl;
  wire[0:0] mux_1327_nl;
  wire[0:0] or_1517_nl;
  wire[0:0] mux_1326_nl;
  wire[0:0] mux_1325_nl;
  wire[0:0] or_1514_nl;
  wire[0:0] or_1512_nl;
  wire[0:0] mux_1324_nl;
  wire[0:0] or_1511_nl;
  wire[0:0] or_1509_nl;
  wire[0:0] mux_1323_nl;
  wire[0:0] nor_354_nl;
  wire[0:0] mux_1322_nl;
  wire[0:0] mux_1321_nl;
  wire[0:0] or_1507_nl;
  wire[0:0] or_1505_nl;
  wire[0:0] or_1504_nl;
  wire[0:0] nor_355_nl;
  wire[0:0] mux_1320_nl;
  wire[0:0] mux_1319_nl;
  wire[0:0] nor_356_nl;
  wire[0:0] and_304_nl;
  wire[0:0] mux_1318_nl;
  wire[0:0] nor_357_nl;
  wire[0:0] mux_1317_nl;
  wire[0:0] nor_358_nl;
  wire[0:0] nor_359_nl;
  wire[0:0] and_305_nl;
  wire[0:0] mux_1316_nl;
  wire[0:0] mux_1315_nl;
  wire[0:0] mux_1314_nl;
  wire[0:0] nor_360_nl;
  wire[0:0] nor_361_nl;
  wire[0:0] mux_1313_nl;
  wire[0:0] nor_363_nl;
  wire[0:0] mux_1312_nl;
  wire[0:0] mux_1311_nl;
  wire[0:0] nor_364_nl;
  wire[0:0] nor_365_nl;
  wire[0:0] nor_366_nl;
  wire[0:0] nor_367_nl;
  wire[0:0] mux_1310_nl;
  wire[0:0] nand_83_nl;
  wire[0:0] mux_1309_nl;
  wire[0:0] mux_1308_nl;
  wire[0:0] mux_1307_nl;
  wire[0:0] nor_369_nl;
  wire[0:0] mux_1306_nl;
  wire[0:0] nor_370_nl;
  wire[0:0] nor_371_nl;
  wire[0:0] nor_372_nl;
  wire[0:0] or_1475_nl;
  wire[0:0] mux_1305_nl;
  wire[0:0] or_1474_nl;
  wire[0:0] mux_1304_nl;
  wire[0:0] mux_1303_nl;
  wire[0:0] or_1472_nl;
  wire[0:0] or_1471_nl;
  wire[0:0] mux_1302_nl;
  wire[0:0] or_1468_nl;
  wire[0:0] mux_1362_nl;
  wire[0:0] mux_1361_nl;
  wire[0:0] mux_1360_nl;
  wire[0:0] nor_346_nl;
  wire[0:0] mux_1359_nl;
  wire[0:0] mux_1358_nl;
  wire[0:0] or_1565_nl;
  wire[0:0] mux_1357_nl;
  wire[0:0] or_1564_nl;
  wire[0:0] and_302_nl;
  wire[0:0] mux_1356_nl;
  wire[0:0] nand_230_nl;
  wire[0:0] mux_1355_nl;
  wire[0:0] mux_1354_nl;
  wire[0:0] or_1561_nl;
  wire[0:0] mux_1353_nl;
  wire[0:0] or_1560_nl;
  wire[0:0] nor_347_nl;
  wire[0:0] mux_1352_nl;
  wire[0:0] or_1557_nl;
  wire[0:0] nor_348_nl;
  wire[0:0] mux_1351_nl;
  wire[0:0] mux_1350_nl;
  wire[0:0] or_1554_nl;
  wire[0:0] nand_231_nl;
  wire[0:0] nand_86_nl;
  wire[0:0] mux_1349_nl;
  wire[0:0] or_1551_nl;
  wire[0:0] mux_1348_nl;
  wire[0:0] or_1550_nl;
  wire[0:0] mux_1347_nl;
  wire[0:0] mux_1346_nl;
  wire[0:0] nor_349_nl;
  wire[0:0] mux_1345_nl;
  wire[0:0] and_303_nl;
  wire[0:0] nor_350_nl;
  wire[0:0] mux_1344_nl;
  wire[0:0] or_1544_nl;
  wire[0:0] mux_1343_nl;
  wire[0:0] or_1543_nl;
  wire[0:0] mux_1342_nl;
  wire[0:0] nor_351_nl;
  wire[0:0] mux_1341_nl;
  wire[0:0] nand_232_nl;
  wire[0:0] mux_1340_nl;
  wire[0:0] mux_1339_nl;
  wire[0:0] or_1537_nl;
  wire[0:0] mux_1338_nl;
  wire[0:0] or_1536_nl;
  wire[0:0] nor_352_nl;
  wire[0:0] mux_1337_nl;
  wire[0:0] mux_1336_nl;
  wire[0:0] mux_1335_nl;
  wire[0:0] or_1532_nl;
  wire[0:0] mux_1334_nl;
  wire[0:0] or_1527_nl;
  wire[0:0] or_1525_nl;
  wire[0:0] mux_1333_nl;
  wire[0:0] or_1524_nl;
  wire[0:0] mux_1393_nl;
  wire[0:0] mux_1392_nl;
  wire[0:0] nor_327_nl;
  wire[0:0] mux_1391_nl;
  wire[0:0] mux_1390_nl;
  wire[0:0] nand_216_nl;
  wire[0:0] mux_1389_nl;
  wire[0:0] or_1615_nl;
  wire[0:0] mux_1388_nl;
  wire[0:0] mux_1387_nl;
  wire[0:0] or_1612_nl;
  wire[0:0] or_1611_nl;
  wire[0:0] mux_1386_nl;
  wire[0:0] nand_368_nl;
  wire[0:0] or_1608_nl;
  wire[0:0] mux_1385_nl;
  wire[0:0] nor_328_nl;
  wire[0:0] mux_1384_nl;
  wire[0:0] mux_1383_nl;
  wire[0:0] or_1606_nl;
  wire[0:0] or_1604_nl;
  wire[0:0] or_1603_nl;
  wire[0:0] nor_329_nl;
  wire[0:0] mux_1382_nl;
  wire[0:0] mux_1381_nl;
  wire[0:0] nor_330_nl;
  wire[0:0] and_299_nl;
  wire[0:0] mux_1380_nl;
  wire[0:0] nor_331_nl;
  wire[0:0] mux_1379_nl;
  wire[0:0] and_300_nl;
  wire[0:0] nor_332_nl;
  wire[0:0] and_301_nl;
  wire[0:0] mux_1378_nl;
  wire[0:0] mux_1377_nl;
  wire[0:0] mux_1376_nl;
  wire[0:0] nor_333_nl;
  wire[0:0] nor_334_nl;
  wire[0:0] mux_1375_nl;
  wire[0:0] nor_336_nl;
  wire[0:0] mux_1374_nl;
  wire[0:0] mux_1373_nl;
  wire[0:0] nor_337_nl;
  wire[0:0] and_430_nl;
  wire[0:0] nor_339_nl;
  wire[0:0] nor_340_nl;
  wire[0:0] mux_1372_nl;
  wire[0:0] nand_89_nl;
  wire[0:0] mux_1371_nl;
  wire[0:0] mux_1370_nl;
  wire[0:0] mux_1369_nl;
  wire[0:0] nor_342_nl;
  wire[0:0] mux_1368_nl;
  wire[0:0] nor_343_nl;
  wire[0:0] nor_344_nl;
  wire[0:0] nor_345_nl;
  wire[0:0] or_1574_nl;
  wire[0:0] mux_1367_nl;
  wire[0:0] or_1573_nl;
  wire[0:0] mux_1366_nl;
  wire[0:0] mux_1365_nl;
  wire[0:0] nand_224_nl;
  wire[0:0] or_1570_nl;
  wire[0:0] mux_1364_nl;
  wire[0:0] nand_351_nl;
  wire[0:0] mux_1424_nl;
  wire[0:0] mux_1423_nl;
  wire[0:0] nor_321_nl;
  wire[0:0] mux_1422_nl;
  wire[0:0] nand_94_nl;
  wire[0:0] mux_1421_nl;
  wire[0:0] mux_1420_nl;
  wire[0:0] or_1662_nl;
  wire[0:0] mux_1419_nl;
  wire[0:0] or_1661_nl;
  wire[0:0] or_1660_nl;
  wire[0:0] mux_1418_nl;
  wire[0:0] and_435_nl;
  wire[0:0] nor_323_nl;
  wire[0:0] mux_1417_nl;
  wire[0:0] or_1655_nl;
  wire[0:0] mux_1416_nl;
  wire[0:0] and_298_nl;
  wire[0:0] mux_1415_nl;
  wire[0:0] nand_375_nl;
  wire[0:0] mux_1414_nl;
  wire[0:0] mux_1413_nl;
  wire[0:0] mux_1412_nl;
  wire[0:0] or_1650_nl;
  wire[0:0] mux_1411_nl;
  wire[0:0] or_1648_nl;
  wire[0:0] or_1647_nl;
  wire[0:0] mux_1410_nl;
  wire[0:0] or_1646_nl;
  wire[0:0] nor_324_nl;
  wire[0:0] mux_1409_nl;
  wire[0:0] nor_325_nl;
  wire[0:0] mux_1408_nl;
  wire[0:0] mux_1407_nl;
  wire[0:0] nand_367_nl;
  wire[0:0] mux_1406_nl;
  wire[0:0] mux_1405_nl;
  wire[0:0] or_1640_nl;
  wire[0:0] mux_1404_nl;
  wire[0:0] or_1638_nl;
  wire[0:0] mux_1403_nl;
  wire[0:0] or_1637_nl;
  wire[0:0] mux_1402_nl;
  wire[0:0] or_1636_nl;
  wire[0:0] nor_326_nl;
  wire[0:0] mux_1401_nl;
  wire[0:0] nand_92_nl;
  wire[0:0] mux_1400_nl;
  wire[0:0] nand_359_nl;
  wire[0:0] mux_1399_nl;
  wire[0:0] mux_1398_nl;
  wire[0:0] or_1631_nl;
  wire[0:0] mux_1397_nl;
  wire[0:0] or_1625_nl;
  wire[0:0] or_1624_nl;
  wire[0:0] mux_1396_nl;
  wire[0:0] or_1623_nl;
  wire[0:0] mux_1395_nl;
  wire[0:0] or_1622_nl;
  wire[0:0] mux_1455_nl;
  wire[0:0] mux_1454_nl;
  wire[0:0] nor_302_nl;
  wire[0:0] mux_1453_nl;
  wire[0:0] mux_1452_nl;
  wire[0:0] nand_196_nl;
  wire[0:0] mux_1451_nl;
  wire[0:0] or_1712_nl;
  wire[0:0] mux_1450_nl;
  wire[0:0] mux_1449_nl;
  wire[0:0] or_1709_nl;
  wire[0:0] or_1707_nl;
  wire[0:0] mux_1448_nl;
  wire[0:0] nand_366_nl;
  wire[0:0] or_1704_nl;
  wire[0:0] mux_1447_nl;
  wire[0:0] nor_303_nl;
  wire[0:0] mux_1446_nl;
  wire[0:0] mux_1445_nl;
  wire[0:0] or_1702_nl;
  wire[0:0] or_1700_nl;
  wire[0:0] or_1699_nl;
  wire[0:0] nor_304_nl;
  wire[0:0] mux_1444_nl;
  wire[0:0] mux_1443_nl;
  wire[0:0] nor_305_nl;
  wire[0:0] and_295_nl;
  wire[0:0] mux_1442_nl;
  wire[0:0] nor_306_nl;
  wire[0:0] mux_1441_nl;
  wire[0:0] and_296_nl;
  wire[0:0] nor_307_nl;
  wire[0:0] and_297_nl;
  wire[0:0] mux_1440_nl;
  wire[0:0] mux_1439_nl;
  wire[0:0] mux_1438_nl;
  wire[0:0] nor_308_nl;
  wire[0:0] nor_309_nl;
  wire[0:0] mux_1437_nl;
  wire[0:0] nor_311_nl;
  wire[0:0] mux_1436_nl;
  wire[0:0] mux_1435_nl;
  wire[0:0] nor_312_nl;
  wire[0:0] and_429_nl;
  wire[0:0] nor_314_nl;
  wire[0:0] nor_315_nl;
  wire[0:0] mux_1434_nl;
  wire[0:0] nand_95_nl;
  wire[0:0] mux_1433_nl;
  wire[0:0] mux_1432_nl;
  wire[0:0] mux_1431_nl;
  wire[0:0] nor_317_nl;
  wire[0:0] mux_1430_nl;
  wire[0:0] nor_318_nl;
  wire[0:0] nor_319_nl;
  wire[0:0] nor_320_nl;
  wire[0:0] or_1671_nl;
  wire[0:0] mux_1429_nl;
  wire[0:0] or_1670_nl;
  wire[0:0] mux_1428_nl;
  wire[0:0] mux_1427_nl;
  wire[0:0] nand_204_nl;
  wire[0:0] or_1667_nl;
  wire[0:0] mux_1426_nl;
  wire[0:0] nand_350_nl;
  wire[0:0] mux_1486_nl;
  wire[0:0] mux_1485_nl;
  wire[0:0] nor_296_nl;
  wire[0:0] mux_1484_nl;
  wire[0:0] nand_100_nl;
  wire[0:0] mux_1483_nl;
  wire[0:0] mux_1482_nl;
  wire[0:0] or_1756_nl;
  wire[0:0] mux_1481_nl;
  wire[0:0] nand_178_nl;
  wire[0:0] or_1754_nl;
  wire[0:0] mux_1480_nl;
  wire[0:0] and_434_nl;
  wire[0:0] nor_298_nl;
  wire[0:0] mux_1479_nl;
  wire[0:0] nand_377_nl;
  wire[0:0] mux_1478_nl;
  wire[0:0] and_294_nl;
  wire[0:0] mux_1477_nl;
  wire[0:0] nand_374_nl;
  wire[0:0] mux_1476_nl;
  wire[0:0] mux_1475_nl;
  wire[0:0] mux_1474_nl;
  wire[0:0] nand_372_nl;
  wire[0:0] mux_1473_nl;
  wire[0:0] nand_183_nl;
  wire[0:0] or_1741_nl;
  wire[0:0] mux_1472_nl;
  wire[0:0] nand_184_nl;
  wire[0:0] nor_299_nl;
  wire[0:0] mux_1471_nl;
  wire[0:0] nor_300_nl;
  wire[0:0] mux_1470_nl;
  wire[0:0] mux_1469_nl;
  wire[0:0] nand_365_nl;
  wire[0:0] mux_1468_nl;
  wire[0:0] mux_1467_nl;
  wire[0:0] nand_362_nl;
  wire[0:0] mux_1466_nl;
  wire[0:0] nand_187_nl;
  wire[0:0] mux_1465_nl;
  wire[0:0] or_1731_nl;
  wire[0:0] mux_1464_nl;
  wire[0:0] nand_188_nl;
  wire[0:0] nor_301_nl;
  wire[0:0] mux_1463_nl;
  wire[0:0] nand_98_nl;
  wire[0:0] mux_1462_nl;
  wire[0:0] nand_358_nl;
  wire[0:0] mux_1461_nl;
  wire[0:0] mux_1460_nl;
  wire[0:0] nand_349_nl;
  wire[0:0] mux_1459_nl;
  wire[0:0] nand_191_nl;
  wire[0:0] or_1721_nl;
  wire[0:0] mux_1458_nl;
  wire[0:0] or_1720_nl;
  wire[0:0] mux_1457_nl;
  wire[0:0] nand_192_nl;
  wire[0:0] mux_1517_nl;
  wire[0:0] mux_1516_nl;
  wire[0:0] nor_282_nl;
  wire[0:0] mux_1515_nl;
  wire[0:0] mux_1514_nl;
  wire[0:0] nand_158_nl;
  wire[0:0] mux_1513_nl;
  wire[0:0] or_1802_nl;
  wire[0:0] mux_1512_nl;
  wire[0:0] mux_1511_nl;
  wire[0:0] nand_162_nl;
  wire[0:0] mux_1510_nl;
  wire[0:0] nand_364_nl;
  wire[0:0] or_1796_nl;
  wire[0:0] mux_1509_nl;
  wire[0:0] nor_283_nl;
  wire[0:0] mux_1508_nl;
  wire[0:0] mux_1507_nl;
  wire[0:0] nand_361_nl;
  wire[0:0] nand_164_nl;
  wire[0:0] or_1791_nl;
  wire[0:0] nor_284_nl;
  wire[0:0] mux_1506_nl;
  wire[0:0] mux_1505_nl;
  wire[0:0] nor_285_nl;
  wire[0:0] and_286_nl;
  wire[0:0] mux_1504_nl;
  wire[0:0] nor_286_nl;
  wire[0:0] mux_1503_nl;
  wire[0:0] and_287_nl;
  wire[0:0] and_288_nl;
  wire[0:0] and_289_nl;
  wire[0:0] mux_1502_nl;
  wire[0:0] mux_1501_nl;
  wire[0:0] mux_1500_nl;
  wire[0:0] and_290_nl;
  wire[0:0] nor_287_nl;
  wire[0:0] mux_1499_nl;
  wire[0:0] and_427_nl;
  wire[0:0] mux_1498_nl;
  wire[0:0] mux_1497_nl;
  wire[0:0] and_292_nl;
  wire[0:0] and_428_nl;
  wire[0:0] nor_290_nl;
  wire[0:0] nor_291_nl;
  wire[0:0] mux_1496_nl;
  wire[0:0] nand_101_nl;
  wire[0:0] mux_1495_nl;
  wire[0:0] mux_1494_nl;
  wire[0:0] mux_1493_nl;
  wire[0:0] and_433_nl;
  wire[0:0] mux_1492_nl;
  wire[0:0] nor_293_nl;
  wire[0:0] and_440_nl;
  wire[0:0] nor_295_nl;
  wire[0:0] or_1764_nl;
  wire[0:0] mux_1491_nl;
  wire[0:0] or_1763_nl;
  wire[0:0] mux_1490_nl;
  wire[0:0] mux_1489_nl;
  wire[0:0] nand_172_nl;
  wire[0:0] mux_1488_nl;
  wire[0:0] nand_348_nl;
  wire[0:0] or_2213_nl;
  wire[0:0] mux_2057_nl;
  wire[0:0] mux_2065_nl;
  wire[0:0] mux_2064_nl;
  wire[0:0] or_2219_nl;
  wire[0:0] mux_2063_nl;
  wire[0:0] or_2218_nl;
  wire[0:0] mux_2062_nl;
  wire[0:0] mux_2061_nl;
  wire[0:0] or_2214_nl;
  wire[0:0] mux_2060_nl;
  wire[0:0] mux_2059_nl;
  wire[0:0] or_2209_nl;
  wire[0:0] or_2208_nl;
  wire[0:0] mux_2056_nl;
  wire[0:0] or_2207_nl;
  wire[0:0] mux_2055_nl;
  wire[0:0] or_2261_nl;
  wire[0:0] or_2267_nl;
  wire[0:0] or_2266_nl;
  wire[0:0] mux_2097_nl;
  wire[0:0] or_2271_nl;
  wire[0:0] or_2270_nl;
  wire[0:0] nand_388_nl;
  wire[0:0] mux_2103_nl;
  wire[0:0] nand_389_nl;
  wire[0:0] mux_2102_nl;
  wire[0:0] mux_2101_nl;
  wire[0:0] or_2272_nl;
  wire[0:0] or_2282_nl;
  wire[0:0] mux_2123_nl;
  wire[0:0] or_2302_nl;
  wire[0:0] mux_2134_nl;
  wire[0:0] mux_2132_nl;
  wire[0:0] mux_2131_nl;
  wire[0:0] mux_2163_nl;
  wire[0:0] mux_2170_nl;
  wire[0:0] mux_2169_nl;
  wire[0:0] mux_2167_nl;
  wire[0:0] mux_2166_nl;
  wire[0:0] mux_2175_nl;
  wire[0:0] mux_2179_nl;
  wire[0:0] or_2346_nl;
  wire[0:0] mux_2215_nl;
  wire[0:0] mux_2220_nl;
  wire[0:0] or_2350_nl;
  wire[0:0] nand_399_nl;
  wire[0:0] or_2360_nl;
  wire[10:0] acc_nl;
  wire[11:0] nl_acc_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_3_nl;
  wire[8:0] COMP_LOOP_COMP_LOOP_mux_15_nl;
  wire[0:0] COMP_LOOP_or_52_nl;
  wire[0:0] COMP_LOOP_or_53_nl;
  wire[3:0] COMP_LOOP_mux1h_271_nl;
  wire[0:0] COMP_LOOP_or_54_nl;
  wire[8:0] acc_1_nl;
  wire[9:0] nl_acc_1_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_4_nl;
  wire[6:0] COMP_LOOP_COMP_LOOP_mux_16_nl;
  wire[0:0] COMP_LOOP_or_55_nl;
  wire[0:0] COMP_LOOP_or_56_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_5_nl;
  wire[4:0] operator_64_false_1_mux_1_nl;
  wire[6:0] acc_3_nl;
  wire[7:0] nl_acc_3_nl;
  wire[5:0] COMP_LOOP_mux_35_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_nand_1_nl;
  wire[7:0] acc_4_nl;
  wire[8:0] nl_acc_4_nl;
  wire[6:0] COMP_LOOP_mux_36_nl;
  wire[0:0] COMP_LOOP_or_57_nl;
  wire[10:0] acc_5_nl;
  wire[12:0] nl_acc_5_nl;
  wire[3:0] COMP_LOOP_or_58_nl;
  wire[3:0] COMP_LOOP_COMP_LOOP_nor_63_nl;
  wire[3:0] COMP_LOOP_mux1h_272_nl;
  wire[0:0] and_706_nl;
  wire[0:0] and_707_nl;
  wire[0:0] and_708_nl;
  wire[0:0] and_709_nl;
  wire[0:0] and_710_nl;
  wire[0:0] and_711_nl;
  wire[0:0] and_712_nl;
  wire[0:0] and_713_nl;
  wire[0:0] and_714_nl;
  wire[0:0] and_715_nl;
  wire[0:0] and_716_nl;
  wire[0:0] and_717_nl;
  wire[0:0] and_718_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_or_1_nl;
  wire[63:0] STAGE_LOOP_STAGE_LOOP_mux_2_nl;
  wire[0:0] STAGE_LOOP_or_2_nl;
  wire[64:0] operator_64_false_acc_nl;
  wire[65:0] nl_operator_64_false_acc_nl;
  wire[60:0] operator_64_false_operator_64_false_operator_64_false_nor_1_nl;
  wire[2:0] operator_64_false_mux_1_nl;
  wire[63:0] operator_64_false_mux1h_1_nl;
  wire[0:0] and_719_nl;
  wire[0:0] and_720_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[63:0] COMP_LOOP_1_acc_5_nl;
  wire[64:0] nl_COMP_LOOP_1_acc_5_nl;
  wire[0:0] mux_1600_nl;
  wire[0:0] mux_1599_nl;
  wire[0:0] mux_1598_nl;
  wire[0:0] and_275_nl;
  wire[0:0] mux_1597_nl;
  wire[0:0] mux_1596_nl;
  wire[0:0] nor_277_nl;
  wire[0:0] mux_1595_nl;
  wire[0:0] mux_1594_nl;
  wire[0:0] mux_1593_nl;
  wire[0:0] nor_278_nl;
  wire[0:0] and_276_nl;
  wire[0:0] mux_1592_nl;
  wire[0:0] and_277_nl;
  wire[0:0] mux_1591_nl;
  wire[0:0] mux_1590_nl;
  wire[0:0] mux_1589_nl;
  wire[0:0] nor_279_nl;
  wire[0:0] mux_1586_nl;
  wire[0:0] mux_1582_nl;
  wire[0:0] or_1816_nl;
  wire[0:0] COMP_LOOP_or_22_nl;
  wire [63:0] nl_modulo_dev_cmp_base_rsc_dat;
  assign nl_COMP_LOOP_1_acc_5_nl = tmp_10_lpi_4_dfm + modulo_dev_cmp_return_rsc_z;
  assign COMP_LOOP_1_acc_5_nl = nl_COMP_LOOP_1_acc_5_nl[63:0];
  assign mux_1596_nl = MUX_s_1_2_2(or_tmp_1794, or_tmp_1793, fsm_output[6]);
  assign mux_1597_nl = MUX_s_1_2_2(or_tmp_1799, mux_1596_nl, fsm_output[2]);
  assign and_275_nl = (fsm_output[4]) & (~ mux_1597_nl);
  assign mux_1594_nl = MUX_s_1_2_2(or_tmp_1788, or_tmp_1796, fsm_output[6]);
  assign mux_1595_nl = MUX_s_1_2_2(or_2306_cse, mux_1594_nl, fsm_output[2]);
  assign nor_277_nl = ~((fsm_output[4]) | mux_1595_nl);
  assign mux_1598_nl = MUX_s_1_2_2(and_275_nl, nor_277_nl, fsm_output[5]);
  assign nor_278_nl = ~((fsm_output[4]) | mux_tmp_1537);
  assign and_276_nl = (fsm_output[4]) & (~ mux_tmp_1534);
  assign mux_1593_nl = MUX_s_1_2_2(nor_278_nl, and_276_nl, fsm_output[5]);
  assign mux_1599_nl = MUX_s_1_2_2(mux_1598_nl, mux_1593_nl, fsm_output[1]);
  assign mux_1589_nl = MUX_s_1_2_2(or_tmp_1799, or_tmp_1794, fsm_output[6]);
  assign mux_1590_nl = MUX_s_1_2_2(mux_1589_nl, or_tmp_1793, fsm_output[2]);
  assign mux_1591_nl = MUX_s_1_2_2(mux_1590_nl, mux_tmp_1537, fsm_output[4]);
  assign and_277_nl = (fsm_output[5]) & (~ mux_1591_nl);
  assign or_1816_nl = (fsm_output[6]) | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9])
      | (fsm_output[8]);
  assign mux_1582_nl = MUX_s_1_2_2(or_tmp_1788, or_1816_nl, fsm_output[2]);
  assign mux_1586_nl = MUX_s_1_2_2(mux_tmp_1534, mux_1582_nl, fsm_output[4]);
  assign nor_279_nl = ~((fsm_output[5]) | mux_1586_nl);
  assign mux_1592_nl = MUX_s_1_2_2(and_277_nl, nor_279_nl, fsm_output[1]);
  assign mux_1600_nl = MUX_s_1_2_2(mux_1599_nl, mux_1592_nl, fsm_output[0]);
  assign COMP_LOOP_or_22_nl = (and_dcpl_35 & and_dcpl_122) | (and_dcpl_30 & and_dcpl_65)
      | (and_dcpl_51 & and_dcpl_28) | (and_dcpl_57 & and_dcpl_28) | (and_dcpl_55
      & and_dcpl_39) | (and_dcpl_30 & and_dcpl_91) | (and_dcpl_40 & and_dcpl_130)
      | (and_dcpl_45 & and_dcpl_130) | (and_dcpl_89 & and_dcpl_73) | (and_dcpl_87
      & and_dcpl_83) | (and_dcpl_68 & and_dcpl_79) | (and_dcpl_75 & and_dcpl_136)
      | (and_dcpl_81 & and_dcpl_138) | (and_dcpl_87 & and_dcpl_101) | (and_dcpl_68
      & and_dcpl_99) | (and_dcpl_95 & and_dcpl_103);
  assign nl_modulo_dev_cmp_base_rsc_dat = MUX1HOT_v_64_3_2(operator_64_false_acc_mut_63_0,
      COMP_LOOP_1_mul_itm, COMP_LOOP_1_acc_5_nl, {mux_1600_nl , COMP_LOOP_or_22_nl
      , not_tmp_370});
  wire [63:0] nl_modulo_dev_cmp_m_rsc_dat;
  assign nl_modulo_dev_cmp_m_rsc_dat = p_sva;
  wire[0:0] mux_1659_nl;
  wire[0:0] mux_1658_nl;
  wire[0:0] mux_1657_nl;
  wire[0:0] mux_1656_nl;
  wire[0:0] mux_1655_nl;
  wire[0:0] or_1873_nl;
  wire[0:0] mux_1654_nl;
  wire[0:0] mux_1653_nl;
  wire[0:0] mux_1652_nl;
  wire[0:0] mux_1651_nl;
  wire[0:0] nand_154_nl;
  wire[0:0] or_1871_nl;
  wire[0:0] mux_1650_nl;
  wire[0:0] mux_1649_nl;
  wire[0:0] mux_1648_nl;
  wire[0:0] mux_1647_nl;
  wire[0:0] mux_1646_nl;
  wire[0:0] mux_1645_nl;
  wire[0:0] mux_1644_nl;
  wire[0:0] mux_1643_nl;
  wire[0:0] mux_1642_nl;
  wire[0:0] mux_1641_nl;
  wire[0:0] mux_1640_nl;
  wire[0:0] mux_1639_nl;
  wire[0:0] mux_1638_nl;
  wire[0:0] mux_1637_nl;
  wire[0:0] mux_1636_nl;
  wire[0:0] mux_1635_nl;
  wire[0:0] mux_1634_nl;
  wire[0:0] mux_1633_nl;
  wire[0:0] mux_1632_nl;
  wire[0:0] mux_1631_nl;
  wire[0:0] or_1866_nl;
  wire[0:0] mux_1629_nl;
  wire[0:0] mux_1628_nl;
  wire[0:0] mux_1627_nl;
  wire[0:0] or_1862_nl;
  wire[0:0] or_1861_nl;
  wire[0:0] mux_1626_nl;
  wire[0:0] mux_1625_nl;
  wire[0:0] mux_1623_nl;
  wire[0:0] mux_1622_nl;
  wire[0:0] mux_1621_nl;
  wire[0:0] or_1857_nl;
  wire[0:0] mux_1620_nl;
  wire[0:0] mux_1619_nl;
  wire[0:0] mux_1618_nl;
  wire[0:0] or_1855_nl;
  wire[0:0] mux_1616_nl;
  wire[0:0] mux_1615_nl;
  wire[0:0] or_1851_nl;
  wire [0:0] nl_modulo_dev_cmp_ccs_ccore_start_rsc_dat;
  assign or_1873_nl = (~ (fsm_output[1])) | (~ (fsm_output[6])) | (fsm_output[5])
      | (fsm_output[9]) | (fsm_output[8]);
  assign mux_1655_nl = MUX_s_1_2_2(mux_tmp_1563, or_1873_nl, fsm_output[7]);
  assign mux_1653_nl = MUX_s_1_2_2(or_tmp_1835, or_tmp_1825, fsm_output[1]);
  assign mux_1654_nl = MUX_s_1_2_2(mux_tmp_1562, mux_1653_nl, fsm_output[7]);
  assign mux_1656_nl = MUX_s_1_2_2(mux_1655_nl, mux_1654_nl, fsm_output[4]);
  assign nand_154_nl = ~((fsm_output[1]) & (fsm_output[5]) & (fsm_output[9]) & (~
      (fsm_output[8])));
  assign or_1871_nl = (fsm_output[1]) | (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[8]);
  assign mux_1651_nl = MUX_s_1_2_2(nand_154_nl, or_1871_nl, fsm_output[7]);
  assign mux_1652_nl = MUX_s_1_2_2(mux_tmp_1566, mux_1651_nl, fsm_output[4]);
  assign mux_1657_nl = MUX_s_1_2_2(mux_1656_nl, mux_1652_nl, fsm_output[3]);
  assign mux_1647_nl = MUX_s_1_2_2(or_tmp_1841, or_tmp_1827, fsm_output[1]);
  assign mux_1648_nl = MUX_s_1_2_2(mux_tmp_1579, mux_1647_nl, fsm_output[7]);
  assign mux_1645_nl = MUX_s_1_2_2(or_tmp_1841, or_tmp_1838, fsm_output[1]);
  assign mux_1644_nl = MUX_s_1_2_2(or_tmp_1841, or_tmp_1824, fsm_output[1]);
  assign mux_1646_nl = MUX_s_1_2_2(mux_1645_nl, mux_1644_nl, fsm_output[7]);
  assign mux_1649_nl = MUX_s_1_2_2(mux_1648_nl, mux_1646_nl, fsm_output[4]);
  assign mux_1641_nl = MUX_s_1_2_2(or_tmp_1840, or_tmp_1830, fsm_output[1]);
  assign mux_1642_nl = MUX_s_1_2_2(mux_tmp_1573, mux_1641_nl, fsm_output[7]);
  assign mux_1639_nl = MUX_s_1_2_2(or_tmp_1823, or_tmp_1818, fsm_output[1]);
  assign mux_1638_nl = MUX_s_1_2_2(or_tmp_1830, or_tmp_1840, fsm_output[1]);
  assign mux_1640_nl = MUX_s_1_2_2(mux_1639_nl, mux_1638_nl, fsm_output[7]);
  assign mux_1643_nl = MUX_s_1_2_2(mux_1642_nl, mux_1640_nl, fsm_output[4]);
  assign mux_1650_nl = MUX_s_1_2_2(mux_1649_nl, mux_1643_nl, fsm_output[3]);
  assign mux_1658_nl = MUX_s_1_2_2(mux_1657_nl, mux_1650_nl, fsm_output[2]);
  assign mux_1633_nl = MUX_s_1_2_2(or_tmp_1830, or_tmp_1835, fsm_output[1]);
  assign mux_1632_nl = MUX_s_1_2_2(or_tmp_1838, or_tmp_1835, fsm_output[1]);
  assign mux_1634_nl = MUX_s_1_2_2(mux_1633_nl, mux_1632_nl, fsm_output[7]);
  assign or_1866_nl = (fsm_output[1]) | (fsm_output[6]) | (~ (fsm_output[5])) | (fsm_output[9])
      | (~ (fsm_output[8]));
  assign mux_1631_nl = MUX_s_1_2_2(or_1866_nl, mux_tmp_1579, fsm_output[7]);
  assign mux_1635_nl = MUX_s_1_2_2(mux_1634_nl, mux_1631_nl, fsm_output[4]);
  assign or_1862_nl = (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[8]);
  assign mux_1627_nl = MUX_s_1_2_2(or_tmp_1824, or_1862_nl, fsm_output[1]);
  assign or_1861_nl = (fsm_output[1]) | (fsm_output[6]) | (~ (fsm_output[5])) | (~
      (fsm_output[9])) | (fsm_output[8]);
  assign mux_1628_nl = MUX_s_1_2_2(mux_1627_nl, or_1861_nl, fsm_output[7]);
  assign mux_1625_nl = MUX_s_1_2_2(or_tmp_1831, or_tmp_1827, fsm_output[1]);
  assign mux_1626_nl = MUX_s_1_2_2(mux_1625_nl, mux_tmp_1573, fsm_output[7]);
  assign mux_1629_nl = MUX_s_1_2_2(mux_1628_nl, mux_1626_nl, fsm_output[4]);
  assign mux_1636_nl = MUX_s_1_2_2(mux_1635_nl, mux_1629_nl, fsm_output[3]);
  assign or_1857_nl = (~ (fsm_output[1])) | (fsm_output[6]) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (fsm_output[8]);
  assign mux_1620_nl = MUX_s_1_2_2(or_tmp_1825, or_tmp_1827, fsm_output[1]);
  assign mux_1621_nl = MUX_s_1_2_2(or_1857_nl, mux_1620_nl, fsm_output[7]);
  assign or_1855_nl = (~ (fsm_output[5])) | (fsm_output[9]) | (fsm_output[8]);
  assign mux_1618_nl = MUX_s_1_2_2(or_1855_nl, or_tmp_1825, fsm_output[1]);
  assign mux_1619_nl = MUX_s_1_2_2(mux_1618_nl, mux_tmp_1566, fsm_output[7]);
  assign mux_1622_nl = MUX_s_1_2_2(mux_1621_nl, mux_1619_nl, fsm_output[4]);
  assign or_1851_nl = (~ (fsm_output[1])) | (~ (fsm_output[6])) | (fsm_output[5])
      | (fsm_output[9]) | (~ (fsm_output[8]));
  assign mux_1615_nl = MUX_s_1_2_2(or_1851_nl, mux_tmp_1563, fsm_output[7]);
  assign mux_1616_nl = MUX_s_1_2_2(mux_1615_nl, mux_tmp_1562, fsm_output[4]);
  assign mux_1623_nl = MUX_s_1_2_2(mux_1622_nl, mux_1616_nl, fsm_output[3]);
  assign mux_1637_nl = MUX_s_1_2_2(mux_1636_nl, mux_1623_nl, fsm_output[2]);
  assign mux_1659_nl = MUX_s_1_2_2(mux_1658_nl, mux_1637_nl, fsm_output[0]);
  assign nl_modulo_dev_cmp_ccs_ccore_start_rsc_dat = ~ mux_1659_nl;
  wire [10:0] nl_operator_66_true_div_cmp_b;
  assign nl_operator_66_true_div_cmp_b = {1'b0, operator_66_true_div_cmp_b_9_0};
  wire [0:0] nl_inPlaceNTT_DIT_core_wait_dp_inst_ensig_cgo_iro;
  assign nl_inPlaceNTT_DIT_core_wait_dp_inst_ensig_cgo_iro = ~ mux_1581_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_3_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_3_tr0 = ~ (z_out_8_64_2[62]);
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0 = ~ COMP_LOOP_nor_11_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_32_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_32_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_64_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_64_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_96_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_96_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_128_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_128_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_160_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_160_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_192_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_192_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_224_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_224_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_256_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_256_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_288_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_288_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_320_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_320_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_352_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_352_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_384_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_384_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_416_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_416_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_448_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_448_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_480_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_480_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 = VEC_LOOP_acc_1_psp_1[10];
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_4_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_4_tr0 = ~ (z_out_8_64_2[0]);
  ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd64)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd64)) r_rsci (
      .dat(r_rsc_dat),
      .idat(r_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_15_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_14_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_13_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_12_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_11_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_10_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_9_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_8_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_7_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_6_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_5_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_4_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_3_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_2_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_1_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  modulo_dev  modulo_dev_cmp (
      .base_rsc_dat(nl_modulo_dev_cmp_base_rsc_dat[63:0]),
      .m_rsc_dat(nl_modulo_dev_cmp_m_rsc_dat[63:0]),
      .return_rsc_z(modulo_dev_cmp_return_rsc_z),
      .ccs_ccore_start_rsc_dat(nl_modulo_dev_cmp_ccs_ccore_start_rsc_dat[0:0]),
      .ccs_ccore_clk(clk),
      .ccs_ccore_srst(rst),
      .ccs_ccore_en(modulo_dev_cmp_ccs_ccore_en)
    );
  mgc_div #(.width_a(32'sd65),
  .width_b(32'sd11),
  .signd(32'sd1)) operator_66_true_div_cmp (
      .a(operator_66_true_div_cmp_a),
      .b(nl_operator_66_true_div_cmp_b[10:0]),
      .z(operator_66_true_div_cmp_z)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd10)) STAGE_LOOP_lshift_rg (
      .a(1'b1),
      .s(STAGE_LOOP_i_3_0_sva),
      .z(STAGE_LOOP_lshift_psp_sva_mx0w0)
    );
  inPlaceNTT_DIT_core_wait_dp inPlaceNTT_DIT_core_wait_dp_inst (
      .ensig_cgo_iro(nl_inPlaceNTT_DIT_core_wait_dp_inst_ensig_cgo_iro[0:0]),
      .ensig_cgo(reg_ensig_cgo_cse),
      .modulo_dev_cmp_ccs_ccore_en(modulo_dev_cmp_ccs_ccore_en)
    );
  inPlaceNTT_DIT_core_core_fsm inPlaceNTT_DIT_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .STAGE_LOOP_C_3_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_3_tr0[0:0]),
      .modExp_dev_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_1_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0[0:0]),
      .COMP_LOOP_1_modExp_dev_1_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_32_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_32_tr0[0:0]),
      .COMP_LOOP_2_modExp_dev_1_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_64_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_64_tr0[0:0]),
      .COMP_LOOP_3_modExp_dev_1_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_96_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_96_tr0[0:0]),
      .COMP_LOOP_4_modExp_dev_1_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_128_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_128_tr0[0:0]),
      .COMP_LOOP_5_modExp_dev_1_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_160_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_160_tr0[0:0]),
      .COMP_LOOP_6_modExp_dev_1_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_192_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_192_tr0[0:0]),
      .COMP_LOOP_7_modExp_dev_1_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_224_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_224_tr0[0:0]),
      .COMP_LOOP_8_modExp_dev_1_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_256_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_256_tr0[0:0]),
      .COMP_LOOP_9_modExp_dev_1_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_288_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_288_tr0[0:0]),
      .COMP_LOOP_10_modExp_dev_1_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_320_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_320_tr0[0:0]),
      .COMP_LOOP_11_modExp_dev_1_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_352_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_352_tr0[0:0]),
      .COMP_LOOP_12_modExp_dev_1_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_384_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_384_tr0[0:0]),
      .COMP_LOOP_13_modExp_dev_1_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_416_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_416_tr0[0:0]),
      .COMP_LOOP_14_modExp_dev_1_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_448_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_448_tr0[0:0]),
      .COMP_LOOP_15_modExp_dev_1_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_480_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_480_tr0[0:0]),
      .COMP_LOOP_16_modExp_dev_1_while_C_14_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_512_tr0(COMP_LOOP_COMP_LOOP_and_10_itm),
      .VEC_LOOP_C_0_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0[0:0]),
      .STAGE_LOOP_C_4_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_4_tr0[0:0])
    );
  assign nand_308_cse = ~((z_out_6_10_1[0]) & (fsm_output[5]) & (fsm_output[7]) &
      (fsm_output[4]));
  assign nand_270_cse_1 = ~((z_out_6_10_1[3]) & (fsm_output[5]) & (fsm_output[7])
      & (fsm_output[4]));
  assign nand_264_cse = ~((z_out_6_10_1[3]) & (z_out_6_10_1[0]) & (fsm_output[5])
      & (fsm_output[7]) & (fsm_output[4]));
  assign nand_260_cse_1 = ~((z_out_6_10_1[1]) & (z_out_6_10_1[3]) & (fsm_output[5])
      & (fsm_output[7]) & (fsm_output[4]));
  assign or_2146_cse = (fsm_output[3:2]!=2'b00);
  assign and_357_cse = (fsm_output[0]) & (fsm_output[2]) & (fsm_output[3]);
  assign mux_1575_nl = MUX_s_1_2_2((~ (fsm_output[9])), nor_tmp_14, fsm_output[3]);
  assign mux_1576_nl = MUX_s_1_2_2(mux_1575_nl, mux_461_cse, fsm_output[2]);
  assign mux_1574_nl = MUX_s_1_2_2(mux_tmp_1514, mux_tmp_1488, fsm_output[0]);
  assign mux_1577_nl = MUX_s_1_2_2(mux_1576_nl, mux_1574_nl, fsm_output[6]);
  assign mux_1578_nl = MUX_s_1_2_2(mux_1577_nl, mux_tmp_1498, fsm_output[7]);
  assign mux_1570_nl = MUX_s_1_2_2(mux_424_cse, nor_tmp_14, or_214_cse);
  assign mux_1571_nl = MUX_s_1_2_2(mux_1570_nl, mux_tmp_1496, fsm_output[0]);
  assign and_278_nl = (and_357_cse | (fsm_output[9])) & (fsm_output[8]);
  assign mux_1572_nl = MUX_s_1_2_2(mux_1571_nl, and_278_nl, fsm_output[6]);
  assign mux_1569_nl = MUX_s_1_2_2(mux_tmp_1503, mux_tmp_1501, fsm_output[6]);
  assign mux_1573_nl = MUX_s_1_2_2(mux_1572_nl, mux_1569_nl, fsm_output[7]);
  assign mux_1579_nl = MUX_s_1_2_2(mux_1578_nl, mux_1573_nl, fsm_output[5]);
  assign mux_1566_nl = MUX_s_1_2_2(mux_tmp_1514, mux_tmp_1496, fsm_output[6]);
  assign mux_1567_nl = MUX_s_1_2_2(mux_1566_nl, mux_tmp_1477, fsm_output[7]);
  assign and_280_nl = ((~((fsm_output[0]) | (fsm_output[2]) | (fsm_output[3]))) |
      (fsm_output[9])) & (fsm_output[8]);
  assign mux_1562_nl = MUX_s_1_2_2(and_280_nl, mux_tmp_1489, fsm_output[6]);
  assign mux_1561_nl = MUX_s_1_2_2(mux_tmp_1485, nor_tmp_190, fsm_output[6]);
  assign mux_1563_nl = MUX_s_1_2_2(mux_1562_nl, mux_1561_nl, fsm_output[7]);
  assign mux_1568_nl = MUX_s_1_2_2(mux_1567_nl, mux_1563_nl, fsm_output[5]);
  assign mux_1580_nl = MUX_s_1_2_2(mux_1579_nl, mux_1568_nl, fsm_output[4]);
  assign mux_1555_nl = MUX_s_1_2_2(nor_697_cse, nor_tmp_14, or_2146_cse);
  assign mux_1556_nl = MUX_s_1_2_2(mux_1555_nl, mux_tmp_1482, fsm_output[0]);
  assign mux_1557_nl = MUX_s_1_2_2(mux_1556_nl, mux_tmp_1503, fsm_output[6]);
  assign mux_1551_nl = MUX_s_1_2_2(nor_tmp_14, mux_tmp_1470, fsm_output[0]);
  assign mux_1553_nl = MUX_s_1_2_2(mux_tmp_1501, mux_1551_nl, fsm_output[6]);
  assign mux_1558_nl = MUX_s_1_2_2(mux_1557_nl, mux_1553_nl, fsm_output[7]);
  assign mux_1544_nl = MUX_s_1_2_2(nor_tmp_186, mux_tmp_1471, fsm_output[2]);
  assign mux_1545_nl = MUX_s_1_2_2(mux_tmp_1473, mux_1544_nl, fsm_output[0]);
  assign mux_1546_nl = MUX_s_1_2_2(mux_tmp_1476, mux_1545_nl, fsm_output[6]);
  assign mux_1550_nl = MUX_s_1_2_2(mux_tmp_1498, mux_1546_nl, fsm_output[7]);
  assign mux_1559_nl = MUX_s_1_2_2(mux_1558_nl, mux_1550_nl, fsm_output[5]);
  assign mux_1541_nl = MUX_s_1_2_2(mux_tmp_1489, mux_tmp_1485, fsm_output[6]);
  assign mux_1530_nl = MUX_s_1_2_2((fsm_output[9]), nor_tmp_14, or_214_cse);
  assign mux_1531_nl = MUX_s_1_2_2(mux_tmp_1476, mux_1530_nl, fsm_output[0]);
  assign mux_1532_nl = MUX_s_1_2_2(nor_tmp_190, mux_1531_nl, fsm_output[6]);
  assign mux_1542_nl = MUX_s_1_2_2(mux_1541_nl, mux_1532_nl, fsm_output[7]);
  assign mux_1525_nl = MUX_s_1_2_2(mux_tmp_1473, mux_tmp_1470, fsm_output[6]);
  assign mux_1529_nl = MUX_s_1_2_2(mux_tmp_1477, mux_1525_nl, fsm_output[7]);
  assign mux_1543_nl = MUX_s_1_2_2(mux_1542_nl, mux_1529_nl, fsm_output[5]);
  assign mux_1560_nl = MUX_s_1_2_2(mux_1559_nl, mux_1543_nl, fsm_output[4]);
  assign mux_1581_itm = MUX_s_1_2_2(mux_1580_nl, mux_1560_nl, fsm_output[1]);
  assign or_1973_cse = (fsm_output[6]) | (fsm_output[2]) | (~ (fsm_output[7])) |
      (fsm_output[9]) | (fsm_output[3]) | (fsm_output[8]);
  assign nor_256_cse = ~((fsm_output[4]) | (fsm_output[6]) | (fsm_output[2]) | (~
      (fsm_output[7])) | (fsm_output[9]) | (fsm_output[3]) | (fsm_output[8]));
  assign or_1916_cse = (~ (fsm_output[8])) | (fsm_output[9]) | (fsm_output[3]);
  assign or_1982_cse = (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[8]));
  assign or_1967_cse = (~ (fsm_output[6])) | (fsm_output[2]) | (fsm_output[7]) |
      (fsm_output[9]) | (fsm_output[3]) | (fsm_output[8]);
  assign or_1977_cse = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) |
      (fsm_output[3]) | (fsm_output[8]);
  assign or_1976_cse = (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9]) |
      (fsm_output[3]) | (fsm_output[8]);
  assign mux_1788_cse = MUX_s_1_2_2(or_1977_cse, or_1976_cse, fsm_output[6]);
  assign or_1995_cse = (fsm_output[2]) | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9])
      | (~ (fsm_output[8]));
  assign mux_1802_cse = MUX_s_1_2_2(or_1995_cse, or_1977_cse, fsm_output[6]);
  assign mux_1797_cse = MUX_s_1_2_2(nand_357_cse, or_279_cse, fsm_output[6]);
  assign or_1980_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[9])
      | nand_321_cse;
  assign mux_1789_cse = MUX_s_1_2_2(or_1980_nl, or_279_cse, fsm_output[6]);
  assign mux_1784_cse = MUX_s_1_2_2(or_279_cse, nand_tmp_106, fsm_output[6]);
  assign mux_1785_cse = MUX_s_1_2_2(mux_1784_cse, or_1973_cse, fsm_output[4]);
  assign and_259_cse = (fsm_output[4]) & (~ mux_1602_cse);
  assign mux_1725_nl = MUX_s_1_2_2(or_2306_cse, mux_tmp_1610, fsm_output[2]);
  assign mux_1726_cse = MUX_s_1_2_2(mux_1725_nl, mux_tmp_1623, fsm_output[1]);
  assign modExp_dev_while_mux_2_nl = MUX_v_64_2_2(operator_64_false_acc_mut_63_0,
      modExp_dev_result_sva, mux_2066_cse);
  assign modExp_dev_while_mux_3_nl = MUX_v_64_2_2(modExp_dev_result_sva, r_sva, mux_2066_cse);
  assign nl_mul_nl = modExp_dev_while_mux_2_nl * modExp_dev_while_mux_3_nl;
  assign mul_nl = nl_mul_nl[63:0];
  assign nl_COMP_LOOP_1_acc_8_nl = tmp_10_lpi_4_dfm - modulo_dev_cmp_return_rsc_z;
  assign COMP_LOOP_1_acc_8_nl = nl_COMP_LOOP_1_acc_8_nl[63:0];
  assign modExp_dev_while_or_1_nl = and_dcpl_183 | not_tmp_402;
  assign and_258_nl = (fsm_output[4]) & (~ mux_1789_cse);
  assign nor_255_nl = ~((fsm_output[4]) | mux_1788_cse);
  assign mux_1790_nl = MUX_s_1_2_2(and_258_nl, nor_255_nl, fsm_output[5]);
  assign mux_1787_nl = MUX_s_1_2_2(nor_256_cse, and_259_cse, fsm_output[5]);
  assign mux_1791_nl = MUX_s_1_2_2(mux_1790_nl, mux_1787_nl, fsm_output[1]);
  assign and_260_nl = (fsm_output[5]) & (~ mux_1785_cse);
  assign mux_1783_nl = MUX_s_1_2_2(mux_1602_cse, or_1967_cse, fsm_output[4]);
  assign nor_257_nl = ~((fsm_output[5]) | mux_1783_nl);
  assign mux_1786_nl = MUX_s_1_2_2(and_260_nl, nor_257_nl, fsm_output[1]);
  assign mux_1792_nl = MUX_s_1_2_2(mux_1791_nl, mux_1786_nl, fsm_output[0]);
  assign modExp_dev_while_mux1h_nl = MUX1HOT_v_64_4_2(mul_nl, 64'b0000000000000000000000000000000000000000000000000000000000000001,
      modulo_dev_cmp_return_rsc_z, COMP_LOOP_1_acc_8_nl, {modExp_dev_while_or_1_nl
      , mux_1911_cse , mux_1792_nl , not_tmp_370});
  assign mux_1693_nl = MUX_s_1_2_2(or_1916_cse, or_tmp_1854, fsm_output[7]);
  assign or_1896_nl = (fsm_output[2]) | mux_1693_nl;
  assign mux_1694_nl = MUX_s_1_2_2(or_1896_nl, mux_tmp_1618, fsm_output[1]);
  assign mux_1691_nl = MUX_s_1_2_2(or_tmp_1799, mux_tmp_1610, fsm_output[2]);
  assign mux_1692_nl = MUX_s_1_2_2(mux_1691_nl, or_tmp_1855, fsm_output[1]);
  assign mux_1695_nl = MUX_s_1_2_2(mux_1694_nl, mux_1692_nl, fsm_output[5]);
  assign mux_1696_nl = MUX_s_1_2_2(mux_1695_nl, mux_tmp_1621, fsm_output[6]);
  assign mux_1727_nl = MUX_s_1_2_2(or_2306_cse, or_tmp_1793, fsm_output[2]);
  assign mux_1688_nl = MUX_s_1_2_2(mux_1727_nl, mux_tmp_1625, fsm_output[1]);
  assign mux_1689_nl = MUX_s_1_2_2(mux_1688_nl, mux_1726_cse, fsm_output[5]);
  assign mux_1686_nl = MUX_s_1_2_2(mux_tmp_1629, mux_tmp_1626, fsm_output[5]);
  assign mux_1690_nl = MUX_s_1_2_2(mux_1689_nl, mux_1686_nl, fsm_output[6]);
  assign mux_1697_nl = MUX_s_1_2_2(mux_1696_nl, mux_1690_nl, fsm_output[4]);
  assign mux_1683_nl = MUX_s_1_2_2(mux_1726_cse, mux_tmp_1629, fsm_output[5]);
  assign mux_1713_nl = MUX_s_1_2_2(mux_tmp_1623, or_1880_cse, fsm_output[1]);
  assign mux_1678_nl = MUX_s_1_2_2(mux_tmp_1626, mux_1713_nl, fsm_output[5]);
  assign mux_1684_nl = MUX_s_1_2_2(mux_1683_nl, mux_1678_nl, fsm_output[6]);
  assign mux_1703_nl = MUX_s_1_2_2(mux_tmp_1610, mux_1583_cse, fsm_output[2]);
  assign mux_1667_nl = MUX_s_1_2_2(or_tmp_1855, mux_1703_nl, fsm_output[1]);
  assign mux_1664_nl = MUX_s_1_2_2(mux_tmp_1612, or_1880_cse, fsm_output[1]);
  assign mux_1668_nl = MUX_s_1_2_2(mux_1667_nl, mux_1664_nl, fsm_output[5]);
  assign mux_1673_nl = MUX_s_1_2_2(mux_tmp_1621, mux_1668_nl, fsm_output[6]);
  assign mux_1685_nl = MUX_s_1_2_2(mux_1684_nl, mux_1673_nl, fsm_output[4]);
  assign mux_1698_nl = MUX_s_1_2_2(mux_1697_nl, mux_1685_nl, fsm_output[0]);
  assign operator_64_false_operator_64_false_mux_rgt = MUX_v_65_2_2(({1'b0 , modExp_dev_while_mux1h_nl}),
      z_out_9, mux_1698_nl);
  assign or_2306_cse = (fsm_output[7]) | (~ (fsm_output[8])) | (fsm_output[3]) |
      (fsm_output[9]);
  assign nor_810_cse = ~((~ (fsm_output[0])) | (fsm_output[4]));
  assign and_418_cse = (fsm_output[2:1]==2'b11);
  assign and_267_cse = (fsm_output[1:0]==2'b11);
  assign and_195_rgt = and_dcpl_132 & and_dcpl_48;
  assign or_2012_cse = (fsm_output[3]) | (fsm_output[9]) | (fsm_output[8]);
  assign modExp_dev_while_or_2_cse = and_dcpl_36 | and_dcpl_44 | and_dcpl_52 | and_dcpl_58
      | and_dcpl_63 | and_dcpl_72 | and_dcpl_78 | and_dcpl_84 | and_dcpl_90 | and_dcpl_93
      | and_dcpl_97 | and_dcpl_102 | and_dcpl_106 | and_dcpl_110 | and_dcpl_115 |
      and_dcpl_119;
  assign or_2186_cse = (fsm_output[1:0]!=2'b00);
  assign or_2040_cse = (fsm_output[4:3]!=2'b00);
  assign or_103_cse = (fsm_output[5]) | (fsm_output[4]) | (fsm_output[7]);
  assign and_375_cse = (fsm_output[4:3]==2'b11);
  assign and_376_cse = (fsm_output[3:2]==2'b11);
  assign and_247_cse = (fsm_output[2:0]==3'b111);
  assign mux_424_cse = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), fsm_output[9]);
  assign or_214_cse = (fsm_output[3:2]!=2'b01);
  assign or_212_cse = (fsm_output[9:8]!=2'b01);
  assign mux_461_cse = MUX_s_1_2_2(mux_424_cse, nor_tmp_14, fsm_output[3]);
  assign mux_459_nl = MUX_s_1_2_2(mux_424_cse, (fsm_output[9]), fsm_output[3]);
  assign mux_460_cse = MUX_s_1_2_2(mux_459_nl, nor_tmp_14, fsm_output[2]);
  assign nor_697_cse = ~((fsm_output[9:8]!=2'b00));
  assign mux_1904_nl = MUX_s_1_2_2(mux_1797_cse, mux_1788_cse, fsm_output[4]);
  assign nor_760_cse = ~((fsm_output[5]) | mux_1904_nl);
  assign nor_758_nl = ~((fsm_output[4]) | mux_1802_cse);
  assign and_256_nl = (fsm_output[4]) & (~ mux_1797_cse);
  assign mux_1909_cse = MUX_s_1_2_2(nor_758_nl, and_256_nl, fsm_output[5]);
  assign mux_1800_nl = MUX_s_1_2_2(or_279_cse, nand_tmp, fsm_output[6]);
  assign and_445_nl = (fsm_output[4]) & (~ mux_1800_nl);
  assign mux_1907_nl = MUX_s_1_2_2(and_445_nl, nor_256_cse, fsm_output[5]);
  assign mux_1910_nl = MUX_s_1_2_2(mux_1909_cse, mux_1907_nl, fsm_output[1]);
  assign mux_1794_nl = MUX_s_1_2_2(nand_tmp, or_1982_cse, fsm_output[6]);
  assign mux_1901_nl = MUX_s_1_2_2(mux_1794_nl, or_1967_cse, fsm_output[4]);
  assign and_446_nl = (fsm_output[5]) & (~ mux_1901_nl);
  assign mux_1905_nl = MUX_s_1_2_2(nor_760_cse, and_446_nl, fsm_output[1]);
  assign mux_1911_cse = MUX_s_1_2_2(mux_1910_nl, mux_1905_nl, fsm_output[0]);
  assign mux_1949_cse = MUX_s_1_2_2((fsm_output[8]), or_tmp_2044, fsm_output[3]);
  assign or_2336_cse = (~((fsm_output[3]) | (~ (fsm_output[9])))) | (fsm_output[8]);
  assign COMP_LOOP_k_COMP_LOOP_k_mux_nl = MUX_v_5_2_2(COMP_LOOP_k_9_4_sva_4_0, (z_out_9[8:4]),
      not_tmp_402);
  assign COMP_LOOP_mux1h_192_rgt = MUX_v_10_2_2(({5'b00000 , COMP_LOOP_k_COMP_LOOP_k_mux_nl}),
      z_out_6_10_1, modExp_dev_while_or_2_cse);
  assign or_2348_cse = (fsm_output[4]) | (fsm_output[0]) | (fsm_output[1]);
  assign or_279_cse = (fsm_output[2]) | (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (~ (fsm_output[3]));
  assign nl_COMP_LOOP_acc_13_psp_sva_1 = (VEC_LOOP_j_sva_9_0[9:2]) + conv_u2u_7_8({COMP_LOOP_k_9_4_sva_4_0
      , 2'b01});
  assign COMP_LOOP_acc_13_psp_sva_1 = nl_COMP_LOOP_acc_13_psp_sva_1[7:0];
  assign nl_COMP_LOOP_acc_1_cse_2_sva_1 = VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0001});
  assign COMP_LOOP_acc_1_cse_2_sva_1 = nl_COMP_LOOP_acc_1_cse_2_sva_1[9:0];
  assign nl_VEC_LOOP_acc_1_psp_1 = conv_u2u_10_11(VEC_LOOP_j_sva_9_0) + conv_u2u_10_11(STAGE_LOOP_lshift_psp_sva);
  assign VEC_LOOP_acc_1_psp_1 = nl_VEC_LOOP_acc_1_psp_1[10:0];
  assign nor_728_cse = ~((fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[8]));
  assign nor_727_nl = ~((~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[8])));
  assign mux_51_nl = MUX_s_1_2_2(nor_727_nl, nor_728_cse, fsm_output[7]);
  assign nand_tmp = ~((fsm_output[2]) & mux_51_nl);
  assign nand_357_cse = ~((fsm_output[2]) & (fsm_output[7]) & (fsm_output[3]) & (~
      (fsm_output[9])) & (fsm_output[8]));
  assign or_tmp_20 = (fsm_output[5]) | and_375_cse;
  assign nor_tmp_14 = (fsm_output[9:8]==2'b11);
  assign or_tmp_74 = (fsm_output[5]) | (fsm_output[7]);
  assign nor_tmp_40 = (fsm_output[5]) & (fsm_output[7]);
  assign nand_321_cse = ~((fsm_output[3]) & (fsm_output[8]));
  assign and_dcpl_13 = ~((fsm_output[2:1]!=2'b00));
  assign and_dcpl_14 = and_dcpl_13 & (~ (fsm_output[6]));
  assign and_dcpl_15 = and_dcpl_14 & nor_697_cse;
  assign and_dcpl_16 = ~((fsm_output[4]) | (fsm_output[0]));
  assign and_dcpl_17 = ~((fsm_output[5]) | (fsm_output[7]));
  assign and_dcpl_18 = and_dcpl_17 & (~ (fsm_output[3]));
  assign and_dcpl_19 = and_dcpl_18 & and_dcpl_16;
  assign and_dcpl_23 = and_418_cse & (~ (fsm_output[6]));
  assign or_2152_nl = (fsm_output[9]) | (fsm_output[6]) | (fsm_output[2]) | (fsm_output[1])
      | (fsm_output[0]) | (fsm_output[4]) | (fsm_output[3]) | (fsm_output[7]) | (fsm_output[5]);
  assign nand_314_nl = ~((fsm_output[9]) & ((fsm_output[6]) | and_247_cse | (fsm_output[5])
      | (fsm_output[4]) | (fsm_output[3]) | (fsm_output[7])));
  assign not_tmp_121 = MUX_s_1_2_2(or_2152_nl, nand_314_nl, fsm_output[8]);
  assign and_dcpl_26 = (fsm_output[2:1]==2'b10);
  assign and_dcpl_27 = and_dcpl_26 & (~ (fsm_output[6]));
  assign and_dcpl_28 = and_dcpl_27 & nor_697_cse;
  assign and_dcpl_29 = (fsm_output[4]) & (~ (fsm_output[0]));
  assign and_dcpl_30 = and_dcpl_18 & and_dcpl_29;
  assign and_dcpl_32 = (~ (fsm_output[4])) & (fsm_output[0]);
  assign and_dcpl_33 = (fsm_output[5]) & (~ (fsm_output[7]));
  assign and_dcpl_34 = and_dcpl_33 & (~ (fsm_output[3]));
  assign and_dcpl_35 = and_dcpl_34 & and_dcpl_32;
  assign and_dcpl_36 = and_dcpl_35 & and_dcpl_28;
  assign and_dcpl_37 = (fsm_output[2:1]==2'b01);
  assign and_dcpl_38 = and_dcpl_37 & (fsm_output[6]);
  assign and_dcpl_39 = and_dcpl_38 & nor_697_cse;
  assign and_dcpl_40 = and_dcpl_18 & and_dcpl_32;
  assign and_dcpl_42 = and_dcpl_26 & (fsm_output[6]);
  assign and_dcpl_43 = and_dcpl_42 & nor_697_cse;
  assign and_dcpl_44 = and_dcpl_30 & and_dcpl_43;
  assign and_dcpl_45 = and_dcpl_34 & and_dcpl_29;
  assign and_dcpl_47 = and_dcpl_37 & (~ (fsm_output[6]));
  assign and_dcpl_48 = and_dcpl_47 & nor_697_cse;
  assign and_dcpl_49 = (~ (fsm_output[5])) & (fsm_output[7]);
  assign and_dcpl_50 = and_dcpl_49 & (~ (fsm_output[3]));
  assign and_dcpl_51 = and_dcpl_50 & and_dcpl_32;
  assign and_dcpl_52 = and_dcpl_51 & and_dcpl_48;
  assign and_dcpl_54 = nor_tmp_40 & (~ (fsm_output[3]));
  assign and_dcpl_55 = and_dcpl_54 & and_dcpl_32;
  assign and_dcpl_57 = and_dcpl_54 & and_dcpl_29;
  assign and_dcpl_58 = and_dcpl_57 & and_dcpl_48;
  assign and_dcpl_59 = and_dcpl_13 & (fsm_output[6]);
  assign and_dcpl_60 = and_dcpl_59 & nor_697_cse;
  assign and_dcpl_61 = and_dcpl_50 & and_dcpl_29;
  assign and_dcpl_63 = and_dcpl_55 & and_dcpl_60;
  assign and_dcpl_64 = and_418_cse & (fsm_output[6]);
  assign and_dcpl_65 = and_dcpl_64 & nor_697_cse;
  assign and_dcpl_66 = (fsm_output[4]) & (fsm_output[0]);
  assign and_dcpl_67 = nor_tmp_40 & (fsm_output[3]);
  assign and_dcpl_68 = and_dcpl_67 & and_dcpl_66;
  assign and_dcpl_70 = (fsm_output[9:8]==2'b01);
  assign and_dcpl_71 = and_dcpl_14 & and_dcpl_70;
  assign and_dcpl_72 = and_dcpl_30 & and_dcpl_71;
  assign and_dcpl_73 = and_dcpl_23 & and_dcpl_70;
  assign and_dcpl_74 = and_dcpl_33 & (fsm_output[3]);
  assign and_dcpl_75 = and_dcpl_74 & and_dcpl_16;
  assign and_dcpl_78 = and_dcpl_74 & and_dcpl_66 & and_dcpl_73;
  assign and_dcpl_79 = and_dcpl_42 & and_dcpl_70;
  assign and_dcpl_80 = and_dcpl_17 & (fsm_output[3]);
  assign and_dcpl_81 = and_dcpl_80 & and_dcpl_66;
  assign and_dcpl_83 = and_dcpl_64 & and_dcpl_70;
  assign and_dcpl_84 = and_dcpl_75 & and_dcpl_83;
  assign and_dcpl_85 = and_dcpl_27 & and_dcpl_70;
  assign and_dcpl_86 = and_dcpl_49 & (fsm_output[3]);
  assign and_dcpl_87 = and_dcpl_86 & and_dcpl_16;
  assign and_dcpl_89 = and_dcpl_86 & and_dcpl_66;
  assign and_dcpl_90 = and_dcpl_89 & and_dcpl_85;
  assign and_dcpl_91 = and_dcpl_47 & and_dcpl_70;
  assign and_dcpl_93 = and_dcpl_87 & and_dcpl_79;
  assign and_dcpl_94 = and_dcpl_38 & and_dcpl_70;
  assign and_dcpl_95 = and_dcpl_67 & and_dcpl_16;
  assign and_dcpl_97 = and_dcpl_68 & and_dcpl_94;
  assign and_dcpl_98 = (fsm_output[9:8]==2'b10);
  assign and_dcpl_99 = and_dcpl_14 & and_dcpl_98;
  assign and_dcpl_101 = and_dcpl_47 & and_dcpl_98;
  assign and_dcpl_102 = and_dcpl_75 & and_dcpl_101;
  assign and_dcpl_103 = and_dcpl_59 & and_dcpl_98;
  assign and_dcpl_106 = and_dcpl_81 & and_dcpl_103;
  assign and_dcpl_107 = and_dcpl_64 & and_dcpl_98;
  assign and_dcpl_108 = and_dcpl_34 & and_dcpl_66;
  assign and_dcpl_110 = and_dcpl_87 & and_dcpl_99;
  assign and_dcpl_111 = and_dcpl_23 & and_dcpl_98;
  assign and_dcpl_112 = and_dcpl_54 & and_dcpl_16;
  assign and_dcpl_115 = and_dcpl_54 & and_dcpl_66 & and_dcpl_111;
  assign and_dcpl_116 = and_dcpl_42 & and_dcpl_98;
  assign and_dcpl_117 = and_dcpl_50 & and_dcpl_66;
  assign and_dcpl_119 = and_dcpl_112 & and_dcpl_107;
  assign or_tmp_237 = (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[3]);
  assign or_265_nl = (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[3]));
  assign mux_514_nl = MUX_s_1_2_2(or_tmp_237, or_265_nl, fsm_output[7]);
  assign nand_tmp_6 = ~((fsm_output[2]) & (~ mux_514_nl));
  assign or_tmp_239 = (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9]) | nand_321_cse;
  assign or_tmp_241 = (fsm_output[9]) | nand_321_cse;
  assign mux_520_nl = MUX_s_1_2_2(or_tmp_241, or_tmp_237, fsm_output[7]);
  assign nand_tmp_7 = ~((fsm_output[2]) & (~ mux_520_nl));
  assign and_dcpl_122 = and_dcpl_23 & nor_697_cse;
  assign and_dcpl_130 = and_dcpl_59 & and_dcpl_70;
  assign and_dcpl_132 = and_dcpl_18 & and_dcpl_66;
  assign and_dcpl_136 = and_dcpl_27 & and_dcpl_98;
  assign and_dcpl_138 = and_dcpl_38 & and_dcpl_98;
  assign or_tmp_252 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1])
      | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0000);
  assign or_tmp_253 = (~ (fsm_output[5])) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0000);
  assign or_tmp_258 = (~ (fsm_output[5])) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0000);
  assign or_tmp_259 = (fsm_output[5]) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0000);
  assign not_tmp_133 = ~((fsm_output[5]) & (fsm_output[7]) & (fsm_output[4]));
  assign not_tmp_134 = ~((fsm_output[7]) & (fsm_output[4]));
  assign or_tmp_346 = (fsm_output[1]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0001);
  assign or_tmp_352 = (~ (fsm_output[1])) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0001);
  assign or_tmp_353 = (~ (fsm_output[1])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0001);
  assign or_tmp_362 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[5])
      | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0001);
  assign or_tmp_438 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1])
      | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0010);
  assign or_tmp_439 = (~ (fsm_output[5])) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0010);
  assign or_tmp_444 = (~ (fsm_output[5])) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0010);
  assign or_tmp_445 = (fsm_output[5]) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0010);
  assign or_tmp_531 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1])
      | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0011);
  assign or_tmp_532 = (~ (fsm_output[5])) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0011);
  assign or_tmp_537 = (~ (fsm_output[5])) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0011);
  assign or_tmp_538 = (fsm_output[5]) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0011);
  assign or_tmp_624 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1])
      | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0100);
  assign or_tmp_625 = (~ (fsm_output[5])) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0100);
  assign or_tmp_630 = (~ (fsm_output[5])) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0100);
  assign or_tmp_631 = (fsm_output[5]) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0100);
  assign or_tmp_718 = (fsm_output[1]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0101);
  assign or_tmp_724 = (~ (fsm_output[1])) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0101);
  assign or_tmp_725 = (~ (fsm_output[1])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0101);
  assign or_tmp_734 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[5])
      | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0101);
  assign or_tmp_810 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1])
      | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0110);
  assign or_tmp_811 = (~ (fsm_output[5])) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0110);
  assign or_tmp_816 = (~ (fsm_output[5])) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0110);
  assign or_tmp_817 = (fsm_output[5]) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0110);
  assign or_tmp_903 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1])
      | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0111);
  assign or_tmp_904 = (~ (fsm_output[5])) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0111);
  assign or_tmp_909 = ~((fsm_output[5]) & (fsm_output[1]) & (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]==4'b0111));
  assign or_tmp_910 = (fsm_output[5]) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0111);
  assign or_tmp_997 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1])
      | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1000);
  assign or_tmp_999 = (~ (fsm_output[5])) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1000);
  assign or_tmp_1005 = (~ (fsm_output[5])) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1000);
  assign or_tmp_1007 = (fsm_output[5]) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1000);
  assign or_tmp_1097 = (fsm_output[1]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1001);
  assign or_tmp_1104 = (~ (fsm_output[1])) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1001);
  assign or_tmp_1106 = (~ (fsm_output[1])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1001);
  assign or_tmp_1116 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[1]) |
      (fsm_output[5]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1001);
  assign or_tmp_1195 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) |
      (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1010);
  assign or_tmp_1197 = (~ (fsm_output[5])) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1010);
  assign or_tmp_1203 = (~ (fsm_output[5])) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1010);
  assign or_tmp_1205 = (fsm_output[5]) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1010);
  assign or_tmp_1294 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) |
      (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1011);
  assign or_tmp_1296 = (~ (fsm_output[5])) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1011);
  assign or_tmp_1302 = ~((fsm_output[5]) & (fsm_output[1]) & (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]==4'b1011));
  assign or_tmp_1304 = (fsm_output[5]) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1011);
  assign not_tmp_289 = ~((COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:2]==2'b11));
  assign or_tmp_1393 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) |
      (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1:0]!=2'b00) | not_tmp_289;
  assign or_tmp_1395 = (~ (fsm_output[5])) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1:0]!=2'b00)
      | not_tmp_289;
  assign or_tmp_1401 = (~ (fsm_output[5])) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1:0]!=2'b00)
      | not_tmp_289;
  assign or_tmp_1403 = (fsm_output[5]) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1:0]!=2'b00)
      | not_tmp_289;
  assign not_tmp_304 = ~((COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[0]) & (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[2])
      & (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3]));
  assign or_tmp_1493 = (fsm_output[1]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1])
      | not_tmp_304;
  assign or_tmp_1500 = (~ (fsm_output[1])) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1])
      | not_tmp_304;
  assign or_tmp_1502 = (~ (fsm_output[1])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1])
      | not_tmp_304;
  assign or_tmp_1512 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[1]) |
      (fsm_output[5]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1]) | not_tmp_304;
  assign or_tmp_1590 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) |
      (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1:0]!=2'b10) | not_tmp_289;
  assign or_tmp_1592 = (~ (fsm_output[5])) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1:0]!=2'b10)
      | not_tmp_289;
  assign or_tmp_1598 = (~((fsm_output[5]) & (fsm_output[1]) & (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1:0]==2'b10)))
      | not_tmp_289;
  assign or_tmp_1600 = (fsm_output[5]) | (~ (fsm_output[1])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1:0]!=2'b10)
      | not_tmp_289;
  assign not_tmp_335 = ~((COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]==4'b1111));
  assign or_tmp_1687 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) |
      (fsm_output[1]) | not_tmp_335;
  assign or_tmp_1689 = (~ (fsm_output[5])) | (fsm_output[1]) | not_tmp_335;
  assign not_tmp_336 = ~((fsm_output[5]) & (fsm_output[1]) & (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]==4'b1111));
  assign or_tmp_1694 = (fsm_output[5]) | (~((fsm_output[1]) & (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]==4'b1111)));
  assign or_2151_cse = (fsm_output[3]) | (fsm_output[9]);
  assign nor_tmp_186 = or_2151_cse & (fsm_output[8]);
  assign mux_1520_nl = MUX_s_1_2_2(nor_tmp_14, mux_424_cse, fsm_output[3]);
  assign mux_tmp_1470 = MUX_s_1_2_2(nor_tmp_186, mux_1520_nl, fsm_output[2]);
  assign mux_tmp_1471 = MUX_s_1_2_2((fsm_output[9]), nor_tmp_14, fsm_output[3]);
  assign mux_tmp_1472 = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), or_2151_cse);
  assign mux_tmp_1473 = MUX_s_1_2_2(mux_tmp_1472, mux_tmp_1471, fsm_output[2]);
  assign mux_tmp_1476 = MUX_s_1_2_2(mux_461_cse, mux_tmp_1471, fsm_output[2]);
  assign nor_tmp_188 = (and_376_cse | (fsm_output[9])) & (fsm_output[8]);
  assign mux_tmp_1477 = MUX_s_1_2_2(nor_tmp_188, mux_tmp_1476, fsm_output[6]);
  assign nor_tmp_190 = ((~((fsm_output[0]) | (~ (fsm_output[2])) | (~ (fsm_output[3]))))
      | (fsm_output[9])) & (fsm_output[8]);
  assign mux_tmp_1482 = MUX_s_1_2_2(mux_461_cse, nor_tmp_186, fsm_output[2]);
  assign mux_tmp_1483 = MUX_s_1_2_2(nor_tmp_14, (fsm_output[9]), fsm_output[3]);
  assign mux_tmp_1484 = MUX_s_1_2_2(mux_tmp_1483, nor_tmp_186, fsm_output[2]);
  assign mux_tmp_1485 = MUX_s_1_2_2(mux_tmp_1484, mux_tmp_1482, fsm_output[0]);
  assign mux_tmp_1488 = MUX_s_1_2_2(mux_tmp_1483, mux_461_cse, fsm_output[2]);
  assign mux_tmp_1489 = MUX_s_1_2_2(mux_tmp_1488, mux_460_cse, fsm_output[0]);
  assign mux_tmp_1496 = MUX_s_1_2_2(mux_tmp_1483, mux_tmp_1472, fsm_output[2]);
  assign mux_1548_nl = MUX_s_1_2_2(mux_tmp_1496, mux_tmp_1484, fsm_output[0]);
  assign mux_tmp_1498 = MUX_s_1_2_2(mux_1548_nl, nor_tmp_188, fsm_output[6]);
  assign mux_tmp_1501 = MUX_s_1_2_2(mux_tmp_1482, mux_tmp_1473, fsm_output[0]);
  assign mux_tmp_1503 = MUX_s_1_2_2(mux_460_cse, mux_tmp_1476, fsm_output[0]);
  assign mux_1564_nl = MUX_s_1_2_2((fsm_output[8]), (fsm_output[9]), fsm_output[3]);
  assign mux_tmp_1514 = MUX_s_1_2_2(mux_1564_nl, mux_461_cse, fsm_output[2]);
  assign or_tmp_1788 = (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[8]);
  assign or_tmp_1793 = ~((fsm_output[7]) & (fsm_output[3]) & (~ (fsm_output[9]))
      & (fsm_output[8]));
  assign or_tmp_1794 = (fsm_output[7]) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (fsm_output[8]);
  assign or_1820_cse = (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[8]));
  assign mux_1583_cse = MUX_s_1_2_2(or_1820_cse, or_tmp_237, fsm_output[7]);
  assign mux_1584_nl = MUX_s_1_2_2(or_tmp_1793, mux_1583_cse, fsm_output[6]);
  assign mux_tmp_1534 = MUX_s_1_2_2(or_tmp_1794, mux_1584_nl, fsm_output[2]);
  assign or_tmp_1796 = (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[8]);
  assign mux_1587_nl = MUX_s_1_2_2(or_2306_cse, or_tmp_1788, fsm_output[6]);
  assign mux_tmp_1537 = MUX_s_1_2_2(mux_1587_nl, or_tmp_1796, fsm_output[2]);
  assign or_tmp_1799 = ~((fsm_output[7]) & (fsm_output[3]) & (fsm_output[9]) & (~
      (fsm_output[8])));
  assign nor_275_nl = ~((fsm_output[9]) | nand_321_cse);
  assign mux_1601_nl = MUX_s_1_2_2(nor_275_nl, nor_728_cse, fsm_output[7]);
  assign nand_tmp_106 = ~((fsm_output[2]) & mux_1601_nl);
  assign mux_1602_cse = MUX_s_1_2_2(nand_tmp_106, or_tmp_239, fsm_output[6]);
  assign mux_1610_nl = MUX_s_1_2_2(mux_1789_cse, mux_1788_cse, fsm_output[4]);
  assign and_272_nl = (fsm_output[5]) & (~ mux_1610_nl);
  assign nor_272_nl = ~((fsm_output[5]) | mux_1785_cse);
  assign mux_1611_nl = MUX_s_1_2_2(and_272_nl, nor_272_nl, fsm_output[1]);
  assign nor_273_nl = ~((fsm_output[4]) | (~ (fsm_output[6])) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[3]) | (fsm_output[8]));
  assign and_273_nl = (fsm_output[4]) & (~ mux_1784_cse);
  assign mux_1605_nl = MUX_s_1_2_2(nor_273_nl, and_273_nl, fsm_output[5]);
  assign nor_274_nl = ~((fsm_output[4]) | (~ (fsm_output[6])) | (fsm_output[2]) |
      (fsm_output[7]) | (fsm_output[9]) | (fsm_output[3]) | (fsm_output[8]));
  assign mux_1603_nl = MUX_s_1_2_2(and_259_cse, nor_274_nl, fsm_output[5]);
  assign mux_1606_nl = MUX_s_1_2_2(mux_1605_nl, mux_1603_nl, fsm_output[1]);
  assign not_tmp_370 = MUX_s_1_2_2(mux_1611_nl, mux_1606_nl, fsm_output[0]);
  assign or_tmp_1816 = (fsm_output[6]) | (fsm_output[5]) | (fsm_output[9]) | (~ (fsm_output[8]));
  assign or_tmp_1818 = ~((fsm_output[6]) & (fsm_output[5]) & (~ (fsm_output[9]))
      & (fsm_output[8]));
  assign mux_tmp_1562 = MUX_s_1_2_2(or_tmp_1818, or_tmp_1816, fsm_output[1]);
  assign or_1849_nl = (~ (fsm_output[5])) | (fsm_output[9]) | (~ (fsm_output[8]));
  assign mux_tmp_1563 = MUX_s_1_2_2(or_1849_nl, or_tmp_1816, fsm_output[1]);
  assign or_tmp_1823 = (fsm_output[6]) | (fsm_output[5]) | (~ (fsm_output[9])) |
      (fsm_output[8]);
  assign or_tmp_1824 = ~((fsm_output[6]) & (fsm_output[5]) & (fsm_output[9]) & (~
      (fsm_output[8])));
  assign mux_tmp_1566 = MUX_s_1_2_2(or_tmp_1824, or_tmp_1823, fsm_output[1]);
  assign or_tmp_1825 = (fsm_output[6]) | (fsm_output[5]) | (fsm_output[9]) | (fsm_output[8]);
  assign or_tmp_1827 = (~ (fsm_output[6])) | (fsm_output[5]) | (~ (fsm_output[9]))
      | (fsm_output[8]);
  assign or_tmp_1830 = (~ (fsm_output[6])) | (fsm_output[5]) | (fsm_output[9]) |
      (~ (fsm_output[8]));
  assign or_tmp_1831 = (fsm_output[6]) | (~ (fsm_output[5])) | (~ (fsm_output[9]))
      | (fsm_output[8]);
  assign mux_tmp_1573 = MUX_s_1_2_2(or_tmp_1831, or_tmp_1830, fsm_output[1]);
  assign or_tmp_1835 = (~ (fsm_output[6])) | (~ (fsm_output[5])) | (fsm_output[9])
      | (fsm_output[8]);
  assign or_1863_nl = (fsm_output[5]) | (fsm_output[9]) | (fsm_output[8]);
  assign mux_tmp_1579 = MUX_s_1_2_2(or_tmp_1835, or_1863_nl, fsm_output[1]);
  assign or_tmp_1838 = (~ (fsm_output[6])) | (fsm_output[5]) | (fsm_output[9]) |
      (fsm_output[8]);
  assign or_tmp_1840 = (fsm_output[6]) | (~ (fsm_output[5])) | (fsm_output[9]) |
      (~ (fsm_output[8]));
  assign or_tmp_1841 = (fsm_output[6]) | (~ (fsm_output[5])) | (fsm_output[9]) |
      (fsm_output[8]);
  assign and_dcpl_169 = and_dcpl_18 & (~ (fsm_output[4])) & (fsm_output[1]) & (~
      (fsm_output[2])) & (~ (fsm_output[6])) & nor_697_cse;
  assign or_tmp_1845 = and_418_cse | (fsm_output[4]) | (fsm_output[3]) | (fsm_output[7])
      | (fsm_output[5]);
  assign and_tmp_12 = (fsm_output[9]) & ((fsm_output[6]) | or_tmp_1845);
  assign mux_tmp_1610 = MUX_s_1_2_2(or_2012_cse, or_1820_cse, fsm_output[7]);
  assign or_1880_cse = (fsm_output[2]) | mux_tmp_1610;
  assign mux_tmp_1612 = MUX_s_1_2_2(or_tmp_1794, mux_1583_cse, fsm_output[2]);
  assign or_tmp_1854 = (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[8]);
  assign mux_tmp_1615 = MUX_s_1_2_2(or_tmp_1854, or_2012_cse, fsm_output[7]);
  assign or_tmp_1855 = (fsm_output[2]) | mux_tmp_1615;
  assign mux_tmp_1618 = MUX_s_1_2_2(mux_tmp_1615, or_tmp_1793, fsm_output[2]);
  assign nand_111_nl = ~((fsm_output[2]) & (~ mux_tmp_1610));
  assign mux_1671_nl = MUX_s_1_2_2(nand_111_nl, mux_tmp_1612, fsm_output[1]);
  assign nand_110_nl = ~((fsm_output[2]) & (~ mux_1583_cse));
  assign mux_1670_nl = MUX_s_1_2_2(mux_tmp_1618, nand_110_nl, fsm_output[1]);
  assign mux_tmp_1621 = MUX_s_1_2_2(mux_1671_nl, mux_1670_nl, fsm_output[5]);
  assign mux_tmp_1623 = MUX_s_1_2_2(or_tmp_1788, mux_1583_cse, fsm_output[2]);
  assign mux_tmp_1625 = MUX_s_1_2_2(mux_tmp_1615, or_tmp_1796, fsm_output[2]);
  assign mux_tmp_1626 = MUX_s_1_2_2(mux_tmp_1625, or_1982_cse, fsm_output[1]);
  assign mux_1679_nl = MUX_s_1_2_2(or_tmp_1794, or_tmp_1796, fsm_output[2]);
  assign mux_tmp_1629 = MUX_s_1_2_2(mux_1679_nl, mux_tmp_1623, fsm_output[1]);
  assign nand_151_nl = ~((fsm_output[1]) & (fsm_output[0]) & (fsm_output[4]));
  assign mux_tmp_1688 = MUX_s_1_2_2(nand_151_nl, or_2348_cse, fsm_output[2]);
  assign or_tmp_1899 = and_375_cse | (fsm_output[7]) | (fsm_output[5]);
  assign and_dcpl_183 = and_dcpl_40 & and_dcpl_28;
  assign nand_342_nl = ~((fsm_output[2]) & (fsm_output[3]) & (~ (fsm_output[9]))
      & (fsm_output[8]));
  assign or_2000_nl = (~ (fsm_output[2])) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (fsm_output[8]);
  assign mux_1768_cse = MUX_s_1_2_2(nand_342_nl, or_2000_nl, fsm_output[7]);
  assign or_1996_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[8]);
  assign mux_1803_nl = MUX_s_1_2_2(or_1996_nl, nand_357_cse, fsm_output[6]);
  assign mux_1804_nl = MUX_s_1_2_2(mux_1803_nl, mux_1802_cse, fsm_output[4]);
  assign and_261_nl = (fsm_output[5]) & (~ mux_1804_nl);
  assign mux_1779_nl = MUX_s_1_2_2(and_261_nl, nor_760_cse, fsm_output[1]);
  assign mux_1769_nl = MUX_s_1_2_2(or_279_cse, mux_1768_cse, fsm_output[6]);
  assign and_263_nl = (fsm_output[4]) & (~ mux_1769_nl);
  assign mux_1770_nl = MUX_s_1_2_2(and_263_nl, nor_256_cse, fsm_output[5]);
  assign mux_1774_nl = MUX_s_1_2_2(mux_1909_cse, mux_1770_nl, fsm_output[1]);
  assign not_tmp_402 = MUX_s_1_2_2(mux_1779_nl, mux_1774_nl, fsm_output[0]);
  assign nor_tmp_203 = (fsm_output[6]) & (fsm_output[7]) & (fsm_output[9]);
  assign not_tmp_418 = ~((fsm_output[6]) | (fsm_output[7]) | (fsm_output[9]));
  assign nor_248_nl = ~((fsm_output[0]) | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[9]));
  assign mux_1827_nl = MUX_s_1_2_2(nor_248_nl, nor_tmp_203, fsm_output[1]);
  assign mux_1828_nl = MUX_s_1_2_2(not_tmp_418, mux_1827_nl, fsm_output[2]);
  assign mux_1829_nl = MUX_s_1_2_2(mux_1828_nl, nor_tmp_203, fsm_output[3]);
  assign mux_1830_nl = MUX_s_1_2_2(not_tmp_418, mux_1829_nl, fsm_output[4]);
  assign mux_1831_nl = MUX_s_1_2_2(mux_1830_nl, nor_tmp_203, fsm_output[5]);
  assign mux_1832_itm = MUX_s_1_2_2(mux_1831_nl, (fsm_output[9]), fsm_output[8]);
  assign or_tmp_1989 = (fsm_output[5]) | (~ nor_tmp_203);
  assign or_tmp_1990 = (fsm_output[5]) | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[9]);
  assign mux_tmp_1782 = MUX_s_1_2_2(or_tmp_1990, or_tmp_1989, fsm_output[4]);
  assign mux_1834_itm = MUX_s_1_2_2(not_tmp_418, nor_tmp_203, fsm_output[5]);
  assign mux_tmp_1786 = MUX_s_1_2_2((~ mux_1834_itm), or_tmp_1990, fsm_output[4]);
  assign mux_1843_nl = MUX_s_1_2_2(or_tmp_1899, or_103_cse, or_2186_cse);
  assign mux_tmp_1793 = MUX_s_1_2_2(or_tmp_1899, mux_1843_nl, fsm_output[2]);
  assign mux_tmp_1799 = MUX_s_1_2_2((~ (fsm_output[5])), (fsm_output[5]), fsm_output[7]);
  assign mux_tmp_1801 = MUX_s_1_2_2(mux_tmp_1799, nor_tmp_40, fsm_output[4]);
  assign mux_tmp_1803 = MUX_s_1_2_2(mux_tmp_1799, nor_tmp_40, and_375_cse);
  assign mux_tmp_1808 = MUX_s_1_2_2(nor_tmp_40, (fsm_output[7]), or_2040_cse);
  assign mux_tmp_1809 = MUX_s_1_2_2(nor_tmp_40, (fsm_output[7]), fsm_output[4]);
  assign not_tmp_431 = ~((fsm_output[6]) | mux_tmp_1793);
  assign nor_tmp_215 = (fsm_output[5]) & (fsm_output[6]) & (fsm_output[9]);
  assign not_tmp_439 = ~((fsm_output[5]) | (fsm_output[6]) | (fsm_output[9]));
  assign nor_244_nl = ~((fsm_output[7]) | (fsm_output[9]));
  assign and_368_nl = (fsm_output[9]) & (fsm_output[7]);
  assign mux_tmp_1839 = MUX_s_1_2_2(nor_244_nl, and_368_nl, fsm_output[6]);
  assign and_dcpl_199 = and_dcpl_132 & and_dcpl_28;
  assign and_dcpl_200 = and_dcpl_19 & and_dcpl_43;
  assign and_dcpl_201 = and_dcpl_108 & and_dcpl_39;
  assign and_dcpl_202 = and_dcpl_112 & and_dcpl_48;
  assign and_dcpl_203 = and_dcpl_117 & and_dcpl_60;
  assign and_dcpl_204 = and_dcpl_19 & and_dcpl_71;
  assign and_dcpl_206 = and_dcpl_74 & and_dcpl_32 & and_dcpl_73;
  assign and_dcpl_207 = and_dcpl_80 & and_dcpl_29;
  assign and_dcpl_208 = and_dcpl_207 & and_dcpl_83;
  assign and_dcpl_210 = and_dcpl_86 & and_dcpl_32 & and_dcpl_85;
  assign and_dcpl_212 = and_dcpl_67 & and_dcpl_29 & and_dcpl_85;
  assign and_dcpl_214 = and_dcpl_67 & and_dcpl_32 & and_dcpl_94;
  assign and_dcpl_215 = and_dcpl_207 & and_dcpl_101;
  assign and_dcpl_217 = and_dcpl_80 & and_dcpl_32 & and_dcpl_103;
  assign and_dcpl_219 = and_dcpl_74 & and_dcpl_29 & and_dcpl_103;
  assign and_dcpl_220 = and_dcpl_55 & and_dcpl_111;
  assign and_dcpl_221 = and_dcpl_61 & and_dcpl_107;
  assign or_tmp_2035 = (~ (fsm_output[2])) | (fsm_output[9]) | (fsm_output[8]);
  assign mux_tmp_1861 = MUX_s_1_2_2(or_tmp_2035, (fsm_output[8]), fsm_output[3]);
  assign or_tmp_2037 = and_376_cse | (fsm_output[9:8]!=2'b01);
  assign mux_tmp_1863 = MUX_s_1_2_2(mux_tmp_1861, or_tmp_2037, fsm_output[7]);
  assign or_tmp_2040 = (~((~ (fsm_output[2])) | (fsm_output[9]))) | (fsm_output[8]);
  assign or_tmp_2041 = (fsm_output[3]) | or_tmp_2040;
  assign mux_tmp_1866 = MUX_s_1_2_2(or_tmp_2041, mux_tmp_1861, fsm_output[7]);
  assign or_tmp_2043 = (~ (fsm_output[2])) | (fsm_output[9]) | (~ (fsm_output[8]));
  assign or_tmp_2044 = (fsm_output[2]) | (~ (fsm_output[9])) | (fsm_output[8]);
  assign mux_1920_cse = MUX_s_1_2_2(or_tmp_2044, or_tmp_2043, fsm_output[3]);
  assign mux_tmp_1870 = MUX_s_1_2_2(or_tmp_2037, mux_1920_cse, fsm_output[7]);
  assign or_2086_cse = (fsm_output[9:8]!=2'b10);
  assign mux_1922_cse = MUX_s_1_2_2(or_2086_cse, or_tmp_2043, fsm_output[3]);
  assign mux_tmp_1872 = MUX_s_1_2_2(or_212_cse, mux_1922_cse, fsm_output[7]);
  assign or_tmp_2047 = (~((fsm_output[2]) | (~ (fsm_output[9])))) | (fsm_output[8]);
  assign mux_tmp_1874 = MUX_s_1_2_2(or_tmp_2035, or_tmp_2047, fsm_output[3]);
  assign mux_tmp_1875 = MUX_s_1_2_2(mux_tmp_1874, or_tmp_2037, fsm_output[7]);
  assign nand_tmp_134 = ~((fsm_output[3]) & (~ or_tmp_2047));
  assign mux_tmp_1876 = MUX_s_1_2_2(nand_tmp_134, or_tmp_2037, fsm_output[7]);
  assign mux_tmp_1877 = MUX_s_1_2_2(mux_tmp_1876, mux_tmp_1875, fsm_output[0]);
  assign mux_tmp_1882 = MUX_s_1_2_2(or_212_cse, or_tmp_2041, fsm_output[7]);
  assign mux_tmp_1883 = MUX_s_1_2_2(mux_tmp_1882, mux_tmp_1872, fsm_output[0]);
  assign mux_1938_cse = MUX_s_1_2_2(or_tmp_2040, or_tmp_2044, fsm_output[3]);
  assign mux_tmp_1888 = MUX_s_1_2_2(mux_1938_cse, mux_tmp_1861, fsm_output[7]);
  assign or_2091_nl = (~((fsm_output[3:2]!=2'b00))) | (fsm_output[9:8]!=2'b01);
  assign mux_tmp_1891 = MUX_s_1_2_2(or_2091_nl, or_tmp_2041, fsm_output[7]);
  assign STAGE_LOOP_i_3_0_sva_mx0c1 = and_dcpl_19 & and_dcpl_23 & nor_tmp_14;
  assign VEC_LOOP_j_sva_9_0_mx0c1 = and_dcpl_40 & and_dcpl_27 & nor_tmp_14;
  assign vec_rsc_0_0_i_d_d_pff = modulo_dev_cmp_return_rsc_z;
  assign and_42_nl = and_dcpl_30 & and_dcpl_28;
  assign and_52_nl = and_dcpl_40 & and_dcpl_39;
  assign and_57_nl = and_dcpl_45 & and_dcpl_39;
  assign and_67_nl = and_dcpl_55 & and_dcpl_15;
  assign and_73_nl = and_dcpl_61 & and_dcpl_60;
  assign and_80_nl = and_dcpl_68 & and_dcpl_65;
  assign and_87_nl = and_dcpl_75 & and_dcpl_73;
  assign and_93_nl = and_dcpl_81 & and_dcpl_79;
  assign and_99_nl = and_dcpl_87 & and_dcpl_85;
  assign and_103_nl = and_dcpl_68 & and_dcpl_91;
  assign and_107_nl = and_dcpl_95 & and_dcpl_94;
  assign and_111_nl = and_dcpl_81 & and_dcpl_99;
  assign and_116_nl = and_dcpl_80 & and_dcpl_16 & and_dcpl_103;
  assign and_120_nl = and_dcpl_108 & and_dcpl_107;
  assign and_124_nl = and_dcpl_112 & and_dcpl_111;
  assign and_129_nl = and_dcpl_117 & and_dcpl_116;
  assign vec_rsc_0_0_i_radr_d_pff = MUX1HOT_v_6_17_2(z_out_4, (z_out_6_10_1[9:4]),
      (COMP_LOOP_acc_1_cse_2_sva[9:4]), (COMP_LOOP_acc_11_psp_sva[8:3]), (COMP_LOOP_acc_1_cse_4_sva[9:4]),
      (COMP_LOOP_acc_13_psp_sva[7:2]), (COMP_LOOP_acc_1_cse_6_sva[9:4]), (COMP_LOOP_acc_14_psp_sva[8:3]),
      (COMP_LOOP_acc_1_cse_8_sva[9:4]), (COMP_LOOP_acc_16_psp_sva[6:1]), (COMP_LOOP_acc_1_cse_10_sva[9:4]),
      (COMP_LOOP_acc_17_psp_sva[8:3]), (COMP_LOOP_acc_1_cse_12_sva[9:4]), (COMP_LOOP_acc_19_psp_sva[7:2]),
      (COMP_LOOP_acc_1_cse_14_sva[9:4]), (COMP_LOOP_acc_20_psp_sva[8:3]), (COMP_LOOP_acc_1_cse_sva[9:4]),
      {and_42_nl , modExp_dev_while_or_2_cse , and_52_nl , and_57_nl , and_67_nl
      , and_73_nl , and_80_nl , and_87_nl , and_93_nl , and_99_nl , and_103_nl ,
      and_107_nl , and_111_nl , and_116_nl , and_120_nl , and_124_nl , and_129_nl});
  assign and_131_nl = and_dcpl_40 & and_dcpl_60;
  assign mux_524_nl = MUX_s_1_2_2(or_279_cse, nand_tmp_7, fsm_output[6]);
  assign or_280_nl = (~ (fsm_output[4])) | (fsm_output[0]) | mux_524_nl;
  assign mux_521_nl = MUX_s_1_2_2(nand_tmp_7, or_tmp_239, fsm_output[6]);
  assign mux_522_nl = MUX_s_1_2_2(or_1973_cse, mux_521_nl, fsm_output[0]);
  assign or_275_nl = (~ (fsm_output[0])) | (~ (fsm_output[6])) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[3]);
  assign mux_523_nl = MUX_s_1_2_2(mux_522_nl, or_275_nl, fsm_output[4]);
  assign mux_525_nl = MUX_s_1_2_2(or_280_nl, mux_523_nl, fsm_output[5]);
  assign or_271_nl = (~ (fsm_output[9])) | (~ (fsm_output[8])) | (fsm_output[3]);
  assign mux_516_nl = MUX_s_1_2_2(or_271_nl, or_tmp_241, fsm_output[7]);
  assign or_272_nl = (fsm_output[2]) | mux_516_nl;
  assign mux_517_nl = MUX_s_1_2_2(or_272_nl, nand_tmp_6, fsm_output[6]);
  assign mux_518_nl = MUX_s_1_2_2(or_1967_cse, mux_517_nl, fsm_output[0]);
  assign or_274_nl = (fsm_output[4]) | mux_518_nl;
  assign mux_515_nl = MUX_s_1_2_2(or_tmp_239, nand_tmp_6, fsm_output[6]);
  assign or_269_nl = (~ (fsm_output[4])) | (fsm_output[0]) | mux_515_nl;
  assign mux_519_nl = MUX_s_1_2_2(or_274_nl, or_269_nl, fsm_output[5]);
  assign mux_526_nl = MUX_s_1_2_2(mux_525_nl, mux_519_nl, fsm_output[1]);
  assign and_132_nl = and_dcpl_45 & and_dcpl_60;
  assign and_134_nl = and_dcpl_89 & and_dcpl_122;
  assign and_135_nl = and_dcpl_87 & and_dcpl_65;
  assign and_136_nl = and_dcpl_68 & and_dcpl_43;
  assign and_137_nl = and_dcpl_75 & and_dcpl_85;
  assign and_138_nl = and_dcpl_81 & and_dcpl_94;
  assign and_139_nl = and_dcpl_87 & and_dcpl_91;
  assign and_140_nl = and_dcpl_68 & and_dcpl_71;
  assign and_142_nl = and_dcpl_95 & and_dcpl_130;
  assign and_144_nl = and_dcpl_132 & and_dcpl_111;
  assign and_145_nl = and_dcpl_19 & and_dcpl_107;
  assign and_146_nl = and_dcpl_108 & and_dcpl_116;
  assign and_148_nl = and_dcpl_112 & and_dcpl_136;
  assign and_150_nl = and_dcpl_117 & and_dcpl_138;
  assign and_152_nl = and_dcpl_19 & and_dcpl_47 & nor_tmp_14;
  assign vec_rsc_0_0_i_wadr_d_pff = MUX1HOT_v_6_17_2(COMP_LOOP_acc_psp_sva, ({COMP_LOOP_acc_10_cse_10_1_1_sva_9_5
      , (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[4])}), (COMP_LOOP_acc_1_cse_2_sva[9:4]),
      (COMP_LOOP_acc_11_psp_sva[8:3]), (COMP_LOOP_acc_1_cse_4_sva[9:4]), (COMP_LOOP_acc_13_psp_sva[7:2]),
      (COMP_LOOP_acc_1_cse_6_sva[9:4]), (COMP_LOOP_acc_14_psp_sva[8:3]), (COMP_LOOP_acc_1_cse_8_sva[9:4]),
      (COMP_LOOP_acc_16_psp_sva[6:1]), (COMP_LOOP_acc_1_cse_10_sva[9:4]), (COMP_LOOP_acc_17_psp_sva[8:3]),
      (COMP_LOOP_acc_1_cse_12_sva[9:4]), (COMP_LOOP_acc_19_psp_sva[7:2]), (COMP_LOOP_acc_1_cse_14_sva[9:4]),
      (COMP_LOOP_acc_20_psp_sva[8:3]), (COMP_LOOP_acc_1_cse_sva[9:4]), {and_131_nl
      , (~ mux_526_nl) , and_132_nl , and_134_nl , and_135_nl , and_136_nl , and_137_nl
      , and_138_nl , and_139_nl , and_140_nl , and_142_nl , and_144_nl , and_145_nl
      , and_146_nl , and_148_nl , and_150_nl , and_152_nl});
  assign or_319_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b0000) | (fsm_output[5]) | (fsm_output[1]);
  assign mux_552_nl = MUX_s_1_2_2(or_tmp_259, or_319_nl, fsm_output[0]);
  assign or_318_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0000) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_551_nl = MUX_s_1_2_2(or_318_nl, or_tmp_253, fsm_output[0]);
  assign mux_553_nl = MUX_s_1_2_2(mux_552_nl, mux_551_nl, fsm_output[4]);
  assign nand_10_nl = ~((fsm_output[6]) & (~ mux_553_nl));
  assign or_317_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0000);
  assign mux_554_nl = MUX_s_1_2_2(nand_10_nl, or_317_nl, fsm_output[7]);
  assign nor_689_nl = ~((fsm_output[8]) | mux_554_nl);
  assign nor_690_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000) | (~ (fsm_output[7]))
      | (~ (fsm_output[6])) | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[5]) | (~ (fsm_output[1])));
  assign or_313_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0000) | (fsm_output[5]) |
      (~ (fsm_output[1]));
  assign mux_549_nl = MUX_s_1_2_2(or_313_nl, or_tmp_259, fsm_output[0]);
  assign nor_691_nl = ~((fsm_output[7]) | (fsm_output[6]) | (fsm_output[4]) | mux_549_nl);
  assign mux_550_nl = MUX_s_1_2_2(nor_690_nl, nor_691_nl, fsm_output[8]);
  assign mux_555_nl = MUX_s_1_2_2(nor_689_nl, mux_550_nl, fsm_output[9]);
  assign or_310_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign or_308_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0000) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_544_nl = MUX_s_1_2_2(or_308_nl, or_tmp_259, fsm_output[0]);
  assign or_306_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b000)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_543_nl = MUX_s_1_2_2(or_tmp_258, or_306_nl, fsm_output[0]);
  assign mux_545_nl = MUX_s_1_2_2(mux_544_nl, mux_543_nl, fsm_output[4]);
  assign or_304_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0000) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_542_nl = MUX_s_1_2_2(or_304_nl, or_tmp_253, fsm_output[0]);
  assign or_305_nl = (fsm_output[4]) | mux_542_nl;
  assign mux_546_nl = MUX_s_1_2_2(mux_545_nl, or_305_nl, fsm_output[6]);
  assign mux_547_nl = MUX_s_1_2_2(or_310_nl, mux_546_nl, fsm_output[7]);
  assign and_344_nl = (fsm_output[8]) & (~ mux_547_nl);
  assign nor_692_nl = ~((fsm_output[8]) | (fsm_output[7]) | (fsm_output[6]) | (~
      (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0000));
  assign mux_548_nl = MUX_s_1_2_2(and_344_nl, nor_692_nl, fsm_output[9]);
  assign mux_556_nl = MUX_s_1_2_2(mux_555_nl, mux_548_nl, fsm_output[3]);
  assign or_301_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b000) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5]) | (~ (fsm_output[1]));
  assign or_299_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0000) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_537_nl = MUX_s_1_2_2(or_299_nl, or_tmp_259, fsm_output[0]);
  assign or_297_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_536_nl = MUX_s_1_2_2(or_tmp_258, or_297_nl, fsm_output[0]);
  assign mux_538_nl = MUX_s_1_2_2(mux_537_nl, mux_536_nl, fsm_output[4]);
  assign mux_539_nl = MUX_s_1_2_2(or_301_nl, mux_538_nl, fsm_output[6]);
  assign or_295_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0000) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_534_nl = MUX_s_1_2_2(or_295_nl, or_tmp_253, fsm_output[0]);
  assign or_296_nl = (fsm_output[4]) | mux_534_nl;
  assign mux_535_nl = MUX_s_1_2_2(or_296_nl, or_tmp_252, fsm_output[6]);
  assign mux_540_nl = MUX_s_1_2_2(mux_539_nl, mux_535_nl, fsm_output[7]);
  assign nor_693_nl = ~((fsm_output[9:8]!=2'b10) | mux_540_nl);
  assign or_292_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000)
      | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5]) | (~ (fsm_output[1]));
  assign or_290_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0000) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_530_nl = MUX_s_1_2_2(or_290_nl, or_tmp_259, fsm_output[0]);
  assign or_286_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_529_nl = MUX_s_1_2_2(or_tmp_258, or_286_nl, fsm_output[0]);
  assign mux_531_nl = MUX_s_1_2_2(mux_530_nl, mux_529_nl, fsm_output[4]);
  assign mux_532_nl = MUX_s_1_2_2(or_292_nl, mux_531_nl, fsm_output[6]);
  assign nand_8_nl = ~((fsm_output[7]) & (~ mux_532_nl));
  assign or_283_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0000) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_527_nl = MUX_s_1_2_2(or_283_nl, or_tmp_253, fsm_output[0]);
  assign or_284_nl = (fsm_output[4]) | mux_527_nl;
  assign mux_528_nl = MUX_s_1_2_2(or_284_nl, or_tmp_252, fsm_output[6]);
  assign or_285_nl = (fsm_output[7]) | mux_528_nl;
  assign mux_533_nl = MUX_s_1_2_2(nand_8_nl, or_285_nl, fsm_output[8]);
  assign nor_694_nl = ~((fsm_output[9]) | mux_533_nl);
  assign mux_541_nl = MUX_s_1_2_2(nor_693_nl, nor_694_nl, fsm_output[3]);
  assign vec_rsc_0_0_i_we_d_pff = MUX_s_1_2_2(mux_556_nl, mux_541_nl, fsm_output[2]);
  assign nor_678_cse = ~((z_out_6_10_1[3:0]!=4'b0000) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign or_368_cse = (z_out_6_10_1[3:0]!=4'b0000) | not_tmp_133;
  assign or_369_cse = (z_out_6_10_1[3:0]!=4'b0000) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_372_nl = (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0000) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_371_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | not_tmp_134;
  assign mux_583_nl = MUX_s_1_2_2(or_371_nl, or_369_cse, fsm_output[0]);
  assign mux_584_nl = MUX_s_1_2_2(or_372_nl, mux_583_nl, fsm_output[6]);
  assign or_366_nl = (z_out_6_10_1[3:0]!=4'b0000) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_581_nl = MUX_s_1_2_2(or_368_cse, or_366_nl, fsm_output[0]);
  assign or_365_nl = (VEC_LOOP_j_sva_9_0[0]) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_363_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0000) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_580_nl = MUX_s_1_2_2(or_365_nl, or_363_nl, fsm_output[0]);
  assign mux_582_nl = MUX_s_1_2_2(mux_581_nl, mux_580_nl, fsm_output[6]);
  assign mux_585_nl = MUX_s_1_2_2(mux_584_nl, mux_582_nl, fsm_output[1]);
  assign nor_669_nl = ~((fsm_output[3]) | mux_585_nl);
  assign or_361_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b0000) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_359_nl = (z_out_6_10_1[3:0]!=4'b0000) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]);
  assign mux_577_nl = MUX_s_1_2_2(or_361_nl, or_359_nl, fsm_output[0]);
  assign or_358_nl = (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b0000) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_578_nl = MUX_s_1_2_2(mux_577_nl, or_358_nl, fsm_output[6]);
  assign nor_670_nl = ~((fsm_output[1]) | mux_578_nl);
  assign nor_671_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0000) | (~ (fsm_output[1]))
      | (~ (fsm_output[6])) | (~ (fsm_output[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | not_tmp_133);
  assign mux_579_nl = MUX_s_1_2_2(nor_670_nl, nor_671_nl, fsm_output[3]);
  assign mux_586_nl = MUX_s_1_2_2(nor_669_nl, mux_579_nl, fsm_output[2]);
  assign nor_672_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b0000)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign nor_673_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0000) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | not_tmp_133);
  assign nor_674_nl = ~((VEC_LOOP_j_sva_9_0[0]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b000)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_675_nl = ~((z_out_6_10_1[3:0]!=4'b0000) | not_tmp_133);
  assign mux_573_nl = MUX_s_1_2_2(nor_674_nl, nor_675_nl, fsm_output[0]);
  assign mux_574_nl = MUX_s_1_2_2(nor_673_nl, mux_573_nl, fsm_output[6]);
  assign and_342_nl = (fsm_output[1]) & mux_574_nl;
  assign mux_575_nl = MUX_s_1_2_2(nor_672_nl, and_342_nl, fsm_output[3]);
  assign nor_676_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b000)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_677_nl = ~((z_out_6_10_1[3:0]!=4'b0000) | (fsm_output[5]) | not_tmp_134);
  assign mux_570_nl = MUX_s_1_2_2(nor_676_nl, nor_677_nl, fsm_output[0]);
  assign nor_679_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_569_nl = MUX_s_1_2_2(nor_678_cse, nor_679_nl, fsm_output[0]);
  assign mux_571_nl = MUX_s_1_2_2(mux_570_nl, mux_569_nl, fsm_output[6]);
  assign nor_680_nl = ~((VEC_LOOP_j_sva_9_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_681_nl = ~((z_out_6_10_1[3:0]!=4'b0000) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_567_nl = MUX_s_1_2_2(nor_680_nl, nor_681_nl, fsm_output[0]);
  assign nor_682_nl = ~((z_out_6_10_1[3:0]!=4'b0000) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[4]));
  assign mux_568_nl = MUX_s_1_2_2(mux_567_nl, nor_682_nl, fsm_output[6]);
  assign mux_572_nl = MUX_s_1_2_2(mux_571_nl, mux_568_nl, fsm_output[1]);
  assign and_343_nl = (fsm_output[3]) & mux_572_nl;
  assign mux_576_nl = MUX_s_1_2_2(mux_575_nl, and_343_nl, fsm_output[2]);
  assign mux_587_nl = MUX_s_1_2_2(mux_586_nl, mux_576_nl, fsm_output[8]);
  assign nor_685_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_563_nl = MUX_s_1_2_2(nor_678_cse, nor_685_nl, fsm_output[0]);
  assign nor_686_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_687_nl = ~((z_out_6_10_1[3:0]!=4'b0000) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_562_nl = MUX_s_1_2_2(nor_686_nl, nor_687_nl, fsm_output[0]);
  assign mux_564_nl = MUX_s_1_2_2(mux_563_nl, mux_562_nl, fsm_output[6]);
  assign nor_688_nl = ~((z_out_6_10_1[3:0]!=4'b0000) | (fsm_output[6]) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_565_nl = MUX_s_1_2_2(mux_564_nl, nor_688_nl, fsm_output[1]);
  assign nand_11_nl = ~((fsm_output[3]) & mux_565_nl);
  assign or_328_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0000) | (~ (fsm_output[6]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[5])
      | not_tmp_134;
  assign or_326_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_559_nl = MUX_s_1_2_2(or_326_nl, or_368_cse, fsm_output[0]);
  assign or_322_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0000) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_558_nl = MUX_s_1_2_2(or_369_cse, or_322_nl, fsm_output[0]);
  assign mux_560_nl = MUX_s_1_2_2(mux_559_nl, mux_558_nl, fsm_output[6]);
  assign mux_561_nl = MUX_s_1_2_2(or_328_nl, mux_560_nl, fsm_output[1]);
  assign or_329_nl = (fsm_output[3]) | mux_561_nl;
  assign mux_566_nl = MUX_s_1_2_2(nand_11_nl, or_329_nl, fsm_output[2]);
  assign nor_683_nl = ~((fsm_output[8]) | mux_566_nl);
  assign vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_587_nl,
      nor_683_nl, fsm_output[9]);
  assign or_413_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b0001) | (fsm_output[1]) | (fsm_output[5]);
  assign mux_614_nl = MUX_s_1_2_2(or_tmp_353, or_413_nl, fsm_output[0]);
  assign or_412_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0001) | (fsm_output[1])
      | (~ (fsm_output[5]));
  assign mux_613_nl = MUX_s_1_2_2(or_412_nl, or_tmp_346, fsm_output[0]);
  assign mux_615_nl = MUX_s_1_2_2(mux_614_nl, mux_613_nl, fsm_output[4]);
  assign nor_661_nl = ~((fsm_output[9]) | (~ (fsm_output[6])) | mux_615_nl);
  assign or_410_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b000) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_9_0[0])) | (~ (fsm_output[1])) |
      (fsm_output[5]);
  assign or_409_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0001) | (~ (fsm_output[1]))
      | (fsm_output[5]);
  assign mux_610_nl = MUX_s_1_2_2(or_409_nl, or_tmp_353, fsm_output[0]);
  assign or_408_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (fsm_output[1]) | (~ (fsm_output[5]));
  assign mux_609_nl = MUX_s_1_2_2(or_tmp_352, or_408_nl, fsm_output[0]);
  assign mux_611_nl = MUX_s_1_2_2(mux_610_nl, mux_609_nl, fsm_output[4]);
  assign mux_612_nl = MUX_s_1_2_2(or_410_nl, mux_611_nl, fsm_output[6]);
  assign and_341_nl = (fsm_output[9]) & (~ mux_612_nl);
  assign mux_616_nl = MUX_s_1_2_2(nor_661_nl, and_341_nl, fsm_output[2]);
  assign or_405_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0001) | (~ (fsm_output[1]))
      | (fsm_output[5]);
  assign mux_608_nl = MUX_s_1_2_2(or_405_nl, or_tmp_353, fsm_output[0]);
  assign nor_662_nl = ~((fsm_output[2]) | (~ (fsm_output[9])) | (fsm_output[6]) |
      (fsm_output[4]) | mux_608_nl);
  assign mux_617_nl = MUX_s_1_2_2(mux_616_nl, nor_662_nl, fsm_output[8]);
  assign or_402_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (fsm_output[1])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0001);
  assign or_401_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_9_0[0])) |
      (~ (fsm_output[1])) | (fsm_output[5]);
  assign mux_606_nl = MUX_s_1_2_2(or_402_nl, or_401_nl, fsm_output[9]);
  assign or_399_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0001) | (fsm_output[1])
      | (~ (fsm_output[5]));
  assign mux_604_nl = MUX_s_1_2_2(or_399_nl, or_tmp_346, fsm_output[0]);
  assign or_400_nl = (fsm_output[4]) | mux_604_nl;
  assign mux_605_nl = MUX_s_1_2_2(or_400_nl, or_tmp_362, fsm_output[6]);
  assign nand_14_nl = ~((fsm_output[9]) & (~ mux_605_nl));
  assign mux_607_nl = MUX_s_1_2_2(mux_606_nl, nand_14_nl, fsm_output[2]);
  assign nor_663_nl = ~((fsm_output[8]) | mux_607_nl);
  assign mux_618_nl = MUX_s_1_2_2(mux_617_nl, nor_663_nl, fsm_output[7]);
  assign nor_664_nl = ~((fsm_output[2]) | (~ (fsm_output[9])) | (fsm_output[6]) |
      (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[5]) |
      (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0001));
  assign nor_665_nl = ~((fsm_output[9]) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000)
      | (~ (fsm_output[6])) | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_9_0[0]))
      | (~ (fsm_output[1])) | (fsm_output[5]));
  assign or_393_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0001) | (fsm_output[1])
      | (~ (fsm_output[5]));
  assign mux_599_nl = MUX_s_1_2_2(or_393_nl, or_tmp_346, fsm_output[0]);
  assign or_394_nl = (fsm_output[4]) | mux_599_nl;
  assign mux_600_nl = MUX_s_1_2_2(or_394_nl, or_tmp_362, fsm_output[6]);
  assign nor_666_nl = ~((fsm_output[9]) | mux_600_nl);
  assign mux_601_nl = MUX_s_1_2_2(nor_665_nl, nor_666_nl, fsm_output[2]);
  assign mux_602_nl = MUX_s_1_2_2(nor_664_nl, mux_601_nl, fsm_output[8]);
  assign or_389_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000)
      | (~ (VEC_LOOP_j_sva_9_0[0])) | (~ (fsm_output[1])) | (fsm_output[5]);
  assign or_388_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0001) | (~ (fsm_output[1]))
      | (fsm_output[5]);
  assign mux_595_nl = MUX_s_1_2_2(or_388_nl, or_tmp_353, fsm_output[0]);
  assign or_387_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (fsm_output[1]) | (~ (fsm_output[5]));
  assign mux_594_nl = MUX_s_1_2_2(or_tmp_352, or_387_nl, fsm_output[0]);
  assign mux_596_nl = MUX_s_1_2_2(mux_595_nl, mux_594_nl, fsm_output[4]);
  assign mux_597_nl = MUX_s_1_2_2(or_389_nl, mux_596_nl, fsm_output[6]);
  assign nor_667_nl = ~((~ (fsm_output[2])) | (fsm_output[9]) | mux_597_nl);
  assign or_383_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0001) | (~ (fsm_output[1]))
      | (fsm_output[5]);
  assign mux_591_nl = MUX_s_1_2_2(or_383_nl, or_tmp_353, fsm_output[0]);
  assign or_380_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b001)
      | (fsm_output[1]) | (~ (fsm_output[5]));
  assign mux_590_nl = MUX_s_1_2_2(or_tmp_352, or_380_nl, fsm_output[0]);
  assign mux_592_nl = MUX_s_1_2_2(mux_591_nl, mux_590_nl, fsm_output[4]);
  assign or_377_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0001) | (fsm_output[1])
      | (~ (fsm_output[5]));
  assign mux_589_nl = MUX_s_1_2_2(or_377_nl, or_tmp_346, fsm_output[0]);
  assign or_378_nl = (fsm_output[4]) | mux_589_nl;
  assign mux_593_nl = MUX_s_1_2_2(mux_592_nl, or_378_nl, fsm_output[6]);
  assign nor_668_nl = ~((fsm_output[2]) | (fsm_output[9]) | mux_593_nl);
  assign mux_598_nl = MUX_s_1_2_2(nor_667_nl, nor_668_nl, fsm_output[8]);
  assign mux_603_nl = MUX_s_1_2_2(mux_602_nl, mux_598_nl, fsm_output[7]);
  assign vec_rsc_0_1_i_we_d_pff = MUX_s_1_2_2(mux_618_nl, mux_603_nl, fsm_output[3]);
  assign nor_650_cse = ~((z_out_6_10_1[3:0]!=4'b0001) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign or_462_cse = (z_out_6_10_1[3:0]!=4'b0001) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_465_nl = (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0001) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_464_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | not_tmp_134;
  assign mux_645_nl = MUX_s_1_2_2(or_464_nl, or_462_cse, fsm_output[0]);
  assign mux_646_nl = MUX_s_1_2_2(or_465_nl, mux_645_nl, fsm_output[6]);
  assign or_461_nl = (z_out_6_10_1[3:1]!=3'b000) | nand_308_cse;
  assign or_459_nl = (z_out_6_10_1[3:0]!=4'b0001) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_643_nl = MUX_s_1_2_2(or_461_nl, or_459_nl, fsm_output[0]);
  assign or_458_nl = (~ (VEC_LOOP_j_sva_9_0[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_456_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0001) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_642_nl = MUX_s_1_2_2(or_458_nl, or_456_nl, fsm_output[0]);
  assign mux_644_nl = MUX_s_1_2_2(mux_643_nl, mux_642_nl, fsm_output[6]);
  assign mux_647_nl = MUX_s_1_2_2(mux_646_nl, mux_644_nl, fsm_output[1]);
  assign nor_641_nl = ~((fsm_output[3]) | mux_647_nl);
  assign or_454_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b0001) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_452_nl = (z_out_6_10_1[3:0]!=4'b0001) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]);
  assign mux_639_nl = MUX_s_1_2_2(or_454_nl, or_452_nl, fsm_output[0]);
  assign or_451_nl = (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b0001) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_640_nl = MUX_s_1_2_2(mux_639_nl, or_451_nl, fsm_output[6]);
  assign nor_642_nl = ~((fsm_output[1]) | mux_640_nl);
  assign nor_643_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0001) | (~ (fsm_output[1]))
      | (~ (fsm_output[6])) | (~ (fsm_output[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | not_tmp_133);
  assign mux_641_nl = MUX_s_1_2_2(nor_642_nl, nor_643_nl, fsm_output[3]);
  assign mux_648_nl = MUX_s_1_2_2(nor_641_nl, mux_641_nl, fsm_output[2]);
  assign nor_644_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b0001)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign nor_645_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0001) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | not_tmp_133);
  assign nor_646_nl = ~((~ (VEC_LOOP_j_sva_9_0[0])) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b000)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_647_nl = ~((z_out_6_10_1[3:0]!=4'b0001) | not_tmp_133);
  assign mux_635_nl = MUX_s_1_2_2(nor_646_nl, nor_647_nl, fsm_output[0]);
  assign mux_636_nl = MUX_s_1_2_2(nor_645_nl, mux_635_nl, fsm_output[6]);
  assign and_339_nl = (fsm_output[1]) & mux_636_nl;
  assign mux_637_nl = MUX_s_1_2_2(nor_644_nl, and_339_nl, fsm_output[3]);
  assign nor_648_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b001)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_649_nl = ~((z_out_6_10_1[3:0]!=4'b0001) | (fsm_output[5]) | not_tmp_134);
  assign mux_632_nl = MUX_s_1_2_2(nor_648_nl, nor_649_nl, fsm_output[0]);
  assign nor_651_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_631_nl = MUX_s_1_2_2(nor_650_cse, nor_651_nl, fsm_output[0]);
  assign mux_633_nl = MUX_s_1_2_2(mux_632_nl, mux_631_nl, fsm_output[6]);
  assign nor_652_nl = ~((~ (VEC_LOOP_j_sva_9_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_653_nl = ~((z_out_6_10_1[3:0]!=4'b0001) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_629_nl = MUX_s_1_2_2(nor_652_nl, nor_653_nl, fsm_output[0]);
  assign nor_654_nl = ~((z_out_6_10_1[3:0]!=4'b0001) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[4]));
  assign mux_630_nl = MUX_s_1_2_2(mux_629_nl, nor_654_nl, fsm_output[6]);
  assign mux_634_nl = MUX_s_1_2_2(mux_633_nl, mux_630_nl, fsm_output[1]);
  assign and_340_nl = (fsm_output[3]) & mux_634_nl;
  assign mux_638_nl = MUX_s_1_2_2(mux_637_nl, and_340_nl, fsm_output[2]);
  assign mux_649_nl = MUX_s_1_2_2(mux_648_nl, mux_638_nl, fsm_output[8]);
  assign nor_657_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_625_nl = MUX_s_1_2_2(nor_650_cse, nor_657_nl, fsm_output[0]);
  assign nor_658_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_659_nl = ~((z_out_6_10_1[3:0]!=4'b0001) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_624_nl = MUX_s_1_2_2(nor_658_nl, nor_659_nl, fsm_output[0]);
  assign mux_626_nl = MUX_s_1_2_2(mux_625_nl, mux_624_nl, fsm_output[6]);
  assign nor_660_nl = ~((z_out_6_10_1[3:0]!=4'b0001) | (fsm_output[6]) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_627_nl = MUX_s_1_2_2(mux_626_nl, nor_660_nl, fsm_output[1]);
  assign nand_17_nl = ~((fsm_output[3]) & mux_627_nl);
  assign or_421_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0001) | (~ (fsm_output[6]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[5])
      | not_tmp_134;
  assign or_419_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000) | (~ (VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_418_nl = (z_out_6_10_1[3:0]!=4'b0001) | not_tmp_133;
  assign mux_621_nl = MUX_s_1_2_2(or_419_nl, or_418_nl, fsm_output[0]);
  assign or_415_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0001) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_620_nl = MUX_s_1_2_2(or_462_cse, or_415_nl, fsm_output[0]);
  assign mux_622_nl = MUX_s_1_2_2(mux_621_nl, mux_620_nl, fsm_output[6]);
  assign mux_623_nl = MUX_s_1_2_2(or_421_nl, mux_622_nl, fsm_output[1]);
  assign or_422_nl = (fsm_output[3]) | mux_623_nl;
  assign mux_628_nl = MUX_s_1_2_2(nand_17_nl, or_422_nl, fsm_output[2]);
  assign nor_655_nl = ~((fsm_output[8]) | mux_628_nl);
  assign vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_649_nl,
      nor_655_nl, fsm_output[9]);
  assign or_505_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b0010) | (fsm_output[5]) | (fsm_output[1]);
  assign mux_676_nl = MUX_s_1_2_2(or_tmp_445, or_505_nl, fsm_output[0]);
  assign or_504_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0010) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_675_nl = MUX_s_1_2_2(or_504_nl, or_tmp_439, fsm_output[0]);
  assign mux_677_nl = MUX_s_1_2_2(mux_676_nl, mux_675_nl, fsm_output[4]);
  assign nand_22_nl = ~((fsm_output[6]) & (~ mux_677_nl));
  assign or_503_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0010);
  assign mux_678_nl = MUX_s_1_2_2(nand_22_nl, or_503_nl, fsm_output[7]);
  assign nor_635_nl = ~((fsm_output[8]) | mux_678_nl);
  assign nor_636_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001) | (~ (fsm_output[7]))
      | (~ (fsm_output[6])) | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[5]) | (~ (fsm_output[1])));
  assign or_499_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0010) | (fsm_output[5]) |
      (~ (fsm_output[1]));
  assign mux_673_nl = MUX_s_1_2_2(or_499_nl, or_tmp_445, fsm_output[0]);
  assign nor_637_nl = ~((fsm_output[7]) | (fsm_output[6]) | (fsm_output[4]) | mux_673_nl);
  assign mux_674_nl = MUX_s_1_2_2(nor_636_nl, nor_637_nl, fsm_output[8]);
  assign mux_679_nl = MUX_s_1_2_2(nor_635_nl, mux_674_nl, fsm_output[9]);
  assign or_496_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign or_494_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0010) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_668_nl = MUX_s_1_2_2(or_494_nl, or_tmp_445, fsm_output[0]);
  assign or_492_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b010)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_667_nl = MUX_s_1_2_2(or_tmp_444, or_492_nl, fsm_output[0]);
  assign mux_669_nl = MUX_s_1_2_2(mux_668_nl, mux_667_nl, fsm_output[4]);
  assign or_490_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0010) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_666_nl = MUX_s_1_2_2(or_490_nl, or_tmp_439, fsm_output[0]);
  assign or_491_nl = (fsm_output[4]) | mux_666_nl;
  assign mux_670_nl = MUX_s_1_2_2(mux_669_nl, or_491_nl, fsm_output[6]);
  assign mux_671_nl = MUX_s_1_2_2(or_496_nl, mux_670_nl, fsm_output[7]);
  assign and_338_nl = (fsm_output[8]) & (~ mux_671_nl);
  assign nor_638_nl = ~((fsm_output[8]) | (fsm_output[7]) | (fsm_output[6]) | (~
      (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0010));
  assign mux_672_nl = MUX_s_1_2_2(and_338_nl, nor_638_nl, fsm_output[9]);
  assign mux_680_nl = MUX_s_1_2_2(mux_679_nl, mux_672_nl, fsm_output[3]);
  assign or_487_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b001) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5]) | (~ (fsm_output[1]));
  assign or_485_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0010) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_661_nl = MUX_s_1_2_2(or_485_nl, or_tmp_445, fsm_output[0]);
  assign or_483_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_660_nl = MUX_s_1_2_2(or_tmp_444, or_483_nl, fsm_output[0]);
  assign mux_662_nl = MUX_s_1_2_2(mux_661_nl, mux_660_nl, fsm_output[4]);
  assign mux_663_nl = MUX_s_1_2_2(or_487_nl, mux_662_nl, fsm_output[6]);
  assign or_481_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0010) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_658_nl = MUX_s_1_2_2(or_481_nl, or_tmp_439, fsm_output[0]);
  assign or_482_nl = (fsm_output[4]) | mux_658_nl;
  assign mux_659_nl = MUX_s_1_2_2(or_482_nl, or_tmp_438, fsm_output[6]);
  assign mux_664_nl = MUX_s_1_2_2(mux_663_nl, mux_659_nl, fsm_output[7]);
  assign nor_639_nl = ~((fsm_output[9:8]!=2'b10) | mux_664_nl);
  assign or_478_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001)
      | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5]) | (~ (fsm_output[1]));
  assign or_476_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0010) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_654_nl = MUX_s_1_2_2(or_476_nl, or_tmp_445, fsm_output[0]);
  assign or_472_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_653_nl = MUX_s_1_2_2(or_tmp_444, or_472_nl, fsm_output[0]);
  assign mux_655_nl = MUX_s_1_2_2(mux_654_nl, mux_653_nl, fsm_output[4]);
  assign mux_656_nl = MUX_s_1_2_2(or_478_nl, mux_655_nl, fsm_output[6]);
  assign nand_20_nl = ~((fsm_output[7]) & (~ mux_656_nl));
  assign or_469_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0010) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_651_nl = MUX_s_1_2_2(or_469_nl, or_tmp_439, fsm_output[0]);
  assign or_470_nl = (fsm_output[4]) | mux_651_nl;
  assign mux_652_nl = MUX_s_1_2_2(or_470_nl, or_tmp_438, fsm_output[6]);
  assign or_471_nl = (fsm_output[7]) | mux_652_nl;
  assign mux_657_nl = MUX_s_1_2_2(nand_20_nl, or_471_nl, fsm_output[8]);
  assign nor_640_nl = ~((fsm_output[9]) | mux_657_nl);
  assign mux_665_nl = MUX_s_1_2_2(nor_639_nl, nor_640_nl, fsm_output[3]);
  assign vec_rsc_0_2_i_we_d_pff = MUX_s_1_2_2(mux_680_nl, mux_665_nl, fsm_output[2]);
  assign nor_624_cse = ~((z_out_6_10_1[3:0]!=4'b0010) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign or_554_cse = (z_out_6_10_1[3:0]!=4'b0010) | not_tmp_133;
  assign or_555_cse = (z_out_6_10_1[3:0]!=4'b0010) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_558_nl = (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0010) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_557_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | not_tmp_134;
  assign mux_707_nl = MUX_s_1_2_2(or_557_nl, or_555_cse, fsm_output[0]);
  assign mux_708_nl = MUX_s_1_2_2(or_558_nl, mux_707_nl, fsm_output[6]);
  assign or_552_nl = (z_out_6_10_1[3:0]!=4'b0010) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_705_nl = MUX_s_1_2_2(or_554_cse, or_552_nl, fsm_output[0]);
  assign or_551_nl = (VEC_LOOP_j_sva_9_0[0]) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_549_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0010) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_704_nl = MUX_s_1_2_2(or_551_nl, or_549_nl, fsm_output[0]);
  assign mux_706_nl = MUX_s_1_2_2(mux_705_nl, mux_704_nl, fsm_output[6]);
  assign mux_709_nl = MUX_s_1_2_2(mux_708_nl, mux_706_nl, fsm_output[1]);
  assign nor_615_nl = ~((fsm_output[3]) | mux_709_nl);
  assign or_547_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b0010) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_545_nl = (z_out_6_10_1[3:0]!=4'b0010) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]);
  assign mux_701_nl = MUX_s_1_2_2(or_547_nl, or_545_nl, fsm_output[0]);
  assign or_544_nl = (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b0010) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_702_nl = MUX_s_1_2_2(mux_701_nl, or_544_nl, fsm_output[6]);
  assign nor_616_nl = ~((fsm_output[1]) | mux_702_nl);
  assign nor_617_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0010) | (~ (fsm_output[1]))
      | (~ (fsm_output[6])) | (~ (fsm_output[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | not_tmp_133);
  assign mux_703_nl = MUX_s_1_2_2(nor_616_nl, nor_617_nl, fsm_output[3]);
  assign mux_710_nl = MUX_s_1_2_2(nor_615_nl, mux_703_nl, fsm_output[2]);
  assign nor_618_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b0010)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign nor_619_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0010) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | not_tmp_133);
  assign nor_620_nl = ~((VEC_LOOP_j_sva_9_0[0]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b001)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_621_nl = ~((z_out_6_10_1[3:0]!=4'b0010) | not_tmp_133);
  assign mux_697_nl = MUX_s_1_2_2(nor_620_nl, nor_621_nl, fsm_output[0]);
  assign mux_698_nl = MUX_s_1_2_2(nor_619_nl, mux_697_nl, fsm_output[6]);
  assign and_336_nl = (fsm_output[1]) & mux_698_nl;
  assign mux_699_nl = MUX_s_1_2_2(nor_618_nl, and_336_nl, fsm_output[3]);
  assign nor_622_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b010)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_623_nl = ~((z_out_6_10_1[3:0]!=4'b0010) | (fsm_output[5]) | not_tmp_134);
  assign mux_694_nl = MUX_s_1_2_2(nor_622_nl, nor_623_nl, fsm_output[0]);
  assign nor_625_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_693_nl = MUX_s_1_2_2(nor_624_cse, nor_625_nl, fsm_output[0]);
  assign mux_695_nl = MUX_s_1_2_2(mux_694_nl, mux_693_nl, fsm_output[6]);
  assign nor_626_nl = ~((VEC_LOOP_j_sva_9_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_627_nl = ~((z_out_6_10_1[3:0]!=4'b0010) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_691_nl = MUX_s_1_2_2(nor_626_nl, nor_627_nl, fsm_output[0]);
  assign nor_628_nl = ~((z_out_6_10_1[3:0]!=4'b0010) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[4]));
  assign mux_692_nl = MUX_s_1_2_2(mux_691_nl, nor_628_nl, fsm_output[6]);
  assign mux_696_nl = MUX_s_1_2_2(mux_695_nl, mux_692_nl, fsm_output[1]);
  assign and_337_nl = (fsm_output[3]) & mux_696_nl;
  assign mux_700_nl = MUX_s_1_2_2(mux_699_nl, and_337_nl, fsm_output[2]);
  assign mux_711_nl = MUX_s_1_2_2(mux_710_nl, mux_700_nl, fsm_output[8]);
  assign nor_631_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_687_nl = MUX_s_1_2_2(nor_624_cse, nor_631_nl, fsm_output[0]);
  assign nor_632_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_633_nl = ~((z_out_6_10_1[3:0]!=4'b0010) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_686_nl = MUX_s_1_2_2(nor_632_nl, nor_633_nl, fsm_output[0]);
  assign mux_688_nl = MUX_s_1_2_2(mux_687_nl, mux_686_nl, fsm_output[6]);
  assign nor_634_nl = ~((z_out_6_10_1[3:0]!=4'b0010) | (fsm_output[6]) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_689_nl = MUX_s_1_2_2(mux_688_nl, nor_634_nl, fsm_output[1]);
  assign nand_23_nl = ~((fsm_output[3]) & mux_689_nl);
  assign or_514_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0010) | (~ (fsm_output[6]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[5])
      | not_tmp_134;
  assign or_512_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_683_nl = MUX_s_1_2_2(or_512_nl, or_554_cse, fsm_output[0]);
  assign or_508_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0010) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_682_nl = MUX_s_1_2_2(or_555_cse, or_508_nl, fsm_output[0]);
  assign mux_684_nl = MUX_s_1_2_2(mux_683_nl, mux_682_nl, fsm_output[6]);
  assign mux_685_nl = MUX_s_1_2_2(or_514_nl, mux_684_nl, fsm_output[1]);
  assign or_515_nl = (fsm_output[3]) | mux_685_nl;
  assign mux_690_nl = MUX_s_1_2_2(nand_23_nl, or_515_nl, fsm_output[2]);
  assign nor_629_nl = ~((fsm_output[8]) | mux_690_nl);
  assign vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_711_nl,
      nor_629_nl, fsm_output[9]);
  assign or_598_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b0011) | (fsm_output[5]) | (fsm_output[1]);
  assign mux_738_nl = MUX_s_1_2_2(or_tmp_538, or_598_nl, fsm_output[0]);
  assign or_597_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0011) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_737_nl = MUX_s_1_2_2(or_597_nl, or_tmp_532, fsm_output[0]);
  assign mux_739_nl = MUX_s_1_2_2(mux_738_nl, mux_737_nl, fsm_output[4]);
  assign nand_28_nl = ~((fsm_output[6]) & (~ mux_739_nl));
  assign or_596_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0011);
  assign mux_740_nl = MUX_s_1_2_2(nand_28_nl, or_596_nl, fsm_output[7]);
  assign nor_609_nl = ~((fsm_output[8]) | mux_740_nl);
  assign and_439_nl = (COMP_LOOP_acc_20_psp_sva[2:0]==3'b001) & (fsm_output[7]) &
      (fsm_output[6]) & (fsm_output[4]) & (fsm_output[0]) & (VEC_LOOP_j_sva_9_0[0])
      & (~ (fsm_output[5])) & (fsm_output[1]);
  assign or_592_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0011) | (fsm_output[5]) |
      (~ (fsm_output[1]));
  assign mux_735_nl = MUX_s_1_2_2(or_592_nl, or_tmp_538, fsm_output[0]);
  assign nor_611_nl = ~((fsm_output[7]) | (fsm_output[6]) | (fsm_output[4]) | mux_735_nl);
  assign mux_736_nl = MUX_s_1_2_2(and_439_nl, nor_611_nl, fsm_output[8]);
  assign mux_741_nl = MUX_s_1_2_2(nor_609_nl, mux_736_nl, fsm_output[9]);
  assign or_589_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_9_0[0])) |
      (fsm_output[5]) | (~ (fsm_output[1]));
  assign or_587_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0011) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_730_nl = MUX_s_1_2_2(or_587_nl, or_tmp_538, fsm_output[0]);
  assign or_585_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b011)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_729_nl = MUX_s_1_2_2(or_tmp_537, or_585_nl, fsm_output[0]);
  assign mux_731_nl = MUX_s_1_2_2(mux_730_nl, mux_729_nl, fsm_output[4]);
  assign or_583_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0011) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_728_nl = MUX_s_1_2_2(or_583_nl, or_tmp_532, fsm_output[0]);
  assign or_584_nl = (fsm_output[4]) | mux_728_nl;
  assign mux_732_nl = MUX_s_1_2_2(mux_731_nl, or_584_nl, fsm_output[6]);
  assign mux_733_nl = MUX_s_1_2_2(or_589_nl, mux_732_nl, fsm_output[7]);
  assign and_335_nl = (fsm_output[8]) & (~ mux_733_nl);
  assign nor_612_nl = ~((fsm_output[8]) | (fsm_output[7]) | (fsm_output[6]) | (~
      (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0011));
  assign mux_734_nl = MUX_s_1_2_2(and_335_nl, nor_612_nl, fsm_output[9]);
  assign mux_742_nl = MUX_s_1_2_2(mux_741_nl, mux_734_nl, fsm_output[3]);
  assign or_580_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b001) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_9_0[0])) | (fsm_output[5]) | (~
      (fsm_output[1]));
  assign or_578_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0011) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_723_nl = MUX_s_1_2_2(or_578_nl, or_tmp_538, fsm_output[0]);
  assign or_576_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_722_nl = MUX_s_1_2_2(or_tmp_537, or_576_nl, fsm_output[0]);
  assign mux_724_nl = MUX_s_1_2_2(mux_723_nl, mux_722_nl, fsm_output[4]);
  assign mux_725_nl = MUX_s_1_2_2(or_580_nl, mux_724_nl, fsm_output[6]);
  assign or_574_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0011) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_720_nl = MUX_s_1_2_2(or_574_nl, or_tmp_532, fsm_output[0]);
  assign or_575_nl = (fsm_output[4]) | mux_720_nl;
  assign mux_721_nl = MUX_s_1_2_2(or_575_nl, or_tmp_531, fsm_output[6]);
  assign mux_726_nl = MUX_s_1_2_2(mux_725_nl, mux_721_nl, fsm_output[7]);
  assign nor_613_nl = ~((fsm_output[9:8]!=2'b10) | mux_726_nl);
  assign or_571_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001)
      | (~ (VEC_LOOP_j_sva_9_0[0])) | (fsm_output[5]) | (~ (fsm_output[1]));
  assign or_569_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0011) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_716_nl = MUX_s_1_2_2(or_569_nl, or_tmp_538, fsm_output[0]);
  assign or_565_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_715_nl = MUX_s_1_2_2(or_tmp_537, or_565_nl, fsm_output[0]);
  assign mux_717_nl = MUX_s_1_2_2(mux_716_nl, mux_715_nl, fsm_output[4]);
  assign mux_718_nl = MUX_s_1_2_2(or_571_nl, mux_717_nl, fsm_output[6]);
  assign nand_26_nl = ~((fsm_output[7]) & (~ mux_718_nl));
  assign or_562_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0011) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_713_nl = MUX_s_1_2_2(or_562_nl, or_tmp_532, fsm_output[0]);
  assign or_563_nl = (fsm_output[4]) | mux_713_nl;
  assign mux_714_nl = MUX_s_1_2_2(or_563_nl, or_tmp_531, fsm_output[6]);
  assign or_564_nl = (fsm_output[7]) | mux_714_nl;
  assign mux_719_nl = MUX_s_1_2_2(nand_26_nl, or_564_nl, fsm_output[8]);
  assign nor_614_nl = ~((fsm_output[9]) | mux_719_nl);
  assign mux_727_nl = MUX_s_1_2_2(nor_613_nl, nor_614_nl, fsm_output[3]);
  assign vec_rsc_0_3_i_we_d_pff = MUX_s_1_2_2(mux_742_nl, mux_727_nl, fsm_output[2]);
  assign nor_598_cse = ~((z_out_6_10_1[3:0]!=4'b0011) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign or_648_cse = (z_out_6_10_1[3:0]!=4'b0011) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_651_nl = (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0011) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_650_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | not_tmp_134;
  assign mux_769_nl = MUX_s_1_2_2(or_650_nl, or_648_cse, fsm_output[0]);
  assign mux_770_nl = MUX_s_1_2_2(or_651_nl, mux_769_nl, fsm_output[6]);
  assign or_647_nl = (z_out_6_10_1[3:1]!=3'b001) | nand_308_cse;
  assign or_645_nl = (z_out_6_10_1[3:0]!=4'b0011) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_767_nl = MUX_s_1_2_2(or_647_nl, or_645_nl, fsm_output[0]);
  assign or_644_nl = (~ (VEC_LOOP_j_sva_9_0[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_642_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0011) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_766_nl = MUX_s_1_2_2(or_644_nl, or_642_nl, fsm_output[0]);
  assign mux_768_nl = MUX_s_1_2_2(mux_767_nl, mux_766_nl, fsm_output[6]);
  assign mux_771_nl = MUX_s_1_2_2(mux_770_nl, mux_768_nl, fsm_output[1]);
  assign nor_589_nl = ~((fsm_output[3]) | mux_771_nl);
  assign or_640_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b0011) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_638_nl = (z_out_6_10_1[3:0]!=4'b0011) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]);
  assign mux_763_nl = MUX_s_1_2_2(or_640_nl, or_638_nl, fsm_output[0]);
  assign or_637_nl = (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b0011) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_764_nl = MUX_s_1_2_2(mux_763_nl, or_637_nl, fsm_output[6]);
  assign nor_590_nl = ~((fsm_output[1]) | mux_764_nl);
  assign nor_591_nl = ~((~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b0011) & (fsm_output[1])
      & (fsm_output[6]) & (fsm_output[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      | not_tmp_133);
  assign mux_765_nl = MUX_s_1_2_2(nor_590_nl, nor_591_nl, fsm_output[3]);
  assign mux_772_nl = MUX_s_1_2_2(nor_589_nl, mux_765_nl, fsm_output[2]);
  assign nor_592_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b0011)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign nor_593_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0011) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | not_tmp_133);
  assign nor_594_nl = ~((~ (VEC_LOOP_j_sva_9_0[0])) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b001)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_595_nl = ~((z_out_6_10_1[3:0]!=4'b0011) | not_tmp_133);
  assign mux_759_nl = MUX_s_1_2_2(nor_594_nl, nor_595_nl, fsm_output[0]);
  assign mux_760_nl = MUX_s_1_2_2(nor_593_nl, mux_759_nl, fsm_output[6]);
  assign and_333_nl = (fsm_output[1]) & mux_760_nl;
  assign mux_761_nl = MUX_s_1_2_2(nor_592_nl, and_333_nl, fsm_output[3]);
  assign nor_596_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b011)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_597_nl = ~((z_out_6_10_1[3:0]!=4'b0011) | (fsm_output[5]) | not_tmp_134);
  assign mux_756_nl = MUX_s_1_2_2(nor_596_nl, nor_597_nl, fsm_output[0]);
  assign nor_599_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_755_nl = MUX_s_1_2_2(nor_598_cse, nor_599_nl, fsm_output[0]);
  assign mux_757_nl = MUX_s_1_2_2(mux_756_nl, mux_755_nl, fsm_output[6]);
  assign nor_600_nl = ~((~ (VEC_LOOP_j_sva_9_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_601_nl = ~((z_out_6_10_1[3:0]!=4'b0011) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_753_nl = MUX_s_1_2_2(nor_600_nl, nor_601_nl, fsm_output[0]);
  assign nor_602_nl = ~((z_out_6_10_1[3:0]!=4'b0011) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[4]));
  assign mux_754_nl = MUX_s_1_2_2(mux_753_nl, nor_602_nl, fsm_output[6]);
  assign mux_758_nl = MUX_s_1_2_2(mux_757_nl, mux_754_nl, fsm_output[1]);
  assign and_334_nl = (fsm_output[3]) & mux_758_nl;
  assign mux_762_nl = MUX_s_1_2_2(mux_761_nl, and_334_nl, fsm_output[2]);
  assign mux_773_nl = MUX_s_1_2_2(mux_772_nl, mux_762_nl, fsm_output[8]);
  assign nor_605_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_749_nl = MUX_s_1_2_2(nor_598_cse, nor_605_nl, fsm_output[0]);
  assign nor_606_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_607_nl = ~((z_out_6_10_1[3:0]!=4'b0011) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_748_nl = MUX_s_1_2_2(nor_606_nl, nor_607_nl, fsm_output[0]);
  assign mux_750_nl = MUX_s_1_2_2(mux_749_nl, mux_748_nl, fsm_output[6]);
  assign nor_608_nl = ~((z_out_6_10_1[3:0]!=4'b0011) | (fsm_output[6]) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_751_nl = MUX_s_1_2_2(mux_750_nl, nor_608_nl, fsm_output[1]);
  assign nand_29_nl = ~((fsm_output[3]) & mux_751_nl);
  assign or_607_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0011) | (~ (fsm_output[6]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[5])
      | not_tmp_134;
  assign or_605_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001) | (~ (VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_604_nl = (z_out_6_10_1[3:0]!=4'b0011) | not_tmp_133;
  assign mux_745_nl = MUX_s_1_2_2(or_605_nl, or_604_nl, fsm_output[0]);
  assign or_601_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0011) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_744_nl = MUX_s_1_2_2(or_648_cse, or_601_nl, fsm_output[0]);
  assign mux_746_nl = MUX_s_1_2_2(mux_745_nl, mux_744_nl, fsm_output[6]);
  assign mux_747_nl = MUX_s_1_2_2(or_607_nl, mux_746_nl, fsm_output[1]);
  assign or_608_nl = (fsm_output[3]) | mux_747_nl;
  assign mux_752_nl = MUX_s_1_2_2(nand_29_nl, or_608_nl, fsm_output[2]);
  assign nor_603_nl = ~((fsm_output[8]) | mux_752_nl);
  assign vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_773_nl,
      nor_603_nl, fsm_output[9]);
  assign or_691_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b0100) | (fsm_output[5]) | (fsm_output[1]);
  assign mux_800_nl = MUX_s_1_2_2(or_tmp_631, or_691_nl, fsm_output[0]);
  assign or_690_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0100) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_799_nl = MUX_s_1_2_2(or_690_nl, or_tmp_625, fsm_output[0]);
  assign mux_801_nl = MUX_s_1_2_2(mux_800_nl, mux_799_nl, fsm_output[4]);
  assign nand_34_nl = ~((fsm_output[6]) & (~ mux_801_nl));
  assign or_689_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0100);
  assign mux_802_nl = MUX_s_1_2_2(nand_34_nl, or_689_nl, fsm_output[7]);
  assign nor_583_nl = ~((fsm_output[8]) | mux_802_nl);
  assign nor_584_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010) | (~ (fsm_output[7]))
      | (~ (fsm_output[6])) | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[5]) | (~ (fsm_output[1])));
  assign or_685_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0100) | (fsm_output[5]) |
      (~ (fsm_output[1]));
  assign mux_797_nl = MUX_s_1_2_2(or_685_nl, or_tmp_631, fsm_output[0]);
  assign nor_585_nl = ~((fsm_output[7]) | (fsm_output[6]) | (fsm_output[4]) | mux_797_nl);
  assign mux_798_nl = MUX_s_1_2_2(nor_584_nl, nor_585_nl, fsm_output[8]);
  assign mux_803_nl = MUX_s_1_2_2(nor_583_nl, mux_798_nl, fsm_output[9]);
  assign or_682_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign or_680_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0100) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_792_nl = MUX_s_1_2_2(or_680_nl, or_tmp_631, fsm_output[0]);
  assign or_678_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b100)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_791_nl = MUX_s_1_2_2(or_tmp_630, or_678_nl, fsm_output[0]);
  assign mux_793_nl = MUX_s_1_2_2(mux_792_nl, mux_791_nl, fsm_output[4]);
  assign or_676_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0100) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_790_nl = MUX_s_1_2_2(or_676_nl, or_tmp_625, fsm_output[0]);
  assign or_677_nl = (fsm_output[4]) | mux_790_nl;
  assign mux_794_nl = MUX_s_1_2_2(mux_793_nl, or_677_nl, fsm_output[6]);
  assign mux_795_nl = MUX_s_1_2_2(or_682_nl, mux_794_nl, fsm_output[7]);
  assign and_332_nl = (fsm_output[8]) & (~ mux_795_nl);
  assign nor_586_nl = ~((fsm_output[8]) | (fsm_output[7]) | (fsm_output[6]) | (~
      (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0100));
  assign mux_796_nl = MUX_s_1_2_2(and_332_nl, nor_586_nl, fsm_output[9]);
  assign mux_804_nl = MUX_s_1_2_2(mux_803_nl, mux_796_nl, fsm_output[3]);
  assign or_673_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b010) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5]) | (~ (fsm_output[1]));
  assign or_671_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0100) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_785_nl = MUX_s_1_2_2(or_671_nl, or_tmp_631, fsm_output[0]);
  assign or_669_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_784_nl = MUX_s_1_2_2(or_tmp_630, or_669_nl, fsm_output[0]);
  assign mux_786_nl = MUX_s_1_2_2(mux_785_nl, mux_784_nl, fsm_output[4]);
  assign mux_787_nl = MUX_s_1_2_2(or_673_nl, mux_786_nl, fsm_output[6]);
  assign or_667_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0100) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_782_nl = MUX_s_1_2_2(or_667_nl, or_tmp_625, fsm_output[0]);
  assign or_668_nl = (fsm_output[4]) | mux_782_nl;
  assign mux_783_nl = MUX_s_1_2_2(or_668_nl, or_tmp_624, fsm_output[6]);
  assign mux_788_nl = MUX_s_1_2_2(mux_787_nl, mux_783_nl, fsm_output[7]);
  assign nor_587_nl = ~((fsm_output[9:8]!=2'b10) | mux_788_nl);
  assign or_664_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010)
      | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5]) | (~ (fsm_output[1]));
  assign or_662_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0100) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_778_nl = MUX_s_1_2_2(or_662_nl, or_tmp_631, fsm_output[0]);
  assign or_658_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_777_nl = MUX_s_1_2_2(or_tmp_630, or_658_nl, fsm_output[0]);
  assign mux_779_nl = MUX_s_1_2_2(mux_778_nl, mux_777_nl, fsm_output[4]);
  assign mux_780_nl = MUX_s_1_2_2(or_664_nl, mux_779_nl, fsm_output[6]);
  assign nand_32_nl = ~((fsm_output[7]) & (~ mux_780_nl));
  assign or_655_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0100) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_775_nl = MUX_s_1_2_2(or_655_nl, or_tmp_625, fsm_output[0]);
  assign or_656_nl = (fsm_output[4]) | mux_775_nl;
  assign mux_776_nl = MUX_s_1_2_2(or_656_nl, or_tmp_624, fsm_output[6]);
  assign or_657_nl = (fsm_output[7]) | mux_776_nl;
  assign mux_781_nl = MUX_s_1_2_2(nand_32_nl, or_657_nl, fsm_output[8]);
  assign nor_588_nl = ~((fsm_output[9]) | mux_781_nl);
  assign mux_789_nl = MUX_s_1_2_2(nor_587_nl, nor_588_nl, fsm_output[3]);
  assign vec_rsc_0_4_i_we_d_pff = MUX_s_1_2_2(mux_804_nl, mux_789_nl, fsm_output[2]);
  assign nor_572_cse = ~((z_out_6_10_1[3:0]!=4'b0100) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign or_740_cse = (z_out_6_10_1[3:0]!=4'b0100) | not_tmp_133;
  assign or_741_cse = (z_out_6_10_1[3:0]!=4'b0100) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_744_nl = (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0100) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_743_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | not_tmp_134;
  assign mux_831_nl = MUX_s_1_2_2(or_743_nl, or_741_cse, fsm_output[0]);
  assign mux_832_nl = MUX_s_1_2_2(or_744_nl, mux_831_nl, fsm_output[6]);
  assign or_738_nl = (z_out_6_10_1[3:0]!=4'b0100) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_829_nl = MUX_s_1_2_2(or_740_cse, or_738_nl, fsm_output[0]);
  assign or_737_nl = (VEC_LOOP_j_sva_9_0[0]) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_735_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0100) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_828_nl = MUX_s_1_2_2(or_737_nl, or_735_nl, fsm_output[0]);
  assign mux_830_nl = MUX_s_1_2_2(mux_829_nl, mux_828_nl, fsm_output[6]);
  assign mux_833_nl = MUX_s_1_2_2(mux_832_nl, mux_830_nl, fsm_output[1]);
  assign nor_563_nl = ~((fsm_output[3]) | mux_833_nl);
  assign or_733_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b0100) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_731_nl = (z_out_6_10_1[3:0]!=4'b0100) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]);
  assign mux_825_nl = MUX_s_1_2_2(or_733_nl, or_731_nl, fsm_output[0]);
  assign or_730_nl = (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b0100) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_826_nl = MUX_s_1_2_2(mux_825_nl, or_730_nl, fsm_output[6]);
  assign nor_564_nl = ~((fsm_output[1]) | mux_826_nl);
  assign nor_565_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0100) | (~ (fsm_output[1]))
      | (~ (fsm_output[6])) | (~ (fsm_output[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | not_tmp_133);
  assign mux_827_nl = MUX_s_1_2_2(nor_564_nl, nor_565_nl, fsm_output[3]);
  assign mux_834_nl = MUX_s_1_2_2(nor_563_nl, mux_827_nl, fsm_output[2]);
  assign nor_566_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b0100)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign nor_567_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0100) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | not_tmp_133);
  assign nor_568_nl = ~((VEC_LOOP_j_sva_9_0[0]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b010)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_569_nl = ~((z_out_6_10_1[3:0]!=4'b0100) | not_tmp_133);
  assign mux_821_nl = MUX_s_1_2_2(nor_568_nl, nor_569_nl, fsm_output[0]);
  assign mux_822_nl = MUX_s_1_2_2(nor_567_nl, mux_821_nl, fsm_output[6]);
  assign and_330_nl = (fsm_output[1]) & mux_822_nl;
  assign mux_823_nl = MUX_s_1_2_2(nor_566_nl, and_330_nl, fsm_output[3]);
  assign nor_570_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b100)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_571_nl = ~((z_out_6_10_1[3:0]!=4'b0100) | (fsm_output[5]) | not_tmp_134);
  assign mux_818_nl = MUX_s_1_2_2(nor_570_nl, nor_571_nl, fsm_output[0]);
  assign nor_573_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_817_nl = MUX_s_1_2_2(nor_572_cse, nor_573_nl, fsm_output[0]);
  assign mux_819_nl = MUX_s_1_2_2(mux_818_nl, mux_817_nl, fsm_output[6]);
  assign nor_574_nl = ~((VEC_LOOP_j_sva_9_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_575_nl = ~((z_out_6_10_1[3:0]!=4'b0100) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_815_nl = MUX_s_1_2_2(nor_574_nl, nor_575_nl, fsm_output[0]);
  assign nor_576_nl = ~((z_out_6_10_1[3:0]!=4'b0100) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[4]));
  assign mux_816_nl = MUX_s_1_2_2(mux_815_nl, nor_576_nl, fsm_output[6]);
  assign mux_820_nl = MUX_s_1_2_2(mux_819_nl, mux_816_nl, fsm_output[1]);
  assign and_331_nl = (fsm_output[3]) & mux_820_nl;
  assign mux_824_nl = MUX_s_1_2_2(mux_823_nl, and_331_nl, fsm_output[2]);
  assign mux_835_nl = MUX_s_1_2_2(mux_834_nl, mux_824_nl, fsm_output[8]);
  assign nor_579_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_811_nl = MUX_s_1_2_2(nor_572_cse, nor_579_nl, fsm_output[0]);
  assign nor_580_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_581_nl = ~((z_out_6_10_1[3:0]!=4'b0100) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_810_nl = MUX_s_1_2_2(nor_580_nl, nor_581_nl, fsm_output[0]);
  assign mux_812_nl = MUX_s_1_2_2(mux_811_nl, mux_810_nl, fsm_output[6]);
  assign nor_582_nl = ~((z_out_6_10_1[3:0]!=4'b0100) | (fsm_output[6]) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_813_nl = MUX_s_1_2_2(mux_812_nl, nor_582_nl, fsm_output[1]);
  assign nand_35_nl = ~((fsm_output[3]) & mux_813_nl);
  assign or_700_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0100) | (~ (fsm_output[6]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[5])
      | not_tmp_134;
  assign or_698_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_807_nl = MUX_s_1_2_2(or_698_nl, or_740_cse, fsm_output[0]);
  assign or_694_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0100) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_806_nl = MUX_s_1_2_2(or_741_cse, or_694_nl, fsm_output[0]);
  assign mux_808_nl = MUX_s_1_2_2(mux_807_nl, mux_806_nl, fsm_output[6]);
  assign mux_809_nl = MUX_s_1_2_2(or_700_nl, mux_808_nl, fsm_output[1]);
  assign or_701_nl = (fsm_output[3]) | mux_809_nl;
  assign mux_814_nl = MUX_s_1_2_2(nand_35_nl, or_701_nl, fsm_output[2]);
  assign nor_577_nl = ~((fsm_output[8]) | mux_814_nl);
  assign vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_835_nl,
      nor_577_nl, fsm_output[9]);
  assign or_785_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b0101) | (fsm_output[1]) | (fsm_output[5]);
  assign mux_862_nl = MUX_s_1_2_2(or_tmp_725, or_785_nl, fsm_output[0]);
  assign or_784_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0101) | (fsm_output[1])
      | (~ (fsm_output[5]));
  assign mux_861_nl = MUX_s_1_2_2(or_784_nl, or_tmp_718, fsm_output[0]);
  assign mux_863_nl = MUX_s_1_2_2(mux_862_nl, mux_861_nl, fsm_output[4]);
  assign nor_555_nl = ~((fsm_output[9]) | (~ (fsm_output[6])) | mux_863_nl);
  assign or_782_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b010) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_9_0[0])) | (~ (fsm_output[1])) |
      (fsm_output[5]);
  assign or_781_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0101) | (~ (fsm_output[1]))
      | (fsm_output[5]);
  assign mux_858_nl = MUX_s_1_2_2(or_781_nl, or_tmp_725, fsm_output[0]);
  assign or_780_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (fsm_output[1]) | (~ (fsm_output[5]));
  assign mux_857_nl = MUX_s_1_2_2(or_tmp_724, or_780_nl, fsm_output[0]);
  assign mux_859_nl = MUX_s_1_2_2(mux_858_nl, mux_857_nl, fsm_output[4]);
  assign mux_860_nl = MUX_s_1_2_2(or_782_nl, mux_859_nl, fsm_output[6]);
  assign and_329_nl = (fsm_output[9]) & (~ mux_860_nl);
  assign mux_864_nl = MUX_s_1_2_2(nor_555_nl, and_329_nl, fsm_output[2]);
  assign or_777_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0101) | (~ (fsm_output[1]))
      | (fsm_output[5]);
  assign mux_856_nl = MUX_s_1_2_2(or_777_nl, or_tmp_725, fsm_output[0]);
  assign nor_556_nl = ~((fsm_output[2]) | (~ (fsm_output[9])) | (fsm_output[6]) |
      (fsm_output[4]) | mux_856_nl);
  assign mux_865_nl = MUX_s_1_2_2(mux_864_nl, nor_556_nl, fsm_output[8]);
  assign or_774_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (fsm_output[1])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0101);
  assign or_773_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_9_0[0])) |
      (~ (fsm_output[1])) | (fsm_output[5]);
  assign mux_854_nl = MUX_s_1_2_2(or_774_nl, or_773_nl, fsm_output[9]);
  assign or_771_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0101) | (fsm_output[1])
      | (~ (fsm_output[5]));
  assign mux_852_nl = MUX_s_1_2_2(or_771_nl, or_tmp_718, fsm_output[0]);
  assign or_772_nl = (fsm_output[4]) | mux_852_nl;
  assign mux_853_nl = MUX_s_1_2_2(or_772_nl, or_tmp_734, fsm_output[6]);
  assign nand_38_nl = ~((fsm_output[9]) & (~ mux_853_nl));
  assign mux_855_nl = MUX_s_1_2_2(mux_854_nl, nand_38_nl, fsm_output[2]);
  assign nor_557_nl = ~((fsm_output[8]) | mux_855_nl);
  assign mux_866_nl = MUX_s_1_2_2(mux_865_nl, nor_557_nl, fsm_output[7]);
  assign nor_558_nl = ~((fsm_output[2]) | (~ (fsm_output[9])) | (fsm_output[6]) |
      (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[5]) |
      (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0101));
  assign nor_559_nl = ~((fsm_output[9]) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010)
      | (~ (fsm_output[6])) | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_9_0[0]))
      | (~ (fsm_output[1])) | (fsm_output[5]));
  assign or_765_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0101) | (fsm_output[1])
      | (~ (fsm_output[5]));
  assign mux_847_nl = MUX_s_1_2_2(or_765_nl, or_tmp_718, fsm_output[0]);
  assign or_766_nl = (fsm_output[4]) | mux_847_nl;
  assign mux_848_nl = MUX_s_1_2_2(or_766_nl, or_tmp_734, fsm_output[6]);
  assign nor_560_nl = ~((fsm_output[9]) | mux_848_nl);
  assign mux_849_nl = MUX_s_1_2_2(nor_559_nl, nor_560_nl, fsm_output[2]);
  assign mux_850_nl = MUX_s_1_2_2(nor_558_nl, mux_849_nl, fsm_output[8]);
  assign or_761_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010)
      | (~ (VEC_LOOP_j_sva_9_0[0])) | (~ (fsm_output[1])) | (fsm_output[5]);
  assign or_760_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0101) | (~ (fsm_output[1]))
      | (fsm_output[5]);
  assign mux_843_nl = MUX_s_1_2_2(or_760_nl, or_tmp_725, fsm_output[0]);
  assign or_759_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (fsm_output[1]) | (~ (fsm_output[5]));
  assign mux_842_nl = MUX_s_1_2_2(or_tmp_724, or_759_nl, fsm_output[0]);
  assign mux_844_nl = MUX_s_1_2_2(mux_843_nl, mux_842_nl, fsm_output[4]);
  assign mux_845_nl = MUX_s_1_2_2(or_761_nl, mux_844_nl, fsm_output[6]);
  assign nor_561_nl = ~((~ (fsm_output[2])) | (fsm_output[9]) | mux_845_nl);
  assign or_755_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0101) | (~ (fsm_output[1]))
      | (fsm_output[5]);
  assign mux_839_nl = MUX_s_1_2_2(or_755_nl, or_tmp_725, fsm_output[0]);
  assign or_752_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b101)
      | (fsm_output[1]) | (~ (fsm_output[5]));
  assign mux_838_nl = MUX_s_1_2_2(or_tmp_724, or_752_nl, fsm_output[0]);
  assign mux_840_nl = MUX_s_1_2_2(mux_839_nl, mux_838_nl, fsm_output[4]);
  assign or_749_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0101) | (fsm_output[1])
      | (~ (fsm_output[5]));
  assign mux_837_nl = MUX_s_1_2_2(or_749_nl, or_tmp_718, fsm_output[0]);
  assign or_750_nl = (fsm_output[4]) | mux_837_nl;
  assign mux_841_nl = MUX_s_1_2_2(mux_840_nl, or_750_nl, fsm_output[6]);
  assign nor_562_nl = ~((fsm_output[2]) | (fsm_output[9]) | mux_841_nl);
  assign mux_846_nl = MUX_s_1_2_2(nor_561_nl, nor_562_nl, fsm_output[8]);
  assign mux_851_nl = MUX_s_1_2_2(mux_850_nl, mux_846_nl, fsm_output[7]);
  assign vec_rsc_0_5_i_we_d_pff = MUX_s_1_2_2(mux_866_nl, mux_851_nl, fsm_output[3]);
  assign nor_544_cse = ~((z_out_6_10_1[3:0]!=4'b0101) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign or_834_cse = (z_out_6_10_1[3:0]!=4'b0101) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_837_nl = (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0101) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_836_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | not_tmp_134;
  assign mux_893_nl = MUX_s_1_2_2(or_836_nl, or_834_cse, fsm_output[0]);
  assign mux_894_nl = MUX_s_1_2_2(or_837_nl, mux_893_nl, fsm_output[6]);
  assign or_833_nl = (z_out_6_10_1[3:1]!=3'b010) | nand_308_cse;
  assign or_831_nl = (z_out_6_10_1[3:0]!=4'b0101) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_891_nl = MUX_s_1_2_2(or_833_nl, or_831_nl, fsm_output[0]);
  assign or_830_nl = (~ (VEC_LOOP_j_sva_9_0[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_828_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0101) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_890_nl = MUX_s_1_2_2(or_830_nl, or_828_nl, fsm_output[0]);
  assign mux_892_nl = MUX_s_1_2_2(mux_891_nl, mux_890_nl, fsm_output[6]);
  assign mux_895_nl = MUX_s_1_2_2(mux_894_nl, mux_892_nl, fsm_output[1]);
  assign nor_535_nl = ~((fsm_output[3]) | mux_895_nl);
  assign or_826_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b0101) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_824_nl = (z_out_6_10_1[3:0]!=4'b0101) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]);
  assign mux_887_nl = MUX_s_1_2_2(or_826_nl, or_824_nl, fsm_output[0]);
  assign or_823_nl = (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b0101) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_888_nl = MUX_s_1_2_2(mux_887_nl, or_823_nl, fsm_output[6]);
  assign nor_536_nl = ~((fsm_output[1]) | mux_888_nl);
  assign nor_537_nl = ~((~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b0101) & (fsm_output[1])
      & (fsm_output[6]) & (fsm_output[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      | not_tmp_133);
  assign mux_889_nl = MUX_s_1_2_2(nor_536_nl, nor_537_nl, fsm_output[3]);
  assign mux_896_nl = MUX_s_1_2_2(nor_535_nl, mux_889_nl, fsm_output[2]);
  assign nor_538_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b0101)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign nor_539_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0101) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | not_tmp_133);
  assign nor_540_nl = ~((~ (VEC_LOOP_j_sva_9_0[0])) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b010)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_541_nl = ~((z_out_6_10_1[3:0]!=4'b0101) | not_tmp_133);
  assign mux_883_nl = MUX_s_1_2_2(nor_540_nl, nor_541_nl, fsm_output[0]);
  assign mux_884_nl = MUX_s_1_2_2(nor_539_nl, mux_883_nl, fsm_output[6]);
  assign and_327_nl = (fsm_output[1]) & mux_884_nl;
  assign mux_885_nl = MUX_s_1_2_2(nor_538_nl, and_327_nl, fsm_output[3]);
  assign nor_542_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b101)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_543_nl = ~((z_out_6_10_1[3:0]!=4'b0101) | (fsm_output[5]) | not_tmp_134);
  assign mux_880_nl = MUX_s_1_2_2(nor_542_nl, nor_543_nl, fsm_output[0]);
  assign nor_545_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_879_nl = MUX_s_1_2_2(nor_544_cse, nor_545_nl, fsm_output[0]);
  assign mux_881_nl = MUX_s_1_2_2(mux_880_nl, mux_879_nl, fsm_output[6]);
  assign nor_546_nl = ~((~ (VEC_LOOP_j_sva_9_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_547_nl = ~((z_out_6_10_1[3:0]!=4'b0101) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_877_nl = MUX_s_1_2_2(nor_546_nl, nor_547_nl, fsm_output[0]);
  assign nor_548_nl = ~((z_out_6_10_1[3:0]!=4'b0101) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[4]));
  assign mux_878_nl = MUX_s_1_2_2(mux_877_nl, nor_548_nl, fsm_output[6]);
  assign mux_882_nl = MUX_s_1_2_2(mux_881_nl, mux_878_nl, fsm_output[1]);
  assign and_328_nl = (fsm_output[3]) & mux_882_nl;
  assign mux_886_nl = MUX_s_1_2_2(mux_885_nl, and_328_nl, fsm_output[2]);
  assign mux_897_nl = MUX_s_1_2_2(mux_896_nl, mux_886_nl, fsm_output[8]);
  assign nor_551_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_873_nl = MUX_s_1_2_2(nor_544_cse, nor_551_nl, fsm_output[0]);
  assign nor_552_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_553_nl = ~((z_out_6_10_1[3:0]!=4'b0101) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_872_nl = MUX_s_1_2_2(nor_552_nl, nor_553_nl, fsm_output[0]);
  assign mux_874_nl = MUX_s_1_2_2(mux_873_nl, mux_872_nl, fsm_output[6]);
  assign nor_554_nl = ~((z_out_6_10_1[3:0]!=4'b0101) | (fsm_output[6]) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_875_nl = MUX_s_1_2_2(mux_874_nl, nor_554_nl, fsm_output[1]);
  assign nand_41_nl = ~((fsm_output[3]) & mux_875_nl);
  assign or_793_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0101) | (~ (fsm_output[6]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[5])
      | not_tmp_134;
  assign or_791_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010) | (~ (VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_790_nl = (z_out_6_10_1[3:0]!=4'b0101) | not_tmp_133;
  assign mux_869_nl = MUX_s_1_2_2(or_791_nl, or_790_nl, fsm_output[0]);
  assign or_787_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0101) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_868_nl = MUX_s_1_2_2(or_834_cse, or_787_nl, fsm_output[0]);
  assign mux_870_nl = MUX_s_1_2_2(mux_869_nl, mux_868_nl, fsm_output[6]);
  assign mux_871_nl = MUX_s_1_2_2(or_793_nl, mux_870_nl, fsm_output[1]);
  assign or_794_nl = (fsm_output[3]) | mux_871_nl;
  assign mux_876_nl = MUX_s_1_2_2(nand_41_nl, or_794_nl, fsm_output[2]);
  assign nor_549_nl = ~((fsm_output[8]) | mux_876_nl);
  assign vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_897_nl,
      nor_549_nl, fsm_output[9]);
  assign or_877_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b0110) | (fsm_output[5]) | (fsm_output[1]);
  assign mux_924_nl = MUX_s_1_2_2(or_tmp_817, or_877_nl, fsm_output[0]);
  assign or_876_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0110) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_923_nl = MUX_s_1_2_2(or_876_nl, or_tmp_811, fsm_output[0]);
  assign mux_925_nl = MUX_s_1_2_2(mux_924_nl, mux_923_nl, fsm_output[4]);
  assign nand_46_nl = ~((fsm_output[6]) & (~ mux_925_nl));
  assign or_875_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0110);
  assign mux_926_nl = MUX_s_1_2_2(nand_46_nl, or_875_nl, fsm_output[7]);
  assign nor_529_nl = ~((fsm_output[8]) | mux_926_nl);
  assign and_438_nl = (COMP_LOOP_acc_20_psp_sva[2:0]==3'b011) & (fsm_output[7]) &
      (fsm_output[6]) & (fsm_output[4]) & (fsm_output[0]) & (~ (VEC_LOOP_j_sva_9_0[0]))
      & (~ (fsm_output[5])) & (fsm_output[1]);
  assign or_871_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0110) | (fsm_output[5]) |
      (~ (fsm_output[1]));
  assign mux_921_nl = MUX_s_1_2_2(or_871_nl, or_tmp_817, fsm_output[0]);
  assign nor_531_nl = ~((fsm_output[7]) | (fsm_output[6]) | (fsm_output[4]) | mux_921_nl);
  assign mux_922_nl = MUX_s_1_2_2(and_438_nl, nor_531_nl, fsm_output[8]);
  assign mux_927_nl = MUX_s_1_2_2(nor_529_nl, mux_922_nl, fsm_output[9]);
  assign or_868_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b011) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign or_866_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0110) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_916_nl = MUX_s_1_2_2(or_866_nl, or_tmp_817, fsm_output[0]);
  assign or_864_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b110)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_915_nl = MUX_s_1_2_2(or_tmp_816, or_864_nl, fsm_output[0]);
  assign mux_917_nl = MUX_s_1_2_2(mux_916_nl, mux_915_nl, fsm_output[4]);
  assign or_862_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0110) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_914_nl = MUX_s_1_2_2(or_862_nl, or_tmp_811, fsm_output[0]);
  assign or_863_nl = (fsm_output[4]) | mux_914_nl;
  assign mux_918_nl = MUX_s_1_2_2(mux_917_nl, or_863_nl, fsm_output[6]);
  assign mux_919_nl = MUX_s_1_2_2(or_868_nl, mux_918_nl, fsm_output[7]);
  assign and_326_nl = (fsm_output[8]) & (~ mux_919_nl);
  assign nor_532_nl = ~((fsm_output[8]) | (fsm_output[7]) | (fsm_output[6]) | (~
      (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0110));
  assign mux_920_nl = MUX_s_1_2_2(and_326_nl, nor_532_nl, fsm_output[9]);
  assign mux_928_nl = MUX_s_1_2_2(mux_927_nl, mux_920_nl, fsm_output[3]);
  assign or_859_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b011) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5]) | (~ (fsm_output[1]));
  assign or_857_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0110) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_909_nl = MUX_s_1_2_2(or_857_nl, or_tmp_817, fsm_output[0]);
  assign or_855_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_908_nl = MUX_s_1_2_2(or_tmp_816, or_855_nl, fsm_output[0]);
  assign mux_910_nl = MUX_s_1_2_2(mux_909_nl, mux_908_nl, fsm_output[4]);
  assign mux_911_nl = MUX_s_1_2_2(or_859_nl, mux_910_nl, fsm_output[6]);
  assign or_853_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0110) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_906_nl = MUX_s_1_2_2(or_853_nl, or_tmp_811, fsm_output[0]);
  assign or_854_nl = (fsm_output[4]) | mux_906_nl;
  assign mux_907_nl = MUX_s_1_2_2(or_854_nl, or_tmp_810, fsm_output[6]);
  assign mux_912_nl = MUX_s_1_2_2(mux_911_nl, mux_907_nl, fsm_output[7]);
  assign nor_533_nl = ~((fsm_output[9:8]!=2'b10) | mux_912_nl);
  assign or_850_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b011)
      | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5]) | (~ (fsm_output[1]));
  assign or_848_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0110) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_902_nl = MUX_s_1_2_2(or_848_nl, or_tmp_817, fsm_output[0]);
  assign or_844_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_901_nl = MUX_s_1_2_2(or_tmp_816, or_844_nl, fsm_output[0]);
  assign mux_903_nl = MUX_s_1_2_2(mux_902_nl, mux_901_nl, fsm_output[4]);
  assign mux_904_nl = MUX_s_1_2_2(or_850_nl, mux_903_nl, fsm_output[6]);
  assign nand_44_nl = ~((fsm_output[7]) & (~ mux_904_nl));
  assign or_841_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0110) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_899_nl = MUX_s_1_2_2(or_841_nl, or_tmp_811, fsm_output[0]);
  assign or_842_nl = (fsm_output[4]) | mux_899_nl;
  assign mux_900_nl = MUX_s_1_2_2(or_842_nl, or_tmp_810, fsm_output[6]);
  assign or_843_nl = (fsm_output[7]) | mux_900_nl;
  assign mux_905_nl = MUX_s_1_2_2(nand_44_nl, or_843_nl, fsm_output[8]);
  assign nor_534_nl = ~((fsm_output[9]) | mux_905_nl);
  assign mux_913_nl = MUX_s_1_2_2(nor_533_nl, nor_534_nl, fsm_output[3]);
  assign vec_rsc_0_6_i_we_d_pff = MUX_s_1_2_2(mux_928_nl, mux_913_nl, fsm_output[2]);
  assign nor_518_cse = ~((z_out_6_10_1[3:0]!=4'b0110) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign or_926_cse = (z_out_6_10_1[3:0]!=4'b0110) | not_tmp_133;
  assign or_927_cse = (z_out_6_10_1[3:0]!=4'b0110) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_930_nl = (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0110) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_929_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | not_tmp_134;
  assign mux_955_nl = MUX_s_1_2_2(or_929_nl, or_927_cse, fsm_output[0]);
  assign mux_956_nl = MUX_s_1_2_2(or_930_nl, mux_955_nl, fsm_output[6]);
  assign or_924_nl = (z_out_6_10_1[3:0]!=4'b0110) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_953_nl = MUX_s_1_2_2(or_926_cse, or_924_nl, fsm_output[0]);
  assign or_923_nl = (VEC_LOOP_j_sva_9_0[0]) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b011)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_921_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0110) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_952_nl = MUX_s_1_2_2(or_923_nl, or_921_nl, fsm_output[0]);
  assign mux_954_nl = MUX_s_1_2_2(mux_953_nl, mux_952_nl, fsm_output[6]);
  assign mux_957_nl = MUX_s_1_2_2(mux_956_nl, mux_954_nl, fsm_output[1]);
  assign nor_509_nl = ~((fsm_output[3]) | mux_957_nl);
  assign or_919_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b0110) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_917_nl = (z_out_6_10_1[3:0]!=4'b0110) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]);
  assign mux_949_nl = MUX_s_1_2_2(or_919_nl, or_917_nl, fsm_output[0]);
  assign or_916_nl = (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b0110) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_950_nl = MUX_s_1_2_2(mux_949_nl, or_916_nl, fsm_output[6]);
  assign nor_510_nl = ~((fsm_output[1]) | mux_950_nl);
  assign nor_511_nl = ~((~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b0110) & (fsm_output[1])
      & (fsm_output[6]) & (fsm_output[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      | not_tmp_133);
  assign mux_951_nl = MUX_s_1_2_2(nor_510_nl, nor_511_nl, fsm_output[3]);
  assign mux_958_nl = MUX_s_1_2_2(nor_509_nl, mux_951_nl, fsm_output[2]);
  assign nor_512_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b0110)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign nor_513_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0110) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | not_tmp_133);
  assign nor_514_nl = ~((VEC_LOOP_j_sva_9_0[0]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b011)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_515_nl = ~((z_out_6_10_1[3:0]!=4'b0110) | not_tmp_133);
  assign mux_945_nl = MUX_s_1_2_2(nor_514_nl, nor_515_nl, fsm_output[0]);
  assign mux_946_nl = MUX_s_1_2_2(nor_513_nl, mux_945_nl, fsm_output[6]);
  assign and_324_nl = (fsm_output[1]) & mux_946_nl;
  assign mux_947_nl = MUX_s_1_2_2(nor_512_nl, and_324_nl, fsm_output[3]);
  assign nor_516_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b110)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_517_nl = ~((z_out_6_10_1[3:0]!=4'b0110) | (fsm_output[5]) | not_tmp_134);
  assign mux_942_nl = MUX_s_1_2_2(nor_516_nl, nor_517_nl, fsm_output[0]);
  assign nor_519_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_941_nl = MUX_s_1_2_2(nor_518_cse, nor_519_nl, fsm_output[0]);
  assign mux_943_nl = MUX_s_1_2_2(mux_942_nl, mux_941_nl, fsm_output[6]);
  assign nor_520_nl = ~((VEC_LOOP_j_sva_9_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b011) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_521_nl = ~((z_out_6_10_1[3:0]!=4'b0110) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_939_nl = MUX_s_1_2_2(nor_520_nl, nor_521_nl, fsm_output[0]);
  assign nor_522_nl = ~((z_out_6_10_1[3:0]!=4'b0110) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[4]));
  assign mux_940_nl = MUX_s_1_2_2(mux_939_nl, nor_522_nl, fsm_output[6]);
  assign mux_944_nl = MUX_s_1_2_2(mux_943_nl, mux_940_nl, fsm_output[1]);
  assign and_325_nl = (fsm_output[3]) & mux_944_nl;
  assign mux_948_nl = MUX_s_1_2_2(mux_947_nl, and_325_nl, fsm_output[2]);
  assign mux_959_nl = MUX_s_1_2_2(mux_958_nl, mux_948_nl, fsm_output[8]);
  assign nor_525_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_935_nl = MUX_s_1_2_2(nor_518_cse, nor_525_nl, fsm_output[0]);
  assign nor_526_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_527_nl = ~((z_out_6_10_1[3:0]!=4'b0110) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_934_nl = MUX_s_1_2_2(nor_526_nl, nor_527_nl, fsm_output[0]);
  assign mux_936_nl = MUX_s_1_2_2(mux_935_nl, mux_934_nl, fsm_output[6]);
  assign nor_528_nl = ~((z_out_6_10_1[3:0]!=4'b0110) | (fsm_output[6]) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_937_nl = MUX_s_1_2_2(mux_936_nl, nor_528_nl, fsm_output[1]);
  assign nand_47_nl = ~((fsm_output[3]) & mux_937_nl);
  assign or_886_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0110) | (~ (fsm_output[6]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[5])
      | not_tmp_134;
  assign or_884_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_931_nl = MUX_s_1_2_2(or_884_nl, or_926_cse, fsm_output[0]);
  assign or_880_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0110) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_930_nl = MUX_s_1_2_2(or_927_cse, or_880_nl, fsm_output[0]);
  assign mux_932_nl = MUX_s_1_2_2(mux_931_nl, mux_930_nl, fsm_output[6]);
  assign mux_933_nl = MUX_s_1_2_2(or_886_nl, mux_932_nl, fsm_output[1]);
  assign or_887_nl = (fsm_output[3]) | mux_933_nl;
  assign mux_938_nl = MUX_s_1_2_2(nand_47_nl, or_887_nl, fsm_output[2]);
  assign nor_523_nl = ~((fsm_output[8]) | mux_938_nl);
  assign vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_959_nl,
      nor_523_nl, fsm_output[9]);
  assign or_970_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b0111) | (fsm_output[5]) | (fsm_output[1]);
  assign mux_986_nl = MUX_s_1_2_2(or_tmp_910, or_970_nl, fsm_output[0]);
  assign or_969_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0111) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_985_nl = MUX_s_1_2_2(or_969_nl, or_tmp_904, fsm_output[0]);
  assign mux_987_nl = MUX_s_1_2_2(mux_986_nl, mux_985_nl, fsm_output[4]);
  assign nand_52_nl = ~((fsm_output[6]) & (~ mux_987_nl));
  assign or_968_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0111);
  assign mux_988_nl = MUX_s_1_2_2(nand_52_nl, or_968_nl, fsm_output[7]);
  assign nor_503_nl = ~((fsm_output[8]) | mux_988_nl);
  assign and_437_nl = (COMP_LOOP_acc_20_psp_sva[2:0]==3'b011) & (fsm_output[7]) &
      (fsm_output[6]) & (fsm_output[4]) & (fsm_output[0]) & (VEC_LOOP_j_sva_9_0[0])
      & (~ (fsm_output[5])) & (fsm_output[1]);
  assign or_964_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0111) | (fsm_output[5]) |
      (~ (fsm_output[1]));
  assign mux_983_nl = MUX_s_1_2_2(or_964_nl, or_tmp_910, fsm_output[0]);
  assign nor_505_nl = ~((fsm_output[7]) | (fsm_output[6]) | (fsm_output[4]) | mux_983_nl);
  assign mux_984_nl = MUX_s_1_2_2(and_437_nl, nor_505_nl, fsm_output[8]);
  assign mux_989_nl = MUX_s_1_2_2(nor_503_nl, mux_984_nl, fsm_output[9]);
  assign nand_376_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]==3'b011) & (fsm_output[6])
      & (fsm_output[4]) & (fsm_output[0]) & (VEC_LOOP_j_sva_9_0[0]) & (~ (fsm_output[5]))
      & (fsm_output[1]));
  assign or_959_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0111) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_978_nl = MUX_s_1_2_2(or_959_nl, or_tmp_910, fsm_output[0]);
  assign or_957_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b111)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_977_nl = MUX_s_1_2_2(or_tmp_909, or_957_nl, fsm_output[0]);
  assign mux_979_nl = MUX_s_1_2_2(mux_978_nl, mux_977_nl, fsm_output[4]);
  assign or_955_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0111) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_976_nl = MUX_s_1_2_2(or_955_nl, or_tmp_904, fsm_output[0]);
  assign or_956_nl = (fsm_output[4]) | mux_976_nl;
  assign mux_980_nl = MUX_s_1_2_2(mux_979_nl, or_956_nl, fsm_output[6]);
  assign mux_981_nl = MUX_s_1_2_2(nand_376_nl, mux_980_nl, fsm_output[7]);
  assign and_323_nl = (fsm_output[8]) & (~ mux_981_nl);
  assign nor_506_nl = ~((fsm_output[8]) | (fsm_output[7]) | (fsm_output[6]) | (~
      (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b0111));
  assign mux_982_nl = MUX_s_1_2_2(and_323_nl, nor_506_nl, fsm_output[9]);
  assign mux_990_nl = MUX_s_1_2_2(mux_989_nl, mux_982_nl, fsm_output[3]);
  assign nand_371_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]==3'b011) & (fsm_output[4])
      & (fsm_output[0]) & (VEC_LOOP_j_sva_9_0[0]) & (~ (fsm_output[5])) & (fsm_output[1]));
  assign or_950_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0111) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_971_nl = MUX_s_1_2_2(or_950_nl, or_tmp_910, fsm_output[0]);
  assign or_948_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_970_nl = MUX_s_1_2_2(or_tmp_909, or_948_nl, fsm_output[0]);
  assign mux_972_nl = MUX_s_1_2_2(mux_971_nl, mux_970_nl, fsm_output[4]);
  assign mux_973_nl = MUX_s_1_2_2(nand_371_nl, mux_972_nl, fsm_output[6]);
  assign or_946_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0111) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_968_nl = MUX_s_1_2_2(or_946_nl, or_tmp_904, fsm_output[0]);
  assign or_947_nl = (fsm_output[4]) | mux_968_nl;
  assign mux_969_nl = MUX_s_1_2_2(or_947_nl, or_tmp_903, fsm_output[6]);
  assign mux_974_nl = MUX_s_1_2_2(mux_973_nl, mux_969_nl, fsm_output[7]);
  assign nor_507_nl = ~((fsm_output[9:8]!=2'b10) | mux_974_nl);
  assign nand_360_nl = ~((fsm_output[4]) & (fsm_output[0]) & (COMP_LOOP_acc_11_psp_sva[2:0]==3'b011)
      & (VEC_LOOP_j_sva_9_0[0]) & (~ (fsm_output[5])) & (fsm_output[1]));
  assign or_941_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0111) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_964_nl = MUX_s_1_2_2(or_941_nl, or_tmp_910, fsm_output[0]);
  assign or_937_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_963_nl = MUX_s_1_2_2(or_tmp_909, or_937_nl, fsm_output[0]);
  assign mux_965_nl = MUX_s_1_2_2(mux_964_nl, mux_963_nl, fsm_output[4]);
  assign mux_966_nl = MUX_s_1_2_2(nand_360_nl, mux_965_nl, fsm_output[6]);
  assign nand_50_nl = ~((fsm_output[7]) & (~ mux_966_nl));
  assign or_934_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0111) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_961_nl = MUX_s_1_2_2(or_934_nl, or_tmp_904, fsm_output[0]);
  assign or_935_nl = (fsm_output[4]) | mux_961_nl;
  assign mux_962_nl = MUX_s_1_2_2(or_935_nl, or_tmp_903, fsm_output[6]);
  assign or_936_nl = (fsm_output[7]) | mux_962_nl;
  assign mux_967_nl = MUX_s_1_2_2(nand_50_nl, or_936_nl, fsm_output[8]);
  assign nor_508_nl = ~((fsm_output[9]) | mux_967_nl);
  assign mux_975_nl = MUX_s_1_2_2(nor_507_nl, nor_508_nl, fsm_output[3]);
  assign vec_rsc_0_7_i_we_d_pff = MUX_s_1_2_2(mux_990_nl, mux_975_nl, fsm_output[2]);
  assign nor_492_cse = ~((z_out_6_10_1[3:0]!=4'b0111) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nand_280_cse = ~((z_out_6_10_1[3:0]==4'b0111));
  assign nand_275_cse = ~((z_out_6_10_1[3:0]==4'b0111) & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4])));
  assign nand_274_nl = ~((fsm_output[0]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm &
      (COMP_LOOP_acc_1_cse_4_sva[3:0]==4'b0111) & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4])));
  assign or_1022_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | not_tmp_134;
  assign mux_1017_nl = MUX_s_1_2_2(or_1022_nl, nand_275_cse, fsm_output[0]);
  assign mux_1018_nl = MUX_s_1_2_2(nand_274_nl, mux_1017_nl, fsm_output[6]);
  assign or_1019_nl = (z_out_6_10_1[3:1]!=3'b011) | nand_308_cse;
  assign or_1017_nl = (z_out_6_10_1[3:0]!=4'b0111) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_1015_nl = MUX_s_1_2_2(or_1019_nl, or_1017_nl, fsm_output[0]);
  assign nand_370_nl = ~((VEC_LOOP_j_sva_9_0[0]) & (COMP_LOOP_acc_11_psp_sva[2:0]==3'b011)
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (~ (fsm_output[7]))
      & (fsm_output[4]));
  assign or_1014_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0111) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_1014_nl = MUX_s_1_2_2(nand_370_nl, or_1014_nl, fsm_output[0]);
  assign mux_1016_nl = MUX_s_1_2_2(mux_1015_nl, mux_1014_nl, fsm_output[6]);
  assign mux_1019_nl = MUX_s_1_2_2(mux_1018_nl, mux_1016_nl, fsm_output[1]);
  assign nor_484_nl = ~((fsm_output[3]) | mux_1019_nl);
  assign or_1012_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b0111) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_1010_nl = (z_out_6_10_1[3:0]!=4'b0111) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]);
  assign mux_1011_nl = MUX_s_1_2_2(or_1012_nl, or_1010_nl, fsm_output[0]);
  assign or_1009_nl = (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b0111) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_1012_nl = MUX_s_1_2_2(mux_1011_nl, or_1009_nl, fsm_output[6]);
  assign nor_485_nl = ~((fsm_output[1]) | mux_1012_nl);
  assign nor_486_nl = ~((~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b0111) & (fsm_output[1])
      & (fsm_output[6]) & (fsm_output[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      | not_tmp_133);
  assign mux_1013_nl = MUX_s_1_2_2(nor_485_nl, nor_486_nl, fsm_output[3]);
  assign mux_1020_nl = MUX_s_1_2_2(nor_484_nl, mux_1013_nl, fsm_output[2]);
  assign nor_487_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b0111)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign nor_488_nl = ~((~((COMP_LOOP_acc_1_cse_10_sva[3:0]==4'b0111) & (fsm_output[0])
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)) | not_tmp_133);
  assign and_321_nl = (VEC_LOOP_j_sva_9_0[0]) & (COMP_LOOP_acc_17_psp_sva[2:0]==3'b011)
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4]));
  assign nor_489_nl = ~(nand_280_cse | not_tmp_133);
  assign mux_1007_nl = MUX_s_1_2_2(and_321_nl, nor_489_nl, fsm_output[0]);
  assign mux_1008_nl = MUX_s_1_2_2(nor_488_nl, mux_1007_nl, fsm_output[6]);
  assign and_320_nl = (fsm_output[1]) & mux_1008_nl;
  assign mux_1009_nl = MUX_s_1_2_2(nor_487_nl, and_320_nl, fsm_output[3]);
  assign nor_490_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b111)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_491_nl = ~((z_out_6_10_1[3:0]!=4'b0111) | (fsm_output[5]) | not_tmp_134);
  assign mux_1004_nl = MUX_s_1_2_2(nor_490_nl, nor_491_nl, fsm_output[0]);
  assign nor_493_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0111) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_1003_nl = MUX_s_1_2_2(nor_492_cse, nor_493_nl, fsm_output[0]);
  assign mux_1005_nl = MUX_s_1_2_2(mux_1004_nl, mux_1003_nl, fsm_output[6]);
  assign nor_494_nl = ~((~ (VEC_LOOP_j_sva_9_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b011) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]));
  assign and_432_nl = (z_out_6_10_1[3:0]==4'b0111) & (fsm_output[5]) & (~ (fsm_output[7]))
      & (fsm_output[4]);
  assign mux_1001_nl = MUX_s_1_2_2(nor_494_nl, and_432_nl, fsm_output[0]);
  assign nor_496_nl = ~((z_out_6_10_1[3:0]!=4'b0111) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1002_nl = MUX_s_1_2_2(mux_1001_nl, nor_496_nl, fsm_output[6]);
  assign mux_1006_nl = MUX_s_1_2_2(mux_1005_nl, mux_1002_nl, fsm_output[1]);
  assign and_322_nl = (fsm_output[3]) & mux_1006_nl;
  assign mux_1010_nl = MUX_s_1_2_2(mux_1009_nl, and_322_nl, fsm_output[2]);
  assign mux_1021_nl = MUX_s_1_2_2(mux_1020_nl, mux_1010_nl, fsm_output[8]);
  assign nor_499_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0111) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_997_nl = MUX_s_1_2_2(nor_492_cse, nor_499_nl, fsm_output[0]);
  assign nor_500_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_501_nl = ~((z_out_6_10_1[3:0]!=4'b0111) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_996_nl = MUX_s_1_2_2(nor_500_nl, nor_501_nl, fsm_output[0]);
  assign mux_998_nl = MUX_s_1_2_2(mux_997_nl, mux_996_nl, fsm_output[6]);
  assign nor_502_nl = ~((z_out_6_10_1[3:0]!=4'b0111) | (fsm_output[6]) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_999_nl = MUX_s_1_2_2(mux_998_nl, nor_502_nl, fsm_output[1]);
  assign nand_53_nl = ~((fsm_output[3]) & mux_999_nl);
  assign or_979_nl = (~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b0111) & (fsm_output[6])
      & (fsm_output[0]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & (~ (fsm_output[5]))))
      | not_tmp_134;
  assign nand_282_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]==3'b011) & (VEC_LOOP_j_sva_9_0[0])
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4])));
  assign or_976_nl = nand_280_cse | not_tmp_133;
  assign mux_993_nl = MUX_s_1_2_2(nand_282_nl, or_976_nl, fsm_output[0]);
  assign nand_354_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b0111) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[5]) & (~ (fsm_output[7])) & (fsm_output[4]));
  assign mux_992_nl = MUX_s_1_2_2(nand_275_cse, nand_354_nl, fsm_output[0]);
  assign mux_994_nl = MUX_s_1_2_2(mux_993_nl, mux_992_nl, fsm_output[6]);
  assign mux_995_nl = MUX_s_1_2_2(or_979_nl, mux_994_nl, fsm_output[1]);
  assign or_980_nl = (fsm_output[3]) | mux_995_nl;
  assign mux_1000_nl = MUX_s_1_2_2(nand_53_nl, or_980_nl, fsm_output[2]);
  assign nor_497_nl = ~((fsm_output[8]) | mux_1000_nl);
  assign vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1021_nl,
      nor_497_nl, fsm_output[9]);
  assign or_1069_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b1000) | (fsm_output[5]) | (fsm_output[1]);
  assign mux_1048_nl = MUX_s_1_2_2(or_tmp_1007, or_1069_nl, fsm_output[0]);
  assign or_1068_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1000) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1047_nl = MUX_s_1_2_2(or_1068_nl, or_tmp_999, fsm_output[0]);
  assign mux_1049_nl = MUX_s_1_2_2(mux_1048_nl, mux_1047_nl, fsm_output[4]);
  assign nand_58_nl = ~((fsm_output[6]) & (~ mux_1049_nl));
  assign or_1067_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1000);
  assign mux_1050_nl = MUX_s_1_2_2(nand_58_nl, or_1067_nl, fsm_output[7]);
  assign nor_478_nl = ~((fsm_output[8]) | mux_1050_nl);
  assign nor_479_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b100) | (~ (fsm_output[7]))
      | (~ (fsm_output[6])) | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0])
      | (fsm_output[5]) | (~ (fsm_output[1])));
  assign or_1062_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1000) | (fsm_output[5]) |
      (~ (fsm_output[1]));
  assign mux_1045_nl = MUX_s_1_2_2(or_1062_nl, or_tmp_1007, fsm_output[0]);
  assign nor_480_nl = ~((fsm_output[7]) | (fsm_output[6]) | (fsm_output[4]) | mux_1045_nl);
  assign mux_1046_nl = MUX_s_1_2_2(nor_479_nl, nor_480_nl, fsm_output[8]);
  assign mux_1051_nl = MUX_s_1_2_2(nor_478_nl, mux_1046_nl, fsm_output[9]);
  assign or_1059_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign or_1057_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1000) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_1040_nl = MUX_s_1_2_2(or_1057_nl, or_tmp_1007, fsm_output[0]);
  assign or_1055_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b000)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_1039_nl = MUX_s_1_2_2(or_tmp_1005, or_1055_nl, fsm_output[0]);
  assign mux_1041_nl = MUX_s_1_2_2(mux_1040_nl, mux_1039_nl, fsm_output[4]);
  assign or_1053_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1000) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1038_nl = MUX_s_1_2_2(or_1053_nl, or_tmp_999, fsm_output[0]);
  assign or_1054_nl = (fsm_output[4]) | mux_1038_nl;
  assign mux_1042_nl = MUX_s_1_2_2(mux_1041_nl, or_1054_nl, fsm_output[6]);
  assign mux_1043_nl = MUX_s_1_2_2(or_1059_nl, mux_1042_nl, fsm_output[7]);
  assign and_319_nl = (fsm_output[8]) & (~ mux_1043_nl);
  assign nor_481_nl = ~((fsm_output[8]) | (fsm_output[7]) | (fsm_output[6]) | (~
      (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1000));
  assign mux_1044_nl = MUX_s_1_2_2(and_319_nl, nor_481_nl, fsm_output[9]);
  assign mux_1052_nl = MUX_s_1_2_2(mux_1051_nl, mux_1044_nl, fsm_output[3]);
  assign or_1049_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b100) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5]) | (~ (fsm_output[1]));
  assign or_1047_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1000) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_1033_nl = MUX_s_1_2_2(or_1047_nl, or_tmp_1007, fsm_output[0]);
  assign or_1045_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_1032_nl = MUX_s_1_2_2(or_tmp_1005, or_1045_nl, fsm_output[0]);
  assign mux_1034_nl = MUX_s_1_2_2(mux_1033_nl, mux_1032_nl, fsm_output[4]);
  assign mux_1035_nl = MUX_s_1_2_2(or_1049_nl, mux_1034_nl, fsm_output[6]);
  assign or_1043_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1000) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1030_nl = MUX_s_1_2_2(or_1043_nl, or_tmp_999, fsm_output[0]);
  assign or_1044_nl = (fsm_output[4]) | mux_1030_nl;
  assign mux_1031_nl = MUX_s_1_2_2(or_1044_nl, or_tmp_997, fsm_output[6]);
  assign mux_1036_nl = MUX_s_1_2_2(mux_1035_nl, mux_1031_nl, fsm_output[7]);
  assign nor_482_nl = ~((fsm_output[9:8]!=2'b10) | mux_1036_nl);
  assign or_1040_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100)
      | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5]) | (~ (fsm_output[1]));
  assign or_1038_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1000) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_1026_nl = MUX_s_1_2_2(or_1038_nl, or_tmp_1007, fsm_output[0]);
  assign or_1032_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_1025_nl = MUX_s_1_2_2(or_tmp_1005, or_1032_nl, fsm_output[0]);
  assign mux_1027_nl = MUX_s_1_2_2(mux_1026_nl, mux_1025_nl, fsm_output[4]);
  assign mux_1028_nl = MUX_s_1_2_2(or_1040_nl, mux_1027_nl, fsm_output[6]);
  assign nand_56_nl = ~((fsm_output[7]) & (~ mux_1028_nl));
  assign or_1029_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1000) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1023_nl = MUX_s_1_2_2(or_1029_nl, or_tmp_999, fsm_output[0]);
  assign or_1030_nl = (fsm_output[4]) | mux_1023_nl;
  assign mux_1024_nl = MUX_s_1_2_2(or_1030_nl, or_tmp_997, fsm_output[6]);
  assign or_1031_nl = (fsm_output[7]) | mux_1024_nl;
  assign mux_1029_nl = MUX_s_1_2_2(nand_56_nl, or_1031_nl, fsm_output[8]);
  assign nor_483_nl = ~((fsm_output[9]) | mux_1029_nl);
  assign mux_1037_nl = MUX_s_1_2_2(nor_482_nl, nor_483_nl, fsm_output[3]);
  assign vec_rsc_0_8_i_we_d_pff = MUX_s_1_2_2(mux_1052_nl, mux_1037_nl, fsm_output[2]);
  assign nor_467_cse = ~((z_out_6_10_1[3:0]!=4'b1000) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign or_1119_cse = (z_out_6_10_1[3:0]!=4'b1000) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_1122_nl = (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1000) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_1121_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | not_tmp_134;
  assign mux_1079_nl = MUX_s_1_2_2(or_1121_nl, or_1119_cse, fsm_output[0]);
  assign mux_1080_nl = MUX_s_1_2_2(or_1122_nl, mux_1079_nl, fsm_output[6]);
  assign or_1118_nl = (z_out_6_10_1[3:0]!=4'b1000) | not_tmp_133;
  assign or_1116_nl = (z_out_6_10_1[3:0]!=4'b1000) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_1077_nl = MUX_s_1_2_2(or_1118_nl, or_1116_nl, fsm_output[0]);
  assign or_1115_nl = (VEC_LOOP_j_sva_9_0[0]) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_1113_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1000) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_1076_nl = MUX_s_1_2_2(or_1115_nl, or_1113_nl, fsm_output[0]);
  assign mux_1078_nl = MUX_s_1_2_2(mux_1077_nl, mux_1076_nl, fsm_output[6]);
  assign mux_1081_nl = MUX_s_1_2_2(mux_1080_nl, mux_1078_nl, fsm_output[1]);
  assign nor_458_nl = ~((fsm_output[3]) | mux_1081_nl);
  assign or_1111_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b1000) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_1109_nl = (z_out_6_10_1[3:0]!=4'b1000) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]);
  assign mux_1073_nl = MUX_s_1_2_2(or_1111_nl, or_1109_nl, fsm_output[0]);
  assign or_1108_nl = (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b1000) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_1074_nl = MUX_s_1_2_2(mux_1073_nl, or_1108_nl, fsm_output[6]);
  assign nor_459_nl = ~((fsm_output[1]) | mux_1074_nl);
  assign nor_460_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1000) | (~ (fsm_output[1]))
      | (~ (fsm_output[6])) | (~ (fsm_output[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | not_tmp_133);
  assign mux_1075_nl = MUX_s_1_2_2(nor_459_nl, nor_460_nl, fsm_output[3]);
  assign mux_1082_nl = MUX_s_1_2_2(nor_458_nl, mux_1075_nl, fsm_output[2]);
  assign nor_461_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b1000)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign nor_462_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1000) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | not_tmp_133);
  assign nor_463_nl = ~((VEC_LOOP_j_sva_9_0[0]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b100)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_464_nl = ~((z_out_6_10_1[2:0]!=3'b000) | nand_270_cse_1);
  assign mux_1069_nl = MUX_s_1_2_2(nor_463_nl, nor_464_nl, fsm_output[0]);
  assign mux_1070_nl = MUX_s_1_2_2(nor_462_nl, mux_1069_nl, fsm_output[6]);
  assign and_317_nl = (fsm_output[1]) & mux_1070_nl;
  assign mux_1071_nl = MUX_s_1_2_2(nor_461_nl, and_317_nl, fsm_output[3]);
  assign nor_465_nl = ~((~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b000)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_466_nl = ~((z_out_6_10_1[3:0]!=4'b1000) | (fsm_output[5]) | not_tmp_134);
  assign mux_1066_nl = MUX_s_1_2_2(nor_465_nl, nor_466_nl, fsm_output[0]);
  assign nor_468_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_1065_nl = MUX_s_1_2_2(nor_467_cse, nor_468_nl, fsm_output[0]);
  assign mux_1067_nl = MUX_s_1_2_2(mux_1066_nl, mux_1065_nl, fsm_output[6]);
  assign nor_469_nl = ~((VEC_LOOP_j_sva_9_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_470_nl = ~((z_out_6_10_1[3:0]!=4'b1000) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_1063_nl = MUX_s_1_2_2(nor_469_nl, nor_470_nl, fsm_output[0]);
  assign nor_471_nl = ~((z_out_6_10_1[3:0]!=4'b1000) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1064_nl = MUX_s_1_2_2(mux_1063_nl, nor_471_nl, fsm_output[6]);
  assign mux_1068_nl = MUX_s_1_2_2(mux_1067_nl, mux_1064_nl, fsm_output[1]);
  assign and_318_nl = (fsm_output[3]) & mux_1068_nl;
  assign mux_1072_nl = MUX_s_1_2_2(mux_1071_nl, and_318_nl, fsm_output[2]);
  assign mux_1083_nl = MUX_s_1_2_2(mux_1082_nl, mux_1072_nl, fsm_output[8]);
  assign nor_474_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_1059_nl = MUX_s_1_2_2(nor_467_cse, nor_474_nl, fsm_output[0]);
  assign nor_475_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_476_nl = ~((z_out_6_10_1[3:0]!=4'b1000) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_1058_nl = MUX_s_1_2_2(nor_475_nl, nor_476_nl, fsm_output[0]);
  assign mux_1060_nl = MUX_s_1_2_2(mux_1059_nl, mux_1058_nl, fsm_output[6]);
  assign nor_477_nl = ~((z_out_6_10_1[3:0]!=4'b1000) | (fsm_output[6]) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1061_nl = MUX_s_1_2_2(mux_1060_nl, nor_477_nl, fsm_output[1]);
  assign nand_59_nl = ~((fsm_output[3]) & mux_1061_nl);
  assign or_1078_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1000) | (~ (fsm_output[6]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[5])
      | not_tmp_134;
  assign or_1076_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_1075_nl = (z_out_6_10_1[2:0]!=3'b000) | nand_270_cse_1;
  assign mux_1055_nl = MUX_s_1_2_2(or_1076_nl, or_1075_nl, fsm_output[0]);
  assign or_1072_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1000) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_1054_nl = MUX_s_1_2_2(or_1119_cse, or_1072_nl, fsm_output[0]);
  assign mux_1056_nl = MUX_s_1_2_2(mux_1055_nl, mux_1054_nl, fsm_output[6]);
  assign mux_1057_nl = MUX_s_1_2_2(or_1078_nl, mux_1056_nl, fsm_output[1]);
  assign or_1079_nl = (fsm_output[3]) | mux_1057_nl;
  assign mux_1062_nl = MUX_s_1_2_2(nand_59_nl, or_1079_nl, fsm_output[2]);
  assign nor_472_nl = ~((fsm_output[8]) | mux_1062_nl);
  assign vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1083_nl,
      nor_472_nl, fsm_output[9]);
  assign or_1169_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b1001) | (fsm_output[1]) | (fsm_output[5]);
  assign mux_1110_nl = MUX_s_1_2_2(or_tmp_1106, or_1169_nl, fsm_output[0]);
  assign or_1168_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1001) | (fsm_output[1])
      | (~ (fsm_output[5]));
  assign mux_1109_nl = MUX_s_1_2_2(or_1168_nl, or_tmp_1097, fsm_output[0]);
  assign mux_1111_nl = MUX_s_1_2_2(mux_1110_nl, mux_1109_nl, fsm_output[4]);
  assign nor_450_nl = ~((fsm_output[9]) | (~ (fsm_output[6])) | mux_1111_nl);
  assign or_1166_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b100) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_9_0[0])) | (~ (fsm_output[1])) |
      (fsm_output[5]);
  assign or_1165_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1001) | (~ (fsm_output[1]))
      | (fsm_output[5]);
  assign mux_1106_nl = MUX_s_1_2_2(or_1165_nl, or_tmp_1106, fsm_output[0]);
  assign or_1164_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (fsm_output[1]) | (~ (fsm_output[5]));
  assign mux_1105_nl = MUX_s_1_2_2(or_tmp_1104, or_1164_nl, fsm_output[0]);
  assign mux_1107_nl = MUX_s_1_2_2(mux_1106_nl, mux_1105_nl, fsm_output[4]);
  assign mux_1108_nl = MUX_s_1_2_2(or_1166_nl, mux_1107_nl, fsm_output[6]);
  assign and_316_nl = (fsm_output[9]) & (~ mux_1108_nl);
  assign mux_1112_nl = MUX_s_1_2_2(nor_450_nl, and_316_nl, fsm_output[2]);
  assign or_1161_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1001) | (~ (fsm_output[1]))
      | (fsm_output[5]);
  assign mux_1104_nl = MUX_s_1_2_2(or_1161_nl, or_tmp_1106, fsm_output[0]);
  assign nor_451_nl = ~((fsm_output[2]) | (~ (fsm_output[9])) | (fsm_output[6]) |
      (fsm_output[4]) | mux_1104_nl);
  assign mux_1113_nl = MUX_s_1_2_2(mux_1112_nl, nor_451_nl, fsm_output[8]);
  assign or_1158_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (fsm_output[1])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1001);
  assign or_1156_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b100) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_9_0[0])) |
      (~ (fsm_output[1])) | (fsm_output[5]);
  assign mux_1102_nl = MUX_s_1_2_2(or_1158_nl, or_1156_nl, fsm_output[9]);
  assign or_1154_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1001) | (fsm_output[1])
      | (~ (fsm_output[5]));
  assign mux_1100_nl = MUX_s_1_2_2(or_1154_nl, or_tmp_1097, fsm_output[0]);
  assign or_1155_nl = (fsm_output[4]) | mux_1100_nl;
  assign mux_1101_nl = MUX_s_1_2_2(or_1155_nl, or_tmp_1116, fsm_output[6]);
  assign nand_62_nl = ~((fsm_output[9]) & (~ mux_1101_nl));
  assign mux_1103_nl = MUX_s_1_2_2(mux_1102_nl, nand_62_nl, fsm_output[2]);
  assign nor_452_nl = ~((fsm_output[8]) | mux_1103_nl);
  assign mux_1114_nl = MUX_s_1_2_2(mux_1113_nl, nor_452_nl, fsm_output[7]);
  assign nor_453_nl = ~((fsm_output[2]) | (~ (fsm_output[9])) | (fsm_output[6]) |
      (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[5]) |
      (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1001));
  assign nor_454_nl = ~((fsm_output[9]) | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100)
      | (~ (fsm_output[6])) | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (~ (VEC_LOOP_j_sva_9_0[0]))
      | (~ (fsm_output[1])) | (fsm_output[5]));
  assign or_1147_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1001) | (fsm_output[1])
      | (~ (fsm_output[5]));
  assign mux_1095_nl = MUX_s_1_2_2(or_1147_nl, or_tmp_1097, fsm_output[0]);
  assign or_1148_nl = (fsm_output[4]) | mux_1095_nl;
  assign mux_1096_nl = MUX_s_1_2_2(or_1148_nl, or_tmp_1116, fsm_output[6]);
  assign nor_455_nl = ~((fsm_output[9]) | mux_1096_nl);
  assign mux_1097_nl = MUX_s_1_2_2(nor_454_nl, nor_455_nl, fsm_output[2]);
  assign mux_1098_nl = MUX_s_1_2_2(nor_453_nl, mux_1097_nl, fsm_output[8]);
  assign or_1142_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100)
      | (~ (VEC_LOOP_j_sva_9_0[0])) | (~ (fsm_output[1])) | (fsm_output[5]);
  assign or_1141_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1001) | (~ (fsm_output[1]))
      | (fsm_output[5]);
  assign mux_1091_nl = MUX_s_1_2_2(or_1141_nl, or_tmp_1106, fsm_output[0]);
  assign or_1140_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (fsm_output[1]) | (~ (fsm_output[5]));
  assign mux_1090_nl = MUX_s_1_2_2(or_tmp_1104, or_1140_nl, fsm_output[0]);
  assign mux_1092_nl = MUX_s_1_2_2(mux_1091_nl, mux_1090_nl, fsm_output[4]);
  assign mux_1093_nl = MUX_s_1_2_2(or_1142_nl, mux_1092_nl, fsm_output[6]);
  assign nor_456_nl = ~((~ (fsm_output[2])) | (fsm_output[9]) | mux_1093_nl);
  assign or_1136_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1001) | (~ (fsm_output[1]))
      | (fsm_output[5]);
  assign mux_1087_nl = MUX_s_1_2_2(or_1136_nl, or_tmp_1106, fsm_output[0]);
  assign or_1131_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b001)
      | (fsm_output[1]) | (~ (fsm_output[5]));
  assign mux_1086_nl = MUX_s_1_2_2(or_tmp_1104, or_1131_nl, fsm_output[0]);
  assign mux_1088_nl = MUX_s_1_2_2(mux_1087_nl, mux_1086_nl, fsm_output[4]);
  assign or_1128_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1001) | (fsm_output[1])
      | (~ (fsm_output[5]));
  assign mux_1085_nl = MUX_s_1_2_2(or_1128_nl, or_tmp_1097, fsm_output[0]);
  assign or_1129_nl = (fsm_output[4]) | mux_1085_nl;
  assign mux_1089_nl = MUX_s_1_2_2(mux_1088_nl, or_1129_nl, fsm_output[6]);
  assign nor_457_nl = ~((fsm_output[2]) | (fsm_output[9]) | mux_1089_nl);
  assign mux_1094_nl = MUX_s_1_2_2(nor_456_nl, nor_457_nl, fsm_output[8]);
  assign mux_1099_nl = MUX_s_1_2_2(mux_1098_nl, mux_1094_nl, fsm_output[7]);
  assign vec_rsc_0_9_i_we_d_pff = MUX_s_1_2_2(mux_1114_nl, mux_1099_nl, fsm_output[3]);
  assign nor_439_cse = ~((z_out_6_10_1[3:0]!=4'b1001) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign or_1218_cse = (z_out_6_10_1[3:0]!=4'b1001) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_1221_nl = (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1001) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_1220_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | not_tmp_134;
  assign mux_1141_nl = MUX_s_1_2_2(or_1220_nl, or_1218_cse, fsm_output[0]);
  assign mux_1142_nl = MUX_s_1_2_2(or_1221_nl, mux_1141_nl, fsm_output[6]);
  assign or_1217_nl = (z_out_6_10_1[2:1]!=2'b00) | nand_264_cse;
  assign or_1215_nl = (z_out_6_10_1[3:0]!=4'b1001) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_1139_nl = MUX_s_1_2_2(or_1217_nl, or_1215_nl, fsm_output[0]);
  assign or_1214_nl = (~ (VEC_LOOP_j_sva_9_0[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_1212_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1001) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_1138_nl = MUX_s_1_2_2(or_1214_nl, or_1212_nl, fsm_output[0]);
  assign mux_1140_nl = MUX_s_1_2_2(mux_1139_nl, mux_1138_nl, fsm_output[6]);
  assign mux_1143_nl = MUX_s_1_2_2(mux_1142_nl, mux_1140_nl, fsm_output[1]);
  assign nor_430_nl = ~((fsm_output[3]) | mux_1143_nl);
  assign or_1210_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b1001) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_1208_nl = (z_out_6_10_1[3:0]!=4'b1001) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]);
  assign mux_1135_nl = MUX_s_1_2_2(or_1210_nl, or_1208_nl, fsm_output[0]);
  assign or_1207_nl = (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b1001) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_1136_nl = MUX_s_1_2_2(mux_1135_nl, or_1207_nl, fsm_output[6]);
  assign nor_431_nl = ~((fsm_output[1]) | mux_1136_nl);
  assign nor_432_nl = ~((~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1001) & (fsm_output[1])
      & (fsm_output[6]) & (fsm_output[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      | not_tmp_133);
  assign mux_1137_nl = MUX_s_1_2_2(nor_431_nl, nor_432_nl, fsm_output[3]);
  assign mux_1144_nl = MUX_s_1_2_2(nor_430_nl, mux_1137_nl, fsm_output[2]);
  assign nor_433_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b1001)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign nor_434_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1001) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | not_tmp_133);
  assign nor_435_nl = ~((~ (VEC_LOOP_j_sva_9_0[0])) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b100)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_436_nl = ~((z_out_6_10_1[2:0]!=3'b001) | nand_270_cse_1);
  assign mux_1131_nl = MUX_s_1_2_2(nor_435_nl, nor_436_nl, fsm_output[0]);
  assign mux_1132_nl = MUX_s_1_2_2(nor_434_nl, mux_1131_nl, fsm_output[6]);
  assign and_314_nl = (fsm_output[1]) & mux_1132_nl;
  assign mux_1133_nl = MUX_s_1_2_2(nor_433_nl, and_314_nl, fsm_output[3]);
  assign nor_437_nl = ~((~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b001)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_438_nl = ~((z_out_6_10_1[3:0]!=4'b1001) | (fsm_output[5]) | not_tmp_134);
  assign mux_1128_nl = MUX_s_1_2_2(nor_437_nl, nor_438_nl, fsm_output[0]);
  assign nor_440_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_1127_nl = MUX_s_1_2_2(nor_439_cse, nor_440_nl, fsm_output[0]);
  assign mux_1129_nl = MUX_s_1_2_2(mux_1128_nl, mux_1127_nl, fsm_output[6]);
  assign nor_441_nl = ~((~ (VEC_LOOP_j_sva_9_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_442_nl = ~((z_out_6_10_1[3:0]!=4'b1001) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_1125_nl = MUX_s_1_2_2(nor_441_nl, nor_442_nl, fsm_output[0]);
  assign nor_443_nl = ~((z_out_6_10_1[3:0]!=4'b1001) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1126_nl = MUX_s_1_2_2(mux_1125_nl, nor_443_nl, fsm_output[6]);
  assign mux_1130_nl = MUX_s_1_2_2(mux_1129_nl, mux_1126_nl, fsm_output[1]);
  assign and_315_nl = (fsm_output[3]) & mux_1130_nl;
  assign mux_1134_nl = MUX_s_1_2_2(mux_1133_nl, and_315_nl, fsm_output[2]);
  assign mux_1145_nl = MUX_s_1_2_2(mux_1144_nl, mux_1134_nl, fsm_output[8]);
  assign nor_446_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_1121_nl = MUX_s_1_2_2(nor_439_cse, nor_446_nl, fsm_output[0]);
  assign nor_447_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_448_nl = ~((z_out_6_10_1[3:0]!=4'b1001) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_1120_nl = MUX_s_1_2_2(nor_447_nl, nor_448_nl, fsm_output[0]);
  assign mux_1122_nl = MUX_s_1_2_2(mux_1121_nl, mux_1120_nl, fsm_output[6]);
  assign nor_449_nl = ~((z_out_6_10_1[3:0]!=4'b1001) | (fsm_output[6]) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1123_nl = MUX_s_1_2_2(mux_1122_nl, nor_449_nl, fsm_output[1]);
  assign nand_65_nl = ~((fsm_output[3]) & mux_1123_nl);
  assign or_1177_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1001) | (~ (fsm_output[6]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[5])
      | not_tmp_134;
  assign or_1175_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b100) | (~ (VEC_LOOP_j_sva_9_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_1174_nl = (z_out_6_10_1[2:0]!=3'b001) | nand_270_cse_1;
  assign mux_1117_nl = MUX_s_1_2_2(or_1175_nl, or_1174_nl, fsm_output[0]);
  assign or_1171_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1001) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_1116_nl = MUX_s_1_2_2(or_1218_cse, or_1171_nl, fsm_output[0]);
  assign mux_1118_nl = MUX_s_1_2_2(mux_1117_nl, mux_1116_nl, fsm_output[6]);
  assign mux_1119_nl = MUX_s_1_2_2(or_1177_nl, mux_1118_nl, fsm_output[1]);
  assign or_1178_nl = (fsm_output[3]) | mux_1119_nl;
  assign mux_1124_nl = MUX_s_1_2_2(nand_65_nl, or_1178_nl, fsm_output[2]);
  assign nor_444_nl = ~((fsm_output[8]) | mux_1124_nl);
  assign vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1145_nl,
      nor_444_nl, fsm_output[9]);
  assign or_1267_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b1010) | (fsm_output[5]) | (fsm_output[1]);
  assign mux_1172_nl = MUX_s_1_2_2(or_tmp_1205, or_1267_nl, fsm_output[0]);
  assign or_1266_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1010) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1171_nl = MUX_s_1_2_2(or_1266_nl, or_tmp_1197, fsm_output[0]);
  assign mux_1173_nl = MUX_s_1_2_2(mux_1172_nl, mux_1171_nl, fsm_output[4]);
  assign nand_70_nl = ~((fsm_output[6]) & (~ mux_1173_nl));
  assign or_1265_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1010);
  assign mux_1174_nl = MUX_s_1_2_2(nand_70_nl, or_1265_nl, fsm_output[7]);
  assign nor_424_nl = ~((fsm_output[8]) | mux_1174_nl);
  assign and_442_nl = (COMP_LOOP_acc_20_psp_sva[2:0]==3'b101) & (fsm_output[7]) &
      (fsm_output[6]) & (fsm_output[4]) & (fsm_output[0]) & (~ (VEC_LOOP_j_sva_9_0[0]))
      & (~ (fsm_output[5])) & (fsm_output[1]);
  assign or_1260_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1010) | (fsm_output[5]) |
      (~ (fsm_output[1]));
  assign mux_1169_nl = MUX_s_1_2_2(or_1260_nl, or_tmp_1205, fsm_output[0]);
  assign nor_426_nl = ~((fsm_output[7]) | (fsm_output[6]) | (fsm_output[4]) | mux_1169_nl);
  assign mux_1170_nl = MUX_s_1_2_2(and_442_nl, nor_426_nl, fsm_output[8]);
  assign mux_1175_nl = MUX_s_1_2_2(nor_424_nl, mux_1170_nl, fsm_output[9]);
  assign or_1257_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b101) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign or_1255_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1010) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_1164_nl = MUX_s_1_2_2(or_1255_nl, or_tmp_1205, fsm_output[0]);
  assign or_1253_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b010)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_1163_nl = MUX_s_1_2_2(or_tmp_1203, or_1253_nl, fsm_output[0]);
  assign mux_1165_nl = MUX_s_1_2_2(mux_1164_nl, mux_1163_nl, fsm_output[4]);
  assign or_1251_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1010) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1162_nl = MUX_s_1_2_2(or_1251_nl, or_tmp_1197, fsm_output[0]);
  assign or_1252_nl = (fsm_output[4]) | mux_1162_nl;
  assign mux_1166_nl = MUX_s_1_2_2(mux_1165_nl, or_1252_nl, fsm_output[6]);
  assign mux_1167_nl = MUX_s_1_2_2(or_1257_nl, mux_1166_nl, fsm_output[7]);
  assign and_313_nl = (fsm_output[8]) & (~ mux_1167_nl);
  assign nor_427_nl = ~((fsm_output[8]) | (fsm_output[7]) | (fsm_output[6]) | (~
      (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1010));
  assign mux_1168_nl = MUX_s_1_2_2(and_313_nl, nor_427_nl, fsm_output[9]);
  assign mux_1176_nl = MUX_s_1_2_2(mux_1175_nl, mux_1168_nl, fsm_output[3]);
  assign or_1247_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b101) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5]) | (~ (fsm_output[1]));
  assign or_1245_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1010) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_1157_nl = MUX_s_1_2_2(or_1245_nl, or_tmp_1205, fsm_output[0]);
  assign or_1243_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_1156_nl = MUX_s_1_2_2(or_tmp_1203, or_1243_nl, fsm_output[0]);
  assign mux_1158_nl = MUX_s_1_2_2(mux_1157_nl, mux_1156_nl, fsm_output[4]);
  assign mux_1159_nl = MUX_s_1_2_2(or_1247_nl, mux_1158_nl, fsm_output[6]);
  assign or_1241_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1010) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1154_nl = MUX_s_1_2_2(or_1241_nl, or_tmp_1197, fsm_output[0]);
  assign or_1242_nl = (fsm_output[4]) | mux_1154_nl;
  assign mux_1155_nl = MUX_s_1_2_2(or_1242_nl, or_tmp_1195, fsm_output[6]);
  assign mux_1160_nl = MUX_s_1_2_2(mux_1159_nl, mux_1155_nl, fsm_output[7]);
  assign nor_428_nl = ~((fsm_output[9:8]!=2'b10) | mux_1160_nl);
  assign or_1238_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b101)
      | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5]) | (~ (fsm_output[1]));
  assign or_1236_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1010) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_1150_nl = MUX_s_1_2_2(or_1236_nl, or_tmp_1205, fsm_output[0]);
  assign or_1230_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_1149_nl = MUX_s_1_2_2(or_tmp_1203, or_1230_nl, fsm_output[0]);
  assign mux_1151_nl = MUX_s_1_2_2(mux_1150_nl, mux_1149_nl, fsm_output[4]);
  assign mux_1152_nl = MUX_s_1_2_2(or_1238_nl, mux_1151_nl, fsm_output[6]);
  assign nand_68_nl = ~((fsm_output[7]) & (~ mux_1152_nl));
  assign or_1227_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1010) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1147_nl = MUX_s_1_2_2(or_1227_nl, or_tmp_1197, fsm_output[0]);
  assign or_1228_nl = (fsm_output[4]) | mux_1147_nl;
  assign mux_1148_nl = MUX_s_1_2_2(or_1228_nl, or_tmp_1195, fsm_output[6]);
  assign or_1229_nl = (fsm_output[7]) | mux_1148_nl;
  assign mux_1153_nl = MUX_s_1_2_2(nand_68_nl, or_1229_nl, fsm_output[8]);
  assign nor_429_nl = ~((fsm_output[9]) | mux_1153_nl);
  assign mux_1161_nl = MUX_s_1_2_2(nor_428_nl, nor_429_nl, fsm_output[3]);
  assign vec_rsc_0_10_i_we_d_pff = MUX_s_1_2_2(mux_1176_nl, mux_1161_nl, fsm_output[2]);
  assign nor_413_cse = ~((z_out_6_10_1[3:0]!=4'b1010) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign or_1317_cse = (z_out_6_10_1[3:0]!=4'b1010) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_1320_nl = (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1010) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_1319_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | not_tmp_134;
  assign mux_1203_nl = MUX_s_1_2_2(or_1319_nl, or_1317_cse, fsm_output[0]);
  assign mux_1204_nl = MUX_s_1_2_2(or_1320_nl, mux_1203_nl, fsm_output[6]);
  assign or_1316_nl = (z_out_6_10_1[3:0]!=4'b1010) | not_tmp_133;
  assign or_1314_nl = (z_out_6_10_1[3:0]!=4'b1010) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_1201_nl = MUX_s_1_2_2(or_1316_nl, or_1314_nl, fsm_output[0]);
  assign or_1313_nl = (VEC_LOOP_j_sva_9_0[0]) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b101)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_1311_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1010) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_1200_nl = MUX_s_1_2_2(or_1313_nl, or_1311_nl, fsm_output[0]);
  assign mux_1202_nl = MUX_s_1_2_2(mux_1201_nl, mux_1200_nl, fsm_output[6]);
  assign mux_1205_nl = MUX_s_1_2_2(mux_1204_nl, mux_1202_nl, fsm_output[1]);
  assign nor_404_nl = ~((fsm_output[3]) | mux_1205_nl);
  assign or_1309_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b1010) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_1307_nl = (z_out_6_10_1[3:0]!=4'b1010) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]);
  assign mux_1197_nl = MUX_s_1_2_2(or_1309_nl, or_1307_nl, fsm_output[0]);
  assign or_1306_nl = (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b1010) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_1198_nl = MUX_s_1_2_2(mux_1197_nl, or_1306_nl, fsm_output[6]);
  assign nor_405_nl = ~((fsm_output[1]) | mux_1198_nl);
  assign nor_406_nl = ~((~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1010) & (fsm_output[1])
      & (fsm_output[6]) & (fsm_output[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      | not_tmp_133);
  assign mux_1199_nl = MUX_s_1_2_2(nor_405_nl, nor_406_nl, fsm_output[3]);
  assign mux_1206_nl = MUX_s_1_2_2(nor_404_nl, mux_1199_nl, fsm_output[2]);
  assign nor_407_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b1010)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign nor_408_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1010) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | not_tmp_133);
  assign nor_409_nl = ~((VEC_LOOP_j_sva_9_0[0]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b101)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_410_nl = ~((z_out_6_10_1[0]) | (z_out_6_10_1[2]) | nand_260_cse_1);
  assign mux_1193_nl = MUX_s_1_2_2(nor_409_nl, nor_410_nl, fsm_output[0]);
  assign mux_1194_nl = MUX_s_1_2_2(nor_408_nl, mux_1193_nl, fsm_output[6]);
  assign and_311_nl = (fsm_output[1]) & mux_1194_nl;
  assign mux_1195_nl = MUX_s_1_2_2(nor_407_nl, and_311_nl, fsm_output[3]);
  assign nor_411_nl = ~((~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b010)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_412_nl = ~((z_out_6_10_1[3:0]!=4'b1010) | (fsm_output[5]) | not_tmp_134);
  assign mux_1190_nl = MUX_s_1_2_2(nor_411_nl, nor_412_nl, fsm_output[0]);
  assign nor_414_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_1189_nl = MUX_s_1_2_2(nor_413_cse, nor_414_nl, fsm_output[0]);
  assign mux_1191_nl = MUX_s_1_2_2(mux_1190_nl, mux_1189_nl, fsm_output[6]);
  assign nor_415_nl = ~((VEC_LOOP_j_sva_9_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b101) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_416_nl = ~((z_out_6_10_1[3:0]!=4'b1010) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_1187_nl = MUX_s_1_2_2(nor_415_nl, nor_416_nl, fsm_output[0]);
  assign nor_417_nl = ~((z_out_6_10_1[3:0]!=4'b1010) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1188_nl = MUX_s_1_2_2(mux_1187_nl, nor_417_nl, fsm_output[6]);
  assign mux_1192_nl = MUX_s_1_2_2(mux_1191_nl, mux_1188_nl, fsm_output[1]);
  assign and_312_nl = (fsm_output[3]) & mux_1192_nl;
  assign mux_1196_nl = MUX_s_1_2_2(mux_1195_nl, and_312_nl, fsm_output[2]);
  assign mux_1207_nl = MUX_s_1_2_2(mux_1206_nl, mux_1196_nl, fsm_output[8]);
  assign nor_420_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_1183_nl = MUX_s_1_2_2(nor_413_cse, nor_420_nl, fsm_output[0]);
  assign nor_421_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_422_nl = ~((z_out_6_10_1[3:0]!=4'b1010) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_1182_nl = MUX_s_1_2_2(nor_421_nl, nor_422_nl, fsm_output[0]);
  assign mux_1184_nl = MUX_s_1_2_2(mux_1183_nl, mux_1182_nl, fsm_output[6]);
  assign nor_423_nl = ~((z_out_6_10_1[3:0]!=4'b1010) | (fsm_output[6]) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1185_nl = MUX_s_1_2_2(mux_1184_nl, nor_423_nl, fsm_output[1]);
  assign nand_71_nl = ~((fsm_output[3]) & mux_1185_nl);
  assign or_1276_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1010) | (~ (fsm_output[6]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[5])
      | not_tmp_134;
  assign or_1274_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_1273_nl = (z_out_6_10_1[0]) | (z_out_6_10_1[2]) | nand_260_cse_1;
  assign mux_1179_nl = MUX_s_1_2_2(or_1274_nl, or_1273_nl, fsm_output[0]);
  assign or_1270_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1010) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_1178_nl = MUX_s_1_2_2(or_1317_cse, or_1270_nl, fsm_output[0]);
  assign mux_1180_nl = MUX_s_1_2_2(mux_1179_nl, mux_1178_nl, fsm_output[6]);
  assign mux_1181_nl = MUX_s_1_2_2(or_1276_nl, mux_1180_nl, fsm_output[1]);
  assign or_1277_nl = (fsm_output[3]) | mux_1181_nl;
  assign mux_1186_nl = MUX_s_1_2_2(nand_71_nl, or_1277_nl, fsm_output[2]);
  assign nor_418_nl = ~((fsm_output[8]) | mux_1186_nl);
  assign vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1207_nl,
      nor_418_nl, fsm_output[9]);
  assign or_1366_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b1011) | (fsm_output[5]) | (fsm_output[1]);
  assign mux_1234_nl = MUX_s_1_2_2(or_tmp_1304, or_1366_nl, fsm_output[0]);
  assign or_1365_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1011) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1233_nl = MUX_s_1_2_2(or_1365_nl, or_tmp_1296, fsm_output[0]);
  assign mux_1235_nl = MUX_s_1_2_2(mux_1234_nl, mux_1233_nl, fsm_output[4]);
  assign nand_76_nl = ~((fsm_output[6]) & (~ mux_1235_nl));
  assign or_1364_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1011);
  assign mux_1236_nl = MUX_s_1_2_2(nand_76_nl, or_1364_nl, fsm_output[7]);
  assign nor_398_nl = ~((fsm_output[8]) | mux_1236_nl);
  assign and_441_nl = (COMP_LOOP_acc_20_psp_sva[2:0]==3'b101) & (fsm_output[7]) &
      (fsm_output[6]) & (fsm_output[4]) & (fsm_output[0]) & (VEC_LOOP_j_sva_9_0[0])
      & (~ (fsm_output[5])) & (fsm_output[1]);
  assign or_1359_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1011) | (fsm_output[5]) |
      (~ (fsm_output[1]));
  assign mux_1231_nl = MUX_s_1_2_2(or_1359_nl, or_tmp_1304, fsm_output[0]);
  assign nor_400_nl = ~((fsm_output[7]) | (fsm_output[6]) | (fsm_output[4]) | mux_1231_nl);
  assign mux_1232_nl = MUX_s_1_2_2(and_441_nl, nor_400_nl, fsm_output[8]);
  assign mux_1237_nl = MUX_s_1_2_2(nor_398_nl, mux_1232_nl, fsm_output[9]);
  assign nand_378_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]==3'b101) & (fsm_output[6])
      & (fsm_output[4]) & (fsm_output[0]) & (VEC_LOOP_j_sva_9_0[0]) & (~ (fsm_output[5]))
      & (fsm_output[1]));
  assign or_1354_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1011) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_1226_nl = MUX_s_1_2_2(or_1354_nl, or_tmp_1304, fsm_output[0]);
  assign or_1352_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b011)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_1225_nl = MUX_s_1_2_2(or_tmp_1302, or_1352_nl, fsm_output[0]);
  assign mux_1227_nl = MUX_s_1_2_2(mux_1226_nl, mux_1225_nl, fsm_output[4]);
  assign or_1350_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1011) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1224_nl = MUX_s_1_2_2(or_1350_nl, or_tmp_1296, fsm_output[0]);
  assign or_1351_nl = (fsm_output[4]) | mux_1224_nl;
  assign mux_1228_nl = MUX_s_1_2_2(mux_1227_nl, or_1351_nl, fsm_output[6]);
  assign mux_1229_nl = MUX_s_1_2_2(nand_378_nl, mux_1228_nl, fsm_output[7]);
  assign and_310_nl = (fsm_output[8]) & (~ mux_1229_nl);
  assign nor_401_nl = ~((fsm_output[8]) | (fsm_output[7]) | (fsm_output[6]) | (~
      (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3:0]!=4'b1011));
  assign mux_1230_nl = MUX_s_1_2_2(and_310_nl, nor_401_nl, fsm_output[9]);
  assign mux_1238_nl = MUX_s_1_2_2(mux_1237_nl, mux_1230_nl, fsm_output[3]);
  assign nand_373_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]==3'b101) & (fsm_output[4])
      & (fsm_output[0]) & (VEC_LOOP_j_sva_9_0[0]) & (~ (fsm_output[5])) & (fsm_output[1]));
  assign or_1344_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1011) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_1219_nl = MUX_s_1_2_2(or_1344_nl, or_tmp_1304, fsm_output[0]);
  assign or_1342_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_1218_nl = MUX_s_1_2_2(or_tmp_1302, or_1342_nl, fsm_output[0]);
  assign mux_1220_nl = MUX_s_1_2_2(mux_1219_nl, mux_1218_nl, fsm_output[4]);
  assign mux_1221_nl = MUX_s_1_2_2(nand_373_nl, mux_1220_nl, fsm_output[6]);
  assign or_1340_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1011) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1216_nl = MUX_s_1_2_2(or_1340_nl, or_tmp_1296, fsm_output[0]);
  assign or_1341_nl = (fsm_output[4]) | mux_1216_nl;
  assign mux_1217_nl = MUX_s_1_2_2(or_1341_nl, or_tmp_1294, fsm_output[6]);
  assign mux_1222_nl = MUX_s_1_2_2(mux_1221_nl, mux_1217_nl, fsm_output[7]);
  assign nor_402_nl = ~((fsm_output[9:8]!=2'b10) | mux_1222_nl);
  assign nand_363_nl = ~((fsm_output[4]) & (fsm_output[0]) & (COMP_LOOP_acc_11_psp_sva[2:0]==3'b101)
      & (VEC_LOOP_j_sva_9_0[0]) & (~ (fsm_output[5])) & (fsm_output[1]));
  assign or_1335_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1011) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_1212_nl = MUX_s_1_2_2(or_1335_nl, or_tmp_1304, fsm_output[0]);
  assign or_1329_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_1211_nl = MUX_s_1_2_2(or_tmp_1302, or_1329_nl, fsm_output[0]);
  assign mux_1213_nl = MUX_s_1_2_2(mux_1212_nl, mux_1211_nl, fsm_output[4]);
  assign mux_1214_nl = MUX_s_1_2_2(nand_363_nl, mux_1213_nl, fsm_output[6]);
  assign nand_74_nl = ~((fsm_output[7]) & (~ mux_1214_nl));
  assign or_1326_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1011) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1209_nl = MUX_s_1_2_2(or_1326_nl, or_tmp_1296, fsm_output[0]);
  assign or_1327_nl = (fsm_output[4]) | mux_1209_nl;
  assign mux_1210_nl = MUX_s_1_2_2(or_1327_nl, or_tmp_1294, fsm_output[6]);
  assign or_1328_nl = (fsm_output[7]) | mux_1210_nl;
  assign mux_1215_nl = MUX_s_1_2_2(nand_74_nl, or_1328_nl, fsm_output[8]);
  assign nor_403_nl = ~((fsm_output[9]) | mux_1215_nl);
  assign mux_1223_nl = MUX_s_1_2_2(nor_402_nl, nor_403_nl, fsm_output[3]);
  assign vec_rsc_0_11_i_we_d_pff = MUX_s_1_2_2(mux_1238_nl, mux_1223_nl, fsm_output[2]);
  assign nor_387_cse = ~((z_out_6_10_1[3:0]!=4'b1011) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nand_241_cse = ~((z_out_6_10_1[3:0]==4'b1011) & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4])));
  assign nand_240_nl = ~((fsm_output[0]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm &
      (COMP_LOOP_acc_1_cse_4_sva[3:0]==4'b1011) & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4])));
  assign or_1418_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | not_tmp_134;
  assign mux_1265_nl = MUX_s_1_2_2(or_1418_nl, nand_241_cse, fsm_output[0]);
  assign mux_1266_nl = MUX_s_1_2_2(nand_240_nl, mux_1265_nl, fsm_output[6]);
  assign or_1415_nl = (z_out_6_10_1[2:1]!=2'b01) | nand_264_cse;
  assign or_1413_nl = (z_out_6_10_1[3:0]!=4'b1011) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_1263_nl = MUX_s_1_2_2(or_1415_nl, or_1413_nl, fsm_output[0]);
  assign nand_369_nl = ~((VEC_LOOP_j_sva_9_0[0]) & (COMP_LOOP_acc_11_psp_sva[2:0]==3'b101)
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (~ (fsm_output[7]))
      & (fsm_output[4]));
  assign or_1410_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1011) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_1262_nl = MUX_s_1_2_2(nand_369_nl, or_1410_nl, fsm_output[0]);
  assign mux_1264_nl = MUX_s_1_2_2(mux_1263_nl, mux_1262_nl, fsm_output[6]);
  assign mux_1267_nl = MUX_s_1_2_2(mux_1266_nl, mux_1264_nl, fsm_output[1]);
  assign nor_379_nl = ~((fsm_output[3]) | mux_1267_nl);
  assign or_1408_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b1011) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_1406_nl = (z_out_6_10_1[3:0]!=4'b1011) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]);
  assign mux_1259_nl = MUX_s_1_2_2(or_1408_nl, or_1406_nl, fsm_output[0]);
  assign or_1405_nl = (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b1011) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_1260_nl = MUX_s_1_2_2(mux_1259_nl, or_1405_nl, fsm_output[6]);
  assign nor_380_nl = ~((fsm_output[1]) | mux_1260_nl);
  assign nor_381_nl = ~((~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1011) & (fsm_output[1])
      & (fsm_output[6]) & (fsm_output[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      | not_tmp_133);
  assign mux_1261_nl = MUX_s_1_2_2(nor_380_nl, nor_381_nl, fsm_output[3]);
  assign mux_1268_nl = MUX_s_1_2_2(nor_379_nl, mux_1261_nl, fsm_output[2]);
  assign nor_382_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b1011)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign nor_383_nl = ~((~((COMP_LOOP_acc_1_cse_10_sva[3:0]==4'b1011) & (fsm_output[0])
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)) | not_tmp_133);
  assign and_308_nl = (VEC_LOOP_j_sva_9_0[0]) & (COMP_LOOP_acc_17_psp_sva[2:0]==3'b101)
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4]));
  assign nor_384_nl = ~((~ (z_out_6_10_1[0])) | (z_out_6_10_1[2]) | nand_260_cse_1);
  assign mux_1255_nl = MUX_s_1_2_2(and_308_nl, nor_384_nl, fsm_output[0]);
  assign mux_1256_nl = MUX_s_1_2_2(nor_383_nl, mux_1255_nl, fsm_output[6]);
  assign and_307_nl = (fsm_output[1]) & mux_1256_nl;
  assign mux_1257_nl = MUX_s_1_2_2(nor_382_nl, and_307_nl, fsm_output[3]);
  assign nor_385_nl = ~((~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b011)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_386_nl = ~((z_out_6_10_1[3:0]!=4'b1011) | (fsm_output[5]) | not_tmp_134);
  assign mux_1252_nl = MUX_s_1_2_2(nor_385_nl, nor_386_nl, fsm_output[0]);
  assign nor_388_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_1251_nl = MUX_s_1_2_2(nor_387_cse, nor_388_nl, fsm_output[0]);
  assign mux_1253_nl = MUX_s_1_2_2(mux_1252_nl, mux_1251_nl, fsm_output[6]);
  assign nor_389_nl = ~((~ (VEC_LOOP_j_sva_9_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b101) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]));
  assign and_431_nl = (z_out_6_10_1[3:0]==4'b1011) & (fsm_output[5]) & (~ (fsm_output[7]))
      & (fsm_output[4]);
  assign mux_1249_nl = MUX_s_1_2_2(nor_389_nl, and_431_nl, fsm_output[0]);
  assign nor_391_nl = ~((z_out_6_10_1[3:0]!=4'b1011) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1250_nl = MUX_s_1_2_2(mux_1249_nl, nor_391_nl, fsm_output[6]);
  assign mux_1254_nl = MUX_s_1_2_2(mux_1253_nl, mux_1250_nl, fsm_output[1]);
  assign and_309_nl = (fsm_output[3]) & mux_1254_nl;
  assign mux_1258_nl = MUX_s_1_2_2(mux_1257_nl, and_309_nl, fsm_output[2]);
  assign mux_1269_nl = MUX_s_1_2_2(mux_1268_nl, mux_1258_nl, fsm_output[8]);
  assign nor_394_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_1245_nl = MUX_s_1_2_2(nor_387_cse, nor_394_nl, fsm_output[0]);
  assign nor_395_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_396_nl = ~((z_out_6_10_1[3:0]!=4'b1011) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_1244_nl = MUX_s_1_2_2(nor_395_nl, nor_396_nl, fsm_output[0]);
  assign mux_1246_nl = MUX_s_1_2_2(mux_1245_nl, mux_1244_nl, fsm_output[6]);
  assign nor_397_nl = ~((z_out_6_10_1[3:0]!=4'b1011) | (fsm_output[6]) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1247_nl = MUX_s_1_2_2(mux_1246_nl, nor_397_nl, fsm_output[1]);
  assign nand_77_nl = ~((fsm_output[3]) & mux_1247_nl);
  assign or_1375_nl = (~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1011) & (fsm_output[6])
      & (fsm_output[0]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & (~ (fsm_output[5]))))
      | not_tmp_134;
  assign nand_248_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]==3'b101) & (VEC_LOOP_j_sva_9_0[0])
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4])));
  assign or_1372_nl = (~ (z_out_6_10_1[0])) | (z_out_6_10_1[2]) | nand_260_cse_1;
  assign mux_1241_nl = MUX_s_1_2_2(nand_248_nl, or_1372_nl, fsm_output[0]);
  assign nand_352_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1011) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[5]) & (~ (fsm_output[7])) & (fsm_output[4]));
  assign mux_1240_nl = MUX_s_1_2_2(nand_241_cse, nand_352_nl, fsm_output[0]);
  assign mux_1242_nl = MUX_s_1_2_2(mux_1241_nl, mux_1240_nl, fsm_output[6]);
  assign mux_1243_nl = MUX_s_1_2_2(or_1375_nl, mux_1242_nl, fsm_output[1]);
  assign or_1376_nl = (fsm_output[3]) | mux_1243_nl;
  assign mux_1248_nl = MUX_s_1_2_2(nand_77_nl, or_1376_nl, fsm_output[2]);
  assign nor_392_nl = ~((fsm_output[8]) | mux_1248_nl);
  assign vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1269_nl,
      nor_392_nl, fsm_output[9]);
  assign or_1465_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b1100) | (fsm_output[5]) | (fsm_output[1]);
  assign mux_1296_nl = MUX_s_1_2_2(or_tmp_1403, or_1465_nl, fsm_output[0]);
  assign or_1464_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1100) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1295_nl = MUX_s_1_2_2(or_1464_nl, or_tmp_1395, fsm_output[0]);
  assign mux_1297_nl = MUX_s_1_2_2(mux_1296_nl, mux_1295_nl, fsm_output[4]);
  assign nand_82_nl = ~((fsm_output[6]) & (~ mux_1297_nl));
  assign or_1463_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1:0]!=2'b00) | not_tmp_289;
  assign mux_1298_nl = MUX_s_1_2_2(nand_82_nl, or_1463_nl, fsm_output[7]);
  assign nor_373_nl = ~((fsm_output[8]) | mux_1298_nl);
  assign and_436_nl = (COMP_LOOP_acc_20_psp_sva[2:0]==3'b110) & (fsm_output[7]) &
      (fsm_output[6]) & (fsm_output[4]) & (fsm_output[0]) & (~ (VEC_LOOP_j_sva_9_0[0]))
      & (~ (fsm_output[5])) & (fsm_output[1]);
  assign or_1458_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1100) | (fsm_output[5]) |
      (~ (fsm_output[1]));
  assign mux_1293_nl = MUX_s_1_2_2(or_1458_nl, or_tmp_1403, fsm_output[0]);
  assign nor_375_nl = ~((fsm_output[7]) | (fsm_output[6]) | (fsm_output[4]) | mux_1293_nl);
  assign mux_1294_nl = MUX_s_1_2_2(and_436_nl, nor_375_nl, fsm_output[8]);
  assign mux_1299_nl = MUX_s_1_2_2(nor_373_nl, mux_1294_nl, fsm_output[9]);
  assign or_1455_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b110) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign or_1453_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1100) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_1288_nl = MUX_s_1_2_2(or_1453_nl, or_tmp_1403, fsm_output[0]);
  assign or_1451_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b100)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_1287_nl = MUX_s_1_2_2(or_tmp_1401, or_1451_nl, fsm_output[0]);
  assign mux_1289_nl = MUX_s_1_2_2(mux_1288_nl, mux_1287_nl, fsm_output[4]);
  assign or_1449_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1100) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1286_nl = MUX_s_1_2_2(or_1449_nl, or_tmp_1395, fsm_output[0]);
  assign or_1450_nl = (fsm_output[4]) | mux_1286_nl;
  assign mux_1290_nl = MUX_s_1_2_2(mux_1289_nl, or_1450_nl, fsm_output[6]);
  assign mux_1291_nl = MUX_s_1_2_2(or_1455_nl, mux_1290_nl, fsm_output[7]);
  assign and_306_nl = (fsm_output[8]) & (~ mux_1291_nl);
  assign nor_376_nl = ~((fsm_output[8]) | (fsm_output[7]) | (fsm_output[6]) | (~
      (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1:0]!=2'b00)
      | not_tmp_289);
  assign mux_1292_nl = MUX_s_1_2_2(and_306_nl, nor_376_nl, fsm_output[9]);
  assign mux_1300_nl = MUX_s_1_2_2(mux_1299_nl, mux_1292_nl, fsm_output[3]);
  assign or_1445_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b110) | (~ (fsm_output[4]))
      | (~ (fsm_output[0])) | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5]) | (~ (fsm_output[1]));
  assign or_1443_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1100) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_1281_nl = MUX_s_1_2_2(or_1443_nl, or_tmp_1403, fsm_output[0]);
  assign or_1441_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_1280_nl = MUX_s_1_2_2(or_tmp_1401, or_1441_nl, fsm_output[0]);
  assign mux_1282_nl = MUX_s_1_2_2(mux_1281_nl, mux_1280_nl, fsm_output[4]);
  assign mux_1283_nl = MUX_s_1_2_2(or_1445_nl, mux_1282_nl, fsm_output[6]);
  assign or_1439_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1100) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1278_nl = MUX_s_1_2_2(or_1439_nl, or_tmp_1395, fsm_output[0]);
  assign or_1440_nl = (fsm_output[4]) | mux_1278_nl;
  assign mux_1279_nl = MUX_s_1_2_2(or_1440_nl, or_tmp_1393, fsm_output[6]);
  assign mux_1284_nl = MUX_s_1_2_2(mux_1283_nl, mux_1279_nl, fsm_output[7]);
  assign nor_377_nl = ~((fsm_output[9:8]!=2'b10) | mux_1284_nl);
  assign or_1436_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b110)
      | (VEC_LOOP_j_sva_9_0[0]) | (fsm_output[5]) | (~ (fsm_output[1]));
  assign or_1434_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1100) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_1274_nl = MUX_s_1_2_2(or_1434_nl, or_tmp_1403, fsm_output[0]);
  assign or_1428_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_1273_nl = MUX_s_1_2_2(or_tmp_1401, or_1428_nl, fsm_output[0]);
  assign mux_1275_nl = MUX_s_1_2_2(mux_1274_nl, mux_1273_nl, fsm_output[4]);
  assign mux_1276_nl = MUX_s_1_2_2(or_1436_nl, mux_1275_nl, fsm_output[6]);
  assign nand_80_nl = ~((fsm_output[7]) & (~ mux_1276_nl));
  assign or_1425_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1100) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1271_nl = MUX_s_1_2_2(or_1425_nl, or_tmp_1395, fsm_output[0]);
  assign or_1426_nl = (fsm_output[4]) | mux_1271_nl;
  assign mux_1272_nl = MUX_s_1_2_2(or_1426_nl, or_tmp_1393, fsm_output[6]);
  assign or_1427_nl = (fsm_output[7]) | mux_1272_nl;
  assign mux_1277_nl = MUX_s_1_2_2(nand_80_nl, or_1427_nl, fsm_output[8]);
  assign nor_378_nl = ~((fsm_output[9]) | mux_1277_nl);
  assign mux_1285_nl = MUX_s_1_2_2(nor_377_nl, nor_378_nl, fsm_output[3]);
  assign vec_rsc_0_12_i_we_d_pff = MUX_s_1_2_2(mux_1300_nl, mux_1285_nl, fsm_output[2]);
  assign nor_362_cse = ~((z_out_6_10_1[3:0]!=4'b1100) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign or_1515_cse = (z_out_6_10_1[3:0]!=4'b1100) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_1518_nl = (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1100) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_1517_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | not_tmp_134;
  assign mux_1327_nl = MUX_s_1_2_2(or_1517_nl, or_1515_cse, fsm_output[0]);
  assign mux_1328_nl = MUX_s_1_2_2(or_1518_nl, mux_1327_nl, fsm_output[6]);
  assign or_1514_nl = (z_out_6_10_1[3:0]!=4'b1100) | not_tmp_133;
  assign or_1512_nl = (z_out_6_10_1[3:0]!=4'b1100) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_1325_nl = MUX_s_1_2_2(or_1514_nl, or_1512_nl, fsm_output[0]);
  assign or_1511_nl = (VEC_LOOP_j_sva_9_0[0]) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b110)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_1509_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1100) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_1324_nl = MUX_s_1_2_2(or_1511_nl, or_1509_nl, fsm_output[0]);
  assign mux_1326_nl = MUX_s_1_2_2(mux_1325_nl, mux_1324_nl, fsm_output[6]);
  assign mux_1329_nl = MUX_s_1_2_2(mux_1328_nl, mux_1326_nl, fsm_output[1]);
  assign nor_353_nl = ~((fsm_output[3]) | mux_1329_nl);
  assign or_1507_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b1100) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_1505_nl = (z_out_6_10_1[3:0]!=4'b1100) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]);
  assign mux_1321_nl = MUX_s_1_2_2(or_1507_nl, or_1505_nl, fsm_output[0]);
  assign or_1504_nl = (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b1100) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_1322_nl = MUX_s_1_2_2(mux_1321_nl, or_1504_nl, fsm_output[6]);
  assign nor_354_nl = ~((fsm_output[1]) | mux_1322_nl);
  assign nor_355_nl = ~((~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1100) & (fsm_output[1])
      & (fsm_output[6]) & (fsm_output[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      | not_tmp_133);
  assign mux_1323_nl = MUX_s_1_2_2(nor_354_nl, nor_355_nl, fsm_output[3]);
  assign mux_1330_nl = MUX_s_1_2_2(nor_353_nl, mux_1323_nl, fsm_output[2]);
  assign nor_356_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b1100)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign nor_357_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1100) | (~ (fsm_output[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | not_tmp_133);
  assign nor_358_nl = ~((VEC_LOOP_j_sva_9_0[0]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b110)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_359_nl = ~((z_out_6_10_1[2:0]!=3'b100) | nand_270_cse_1);
  assign mux_1317_nl = MUX_s_1_2_2(nor_358_nl, nor_359_nl, fsm_output[0]);
  assign mux_1318_nl = MUX_s_1_2_2(nor_357_nl, mux_1317_nl, fsm_output[6]);
  assign and_304_nl = (fsm_output[1]) & mux_1318_nl;
  assign mux_1319_nl = MUX_s_1_2_2(nor_356_nl, and_304_nl, fsm_output[3]);
  assign nor_360_nl = ~((~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b100)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_361_nl = ~((z_out_6_10_1[3:0]!=4'b1100) | (fsm_output[5]) | not_tmp_134);
  assign mux_1314_nl = MUX_s_1_2_2(nor_360_nl, nor_361_nl, fsm_output[0]);
  assign nor_363_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_1313_nl = MUX_s_1_2_2(nor_362_cse, nor_363_nl, fsm_output[0]);
  assign mux_1315_nl = MUX_s_1_2_2(mux_1314_nl, mux_1313_nl, fsm_output[6]);
  assign nor_364_nl = ~((VEC_LOOP_j_sva_9_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b110) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_365_nl = ~((z_out_6_10_1[3:0]!=4'b1100) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_1311_nl = MUX_s_1_2_2(nor_364_nl, nor_365_nl, fsm_output[0]);
  assign nor_366_nl = ~((z_out_6_10_1[3:0]!=4'b1100) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1312_nl = MUX_s_1_2_2(mux_1311_nl, nor_366_nl, fsm_output[6]);
  assign mux_1316_nl = MUX_s_1_2_2(mux_1315_nl, mux_1312_nl, fsm_output[1]);
  assign and_305_nl = (fsm_output[3]) & mux_1316_nl;
  assign mux_1320_nl = MUX_s_1_2_2(mux_1319_nl, and_305_nl, fsm_output[2]);
  assign mux_1331_nl = MUX_s_1_2_2(mux_1330_nl, mux_1320_nl, fsm_output[8]);
  assign nor_369_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_1307_nl = MUX_s_1_2_2(nor_362_cse, nor_369_nl, fsm_output[0]);
  assign nor_370_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b00)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_371_nl = ~((z_out_6_10_1[3:0]!=4'b1100) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_1306_nl = MUX_s_1_2_2(nor_370_nl, nor_371_nl, fsm_output[0]);
  assign mux_1308_nl = MUX_s_1_2_2(mux_1307_nl, mux_1306_nl, fsm_output[6]);
  assign nor_372_nl = ~((z_out_6_10_1[3:0]!=4'b1100) | (fsm_output[6]) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1309_nl = MUX_s_1_2_2(mux_1308_nl, nor_372_nl, fsm_output[1]);
  assign nand_83_nl = ~((fsm_output[3]) & mux_1309_nl);
  assign or_1474_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1100) | (~ (fsm_output[6]))
      | (~ (fsm_output[0])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[5])
      | not_tmp_134;
  assign or_1472_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_sva_9_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign or_1471_nl = (z_out_6_10_1[2:0]!=3'b100) | nand_270_cse_1;
  assign mux_1303_nl = MUX_s_1_2_2(or_1472_nl, or_1471_nl, fsm_output[0]);
  assign or_1468_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1100) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_1302_nl = MUX_s_1_2_2(or_1515_cse, or_1468_nl, fsm_output[0]);
  assign mux_1304_nl = MUX_s_1_2_2(mux_1303_nl, mux_1302_nl, fsm_output[6]);
  assign mux_1305_nl = MUX_s_1_2_2(or_1474_nl, mux_1304_nl, fsm_output[1]);
  assign or_1475_nl = (fsm_output[3]) | mux_1305_nl;
  assign mux_1310_nl = MUX_s_1_2_2(nand_83_nl, or_1475_nl, fsm_output[2]);
  assign nor_367_nl = ~((fsm_output[8]) | mux_1310_nl);
  assign vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1331_nl,
      nor_367_nl, fsm_output[9]);
  assign or_1565_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b1101) | (fsm_output[1]) | (fsm_output[5]);
  assign mux_1358_nl = MUX_s_1_2_2(or_tmp_1502, or_1565_nl, fsm_output[0]);
  assign or_1564_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1101) | (fsm_output[1])
      | (~ (fsm_output[5]));
  assign mux_1357_nl = MUX_s_1_2_2(or_1564_nl, or_tmp_1493, fsm_output[0]);
  assign mux_1359_nl = MUX_s_1_2_2(mux_1358_nl, mux_1357_nl, fsm_output[4]);
  assign nor_346_nl = ~((fsm_output[9]) | (~ (fsm_output[6])) | mux_1359_nl);
  assign nand_230_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]==3'b110) & (fsm_output[4])
      & (fsm_output[0]) & (VEC_LOOP_j_sva_9_0[0]) & (fsm_output[1]) & (~ (fsm_output[5])));
  assign or_1561_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1101) | (~ (fsm_output[1]))
      | (fsm_output[5]);
  assign mux_1354_nl = MUX_s_1_2_2(or_1561_nl, or_tmp_1502, fsm_output[0]);
  assign or_1560_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (fsm_output[1]) | (~ (fsm_output[5]));
  assign mux_1353_nl = MUX_s_1_2_2(or_tmp_1500, or_1560_nl, fsm_output[0]);
  assign mux_1355_nl = MUX_s_1_2_2(mux_1354_nl, mux_1353_nl, fsm_output[4]);
  assign mux_1356_nl = MUX_s_1_2_2(nand_230_nl, mux_1355_nl, fsm_output[6]);
  assign and_302_nl = (fsm_output[9]) & (~ mux_1356_nl);
  assign mux_1360_nl = MUX_s_1_2_2(nor_346_nl, and_302_nl, fsm_output[2]);
  assign or_1557_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1101) | (~ (fsm_output[1]))
      | (fsm_output[5]);
  assign mux_1352_nl = MUX_s_1_2_2(or_1557_nl, or_tmp_1502, fsm_output[0]);
  assign nor_347_nl = ~((fsm_output[2]) | (~ (fsm_output[9])) | (fsm_output[6]) |
      (fsm_output[4]) | mux_1352_nl);
  assign mux_1361_nl = MUX_s_1_2_2(mux_1360_nl, nor_347_nl, fsm_output[8]);
  assign or_1554_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (fsm_output[1])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1]) | not_tmp_304;
  assign nand_231_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]==3'b110) & (fsm_output[6])
      & (fsm_output[4]) & (fsm_output[0]) & (VEC_LOOP_j_sva_9_0[0]) & (fsm_output[1])
      & (~ (fsm_output[5])));
  assign mux_1350_nl = MUX_s_1_2_2(or_1554_nl, nand_231_nl, fsm_output[9]);
  assign or_1550_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1101) | (fsm_output[1])
      | (~ (fsm_output[5]));
  assign mux_1348_nl = MUX_s_1_2_2(or_1550_nl, or_tmp_1493, fsm_output[0]);
  assign or_1551_nl = (fsm_output[4]) | mux_1348_nl;
  assign mux_1349_nl = MUX_s_1_2_2(or_1551_nl, or_tmp_1512, fsm_output[6]);
  assign nand_86_nl = ~((fsm_output[9]) & (~ mux_1349_nl));
  assign mux_1351_nl = MUX_s_1_2_2(mux_1350_nl, nand_86_nl, fsm_output[2]);
  assign nor_348_nl = ~((fsm_output[8]) | mux_1351_nl);
  assign mux_1362_nl = MUX_s_1_2_2(mux_1361_nl, nor_348_nl, fsm_output[7]);
  assign nor_349_nl = ~((fsm_output[2]) | (~ (fsm_output[9])) | (fsm_output[6]) |
      (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[5]) |
      (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1]) | not_tmp_304);
  assign and_303_nl = (~ (fsm_output[9])) & (COMP_LOOP_acc_14_psp_sva[2:0]==3'b110)
      & (fsm_output[6]) & (fsm_output[4]) & (fsm_output[0]) & (VEC_LOOP_j_sva_9_0[0])
      & (fsm_output[1]) & (~ (fsm_output[5]));
  assign or_1543_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1101) | (fsm_output[1])
      | (~ (fsm_output[5]));
  assign mux_1343_nl = MUX_s_1_2_2(or_1543_nl, or_tmp_1493, fsm_output[0]);
  assign or_1544_nl = (fsm_output[4]) | mux_1343_nl;
  assign mux_1344_nl = MUX_s_1_2_2(or_1544_nl, or_tmp_1512, fsm_output[6]);
  assign nor_350_nl = ~((fsm_output[9]) | mux_1344_nl);
  assign mux_1345_nl = MUX_s_1_2_2(and_303_nl, nor_350_nl, fsm_output[2]);
  assign mux_1346_nl = MUX_s_1_2_2(nor_349_nl, mux_1345_nl, fsm_output[8]);
  assign nand_232_nl = ~((fsm_output[4]) & (fsm_output[0]) & (COMP_LOOP_acc_11_psp_sva[2:0]==3'b110)
      & (VEC_LOOP_j_sva_9_0[0]) & (fsm_output[1]) & (~ (fsm_output[5])));
  assign or_1537_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1101) | (~ (fsm_output[1]))
      | (fsm_output[5]);
  assign mux_1339_nl = MUX_s_1_2_2(or_1537_nl, or_tmp_1502, fsm_output[0]);
  assign or_1536_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (fsm_output[1]) | (~ (fsm_output[5]));
  assign mux_1338_nl = MUX_s_1_2_2(or_tmp_1500, or_1536_nl, fsm_output[0]);
  assign mux_1340_nl = MUX_s_1_2_2(mux_1339_nl, mux_1338_nl, fsm_output[4]);
  assign mux_1341_nl = MUX_s_1_2_2(nand_232_nl, mux_1340_nl, fsm_output[6]);
  assign nor_351_nl = ~((~ (fsm_output[2])) | (fsm_output[9]) | mux_1341_nl);
  assign or_1532_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1101) | (~ (fsm_output[1]))
      | (fsm_output[5]);
  assign mux_1335_nl = MUX_s_1_2_2(or_1532_nl, or_tmp_1502, fsm_output[0]);
  assign or_1527_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b101)
      | (fsm_output[1]) | (~ (fsm_output[5]));
  assign mux_1334_nl = MUX_s_1_2_2(or_tmp_1500, or_1527_nl, fsm_output[0]);
  assign mux_1336_nl = MUX_s_1_2_2(mux_1335_nl, mux_1334_nl, fsm_output[4]);
  assign or_1524_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1101) | (fsm_output[1])
      | (~ (fsm_output[5]));
  assign mux_1333_nl = MUX_s_1_2_2(or_1524_nl, or_tmp_1493, fsm_output[0]);
  assign or_1525_nl = (fsm_output[4]) | mux_1333_nl;
  assign mux_1337_nl = MUX_s_1_2_2(mux_1336_nl, or_1525_nl, fsm_output[6]);
  assign nor_352_nl = ~((fsm_output[2]) | (fsm_output[9]) | mux_1337_nl);
  assign mux_1342_nl = MUX_s_1_2_2(nor_351_nl, nor_352_nl, fsm_output[8]);
  assign mux_1347_nl = MUX_s_1_2_2(mux_1346_nl, mux_1342_nl, fsm_output[7]);
  assign vec_rsc_0_13_i_we_d_pff = MUX_s_1_2_2(mux_1362_nl, mux_1347_nl, fsm_output[3]);
  assign nor_335_cse = ~((z_out_6_10_1[3:0]!=4'b1101) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nand_217_cse = ~((z_out_6_10_1[3:0]==4'b1101) & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4])));
  assign nand_216_nl = ~((fsm_output[0]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm &
      (COMP_LOOP_acc_1_cse_4_sva[3:0]==4'b1101) & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4])));
  assign or_1615_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | not_tmp_134;
  assign mux_1389_nl = MUX_s_1_2_2(or_1615_nl, nand_217_cse, fsm_output[0]);
  assign mux_1390_nl = MUX_s_1_2_2(nand_216_nl, mux_1389_nl, fsm_output[6]);
  assign or_1612_nl = (z_out_6_10_1[1]) | (~((z_out_6_10_1[2]) & (z_out_6_10_1[3])
      & (z_out_6_10_1[0]) & (fsm_output[5]) & (fsm_output[7]) & (fsm_output[4])));
  assign or_1611_nl = (z_out_6_10_1[3:0]!=4'b1101) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_1387_nl = MUX_s_1_2_2(or_1612_nl, or_1611_nl, fsm_output[0]);
  assign nand_368_nl = ~((VEC_LOOP_j_sva_9_0[0]) & (COMP_LOOP_acc_11_psp_sva[2:0]==3'b110)
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (~ (fsm_output[7]))
      & (fsm_output[4]));
  assign or_1608_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1101) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_1386_nl = MUX_s_1_2_2(nand_368_nl, or_1608_nl, fsm_output[0]);
  assign mux_1388_nl = MUX_s_1_2_2(mux_1387_nl, mux_1386_nl, fsm_output[6]);
  assign mux_1391_nl = MUX_s_1_2_2(mux_1390_nl, mux_1388_nl, fsm_output[1]);
  assign nor_327_nl = ~((fsm_output[3]) | mux_1391_nl);
  assign or_1606_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b1101) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_1604_nl = (z_out_6_10_1[3:0]!=4'b1101) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]);
  assign mux_1383_nl = MUX_s_1_2_2(or_1606_nl, or_1604_nl, fsm_output[0]);
  assign or_1603_nl = (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b1101) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_1384_nl = MUX_s_1_2_2(mux_1383_nl, or_1603_nl, fsm_output[6]);
  assign nor_328_nl = ~((fsm_output[1]) | mux_1384_nl);
  assign nor_329_nl = ~((~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1101) & (fsm_output[1])
      & (fsm_output[6]) & (fsm_output[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      | not_tmp_133);
  assign mux_1385_nl = MUX_s_1_2_2(nor_328_nl, nor_329_nl, fsm_output[3]);
  assign mux_1392_nl = MUX_s_1_2_2(nor_327_nl, mux_1385_nl, fsm_output[2]);
  assign nor_330_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b1101)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign nor_331_nl = ~((~((COMP_LOOP_acc_1_cse_10_sva[3:0]==4'b1101) & (fsm_output[0])
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)) | not_tmp_133);
  assign and_300_nl = (VEC_LOOP_j_sva_9_0[0]) & (COMP_LOOP_acc_17_psp_sva[2:0]==3'b110)
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4]));
  assign nor_332_nl = ~((z_out_6_10_1[2:0]!=3'b101) | nand_270_cse_1);
  assign mux_1379_nl = MUX_s_1_2_2(and_300_nl, nor_332_nl, fsm_output[0]);
  assign mux_1380_nl = MUX_s_1_2_2(nor_331_nl, mux_1379_nl, fsm_output[6]);
  assign and_299_nl = (fsm_output[1]) & mux_1380_nl;
  assign mux_1381_nl = MUX_s_1_2_2(nor_330_nl, and_299_nl, fsm_output[3]);
  assign nor_333_nl = ~((~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b101)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_334_nl = ~((z_out_6_10_1[3:0]!=4'b1101) | (fsm_output[5]) | not_tmp_134);
  assign mux_1376_nl = MUX_s_1_2_2(nor_333_nl, nor_334_nl, fsm_output[0]);
  assign nor_336_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_1375_nl = MUX_s_1_2_2(nor_335_cse, nor_336_nl, fsm_output[0]);
  assign mux_1377_nl = MUX_s_1_2_2(mux_1376_nl, mux_1375_nl, fsm_output[6]);
  assign nor_337_nl = ~((~ (VEC_LOOP_j_sva_9_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b110) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]));
  assign and_430_nl = (z_out_6_10_1[3:0]==4'b1101) & (fsm_output[5]) & (~ (fsm_output[7]))
      & (fsm_output[4]);
  assign mux_1373_nl = MUX_s_1_2_2(nor_337_nl, and_430_nl, fsm_output[0]);
  assign nor_339_nl = ~((z_out_6_10_1[3:0]!=4'b1101) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1374_nl = MUX_s_1_2_2(mux_1373_nl, nor_339_nl, fsm_output[6]);
  assign mux_1378_nl = MUX_s_1_2_2(mux_1377_nl, mux_1374_nl, fsm_output[1]);
  assign and_301_nl = (fsm_output[3]) & mux_1378_nl;
  assign mux_1382_nl = MUX_s_1_2_2(mux_1381_nl, and_301_nl, fsm_output[2]);
  assign mux_1393_nl = MUX_s_1_2_2(mux_1392_nl, mux_1382_nl, fsm_output[8]);
  assign nor_342_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_1369_nl = MUX_s_1_2_2(nor_335_cse, nor_342_nl, fsm_output[0]);
  assign nor_343_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b01)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_344_nl = ~((z_out_6_10_1[3:0]!=4'b1101) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_1368_nl = MUX_s_1_2_2(nor_343_nl, nor_344_nl, fsm_output[0]);
  assign mux_1370_nl = MUX_s_1_2_2(mux_1369_nl, mux_1368_nl, fsm_output[6]);
  assign nor_345_nl = ~((z_out_6_10_1[3:0]!=4'b1101) | (fsm_output[6]) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1371_nl = MUX_s_1_2_2(mux_1370_nl, nor_345_nl, fsm_output[1]);
  assign nand_89_nl = ~((fsm_output[3]) & mux_1371_nl);
  assign or_1573_nl = (~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1101) & (fsm_output[6])
      & (fsm_output[0]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & (~ (fsm_output[5]))))
      | not_tmp_134;
  assign nand_224_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]==3'b110) & (VEC_LOOP_j_sva_9_0[0])
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4])));
  assign or_1570_nl = (z_out_6_10_1[2:0]!=3'b101) | nand_270_cse_1;
  assign mux_1365_nl = MUX_s_1_2_2(nand_224_nl, or_1570_nl, fsm_output[0]);
  assign nand_351_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1101) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[5]) & (~ (fsm_output[7])) & (fsm_output[4]));
  assign mux_1364_nl = MUX_s_1_2_2(nand_217_cse, nand_351_nl, fsm_output[0]);
  assign mux_1366_nl = MUX_s_1_2_2(mux_1365_nl, mux_1364_nl, fsm_output[6]);
  assign mux_1367_nl = MUX_s_1_2_2(or_1573_nl, mux_1366_nl, fsm_output[1]);
  assign or_1574_nl = (fsm_output[3]) | mux_1367_nl;
  assign mux_1372_nl = MUX_s_1_2_2(nand_89_nl, or_1574_nl, fsm_output[2]);
  assign nor_340_nl = ~((fsm_output[8]) | mux_1372_nl);
  assign vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1393_nl,
      nor_340_nl, fsm_output[9]);
  assign or_1662_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b1110) | (fsm_output[5]) | (fsm_output[1]);
  assign mux_1420_nl = MUX_s_1_2_2(or_tmp_1600, or_1662_nl, fsm_output[0]);
  assign or_1661_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1110) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1419_nl = MUX_s_1_2_2(or_1661_nl, or_tmp_1592, fsm_output[0]);
  assign mux_1421_nl = MUX_s_1_2_2(mux_1420_nl, mux_1419_nl, fsm_output[4]);
  assign nand_94_nl = ~((fsm_output[6]) & (~ mux_1421_nl));
  assign or_1660_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1:0]!=2'b10) | not_tmp_289;
  assign mux_1422_nl = MUX_s_1_2_2(nand_94_nl, or_1660_nl, fsm_output[7]);
  assign nor_321_nl = ~((fsm_output[8]) | mux_1422_nl);
  assign and_435_nl = (COMP_LOOP_acc_20_psp_sva[2:0]==3'b111) & (fsm_output[7]) &
      (fsm_output[6]) & (fsm_output[4]) & (fsm_output[0]) & (~ (VEC_LOOP_j_sva_9_0[0]))
      & (~ (fsm_output[5])) & (fsm_output[1]);
  assign or_1655_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1110) | (fsm_output[5]) |
      (~ (fsm_output[1]));
  assign mux_1417_nl = MUX_s_1_2_2(or_1655_nl, or_tmp_1600, fsm_output[0]);
  assign nor_323_nl = ~((fsm_output[7]) | (fsm_output[6]) | (fsm_output[4]) | mux_1417_nl);
  assign mux_1418_nl = MUX_s_1_2_2(and_435_nl, nor_323_nl, fsm_output[8]);
  assign mux_1423_nl = MUX_s_1_2_2(nor_321_nl, mux_1418_nl, fsm_output[9]);
  assign nand_375_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]==3'b111) & (fsm_output[6])
      & (fsm_output[4]) & (fsm_output[0]) & (~ (VEC_LOOP_j_sva_9_0[0])) & (~ (fsm_output[5]))
      & (fsm_output[1]));
  assign or_1650_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1110) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_1412_nl = MUX_s_1_2_2(or_1650_nl, or_tmp_1600, fsm_output[0]);
  assign or_1648_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b110)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_1411_nl = MUX_s_1_2_2(or_tmp_1598, or_1648_nl, fsm_output[0]);
  assign mux_1413_nl = MUX_s_1_2_2(mux_1412_nl, mux_1411_nl, fsm_output[4]);
  assign or_1646_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1110) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1410_nl = MUX_s_1_2_2(or_1646_nl, or_tmp_1592, fsm_output[0]);
  assign or_1647_nl = (fsm_output[4]) | mux_1410_nl;
  assign mux_1414_nl = MUX_s_1_2_2(mux_1413_nl, or_1647_nl, fsm_output[6]);
  assign mux_1415_nl = MUX_s_1_2_2(nand_375_nl, mux_1414_nl, fsm_output[7]);
  assign and_298_nl = (fsm_output[8]) & (~ mux_1415_nl);
  assign nor_324_nl = ~((fsm_output[8]) | (fsm_output[7]) | (fsm_output[6]) | (~
      (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1]) | (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1:0]!=2'b10)
      | not_tmp_289);
  assign mux_1416_nl = MUX_s_1_2_2(and_298_nl, nor_324_nl, fsm_output[9]);
  assign mux_1424_nl = MUX_s_1_2_2(mux_1423_nl, mux_1416_nl, fsm_output[3]);
  assign nand_367_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]==3'b111) & (fsm_output[4])
      & (fsm_output[0]) & (~ (VEC_LOOP_j_sva_9_0[0])) & (~ (fsm_output[5])) & (fsm_output[1]));
  assign or_1640_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1110) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_1405_nl = MUX_s_1_2_2(or_1640_nl, or_tmp_1600, fsm_output[0]);
  assign or_1638_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_1404_nl = MUX_s_1_2_2(or_tmp_1598, or_1638_nl, fsm_output[0]);
  assign mux_1406_nl = MUX_s_1_2_2(mux_1405_nl, mux_1404_nl, fsm_output[4]);
  assign mux_1407_nl = MUX_s_1_2_2(nand_367_nl, mux_1406_nl, fsm_output[6]);
  assign or_1636_nl = (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1110) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1402_nl = MUX_s_1_2_2(or_1636_nl, or_tmp_1592, fsm_output[0]);
  assign or_1637_nl = (fsm_output[4]) | mux_1402_nl;
  assign mux_1403_nl = MUX_s_1_2_2(or_1637_nl, or_tmp_1590, fsm_output[6]);
  assign mux_1408_nl = MUX_s_1_2_2(mux_1407_nl, mux_1403_nl, fsm_output[7]);
  assign nor_325_nl = ~((fsm_output[9:8]!=2'b10) | mux_1408_nl);
  assign nand_359_nl = ~((fsm_output[4]) & (fsm_output[0]) & (COMP_LOOP_acc_11_psp_sva[2:0]==3'b111)
      & (~ (VEC_LOOP_j_sva_9_0[0])) & (~ (fsm_output[5])) & (fsm_output[1]));
  assign or_1631_nl = (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1110) | (fsm_output[5])
      | (~ (fsm_output[1]));
  assign mux_1398_nl = MUX_s_1_2_2(or_1631_nl, or_tmp_1600, fsm_output[0]);
  assign or_1625_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_1397_nl = MUX_s_1_2_2(or_tmp_1598, or_1625_nl, fsm_output[0]);
  assign mux_1399_nl = MUX_s_1_2_2(mux_1398_nl, mux_1397_nl, fsm_output[4]);
  assign mux_1400_nl = MUX_s_1_2_2(nand_359_nl, mux_1399_nl, fsm_output[6]);
  assign nand_92_nl = ~((fsm_output[7]) & (~ mux_1400_nl));
  assign or_1622_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1110) | (~ (fsm_output[5]))
      | (fsm_output[1]);
  assign mux_1395_nl = MUX_s_1_2_2(or_1622_nl, or_tmp_1592, fsm_output[0]);
  assign or_1623_nl = (fsm_output[4]) | mux_1395_nl;
  assign mux_1396_nl = MUX_s_1_2_2(or_1623_nl, or_tmp_1590, fsm_output[6]);
  assign or_1624_nl = (fsm_output[7]) | mux_1396_nl;
  assign mux_1401_nl = MUX_s_1_2_2(nand_92_nl, or_1624_nl, fsm_output[8]);
  assign nor_326_nl = ~((fsm_output[9]) | mux_1401_nl);
  assign mux_1409_nl = MUX_s_1_2_2(nor_325_nl, nor_326_nl, fsm_output[3]);
  assign vec_rsc_0_14_i_we_d_pff = MUX_s_1_2_2(mux_1424_nl, mux_1409_nl, fsm_output[2]);
  assign nor_310_cse = ~((z_out_6_10_1[3:0]!=4'b1110) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nand_202_cse = ~((z_out_6_10_1[3:1]==3'b111) & (fsm_output[5]) & (fsm_output[7])
      & (fsm_output[4]));
  assign nand_197_cse = ~((z_out_6_10_1[3:0]==4'b1110) & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4])));
  assign nand_196_nl = ~((fsm_output[0]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm &
      (COMP_LOOP_acc_1_cse_4_sva[3:0]==4'b1110) & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4])));
  assign or_1712_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | not_tmp_134;
  assign mux_1451_nl = MUX_s_1_2_2(or_1712_nl, nand_197_cse, fsm_output[0]);
  assign mux_1452_nl = MUX_s_1_2_2(nand_196_nl, mux_1451_nl, fsm_output[6]);
  assign or_1709_nl = (~((z_out_6_10_1[3:0]==4'b1110))) | not_tmp_133;
  assign or_1707_nl = (z_out_6_10_1[3:0]!=4'b1110) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]);
  assign mux_1449_nl = MUX_s_1_2_2(or_1709_nl, or_1707_nl, fsm_output[0]);
  assign nand_366_nl = ~((~ (VEC_LOOP_j_sva_9_0[0])) & (COMP_LOOP_acc_11_psp_sva[2:0]==3'b111)
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (~ (fsm_output[7]))
      & (fsm_output[4]));
  assign or_1704_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1110) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_1448_nl = MUX_s_1_2_2(nand_366_nl, or_1704_nl, fsm_output[0]);
  assign mux_1450_nl = MUX_s_1_2_2(mux_1449_nl, mux_1448_nl, fsm_output[6]);
  assign mux_1453_nl = MUX_s_1_2_2(mux_1452_nl, mux_1450_nl, fsm_output[1]);
  assign nor_302_nl = ~((fsm_output[3]) | mux_1453_nl);
  assign or_1702_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b1110) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign or_1700_nl = (z_out_6_10_1[3:0]!=4'b1110) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]);
  assign mux_1445_nl = MUX_s_1_2_2(or_1702_nl, or_1700_nl, fsm_output[0]);
  assign or_1699_nl = (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b1110) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_1446_nl = MUX_s_1_2_2(mux_1445_nl, or_1699_nl, fsm_output[6]);
  assign nor_303_nl = ~((fsm_output[1]) | mux_1446_nl);
  assign nor_304_nl = ~((~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1110) & (fsm_output[1])
      & (fsm_output[6]) & (fsm_output[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      | not_tmp_133);
  assign mux_1447_nl = MUX_s_1_2_2(nor_303_nl, nor_304_nl, fsm_output[3]);
  assign mux_1454_nl = MUX_s_1_2_2(nor_302_nl, mux_1447_nl, fsm_output[2]);
  assign nor_305_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b1110)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign nor_306_nl = ~((~((COMP_LOOP_acc_1_cse_10_sva[3:0]==4'b1110) & (fsm_output[0])
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)) | not_tmp_133);
  assign and_296_nl = (~ (VEC_LOOP_j_sva_9_0[0])) & (COMP_LOOP_acc_17_psp_sva[2:0]==3'b111)
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4]));
  assign nor_307_nl = ~((z_out_6_10_1[0]) | nand_202_cse);
  assign mux_1441_nl = MUX_s_1_2_2(and_296_nl, nor_307_nl, fsm_output[0]);
  assign mux_1442_nl = MUX_s_1_2_2(nor_306_nl, mux_1441_nl, fsm_output[6]);
  assign and_295_nl = (fsm_output[1]) & mux_1442_nl;
  assign mux_1443_nl = MUX_s_1_2_2(nor_305_nl, and_295_nl, fsm_output[3]);
  assign nor_308_nl = ~((~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_9_0[2:0]!=3'b110)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[4]));
  assign nor_309_nl = ~((z_out_6_10_1[3:0]!=4'b1110) | (fsm_output[5]) | not_tmp_134);
  assign mux_1438_nl = MUX_s_1_2_2(nor_308_nl, nor_309_nl, fsm_output[0]);
  assign nor_311_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_1437_nl = MUX_s_1_2_2(nor_310_cse, nor_311_nl, fsm_output[0]);
  assign mux_1439_nl = MUX_s_1_2_2(mux_1438_nl, mux_1437_nl, fsm_output[6]);
  assign nor_312_nl = ~((VEC_LOOP_j_sva_9_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b111) | (~ (fsm_output[5])) | (fsm_output[7])
      | (fsm_output[4]));
  assign and_429_nl = (z_out_6_10_1[3:0]==4'b1110) & (fsm_output[5]) & (~ (fsm_output[7]))
      & (fsm_output[4]);
  assign mux_1435_nl = MUX_s_1_2_2(nor_312_nl, and_429_nl, fsm_output[0]);
  assign nor_314_nl = ~((z_out_6_10_1[3:0]!=4'b1110) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1436_nl = MUX_s_1_2_2(mux_1435_nl, nor_314_nl, fsm_output[6]);
  assign mux_1440_nl = MUX_s_1_2_2(mux_1439_nl, mux_1436_nl, fsm_output[1]);
  assign and_297_nl = (fsm_output[3]) & mux_1440_nl;
  assign mux_1444_nl = MUX_s_1_2_2(mux_1443_nl, and_297_nl, fsm_output[2]);
  assign mux_1455_nl = MUX_s_1_2_2(mux_1454_nl, mux_1444_nl, fsm_output[8]);
  assign nor_317_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_1431_nl = MUX_s_1_2_2(nor_310_cse, nor_317_nl, fsm_output[0]);
  assign nor_318_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b10)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[4]));
  assign nor_319_nl = ~((z_out_6_10_1[3:0]!=4'b1110) | (fsm_output[5]) | (fsm_output[7])
      | (~ (fsm_output[4])));
  assign mux_1430_nl = MUX_s_1_2_2(nor_318_nl, nor_319_nl, fsm_output[0]);
  assign mux_1432_nl = MUX_s_1_2_2(mux_1431_nl, mux_1430_nl, fsm_output[6]);
  assign nor_320_nl = ~((z_out_6_10_1[3:0]!=4'b1110) | (fsm_output[6]) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1433_nl = MUX_s_1_2_2(mux_1432_nl, nor_320_nl, fsm_output[1]);
  assign nand_95_nl = ~((fsm_output[3]) & mux_1433_nl);
  assign or_1670_nl = (~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1110) & (fsm_output[6])
      & (fsm_output[0]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & (~ (fsm_output[5]))))
      | not_tmp_134;
  assign nand_204_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]==3'b111) & (~ (VEC_LOOP_j_sva_9_0[0]))
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4])));
  assign or_1667_nl = (z_out_6_10_1[0]) | nand_202_cse;
  assign mux_1427_nl = MUX_s_1_2_2(nand_204_nl, or_1667_nl, fsm_output[0]);
  assign nand_350_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1110) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[5]) & (~ (fsm_output[7])) & (fsm_output[4]));
  assign mux_1426_nl = MUX_s_1_2_2(nand_197_cse, nand_350_nl, fsm_output[0]);
  assign mux_1428_nl = MUX_s_1_2_2(mux_1427_nl, mux_1426_nl, fsm_output[6]);
  assign mux_1429_nl = MUX_s_1_2_2(or_1670_nl, mux_1428_nl, fsm_output[1]);
  assign or_1671_nl = (fsm_output[3]) | mux_1429_nl;
  assign mux_1434_nl = MUX_s_1_2_2(nand_95_nl, or_1671_nl, fsm_output[2]);
  assign nor_315_nl = ~((fsm_output[8]) | mux_1434_nl);
  assign vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1455_nl,
      nor_315_nl, fsm_output[9]);
  assign or_1756_nl = (VEC_LOOP_j_sva_9_0[3:0]!=4'b1111) | (fsm_output[5]) | (fsm_output[1]);
  assign mux_1482_nl = MUX_s_1_2_2(or_tmp_1694, or_1756_nl, fsm_output[0]);
  assign nand_178_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]==4'b1111) & (fsm_output[5])
      & (~ (fsm_output[1])));
  assign mux_1481_nl = MUX_s_1_2_2(nand_178_nl, or_tmp_1689, fsm_output[0]);
  assign mux_1483_nl = MUX_s_1_2_2(mux_1482_nl, mux_1481_nl, fsm_output[4]);
  assign nand_100_nl = ~((fsm_output[6]) & (~ mux_1483_nl));
  assign or_1754_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[1]) | not_tmp_335;
  assign mux_1484_nl = MUX_s_1_2_2(nand_100_nl, or_1754_nl, fsm_output[7]);
  assign nor_296_nl = ~((fsm_output[8]) | mux_1484_nl);
  assign and_434_nl = (COMP_LOOP_acc_20_psp_sva[2:0]==3'b111) & (fsm_output[7]) &
      (fsm_output[6]) & (fsm_output[4]) & (fsm_output[0]) & (VEC_LOOP_j_sva_9_0[0])
      & (~ (fsm_output[5])) & (fsm_output[1]);
  assign nand_377_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1111) & (~ (fsm_output[5]))
      & (fsm_output[1]));
  assign mux_1479_nl = MUX_s_1_2_2(nand_377_nl, or_tmp_1694, fsm_output[0]);
  assign nor_298_nl = ~((fsm_output[7]) | (fsm_output[6]) | (fsm_output[4]) | mux_1479_nl);
  assign mux_1480_nl = MUX_s_1_2_2(and_434_nl, nor_298_nl, fsm_output[8]);
  assign mux_1485_nl = MUX_s_1_2_2(nor_296_nl, mux_1480_nl, fsm_output[9]);
  assign nand_374_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]==3'b111) & (fsm_output[6])
      & (fsm_output[4]) & (fsm_output[0]) & (VEC_LOOP_j_sva_9_0[0]) & (~ (fsm_output[5]))
      & (fsm_output[1]));
  assign nand_372_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b1111) & (~ (fsm_output[5]))
      & (fsm_output[1]));
  assign mux_1474_nl = MUX_s_1_2_2(nand_372_nl, or_tmp_1694, fsm_output[0]);
  assign nand_183_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) & (VEC_LOOP_j_sva_9_0[2:0]==3'b111)
      & (fsm_output[5]) & (~ (fsm_output[1])));
  assign mux_1473_nl = MUX_s_1_2_2(not_tmp_336, nand_183_nl, fsm_output[0]);
  assign mux_1475_nl = MUX_s_1_2_2(mux_1474_nl, mux_1473_nl, fsm_output[4]);
  assign nand_184_nl = ~((COMP_LOOP_acc_1_cse_10_sva[3:0]==4'b1111) & (fsm_output[5])
      & (~ (fsm_output[1])));
  assign mux_1472_nl = MUX_s_1_2_2(nand_184_nl, or_tmp_1689, fsm_output[0]);
  assign or_1741_nl = (fsm_output[4]) | mux_1472_nl;
  assign mux_1476_nl = MUX_s_1_2_2(mux_1475_nl, or_1741_nl, fsm_output[6]);
  assign mux_1477_nl = MUX_s_1_2_2(nand_374_nl, mux_1476_nl, fsm_output[7]);
  assign and_294_nl = (fsm_output[8]) & (~ mux_1477_nl);
  assign nor_299_nl = ~((fsm_output[8]) | (fsm_output[7]) | (fsm_output[6]) | (~
      (fsm_output[4])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[1]) | not_tmp_335);
  assign mux_1478_nl = MUX_s_1_2_2(and_294_nl, nor_299_nl, fsm_output[9]);
  assign mux_1486_nl = MUX_s_1_2_2(mux_1485_nl, mux_1478_nl, fsm_output[3]);
  assign nand_365_nl = ~((COMP_LOOP_acc_17_psp_sva[2:0]==3'b111) & (fsm_output[4])
      & (fsm_output[0]) & (VEC_LOOP_j_sva_9_0[0]) & (~ (fsm_output[5])) & (fsm_output[1]));
  assign nand_362_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b1111) & (~ (fsm_output[5]))
      & (fsm_output[1]));
  assign mux_1467_nl = MUX_s_1_2_2(nand_362_nl, or_tmp_1694, fsm_output[0]);
  assign nand_187_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]==2'b11) & (VEC_LOOP_j_sva_9_0[1:0]==2'b11)
      & (fsm_output[5]) & (~ (fsm_output[1])));
  assign mux_1466_nl = MUX_s_1_2_2(not_tmp_336, nand_187_nl, fsm_output[0]);
  assign mux_1468_nl = MUX_s_1_2_2(mux_1467_nl, mux_1466_nl, fsm_output[4]);
  assign mux_1469_nl = MUX_s_1_2_2(nand_365_nl, mux_1468_nl, fsm_output[6]);
  assign nand_188_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1111) & (fsm_output[5])
      & (~ (fsm_output[1])));
  assign mux_1464_nl = MUX_s_1_2_2(nand_188_nl, or_tmp_1689, fsm_output[0]);
  assign or_1731_nl = (fsm_output[4]) | mux_1464_nl;
  assign mux_1465_nl = MUX_s_1_2_2(or_1731_nl, or_tmp_1687, fsm_output[6]);
  assign mux_1470_nl = MUX_s_1_2_2(mux_1469_nl, mux_1465_nl, fsm_output[7]);
  assign nor_300_nl = ~((fsm_output[9:8]!=2'b10) | mux_1470_nl);
  assign nand_358_nl = ~((fsm_output[4]) & (fsm_output[0]) & (COMP_LOOP_acc_11_psp_sva[2:0]==3'b111)
      & (VEC_LOOP_j_sva_9_0[0]) & (~ (fsm_output[5])) & (fsm_output[1]));
  assign nand_349_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]==4'b1111) & (~ (fsm_output[5]))
      & (fsm_output[1]));
  assign mux_1460_nl = MUX_s_1_2_2(nand_349_nl, or_tmp_1694, fsm_output[0]);
  assign nand_191_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]==2'b11) & (VEC_LOOP_j_sva_9_0[1:0]==2'b11)
      & (fsm_output[5]) & (~ (fsm_output[1])));
  assign mux_1459_nl = MUX_s_1_2_2(not_tmp_336, nand_191_nl, fsm_output[0]);
  assign mux_1461_nl = MUX_s_1_2_2(mux_1460_nl, mux_1459_nl, fsm_output[4]);
  assign mux_1462_nl = MUX_s_1_2_2(nand_358_nl, mux_1461_nl, fsm_output[6]);
  assign nand_98_nl = ~((fsm_output[7]) & (~ mux_1462_nl));
  assign nand_192_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1111) & (fsm_output[5])
      & (~ (fsm_output[1])));
  assign mux_1457_nl = MUX_s_1_2_2(nand_192_nl, or_tmp_1689, fsm_output[0]);
  assign or_1720_nl = (fsm_output[4]) | mux_1457_nl;
  assign mux_1458_nl = MUX_s_1_2_2(or_1720_nl, or_tmp_1687, fsm_output[6]);
  assign or_1721_nl = (fsm_output[7]) | mux_1458_nl;
  assign mux_1463_nl = MUX_s_1_2_2(nand_98_nl, or_1721_nl, fsm_output[8]);
  assign nor_301_nl = ~((fsm_output[9]) | mux_1463_nl);
  assign mux_1471_nl = MUX_s_1_2_2(nor_300_nl, nor_301_nl, fsm_output[3]);
  assign vec_rsc_0_15_i_we_d_pff = MUX_s_1_2_2(mux_1486_nl, mux_1471_nl, fsm_output[2]);
  assign and_291_cse = (z_out_6_10_1[3:0]==4'b1111) & (~ (fsm_output[5])) & (fsm_output[7])
      & (~ (fsm_output[4]));
  assign nand_161_cse = ~((z_out_6_10_1[3:0]==4'b1111) & (fsm_output[5]) & (fsm_output[7])
      & (fsm_output[4]));
  assign nand_160_cse = ~((z_out_6_10_1[3:0]==4'b1111) & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4])));
  assign nand_158_nl = ~((fsm_output[0]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm &
      (COMP_LOOP_acc_1_cse_4_sva[3:0]==4'b1111) & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4])));
  assign or_1802_nl = (~((COMP_LOOP_acc_13_psp_sva[1:0]==2'b11) & (VEC_LOOP_j_sva_9_0[1:0]==2'b11)
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (~ (fsm_output[5])))) | not_tmp_134;
  assign mux_1513_nl = MUX_s_1_2_2(or_1802_nl, nand_160_cse, fsm_output[0]);
  assign mux_1514_nl = MUX_s_1_2_2(nand_158_nl, mux_1513_nl, fsm_output[6]);
  assign nand_162_nl = ~((z_out_6_10_1[3:0]==4'b1111) & (~ (fsm_output[5])) & (fsm_output[7])
      & (~ (fsm_output[4])));
  assign mux_1511_nl = MUX_s_1_2_2(nand_161_cse, nand_162_nl, fsm_output[0]);
  assign nand_364_nl = ~((VEC_LOOP_j_sva_9_0[0]) & (COMP_LOOP_acc_11_psp_sva[2:0]==3'b111)
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (~ (fsm_output[7]))
      & (fsm_output[4]));
  assign or_1796_nl = (COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1111) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_1510_nl = MUX_s_1_2_2(nand_364_nl, or_1796_nl, fsm_output[0]);
  assign mux_1512_nl = MUX_s_1_2_2(mux_1511_nl, mux_1510_nl, fsm_output[6]);
  assign mux_1515_nl = MUX_s_1_2_2(mux_1514_nl, mux_1512_nl, fsm_output[1]);
  assign nor_282_nl = ~((fsm_output[3]) | mux_1515_nl);
  assign nand_361_nl = ~((VEC_LOOP_j_sva_9_0[3:0]==4'b1111) & (~ (fsm_output[5]))
      & (~ (fsm_output[7])) & (fsm_output[4]));
  assign nand_164_nl = ~((z_out_6_10_1[3:0]==4'b1111) & (fsm_output[5]) & (~ (fsm_output[7]))
      & (~ (fsm_output[4])));
  assign mux_1507_nl = MUX_s_1_2_2(nand_361_nl, nand_164_nl, fsm_output[0]);
  assign or_1791_nl = (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b1111) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_1508_nl = MUX_s_1_2_2(mux_1507_nl, or_1791_nl, fsm_output[6]);
  assign nor_283_nl = ~((fsm_output[1]) | mux_1508_nl);
  assign nor_284_nl = ~((~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1111) & (fsm_output[1])
      & (fsm_output[6]) & (fsm_output[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      | not_tmp_133);
  assign mux_1509_nl = MUX_s_1_2_2(nor_283_nl, nor_284_nl, fsm_output[3]);
  assign mux_1516_nl = MUX_s_1_2_2(nor_282_nl, mux_1509_nl, fsm_output[2]);
  assign nor_285_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[0]) | (z_out_6_10_1[3:0]!=4'b1111)
      | (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[4])));
  assign nor_286_nl = ~((~((COMP_LOOP_acc_1_cse_10_sva[3:0]==4'b1111) & (fsm_output[0])
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)) | not_tmp_133);
  assign and_287_nl = (VEC_LOOP_j_sva_9_0[0]) & (COMP_LOOP_acc_17_psp_sva[2:0]==3'b111)
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4]));
  assign and_288_nl = (z_out_6_10_1[3:0]==4'b1111) & (fsm_output[5]) & (fsm_output[7])
      & (fsm_output[4]);
  assign mux_1503_nl = MUX_s_1_2_2(and_287_nl, and_288_nl, fsm_output[0]);
  assign mux_1504_nl = MUX_s_1_2_2(nor_286_nl, mux_1503_nl, fsm_output[6]);
  assign and_286_nl = (fsm_output[1]) & mux_1504_nl;
  assign mux_1505_nl = MUX_s_1_2_2(nor_285_nl, and_286_nl, fsm_output[3]);
  assign and_290_nl = (COMP_LOOP_acc_16_psp_sva[0]) & (VEC_LOOP_j_sva_9_0[2:0]==3'b111)
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (~ (fsm_output[5])) & (fsm_output[7])
      & (~ (fsm_output[4]));
  assign nor_287_nl = ~((~((z_out_6_10_1[3:0]==4'b1111) & (~ (fsm_output[5])))) |
      not_tmp_134);
  assign mux_1500_nl = MUX_s_1_2_2(and_290_nl, nor_287_nl, fsm_output[0]);
  assign and_427_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b1111) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      & (~ (fsm_output[5])) & (~ (fsm_output[7])) & (fsm_output[4]);
  assign mux_1499_nl = MUX_s_1_2_2(and_291_cse, and_427_nl, fsm_output[0]);
  assign mux_1501_nl = MUX_s_1_2_2(mux_1500_nl, mux_1499_nl, fsm_output[6]);
  assign and_292_nl = (VEC_LOOP_j_sva_9_0[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (COMP_LOOP_acc_14_psp_sva[2:0]==3'b111) & (fsm_output[5]) & (~ (fsm_output[7]))
      & (~ (fsm_output[4]));
  assign and_428_nl = (z_out_6_10_1[3:0]==4'b1111) & (fsm_output[5]) & (~ (fsm_output[7]))
      & (fsm_output[4]);
  assign mux_1497_nl = MUX_s_1_2_2(and_292_nl, and_428_nl, fsm_output[0]);
  assign nor_290_nl = ~((z_out_6_10_1[3:0]!=4'b1111) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1498_nl = MUX_s_1_2_2(mux_1497_nl, nor_290_nl, fsm_output[6]);
  assign mux_1502_nl = MUX_s_1_2_2(mux_1501_nl, mux_1498_nl, fsm_output[1]);
  assign and_289_nl = (fsm_output[3]) & mux_1502_nl;
  assign mux_1506_nl = MUX_s_1_2_2(mux_1505_nl, and_289_nl, fsm_output[2]);
  assign mux_1517_nl = MUX_s_1_2_2(mux_1516_nl, mux_1506_nl, fsm_output[8]);
  assign and_433_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b1111) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      & (~ (fsm_output[5])) & (~ (fsm_output[7])) & (fsm_output[4]);
  assign mux_1493_nl = MUX_s_1_2_2(and_291_cse, and_433_nl, fsm_output[0]);
  assign nor_293_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_9_0[1:0]!=2'b11)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[4]));
  assign and_440_nl = (z_out_6_10_1[3:0]==4'b1111) & (~ (fsm_output[5])) & (~ (fsm_output[7]))
      & (fsm_output[4]);
  assign mux_1492_nl = MUX_s_1_2_2(nor_293_nl, and_440_nl, fsm_output[0]);
  assign mux_1494_nl = MUX_s_1_2_2(mux_1493_nl, mux_1492_nl, fsm_output[6]);
  assign nor_295_nl = ~((z_out_6_10_1[3:0]!=4'b1111) | (fsm_output[6]) | (fsm_output[0])
      | (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1495_nl = MUX_s_1_2_2(mux_1494_nl, nor_295_nl, fsm_output[1]);
  assign nand_101_nl = ~((fsm_output[3]) & mux_1495_nl);
  assign or_1763_nl = (~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1111) & (fsm_output[6])
      & (fsm_output[0]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & (~ (fsm_output[5]))))
      | not_tmp_134;
  assign nand_172_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]==3'b111) & (VEC_LOOP_j_sva_9_0[0])
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (fsm_output[7])
      & (~ (fsm_output[4])));
  assign mux_1489_nl = MUX_s_1_2_2(nand_172_nl, nand_161_cse, fsm_output[0]);
  assign nand_348_nl = ~((COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1111) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[5]) & (~ (fsm_output[7])) & (fsm_output[4]));
  assign mux_1488_nl = MUX_s_1_2_2(nand_160_cse, nand_348_nl, fsm_output[0]);
  assign mux_1490_nl = MUX_s_1_2_2(mux_1489_nl, mux_1488_nl, fsm_output[6]);
  assign mux_1491_nl = MUX_s_1_2_2(or_1763_nl, mux_1490_nl, fsm_output[1]);
  assign or_1764_nl = (fsm_output[3]) | mux_1491_nl;
  assign mux_1496_nl = MUX_s_1_2_2(nand_101_nl, or_1764_nl, fsm_output[2]);
  assign nor_291_nl = ~((fsm_output[8]) | mux_1496_nl);
  assign vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1517_nl,
      nor_291_nl, fsm_output[9]);
  assign or_2213_nl = (fsm_output[0]) | (~ (fsm_output[7])) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (~ (fsm_output[8])) | (fsm_output[9]);
  assign mux_2057_nl = MUX_s_1_2_2(or_1977_cse, or_279_cse, fsm_output[0]);
  assign mux_tmp_2006 = MUX_s_1_2_2(or_2213_nl, mux_2057_nl, fsm_output[4]);
  assign or_2219_nl = (fsm_output[4]) | (~ (fsm_output[0])) | (fsm_output[7]) | (fsm_output[2])
      | (fsm_output[3]) | (~ (fsm_output[8])) | (fsm_output[9]);
  assign or_2218_nl = (fsm_output[0]) | (~ (fsm_output[7])) | (fsm_output[2]) | (~
      (fsm_output[3])) | (fsm_output[8]) | (~ (fsm_output[9]));
  assign mux_2062_nl = MUX_s_1_2_2(or_1995_cse, nand_357_cse, fsm_output[0]);
  assign mux_2063_nl = MUX_s_1_2_2(or_2218_nl, mux_2062_nl, fsm_output[4]);
  assign mux_2064_nl = MUX_s_1_2_2(or_2219_nl, mux_2063_nl, fsm_output[5]);
  assign or_2214_nl = (fsm_output[4]) | (~ (fsm_output[0])) | (fsm_output[7]) | (~
      (fsm_output[2])) | (fsm_output[3]) | (fsm_output[8]) | (fsm_output[9]);
  assign mux_2061_nl = MUX_s_1_2_2(or_2214_nl, mux_tmp_2006, fsm_output[5]);
  assign mux_2065_nl = MUX_s_1_2_2(mux_2064_nl, mux_2061_nl, fsm_output[6]);
  assign or_2209_nl = (fsm_output[4]) | (~ (fsm_output[0])) | (~ (fsm_output[7]))
      | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[8]) | (fsm_output[9]);
  assign mux_2059_nl = MUX_s_1_2_2(mux_tmp_2006, or_2209_nl, fsm_output[5]);
  assign or_2207_nl = (fsm_output[0]) | (fsm_output[7]) | (fsm_output[2]) | (~ (fsm_output[3]))
      | (fsm_output[8]) | (~ (fsm_output[9]));
  assign mux_2055_nl = MUX_s_1_2_2(or_1976_cse, mux_1768_cse, fsm_output[0]);
  assign mux_2056_nl = MUX_s_1_2_2(or_2207_nl, mux_2055_nl, fsm_output[4]);
  assign or_2208_nl = (fsm_output[5]) | mux_2056_nl;
  assign mux_2060_nl = MUX_s_1_2_2(mux_2059_nl, or_2208_nl, fsm_output[6]);
  assign mux_2066_cse = MUX_s_1_2_2(mux_2065_nl, mux_2060_nl, fsm_output[1]);
  assign and_dcpl_231 = ~((fsm_output[1]) | (fsm_output[6]));
  assign and_dcpl_232 = and_dcpl_231 & (~ (fsm_output[5]));
  assign and_dcpl_233 = and_dcpl_232 & and_dcpl_29;
  assign and_dcpl_234 = (~ (fsm_output[7])) & (fsm_output[2]);
  assign and_dcpl_236 = ~((fsm_output[9]) | (fsm_output[8]) | (fsm_output[3]));
  assign and_dcpl_237 = and_dcpl_236 & and_dcpl_234;
  assign and_dcpl_238 = and_dcpl_237 & and_dcpl_233;
  assign and_dcpl_242 = and_dcpl_237 & and_dcpl_231 & (fsm_output[5]) & and_dcpl_32;
  assign and_dcpl_243 = (~ (fsm_output[1])) & (fsm_output[6]);
  assign and_dcpl_244 = and_dcpl_243 & (~ (fsm_output[5]));
  assign and_dcpl_246 = and_dcpl_237 & and_dcpl_244 & and_dcpl_29;
  assign and_dcpl_248 = (fsm_output[1]) & (~ (fsm_output[6])) & (fsm_output[5]);
  assign and_dcpl_250 = (fsm_output[7]) & (~ (fsm_output[2]));
  assign and_dcpl_251 = and_dcpl_236 & and_dcpl_250;
  assign and_dcpl_252 = and_dcpl_251 & and_dcpl_248 & and_dcpl_29;
  assign and_dcpl_255 = and_dcpl_251 & and_dcpl_243 & (fsm_output[5]) & and_dcpl_32;
  assign and_dcpl_256 = ~((fsm_output[7]) | (fsm_output[2]));
  assign and_dcpl_260 = and_dcpl_70 & (~ (fsm_output[3])) & and_dcpl_256 & and_dcpl_233;
  assign and_dcpl_265 = and_dcpl_70 & (fsm_output[3]);
  assign and_dcpl_267 = and_dcpl_265 & and_dcpl_234 & (fsm_output[1]) & (fsm_output[6])
      & (fsm_output[5]) & and_dcpl_16;
  assign and_dcpl_271 = and_dcpl_265 & (fsm_output[7]) & (fsm_output[2]);
  assign and_dcpl_272 = and_dcpl_271 & and_dcpl_232 & and_dcpl_66;
  assign and_dcpl_274 = and_dcpl_271 & and_dcpl_244 & and_dcpl_16;
  assign and_dcpl_277 = (fsm_output[9]) & (~ (fsm_output[8])) & (fsm_output[3]);
  assign and_dcpl_278 = and_dcpl_277 & and_dcpl_256;
  assign and_dcpl_279 = and_dcpl_278 & and_dcpl_248 & and_dcpl_16;
  assign and_dcpl_281 = and_dcpl_278 & and_dcpl_244 & and_dcpl_66;
  assign and_dcpl_284 = and_dcpl_277 & and_dcpl_250 & and_dcpl_232 & and_dcpl_16;
  assign and_dcpl_293 = and_dcpl_236 & (~ (fsm_output[7])) & (fsm_output[2]) & (~
      (fsm_output[1])) & (~ (fsm_output[6])) & (~ (fsm_output[5])) & (~ (fsm_output[0]))
      & (fsm_output[4]);
  assign and_dcpl_300 = and_dcpl_236 & and_dcpl_250 & (fsm_output[1]) & (~ (fsm_output[6]))
      & (~ (fsm_output[5])) & (fsm_output[0]) & (~ (fsm_output[4]));
  assign and_dcpl_308 = (fsm_output[8]) & (~ (fsm_output[9])) & (fsm_output[3]) &
      and_dcpl_250 & (fsm_output[1]) & (fsm_output[6]) & (fsm_output[5]) & (fsm_output[0])
      & (fsm_output[4]);
  assign and_dcpl_344 = ~((fsm_output!=10'b0000010100));
  assign and_dcpl_361 = (~ (fsm_output[9])) & (fsm_output[8]) & (fsm_output[3]) &
      and_dcpl_234 & (fsm_output[1]) & (~ (fsm_output[6])) & (fsm_output[5]) & (fsm_output[0])
      & (fsm_output[4]);
  assign and_dcpl_376 = (fsm_output[1]) & (~ (fsm_output[6]));
  assign and_dcpl_382 = and_dcpl_376 & (fsm_output[5]);
  assign and_dcpl_396 = and_dcpl_382 & and_dcpl_66;
  assign and_dcpl_398 = and_dcpl_265 & and_dcpl_234;
  assign and_dcpl_402 = (fsm_output[1]) & (fsm_output[6]) & (fsm_output[5]);
  assign and_dcpl_403 = and_dcpl_402 & and_dcpl_16;
  assign and_dcpl_406 = (fsm_output[7]) & (fsm_output[2]);
  assign and_dcpl_407 = and_dcpl_265 & and_dcpl_406;
  assign and_dcpl_416 = and_dcpl_98 & (fsm_output[3]);
  assign and_dcpl_417 = and_dcpl_416 & and_dcpl_256;
  assign and_dcpl_425 = and_dcpl_98 & (~ (fsm_output[3])) & and_dcpl_406;
  assign and_dcpl_444 = ~((fsm_output[9]) | (fsm_output[8]) | (fsm_output[3]) | (~
      and_dcpl_234) | (fsm_output[1]) | (fsm_output[6]) | (fsm_output[5]) | (~ (fsm_output[0]))
      | (fsm_output[4]));
  assign and_dcpl_460 = (fsm_output[8]) & (fsm_output[9]) & (~ (fsm_output[3])) &
      (~ (fsm_output[7])) & (fsm_output[2]) & (fsm_output[1]) & (~ (fsm_output[6]))
      & (~ (fsm_output[5])) & and_dcpl_16;
  assign nor_761_cse = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[5]));
  assign and_dcpl_464 = nor_761_cse & (fsm_output[0]) & (~ (fsm_output[4]));
  assign and_551_ssc = (fsm_output[9]) & (~ (fsm_output[8])) & (~ (fsm_output[3]))
      & (fsm_output[7]) & (fsm_output[2]) & (fsm_output[1]) & (fsm_output[6]) & (fsm_output[5])
      & and_dcpl_16;
  assign nand_tmp_139 = ~((fsm_output[3]) & (~(and_dcpl_16 | (fsm_output[9:8]!=2'b01))));
  assign or_tmp_2154 = (fsm_output[3]) | (~ (fsm_output[0])) | (fsm_output[8]) |
      (fsm_output[9]);
  assign or_2261_nl = (~ (fsm_output[3])) | (fsm_output[4]) | (fsm_output[0]) | (~
      (fsm_output[8])) | (fsm_output[9]);
  assign mux_tmp_2041 = MUX_s_1_2_2(or_tmp_2154, or_2261_nl, fsm_output[2]);
  assign or_tmp_2156 = nor_810_cse | (fsm_output[9:8]!=2'b10);
  assign or_2267_nl = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[8]) | (fsm_output[9]);
  assign or_2266_nl = (~ (fsm_output[0])) | (~ (fsm_output[8])) | (fsm_output[9]);
  assign mux_tmp_2043 = MUX_s_1_2_2(or_2267_nl, or_2266_nl, fsm_output[3]);
  assign or_2271_nl = (~ (fsm_output[4])) | (~ (fsm_output[0])) | (fsm_output[8])
      | (fsm_output[9]);
  assign or_2270_nl = (fsm_output[4]) | (fsm_output[0]) | (fsm_output[8]) | (~ (fsm_output[9]));
  assign mux_2097_nl = MUX_s_1_2_2(or_2271_nl, or_2270_nl, fsm_output[3]);
  assign nand_388_nl = ~((fsm_output[3]) & (~(nor_810_cse | (fsm_output[9:8]!=2'b01))));
  assign mux_tmp_2046 = MUX_s_1_2_2(mux_2097_nl, nand_388_nl, fsm_output[2]);
  assign or_tmp_2166 = (~ (fsm_output[0])) | (fsm_output[8]) | (~ (fsm_output[9]));
  assign or_tmp_2168 = (fsm_output[3]) | and_dcpl_66 | (fsm_output[9:8]!=2'b00);
  assign nand_389_nl = ~((fsm_output[3]) & (~ or_tmp_2156));
  assign mux_2103_nl = MUX_s_1_2_2(nand_389_nl, mux_tmp_2043, fsm_output[2]);
  assign or_2272_nl = (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[8])) | (fsm_output[9]);
  assign mux_2101_nl = MUX_s_1_2_2(or_tmp_2166, or_2272_nl, fsm_output[3]);
  assign mux_2102_nl = MUX_s_1_2_2(or_tmp_2168, mux_2101_nl, fsm_output[2]);
  assign mux_tmp_2052 = MUX_s_1_2_2(mux_2103_nl, mux_2102_nl, fsm_output[7]);
  assign or_tmp_2171 = and_dcpl_16 | (fsm_output[9:8]!=2'b10);
  assign or_2282_nl = (~ (fsm_output[3])) | (fsm_output[4]) | (fsm_output[0]) | (fsm_output[8])
      | (~ (fsm_output[9]));
  assign mux_tmp_2058 = MUX_s_1_2_2(or_2282_nl, nand_tmp_139, fsm_output[2]);
  assign or_tmp_2183 = ~((fsm_output[4]) & (fsm_output[7]) & (fsm_output[8]) & (fsm_output[3])
      & (~ (fsm_output[9])));
  assign mux_2123_nl = MUX_s_1_2_2(mux_tmp_1610, or_tmp_1796, fsm_output[4]);
  assign mux_tmp_2072 = MUX_s_1_2_2(or_tmp_2183, mux_2123_nl, fsm_output[0]);
  assign not_tmp_571 = ~((fsm_output[3]) & (fsm_output[9]));
  assign or_tmp_2191 = (fsm_output[8:7]!=2'b00) | not_tmp_571;
  assign or_tmp_2193 = (~ (fsm_output[4])) | (fsm_output[7]) | (fsm_output[8]) |
      not_tmp_571;
  assign or_2302_nl = (fsm_output[8]) | not_tmp_571;
  assign mux_tmp_2081 = MUX_s_1_2_2(or_2302_nl, or_2012_cse, fsm_output[7]);
  assign mux_2134_nl = MUX_s_1_2_2(mux_tmp_2081, or_tmp_2193, fsm_output[0]);
  assign mux_2131_nl = MUX_s_1_2_2(or_tmp_1793, or_tmp_1796, fsm_output[4]);
  assign mux_2132_nl = MUX_s_1_2_2(mux_2131_nl, mux_1583_cse, fsm_output[0]);
  assign mux_tmp_2083 = MUX_s_1_2_2(mux_2134_nl, mux_2132_nl, fsm_output[2]);
  assign mux_tmp_2108 = MUX_s_1_2_2(mux_tmp_1874, mux_tmp_1861, fsm_output[1]);
  assign or_tmp_2223 = ((fsm_output[3:1]==3'b111)) | (fsm_output[9:8]!=2'b01);
  assign mux_2163_nl = MUX_s_1_2_2(or_tmp_2041, mux_1920_cse, fsm_output[1]);
  assign mux_tmp_2112 = MUX_s_1_2_2(or_tmp_2223, mux_2163_nl, fsm_output[7]);
  assign or_tmp_2227 = (~((fsm_output[3:1]!=3'b000))) | (fsm_output[9:8]!=2'b01);
  assign mux_2169_nl = MUX_s_1_2_2(or_tmp_2041, mux_1922_cse, fsm_output[1]);
  assign mux_2170_nl = MUX_s_1_2_2(or_tmp_2227, mux_2169_nl, fsm_output[7]);
  assign mux_2166_nl = MUX_s_1_2_2(nand_tmp_134, mux_tmp_1861, fsm_output[1]);
  assign mux_2167_nl = MUX_s_1_2_2(mux_2166_nl, or_tmp_2037, fsm_output[7]);
  assign mux_tmp_2119 = MUX_s_1_2_2(mux_2170_nl, mux_2167_nl, fsm_output[6]);
  assign mux_2175_nl = MUX_s_1_2_2(nand_tmp_134, mux_tmp_1874, fsm_output[1]);
  assign mux_tmp_2124 = MUX_s_1_2_2(mux_2175_nl, or_tmp_2037, fsm_output[7]);
  assign mux_2179_nl = MUX_s_1_2_2(mux_1938_cse, or_tmp_2041, fsm_output[1]);
  assign mux_tmp_2128 = MUX_s_1_2_2(mux_2179_nl, mux_tmp_1861, fsm_output[7]);
  assign or_tmp_2236 = (fsm_output[9:8]!=2'b00);
  assign mux_tmp_2150 = MUX_s_1_2_2(or_tmp_2236, (fsm_output[8]), or_2146_cse);
  assign mux_tmp_2153 = MUX_s_1_2_2((fsm_output[8]), or_2086_cse, fsm_output[2]);
  assign mux_tmp_2154 = MUX_s_1_2_2(mux_tmp_2153, or_tmp_2043, fsm_output[3]);
  assign mux_tmp_2156 = MUX_s_1_2_2(or_tmp_2236, (fsm_output[8]), fsm_output[3]);
  assign mux_tmp_2159 = MUX_s_1_2_2(mux_tmp_2154, or_tmp_2037, fsm_output[4]);
  assign or_2346_nl = and_357_cse | (fsm_output[9:8]!=2'b01);
  assign mux_2215_nl = MUX_s_1_2_2(mux_tmp_1861, mux_tmp_2156, fsm_output[0]);
  assign mux_tmp_2164 = MUX_s_1_2_2(or_2346_nl, mux_2215_nl, fsm_output[4]);
  assign mux_tmp_2165 = MUX_s_1_2_2(mux_tmp_1861, mux_tmp_2154, fsm_output[4]);
  assign mux_tmp_2167 = MUX_s_1_2_2(mux_tmp_2153, or_tmp_2044, fsm_output[3]);
  assign mux_2220_nl = MUX_s_1_2_2(mux_tmp_2167, mux_tmp_2154, fsm_output[0]);
  assign mux_tmp_2169 = MUX_s_1_2_2(mux_2220_nl, or_212_cse, fsm_output[4]);
  assign mux_tmp_2170 = MUX_s_1_2_2(or_212_cse, mux_tmp_1861, fsm_output[4]);
  assign mux_tmp_2179 = MUX_s_1_2_2(or_tmp_2236, (fsm_output[8]), fsm_output[2]);
  assign mux_tmp_2180 = MUX_s_1_2_2(or_tmp_2035, mux_tmp_2179, fsm_output[3]);
  assign or_tmp_2243 = (fsm_output[5]) | (fsm_output[1]);
  assign or_tmp_2244 = (fsm_output[5]) | (~ (fsm_output[1]));
  assign mux_tmp_2192 = MUX_s_1_2_2(or_tmp_2244, or_tmp_2243, fsm_output[0]);
  assign or_2350_nl = (~((fsm_output[0]) | (fsm_output[5]))) | (fsm_output[1]);
  assign mux_tmp_2193 = MUX_s_1_2_2(mux_tmp_2192, or_2350_nl, fsm_output[4]);
  assign or_tmp_2245 = (fsm_output[0]) | (~((fsm_output[5]) & (fsm_output[1])));
  assign mux_tmp_2196 = MUX_s_1_2_2(or_tmp_2245, or_tmp_2244, fsm_output[4]);
  assign nand_399_nl = ~((fsm_output[0]) & (fsm_output[5]) & (fsm_output[1]));
  assign mux_2249_itm = MUX_s_1_2_2(nand_399_nl, mux_tmp_2196, fsm_output[6]);
  assign mux_tmp_2199 = MUX_s_1_2_2(or_tmp_2243, or_2186_cse, fsm_output[4]);
  assign or_2360_nl = (~ (fsm_output[0])) | (~ (fsm_output[5])) | (fsm_output[1]);
  assign mux_tmp_2204 = MUX_s_1_2_2(or_2360_nl, mux_tmp_2192, fsm_output[4]);
  always @(posedge clk) begin
    if ( (and_dcpl_19 & and_dcpl_15) | STAGE_LOOP_i_3_0_sva_mx0c1 ) begin
      STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(4'b0001, (z_out_7[3:0]), STAGE_LOOP_i_3_0_sva_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ not_tmp_121 ) begin
      p_sva <= p_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( ~ not_tmp_121 ) begin
      r_sva <= r_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_vec_rsc_triosy_0_15_obj_ld_cse <= 1'b0;
      reg_ensig_cgo_cse <= 1'b0;
      COMP_LOOP_nor_11_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_nor_1_itm <= 1'b0;
      COMP_LOOP_nor_12_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_139_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_140_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_141_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_143_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_144_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_145_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_146_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_147_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_148_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_149_itm <= 1'b0;
      COMP_LOOP_nor_134_itm <= 1'b0;
      COMP_LOOP_nor_137_itm <= 1'b0;
    end
    else begin
      reg_vec_rsc_triosy_0_15_obj_ld_cse <= and_dcpl_18 & and_dcpl_16 & (fsm_output[1])
          & (fsm_output[2]) & (~ (fsm_output[6])) & (fsm_output[9]) & (fsm_output[8])
          & (~ (z_out_8_64_2[0]));
      reg_ensig_cgo_cse <= ~ mux_1581_itm;
      COMP_LOOP_nor_11_itm <= MUX_s_1_2_2((z_out_3[5]), COMP_LOOP_nor_11_nl, modExp_dev_while_or_2_cse);
      COMP_LOOP_COMP_LOOP_nor_1_itm <= ~((z_out_6_10_1[3:0]!=4'b0000));
      COMP_LOOP_nor_12_itm <= ~((z_out_6_10_1[3]) | (z_out_6_10_1[2]) | (z_out_6_10_1[0]));
      COMP_LOOP_COMP_LOOP_and_139_itm <= (z_out_6_10_1[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_140_itm <= (z_out_6_10_1[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_141_itm <= (z_out_6_10_1[3:0]==4'b0111);
      COMP_LOOP_COMP_LOOP_and_143_itm <= (z_out_6_10_1[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_144_itm <= (z_out_6_10_1[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_145_itm <= (z_out_6_10_1[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_146_itm <= (z_out_6_10_1[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_147_itm <= (z_out_6_10_1[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_148_itm <= (z_out_6_10_1[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_149_itm <= (z_out_6_10_1[3:0]==4'b1111);
      COMP_LOOP_nor_134_itm <= ~((z_out_6_10_1[3]) | (z_out_6_10_1[1]) | (z_out_6_10_1[0]));
      COMP_LOOP_nor_137_itm <= ~((z_out_6_10_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    operator_66_true_div_cmp_a <= MUX_v_65_2_2(z_out_9, ({operator_64_false_acc_mut_64
        , operator_64_false_acc_mut_63_0}), and_dcpl_169);
    operator_66_true_div_cmp_b_9_0 <= MUX_v_10_2_2(STAGE_LOOP_lshift_psp_sva_mx0w0,
        STAGE_LOOP_lshift_psp_sva, and_dcpl_169);
    modExp_dev_exp_1_sva_3_0 <= MUX_v_4_2_2(COMP_LOOP_and_nl, 4'b1111, and_dcpl_221);
    COMP_LOOP_1_mul_itm <= nl_COMP_LOOP_1_mul_itm[63:0];
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(nor_271_nl, and_tmp_12, fsm_output[8]) ) begin
      STAGE_LOOP_lshift_psp_sva <= STAGE_LOOP_lshift_psp_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ mux_2121_nl ) begin
      operator_64_false_acc_mut_64 <= operator_64_false_operator_64_false_mux_rgt[64];
    end
  end
  always @(posedge clk) begin
    if ( ~ mux_2153_nl ) begin
      operator_64_false_acc_mut_63_0 <= operator_64_false_operator_64_false_mux_rgt[63:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      VEC_LOOP_j_sva_9_0 <= 10'b0000000000;
    end
    else if ( (~(mux_tmp_1688 | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[3])
        | (fsm_output[6]) | (~ nor_697_cse))) | VEC_LOOP_j_sva_9_0_mx0c1 ) begin
      VEC_LOOP_j_sva_9_0 <= MUX_v_10_2_2(10'b0000000000, (VEC_LOOP_acc_1_psp_1[9:0]),
          VEC_LOOP_j_sva_9_0_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~(mux_2156_nl | (fsm_output[3])) ) begin
      COMP_LOOP_k_9_4_sva_4_0 <= MUX_v_5_2_2(5'b00000, (z_out_3[4:0]), or_nl);
    end
  end
  always @(posedge clk) begin
    if ( mux_1749_nl | and_195_rgt ) begin
      modExp_dev_result_sva <= MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000001,
          modulo_dev_cmp_return_rsc_z, and_195_rgt);
    end
  end
  always @(posedge clk) begin
    if ( mux_1754_nl | (fsm_output[7:5]!=3'b000) | (~ nor_697_cse) ) begin
      modExp_dev_exp_sva <= MUX_v_64_2_2((operator_66_true_div_cmp_z[63:0]), (z_out_9[63:0]),
          and_dcpl_183);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_137_itm <= 1'b0;
    end
    else if ( and_dcpl_183 | not_tmp_402 | and_dcpl_36 | and_dcpl_44 | and_dcpl_52
        | and_dcpl_58 | and_dcpl_63 | and_dcpl_72 | and_dcpl_78 | and_dcpl_84 | and_dcpl_90
        | and_dcpl_93 | and_dcpl_97 | and_dcpl_102 | and_dcpl_106 | and_dcpl_110
        | and_dcpl_115 | and_dcpl_119 ) begin
      COMP_LOOP_COMP_LOOP_and_137_itm <= MUX_s_1_2_2((~ (z_out_7[64])), COMP_LOOP_COMP_LOOP_and_17_nl,
          modExp_dev_while_or_2_cse);
    end
  end
  always @(posedge clk) begin
    if ( ~(or_tmp_74 | (fsm_output[3]) | (~ (fsm_output[4])) | (fsm_output[0]) |
        (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[6]) | (fsm_output[9])
        | (fsm_output[8])) ) begin
      COMP_LOOP_acc_psp_sva <= z_out_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_244_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_62_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_2_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_64_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_4_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_5_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_6_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_68_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_8_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_9_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_11_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_12_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_13_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_14_itm <= 1'b0;
    end
    else if ( mux_1832_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_itm <= ~((VEC_LOOP_j_sva_9_0[3:0]!=4'b0000));
      COMP_LOOP_COMP_LOOP_and_244_itm <= (COMP_LOOP_acc_13_psp_sva_1[0]) & (VEC_LOOP_j_sva_9_0[0])
          & (~((COMP_LOOP_acc_13_psp_sva_1[1]) | (VEC_LOOP_j_sva_9_0[1])));
      COMP_LOOP_COMP_LOOP_and_62_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b0011);
      COMP_LOOP_COMP_LOOP_and_2_itm <= (VEC_LOOP_j_sva_9_0[3:0]==4'b0011);
      COMP_LOOP_COMP_LOOP_and_64_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_4_itm <= (VEC_LOOP_j_sva_9_0[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_5_itm <= (VEC_LOOP_j_sva_9_0[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_6_itm <= (VEC_LOOP_j_sva_9_0[3:0]==4'b0111);
      COMP_LOOP_COMP_LOOP_and_68_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_8_itm <= (VEC_LOOP_j_sva_9_0[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_9_itm <= (VEC_LOOP_j_sva_9_0[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_11_itm <= (VEC_LOOP_j_sva_9_0[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_12_itm <= (VEC_LOOP_j_sva_9_0[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_13_itm <= (VEC_LOOP_j_sva_9_0[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_14_itm <= (VEC_LOOP_j_sva_9_0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_10_itm <= 1'b0;
    end
    else if ( ~ mux_1842_nl ) begin
      COMP_LOOP_COMP_LOOP_and_10_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_10_nl,
          (~ (readslicef_10_1_9(COMP_LOOP_1_acc_nl))), and_dcpl_119);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_13_psp_sva <= 8'b00000000;
    end
    else if ( ~(mux_1845_nl & nor_697_cse) ) begin
      COMP_LOOP_acc_13_psp_sva <= COMP_LOOP_acc_13_psp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_2_sva <= 10'b0000000000;
    end
    else if ( (~ mux_1848_nl) | (fsm_output[9:7]!=3'b000) ) begin
      COMP_LOOP_acc_1_cse_2_sva <= COMP_LOOP_acc_1_cse_2_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_11_psp_sva <= 9'b000000000;
    end
    else if ( ~((~ mux_1858_nl) & nor_697_cse) ) begin
      COMP_LOOP_acc_11_psp_sva <= nl_COMP_LOOP_acc_11_psp_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_4_sva <= 10'b0000000000;
    end
    else if ( ~(mux_1862_nl & nor_697_cse) ) begin
      COMP_LOOP_acc_1_cse_4_sva <= nl_COMP_LOOP_acc_1_cse_4_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_6_sva <= 10'b0000000000;
    end
    else if ( mux_1866_nl | (fsm_output[9]) ) begin
      COMP_LOOP_acc_1_cse_6_sva <= z_out_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_14_psp_sva <= 9'b000000000;
    end
    else if ( mux_1869_nl | (fsm_output[9]) ) begin
      COMP_LOOP_acc_14_psp_sva <= nl_COMP_LOOP_acc_14_psp_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_8_sva <= 10'b0000000000;
    end
    else if ( mux_1872_nl | (fsm_output[9]) ) begin
      COMP_LOOP_acc_1_cse_8_sva <= nl_COMP_LOOP_acc_1_cse_8_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_16_psp_sva <= 7'b0000000;
    end
    else if ( mux_1874_nl | (fsm_output[9]) ) begin
      COMP_LOOP_acc_16_psp_sva <= z_out_5;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_10_sva <= 10'b0000000000;
    end
    else if ( mux_1875_nl | (fsm_output[9]) ) begin
      COMP_LOOP_acc_1_cse_10_sva <= nl_COMP_LOOP_acc_1_cse_10_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_17_psp_sva <= 9'b000000000;
    end
    else if ( MUX_s_1_2_2(mux_1877_nl, (fsm_output[9]), fsm_output[8]) ) begin
      COMP_LOOP_acc_17_psp_sva <= nl_COMP_LOOP_acc_17_psp_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_12_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_1880_nl, (fsm_output[9]), fsm_output[8]) ) begin
      COMP_LOOP_acc_1_cse_12_sva <= nl_COMP_LOOP_acc_1_cse_12_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_19_psp_sva <= 8'b00000000;
    end
    else if ( MUX_s_1_2_2(mux_1885_nl, (fsm_output[9]), or_110_nl) ) begin
      COMP_LOOP_acc_19_psp_sva <= z_out_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_14_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_1888_nl, (fsm_output[9]), fsm_output[8]) ) begin
      COMP_LOOP_acc_1_cse_14_sva <= nl_COMP_LOOP_acc_1_cse_14_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_20_psp_sva <= 9'b000000000;
    end
    else if ( MUX_s_1_2_2(mux_1896_nl, (fsm_output[9]), fsm_output[8]) ) begin
      COMP_LOOP_acc_20_psp_sva <= nl_COMP_LOOP_acc_20_psp_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(nor_nl, and_nl, fsm_output[8]) ) begin
      COMP_LOOP_acc_1_cse_sva <= nl_COMP_LOOP_acc_1_cse_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( and_dcpl_199 | and_dcpl_200 | and_dcpl_201 | and_dcpl_202 | and_dcpl_203
        | and_dcpl_204 | and_dcpl_206 | and_dcpl_208 | and_dcpl_210 | and_dcpl_212
        | and_dcpl_214 | and_dcpl_215 | and_dcpl_217 | and_dcpl_219 | and_dcpl_220
        | and_dcpl_221 ) begin
      tmp_10_lpi_4_dfm <= MUX1HOT_v_64_16_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d,
          vec_rsc_0_2_i_q_d, vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d,
          vec_rsc_0_6_i_q_d, vec_rsc_0_7_i_q_d, vec_rsc_0_8_i_q_d, vec_rsc_0_9_i_q_d,
          vec_rsc_0_10_i_q_d, vec_rsc_0_11_i_q_d, vec_rsc_0_12_i_q_d, vec_rsc_0_13_i_q_d,
          vec_rsc_0_14_i_q_d, vec_rsc_0_15_i_q_d, {COMP_LOOP_or_6_nl , COMP_LOOP_or_7_nl
          , COMP_LOOP_or_8_nl , COMP_LOOP_or_9_nl , COMP_LOOP_or_10_nl , COMP_LOOP_or_11_nl
          , COMP_LOOP_or_12_nl , COMP_LOOP_or_13_nl , COMP_LOOP_or_14_nl , COMP_LOOP_or_15_nl
          , COMP_LOOP_or_16_nl , COMP_LOOP_or_17_nl , COMP_LOOP_or_18_nl , COMP_LOOP_or_19_nl
          , COMP_LOOP_or_20_nl , COMP_LOOP_or_21_nl});
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_2196_nl, mux_2184_nl, fsm_output[4]) ) begin
      modExp_dev_exp_1_sva_63_9 <= MUX_v_55_2_2(55'b0000000000000000000000000000000000000000000000000000000,
          (z_out_9[63:9]), not_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_1_sva_9_5 <= 5'b00000;
    end
    else if ( ~ mux_2243_nl ) begin
      COMP_LOOP_acc_10_cse_10_1_1_sva_9_5 <= COMP_LOOP_mux1h_192_rgt[9:5];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_1_sva_4_0 <= 5'b00000;
    end
    else if ( MUX_s_1_2_2(mux_2262_nl, nor_800_nl, fsm_output[8]) ) begin
      COMP_LOOP_acc_10_cse_10_1_1_sva_4_0 <= COMP_LOOP_mux1h_192_rgt[4:0];
    end
  end
  always @(posedge clk) begin
    if ( and_dcpl_36 | and_dcpl_44 | and_dcpl_58 | and_dcpl_63 | and_dcpl_72 | and_dcpl_84
        | and_dcpl_90 | and_dcpl_93 | and_dcpl_102 | and_dcpl_106 | and_dcpl_110
        ) begin
      COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm <= z_out_1[9];
    end
  end
  always @(posedge clk) begin
    if ( and_dcpl_52 | and_dcpl_78 | and_dcpl_97 | and_dcpl_115 ) begin
      COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= MUX1HOT_s_1_3_2((z_out_2[7]), (z_out_5[6]),
          (z_out_4[5]), {COMP_LOOP_or_27_nl , and_dcpl_78 , and_dcpl_115});
    end
  end
  assign COMP_LOOP_nor_11_nl = ~((z_out_6_10_1[3:1]!=3'b000));
  assign mux_1950_nl = MUX_s_1_2_2(mux_1949_cse, mux_tmp_1874, fsm_output[7]);
  assign mux_1951_nl = MUX_s_1_2_2(mux_1950_nl, mux_tmp_1888, fsm_output[0]);
  assign mux_1952_nl = MUX_s_1_2_2(mux_tmp_1891, mux_1951_nl, fsm_output[5]);
  assign mux_1948_nl = MUX_s_1_2_2(mux_tmp_1876, mux_tmp_1883, fsm_output[5]);
  assign mux_1953_nl = MUX_s_1_2_2(mux_1952_nl, mux_1948_nl, fsm_output[6]);
  assign mux_1944_nl = MUX_s_1_2_2(nand_tmp_134, or_212_cse, fsm_output[7]);
  assign mux_1945_nl = MUX_s_1_2_2(mux_1944_nl, mux_tmp_1876, fsm_output[0]);
  assign mux_1943_nl = MUX_s_1_2_2(mux_tmp_1891, mux_tmp_1882, fsm_output[0]);
  assign mux_1946_nl = MUX_s_1_2_2(mux_1945_nl, mux_1943_nl, fsm_output[5]);
  assign mux_1940_nl = MUX_s_1_2_2(mux_tmp_1888, mux_tmp_1866, fsm_output[0]);
  assign mux_1941_nl = MUX_s_1_2_2(mux_1940_nl, mux_tmp_1877, fsm_output[5]);
  assign mux_1947_nl = MUX_s_1_2_2(mux_1946_nl, mux_1941_nl, fsm_output[6]);
  assign mux_1954_nl = MUX_s_1_2_2(mux_1953_nl, mux_1947_nl, fsm_output[4]);
  assign mux_1935_nl = MUX_s_1_2_2(mux_tmp_1883, mux_tmp_1866, fsm_output[5]);
  assign mux_1931_nl = MUX_s_1_2_2(mux_tmp_1875, mux_tmp_1863, fsm_output[0]);
  assign mux_1932_nl = MUX_s_1_2_2(mux_1931_nl, mux_tmp_1870, fsm_output[5]);
  assign mux_1936_nl = MUX_s_1_2_2(mux_1935_nl, mux_1932_nl, fsm_output[6]);
  assign mux_1924_nl = MUX_s_1_2_2(mux_tmp_1872, mux_tmp_1870, fsm_output[0]);
  assign mux_1929_nl = MUX_s_1_2_2(mux_tmp_1877, mux_1924_nl, fsm_output[5]);
  assign mux_1916_nl = MUX_s_1_2_2(or_tmp_2041, or_2336_cse, fsm_output[7]);
  assign mux_1918_nl = MUX_s_1_2_2(mux_tmp_1866, mux_1916_nl, fsm_output[0]);
  assign mux_1913_nl = MUX_s_1_2_2(mux_tmp_1861, or_1916_cse, fsm_output[7]);
  assign mux_1915_nl = MUX_s_1_2_2(mux_tmp_1863, mux_1913_nl, fsm_output[0]);
  assign mux_1919_nl = MUX_s_1_2_2(mux_1918_nl, mux_1915_nl, fsm_output[5]);
  assign mux_1930_nl = MUX_s_1_2_2(mux_1929_nl, mux_1919_nl, fsm_output[6]);
  assign mux_1937_nl = MUX_s_1_2_2(mux_1936_nl, mux_1930_nl, fsm_output[4]);
  assign mux_1955_nl = MUX_s_1_2_2(mux_1954_nl, mux_1937_nl, fsm_output[1]);
  assign COMP_LOOP_mux1h_186_nl = MUX1HOT_v_4_16_2((z_out_9[3:0]), modExp_dev_exp_1_sva_3_0,
      4'b0001, 4'b0010, 4'b0011, 4'b0100, 4'b0101, 4'b0110, 4'b0111, 4'b1000, 4'b1001,
      4'b1010, 4'b1011, 4'b1100, 4'b1101, 4'b1110, {not_tmp_402 , (~ mux_1955_nl)
      , and_dcpl_200 , and_dcpl_201 , and_dcpl_202 , and_dcpl_203 , and_dcpl_204
      , and_dcpl_206 , and_dcpl_208 , and_dcpl_210 , and_dcpl_212 , and_dcpl_214
      , and_dcpl_215 , and_dcpl_217 , and_dcpl_219 , and_dcpl_220});
  assign not_4628_nl = ~ and_dcpl_199;
  assign COMP_LOOP_and_nl = MUX_v_4_2_2(4'b0000, COMP_LOOP_mux1h_186_nl, not_4628_nl);
  assign COMP_LOOP_COMP_LOOP_and_930_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[0])
      & COMP_LOOP_nor_11_itm;
  assign COMP_LOOP_COMP_LOOP_and_932_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[1])
      & COMP_LOOP_nor_12_itm;
  assign COMP_LOOP_COMP_LOOP_and_934_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[2])
      & COMP_LOOP_nor_134_itm;
  assign COMP_LOOP_COMP_LOOP_and_936_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0[3])
      & COMP_LOOP_nor_137_itm;
  assign COMP_LOOP_mux1h_209_nl = MUX1HOT_v_64_16_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d,
      vec_rsc_0_2_i_q_d, vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d,
      vec_rsc_0_6_i_q_d, vec_rsc_0_7_i_q_d, vec_rsc_0_8_i_q_d, vec_rsc_0_9_i_q_d,
      vec_rsc_0_10_i_q_d, vec_rsc_0_11_i_q_d, vec_rsc_0_12_i_q_d, vec_rsc_0_13_i_q_d,
      vec_rsc_0_14_i_q_d, vec_rsc_0_15_i_q_d, {COMP_LOOP_COMP_LOOP_nor_1_itm , COMP_LOOP_COMP_LOOP_and_930_nl
      , COMP_LOOP_COMP_LOOP_and_932_nl , COMP_LOOP_COMP_LOOP_and_137_itm , COMP_LOOP_COMP_LOOP_and_934_nl
      , COMP_LOOP_COMP_LOOP_and_139_itm , COMP_LOOP_COMP_LOOP_and_140_itm , COMP_LOOP_COMP_LOOP_and_141_itm
      , COMP_LOOP_COMP_LOOP_and_936_nl , COMP_LOOP_COMP_LOOP_and_143_itm , COMP_LOOP_COMP_LOOP_and_144_itm
      , COMP_LOOP_COMP_LOOP_and_145_itm , COMP_LOOP_COMP_LOOP_and_146_itm , COMP_LOOP_COMP_LOOP_and_147_itm
      , COMP_LOOP_COMP_LOOP_and_148_itm , COMP_LOOP_COMP_LOOP_and_149_itm});
  assign nl_COMP_LOOP_1_mul_itm  = $signed(operator_64_false_acc_mut_63_0) * $signed(conv_u2s_64_65(COMP_LOOP_mux1h_209_nl));
  assign nor_271_nl = ~((fsm_output[9]) | (fsm_output[6]) | (fsm_output[2]) | (fsm_output[1])
      | (fsm_output[4]) | (fsm_output[3]) | (fsm_output[7]) | (fsm_output[5]));
  assign or_2286_nl = (~((fsm_output[0]) | (fsm_output[8]))) | (fsm_output[9]);
  assign or_2284_nl = (fsm_output[0]) | (~ (fsm_output[8])) | (fsm_output[9]);
  assign mux_2116_nl = MUX_s_1_2_2(or_2286_nl, or_2284_nl, fsm_output[4]);
  assign or_2287_nl = (fsm_output[3]) | mux_2116_nl;
  assign mux_2117_nl = MUX_s_1_2_2(or_2287_nl, or_tmp_2154, fsm_output[2]);
  assign mux_2118_nl = MUX_s_1_2_2(mux_2117_nl, mux_tmp_2058, fsm_output[7]);
  assign or_2283_nl = (~ (fsm_output[4])) | (fsm_output[0]) | (~ (fsm_output[8]))
      | (fsm_output[9]);
  assign mux_2113_nl = MUX_s_1_2_2(or_2283_nl, or_tmp_2166, fsm_output[3]);
  assign mux_2114_nl = MUX_s_1_2_2(mux_2113_nl, or_tmp_2168, fsm_output[2]);
  assign mux_2115_nl = MUX_s_1_2_2(mux_2114_nl, mux_tmp_2046, fsm_output[7]);
  assign mux_2119_nl = MUX_s_1_2_2(mux_2118_nl, mux_2115_nl, fsm_output[5]);
  assign or_2280_nl = (fsm_output[3]) | or_tmp_2171;
  assign mux_2109_nl = MUX_s_1_2_2(or_tmp_2168, or_2280_nl, fsm_output[2]);
  assign mux_2111_nl = MUX_s_1_2_2(mux_tmp_2058, mux_2109_nl, fsm_output[7]);
  assign mux_2112_nl = MUX_s_1_2_2(mux_tmp_2052, mux_2111_nl, fsm_output[5]);
  assign mux_2120_nl = MUX_s_1_2_2(mux_2119_nl, mux_2112_nl, fsm_output[1]);
  assign nand_390_nl = ~((fsm_output[3]) & (~ or_tmp_2171));
  assign mux_2105_nl = MUX_s_1_2_2(nand_390_nl, or_tmp_2168, fsm_output[2]);
  assign mux_2106_nl = MUX_s_1_2_2(mux_2105_nl, mux_tmp_2041, fsm_output[7]);
  assign mux_2107_nl = MUX_s_1_2_2(mux_2106_nl, mux_tmp_2052, fsm_output[5]);
  assign or_2265_nl = (fsm_output[3]) | or_tmp_2156;
  assign mux_2096_nl = MUX_s_1_2_2(mux_tmp_2043, or_2265_nl, fsm_output[2]);
  assign mux_2099_nl = MUX_s_1_2_2(mux_tmp_2046, mux_2096_nl, fsm_output[7]);
  assign or_2258_nl = (fsm_output[3]) | (fsm_output[4]) | (fsm_output[0]) | (fsm_output[8])
      | (~ (fsm_output[9]));
  assign mux_nl = MUX_s_1_2_2(nand_tmp_139, or_2258_nl, fsm_output[2]);
  assign mux_2094_nl = MUX_s_1_2_2(mux_tmp_2041, mux_nl, fsm_output[7]);
  assign mux_2100_nl = MUX_s_1_2_2(mux_2099_nl, mux_2094_nl, fsm_output[5]);
  assign mux_2108_nl = MUX_s_1_2_2(mux_2107_nl, mux_2100_nl, fsm_output[1]);
  assign mux_2121_nl = MUX_s_1_2_2(mux_2120_nl, mux_2108_nl, fsm_output[6]);
  assign or_2310_nl = (fsm_output[4]) | (fsm_output[7]) | (~ (fsm_output[8])) | (fsm_output[3])
      | (fsm_output[9]);
  assign or_2309_nl = (fsm_output[4]) | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9]);
  assign mux_2149_nl = MUX_s_1_2_2(or_2310_nl, or_2309_nl, fsm_output[0]);
  assign mux_2150_nl = MUX_s_1_2_2(mux_2149_nl, mux_tmp_2072, fsm_output[2]);
  assign or_2308_nl = (fsm_output[8:7]!=2'b01) | not_tmp_571;
  assign mux_2146_nl = MUX_s_1_2_2(or_2308_nl, or_2306_cse, fsm_output[4]);
  assign mux_2145_nl = MUX_s_1_2_2(or_tmp_2191, mux_tmp_2081, fsm_output[4]);
  assign mux_2147_nl = MUX_s_1_2_2(mux_2146_nl, mux_2145_nl, fsm_output[0]);
  assign mux_2144_nl = MUX_s_1_2_2(mux_tmp_1610, or_tmp_2183, fsm_output[0]);
  assign mux_2148_nl = MUX_s_1_2_2(mux_2147_nl, mux_2144_nl, fsm_output[2]);
  assign mux_2151_nl = MUX_s_1_2_2(mux_2150_nl, mux_2148_nl, fsm_output[5]);
  assign or_2305_nl = (fsm_output[4]) | (~ (fsm_output[7])) | (fsm_output[8]) | (fsm_output[3])
      | (fsm_output[9]);
  assign nand_392_nl = ~((fsm_output[4]) & (~ mux_1583_cse));
  assign or_2304_nl = (fsm_output[4]) | mux_1583_cse;
  assign mux_2141_nl = MUX_s_1_2_2(nand_392_nl, or_2304_nl, fsm_output[0]);
  assign mux_2142_nl = MUX_s_1_2_2(or_2305_nl, mux_2141_nl, fsm_output[2]);
  assign mux_2143_nl = MUX_s_1_2_2(mux_tmp_2083, mux_2142_nl, fsm_output[5]);
  assign mux_2152_nl = MUX_s_1_2_2(mux_2151_nl, mux_2143_nl, fsm_output[1]);
  assign mux_2136_nl = MUX_s_1_2_2(mux_tmp_2081, or_tmp_1788, fsm_output[4]);
  assign mux_2137_nl = MUX_s_1_2_2(or_tmp_2193, mux_2136_nl, fsm_output[0]);
  assign or_2303_nl = (fsm_output[4]) | (fsm_output[7]) | (fsm_output[8]) | (fsm_output[3])
      | (fsm_output[9]);
  assign mux_2138_nl = MUX_s_1_2_2(mux_2137_nl, or_2303_nl, fsm_output[2]);
  assign mux_2139_nl = MUX_s_1_2_2(mux_2138_nl, mux_tmp_2083, fsm_output[5]);
  assign mux_2127_nl = MUX_s_1_2_2(or_tmp_2191, or_tmp_1788, fsm_output[4]);
  assign mux_2126_nl = MUX_s_1_2_2(or_tmp_1793, mux_tmp_1610, fsm_output[4]);
  assign mux_2128_nl = MUX_s_1_2_2(mux_2127_nl, mux_2126_nl, fsm_output[0]);
  assign or_2367_nl = nor_810_cse | mux_1583_cse;
  assign mux_2129_nl = MUX_s_1_2_2(mux_2128_nl, or_2367_nl, fsm_output[2]);
  assign or_2292_nl = (fsm_output[2]) | mux_tmp_2072;
  assign mux_2130_nl = MUX_s_1_2_2(mux_2129_nl, or_2292_nl, fsm_output[5]);
  assign mux_2140_nl = MUX_s_1_2_2(mux_2139_nl, mux_2130_nl, fsm_output[1]);
  assign mux_2153_nl = MUX_s_1_2_2(mux_2152_nl, mux_2140_nl, fsm_output[6]);
  assign or_1923_nl = (fsm_output[9]) | mux_tmp_1688;
  assign or_1922_nl = (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[1])
      | (~ (fsm_output[0])) | (fsm_output[4]);
  assign mux_1740_nl = MUX_s_1_2_2(or_1923_nl, or_1922_nl, fsm_output[8]);
  assign or_nl = mux_1740_nl | (~ and_dcpl_17) | (fsm_output[3]) | (fsm_output[6]);
  assign or_2316_nl = (fsm_output[9]) | (fsm_output[1]) | (fsm_output[8]) | (~ (fsm_output[2]))
      | (fsm_output[4]);
  assign or_2315_nl = (~ (fsm_output[1])) | (fsm_output[8]) | (fsm_output[2]) | (~
      (fsm_output[4]));
  assign or_2313_nl = (fsm_output[1]) | (~ (fsm_output[8])) | (~ (fsm_output[2]))
      | (fsm_output[4]);
  assign mux_2154_nl = MUX_s_1_2_2(or_2315_nl, or_2313_nl, fsm_output[9]);
  assign mux_2155_nl = MUX_s_1_2_2(or_2316_nl, mux_2154_nl, fsm_output[0]);
  assign or_2365_nl = (fsm_output[7:6]!=2'b00) | mux_2155_nl;
  assign or_2366_nl = (~ (fsm_output[7])) | (~ (fsm_output[6])) | (fsm_output[0])
      | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[8]) | (~ (fsm_output[2]))
      | (fsm_output[4]);
  assign mux_2156_nl = MUX_s_1_2_2(or_2365_nl, or_2366_nl, fsm_output[5]);
  assign mux_1747_nl = MUX_s_1_2_2(or_tmp_1899, or_103_cse, and_267_cse);
  assign mux_1748_nl = MUX_s_1_2_2(mux_1747_nl, or_103_cse, fsm_output[2]);
  assign nor_269_nl = ~((fsm_output[9]) | (fsm_output[6]) | mux_1748_nl);
  assign mux_1749_nl = MUX_s_1_2_2(nor_269_nl, and_tmp_12, fsm_output[8]);
  assign mux_1753_nl = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), fsm_output[4]);
  assign or_1936_nl = (fsm_output[4:3]!=2'b01);
  assign mux_1752_nl = MUX_s_1_2_2(or_1936_nl, (fsm_output[4]), fsm_output[1]);
  assign mux_1754_nl = MUX_s_1_2_2(mux_1753_nl, mux_1752_nl, fsm_output[2]);
  assign COMP_LOOP_COMP_LOOP_and_17_nl = (z_out_6_10_1[3:0]==4'b0011);
  assign COMP_LOOP_COMP_LOOP_and_10_nl = (VEC_LOOP_j_sva_9_0[3:0]==4'b1011);
  assign nl_COMP_LOOP_1_acc_nl = ({z_out_3 , 4'b0000}) + ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[9:1]))})
      + 10'b0000000001;
  assign COMP_LOOP_1_acc_nl = nl_COMP_LOOP_1_acc_nl[9:0];
  assign mux_1836_nl = MUX_s_1_2_2((~ mux_1834_itm), or_tmp_1989, fsm_output[4]);
  assign mux_1838_nl = MUX_s_1_2_2(mux_tmp_1786, mux_1836_nl, fsm_output[1]);
  assign or_2033_nl = (fsm_output[4]) | (~ mux_1834_itm);
  assign mux_1835_nl = MUX_s_1_2_2(or_2033_nl, mux_tmp_1782, fsm_output[1]);
  assign mux_1839_nl = MUX_s_1_2_2(mux_1838_nl, mux_1835_nl, fsm_output[0]);
  assign mux_1840_nl = MUX_s_1_2_2(mux_tmp_1786, mux_1839_nl, fsm_output[2]);
  assign mux_1841_nl = MUX_s_1_2_2(mux_1840_nl, mux_tmp_1782, fsm_output[3]);
  assign nand_146_nl = ~(((fsm_output[7:2]!=6'b000000)) & (fsm_output[9]));
  assign mux_1842_nl = MUX_s_1_2_2(mux_1841_nl, nand_146_nl, fsm_output[8]);
  assign nand_338_nl = ~((fsm_output[2]) & or_2186_cse & (fsm_output[4]) & (fsm_output[3])
      & (fsm_output[7]) & (fsm_output[5]));
  assign mux_1845_nl = MUX_s_1_2_2(mux_tmp_1793, nand_338_nl, fsm_output[6]);
  assign or_23_nl = (fsm_output[5:4]!=2'b00);
  assign mux_66_nl = MUX_s_1_2_2(or_tmp_20, or_23_nl, or_2186_cse);
  assign mux_67_nl = MUX_s_1_2_2(or_tmp_20, mux_66_nl, fsm_output[2]);
  assign nand_145_nl = ~((fsm_output[5:4]==2'b11));
  assign mux_1848_nl = MUX_s_1_2_2(mux_67_nl, nand_145_nl, fsm_output[6]);
  assign nl_COMP_LOOP_acc_11_psp_sva  = (VEC_LOOP_j_sva_9_0[9:1]) + conv_u2u_8_9({COMP_LOOP_k_9_4_sva_4_0
      , 3'b001});
  assign mux_1855_nl = MUX_s_1_2_2(mux_tmp_1803, mux_tmp_1801, fsm_output[0]);
  assign mux_1849_nl = MUX_s_1_2_2(nor_tmp_40, (fsm_output[7]), fsm_output[3]);
  assign mux_1851_nl = MUX_s_1_2_2(mux_tmp_1799, mux_1849_nl, fsm_output[4]);
  assign mux_1853_nl = MUX_s_1_2_2(mux_tmp_1801, mux_1851_nl, fsm_output[0]);
  assign mux_1856_nl = MUX_s_1_2_2(mux_1855_nl, mux_1853_nl, fsm_output[1]);
  assign mux_1857_nl = MUX_s_1_2_2(mux_tmp_1803, mux_1856_nl, fsm_output[2]);
  assign mux_1858_nl = MUX_s_1_2_2(mux_1857_nl, (fsm_output[7]), fsm_output[6]);
  assign nl_COMP_LOOP_acc_1_cse_4_sva  = VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0011});
  assign mux_1861_nl = MUX_s_1_2_2(mux_tmp_1809, mux_tmp_1808, and_418_cse);
  assign mux_1862_nl = MUX_s_1_2_2(mux_tmp_1793, (~ mux_1861_nl), fsm_output[6]);
  assign mux_1864_nl = MUX_s_1_2_2((fsm_output[7]), or_tmp_74, fsm_output[4]);
  assign mux_1863_nl = MUX_s_1_2_2((fsm_output[7]), or_tmp_74, or_2040_cse);
  assign mux_1865_nl = MUX_s_1_2_2(mux_1864_nl, mux_1863_nl, fsm_output[2]);
  assign or_2041_nl = (fsm_output[6]) | mux_1865_nl;
  assign mux_1866_nl = MUX_s_1_2_2(not_tmp_431, or_2041_nl, fsm_output[8]);
  assign nl_COMP_LOOP_acc_14_psp_sva  = (VEC_LOOP_j_sva_9_0[9:1]) + conv_u2u_8_9({COMP_LOOP_k_9_4_sva_4_0
      , 3'b011});
  assign or_2043_nl = ((fsm_output[1]) & (fsm_output[0]) & (fsm_output[4]) & (fsm_output[3]))
      | (fsm_output[7]) | (fsm_output[5]);
  assign mux_1867_nl = MUX_s_1_2_2(or_2043_nl, or_tmp_1899, fsm_output[2]);
  assign mux_1868_nl = MUX_s_1_2_2((fsm_output[7]), mux_1867_nl, fsm_output[6]);
  assign mux_1869_nl = MUX_s_1_2_2(not_tmp_431, mux_1868_nl, fsm_output[8]);
  assign nl_COMP_LOOP_acc_1_cse_8_sva  = VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0111});
  assign or_2175_nl = (fsm_output[2:1]!=2'b00);
  assign mux_1870_nl = MUX_s_1_2_2(mux_tmp_1809, mux_tmp_1808, or_2175_nl);
  assign mux_1871_nl = MUX_s_1_2_2(mux_1870_nl, (fsm_output[7]), fsm_output[6]);
  assign mux_1872_nl = MUX_s_1_2_2(not_tmp_431, mux_1871_nl, fsm_output[8]);
  assign and_248_nl = ((fsm_output[2:0]!=3'b000)) & (fsm_output[4]) & (fsm_output[3])
      & (fsm_output[7]) & (fsm_output[5]);
  assign mux_1873_nl = MUX_s_1_2_2(and_248_nl, (fsm_output[7]), fsm_output[6]);
  assign mux_1874_nl = MUX_s_1_2_2(not_tmp_431, mux_1873_nl, fsm_output[8]);
  assign nl_COMP_LOOP_acc_1_cse_10_sva  = VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1001});
  assign and_213_nl = (fsm_output[6]) & or_2040_cse & (fsm_output[7]) & (fsm_output[5]);
  assign mux_1875_nl = MUX_s_1_2_2(not_tmp_431, and_213_nl, fsm_output[8]);
  assign nl_COMP_LOOP_acc_17_psp_sva  = (VEC_LOOP_j_sva_9_0[9:1]) + conv_u2u_8_9({COMP_LOOP_k_9_4_sva_4_0
      , 3'b101});
  assign mux_1876_nl = MUX_s_1_2_2(or_tmp_1899, or_103_cse, and_247_cse);
  assign or_2047_nl = (fsm_output[6]) | mux_1876_nl;
  assign mux_1877_nl = MUX_s_1_2_2(not_tmp_431, or_2047_nl, fsm_output[9]);
  assign nl_COMP_LOOP_acc_1_cse_12_sva  = VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1011});
  assign mux_1879_nl = MUX_s_1_2_2((fsm_output[7]), or_tmp_1845, fsm_output[6]);
  assign mux_1880_nl = MUX_s_1_2_2(not_tmp_431, mux_1879_nl, fsm_output[9]);
  assign mux_1882_nl = MUX_s_1_2_2(not_tmp_439, nor_tmp_215, or_2186_cse);
  assign mux_1883_nl = MUX_s_1_2_2(not_tmp_439, mux_1882_nl, fsm_output[2]);
  assign mux_1884_nl = MUX_s_1_2_2(mux_1883_nl, nor_tmp_215, fsm_output[3]);
  assign mux_1885_nl = MUX_s_1_2_2(not_tmp_439, mux_1884_nl, fsm_output[4]);
  assign or_110_nl = (fsm_output[8:7]!=2'b00);
  assign nl_COMP_LOOP_acc_1_cse_14_sva  = VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1101});
  assign and_245_nl = ((fsm_output[4:2]!=3'b000)) & (fsm_output[7]) & (fsm_output[5]);
  assign mux_1887_nl = MUX_s_1_2_2(and_245_nl, (fsm_output[7]), fsm_output[6]);
  assign mux_1888_nl = MUX_s_1_2_2(not_tmp_431, mux_1887_nl, fsm_output[9]);
  assign nl_COMP_LOOP_acc_20_psp_sva  = (VEC_LOOP_j_sva_9_0[9:1]) + conv_u2u_8_9({COMP_LOOP_k_9_4_sva_4_0
      , 3'b111});
  assign mux_1892_nl = MUX_s_1_2_2(not_tmp_418, mux_tmp_1839, and_267_cse);
  assign mux_1891_nl = MUX_s_1_2_2(mux_tmp_1839, nor_tmp_203, or_2186_cse);
  assign mux_1893_nl = MUX_s_1_2_2(mux_1892_nl, mux_1891_nl, fsm_output[2]);
  assign mux_1894_nl = MUX_s_1_2_2(mux_1893_nl, nor_tmp_203, fsm_output[3]);
  assign mux_1895_nl = MUX_s_1_2_2(not_tmp_418, mux_1894_nl, fsm_output[4]);
  assign mux_1896_nl = MUX_s_1_2_2(mux_1895_nl, nor_tmp_203, fsm_output[5]);
  assign nl_COMP_LOOP_acc_1_cse_sva  = VEC_LOOP_j_sva_9_0 + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1111});
  assign nor_nl = ~((fsm_output[9]) | (fsm_output[6]) | mux_tmp_1793);
  assign and_nl = (fsm_output[9]) & ((fsm_output[7:1]!=7'b0000000));
  assign COMP_LOOP_or_6_nl = (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_199) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_200) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_201) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_202) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_dcpl_203) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_204) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_dcpl_206) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_dcpl_208) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_210) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_212) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_dcpl_214) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_dcpl_215) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_217) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_dcpl_219) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_220) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_dcpl_221);
  assign COMP_LOOP_or_7_nl = (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_199) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_200) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_201) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_202) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_203) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_dcpl_204) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_206) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_dcpl_208) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_dcpl_210) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_dcpl_212) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_214) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_dcpl_215) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_dcpl_217) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_dcpl_219) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_dcpl_220) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_221);
  assign COMP_LOOP_or_8_nl = (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_199) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_dcpl_200) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_201) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_202) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_203) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_204) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_dcpl_206) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_208) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_dcpl_210) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_dcpl_212) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_214) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_215) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_dcpl_217) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_dcpl_219) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_220) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_dcpl_221);
  assign COMP_LOOP_or_9_nl = (COMP_LOOP_COMP_LOOP_and_2_itm & and_dcpl_199) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_200) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_201) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_202) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_203) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_204) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_206) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_dcpl_208) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_210) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_dcpl_212) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_dcpl_214) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_dcpl_215) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_217) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_dcpl_219) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_dcpl_220) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_dcpl_221);
  assign COMP_LOOP_or_10_nl = (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_199) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_dcpl_200) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_201) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_dcpl_202) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_203) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_204) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_206) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_208) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_dcpl_210) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_212) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_dcpl_214) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_dcpl_215) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_217) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_219) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_dcpl_220) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_dcpl_221);
  assign COMP_LOOP_or_11_nl = (COMP_LOOP_COMP_LOOP_and_4_itm & and_dcpl_199) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_dcpl_200) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_dcpl_201) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_202) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_203) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_204) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_206) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_208) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_210) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_dcpl_212) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_214) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_dcpl_215) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_dcpl_217) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_dcpl_219) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_220) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_dcpl_221);
  assign COMP_LOOP_or_12_nl = (COMP_LOOP_COMP_LOOP_and_5_itm & and_dcpl_199) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_dcpl_200) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_201) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_dcpl_202) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_203) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_dcpl_204) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_206) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_208) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_210) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_212) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_dcpl_214) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_215) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_dcpl_217) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_dcpl_219) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_220) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_221);
  assign COMP_LOOP_or_13_nl = (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_199) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_dcpl_200) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_dcpl_201) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_dcpl_202) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_dcpl_203) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_204) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_206) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_208) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_210) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_212) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_214) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_dcpl_215) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_217) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_dcpl_219) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_dcpl_220) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_dcpl_221);
  assign COMP_LOOP_or_14_nl = (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_199) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_200) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_dcpl_201) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_dcpl_202) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_203) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_dcpl_204) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_206) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_dcpl_208) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_210) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_212) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_214) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_215) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_dcpl_217) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_219) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_dcpl_220) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_dcpl_221);
  assign COMP_LOOP_or_15_nl = (COMP_LOOP_COMP_LOOP_and_8_itm & and_dcpl_199) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_dcpl_200) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_201) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_dcpl_202) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_dcpl_203) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_dcpl_204) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_dcpl_206) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_208) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_210) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_212) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_214) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_215) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_217) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_dcpl_219) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_220) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_dcpl_221);
  assign COMP_LOOP_or_16_nl = (COMP_LOOP_COMP_LOOP_and_9_itm & and_dcpl_199) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_dcpl_200) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_201) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_202) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_dcpl_203) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_dcpl_204) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_206) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_dcpl_208) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_210) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_dcpl_212) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_214) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_215) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_217) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_219) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_dcpl_220) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_221);
  assign COMP_LOOP_or_17_nl = (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_199) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_dcpl_200) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_dcpl_201) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_dcpl_202) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_203) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_dcpl_204) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_dcpl_206) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_dcpl_208) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_dcpl_210) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_212) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_214) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_215) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_217) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_219) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_220) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_dcpl_221);
  assign COMP_LOOP_or_18_nl = (COMP_LOOP_COMP_LOOP_and_11_itm & and_dcpl_199) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_200) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_dcpl_201) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_dcpl_202) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_203) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_204) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_dcpl_206) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_dcpl_208) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_210) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_dcpl_212) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_214) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_dcpl_215) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_217) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_219) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_220) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_221);
  assign COMP_LOOP_or_19_nl = (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_199) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_dcpl_200) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_201) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_dcpl_202) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_dcpl_203) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_dcpl_204) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_206) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_dcpl_208) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_dcpl_210) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_dcpl_212) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_dcpl_214) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_215) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_217) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_219) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_220) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_221);
  assign COMP_LOOP_or_20_nl = (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_199) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_200) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_dcpl_201) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_202) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_dcpl_203) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_dcpl_204) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_206) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_208) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_dcpl_210) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_dcpl_212) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_214) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_dcpl_215) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_217) | (COMP_LOOP_COMP_LOOP_and_244_itm
      & and_dcpl_219) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_220) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_221);
  assign COMP_LOOP_or_21_nl = (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_199) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_200) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_201) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_dcpl_202) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_203) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_dcpl_204) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_dcpl_206) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_dcpl_208) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_210) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_dcpl_212) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_dcpl_214) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_dcpl_215) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_dcpl_217) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_219) | (COMP_LOOP_COMP_LOOP_and_244_itm & and_dcpl_220) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_221);
  assign not_nl = ~ mux_1911_cse;
  assign mux_2193_nl = MUX_s_1_2_2(or_tmp_2227, or_tmp_2041, fsm_output[7]);
  assign mux_2194_nl = MUX_s_1_2_2(mux_2193_nl, mux_tmp_2124, fsm_output[6]);
  assign mux_2195_nl = MUX_s_1_2_2(mux_2194_nl, mux_tmp_2119, fsm_output[0]);
  assign mux_2189_nl = MUX_s_1_2_2(mux_1949_cse, or_tmp_2041, fsm_output[1]);
  assign mux_2190_nl = MUX_s_1_2_2(mux_2189_nl, mux_tmp_2108, fsm_output[7]);
  assign mux_2191_nl = MUX_s_1_2_2(mux_2190_nl, mux_tmp_2112, fsm_output[6]);
  assign mux_2185_nl = MUX_s_1_2_2(mux_1922_cse, mux_1920_cse, fsm_output[1]);
  assign mux_2186_nl = MUX_s_1_2_2(or_tmp_2223, mux_2185_nl, fsm_output[7]);
  assign mux_2187_nl = MUX_s_1_2_2(mux_tmp_2128, mux_2186_nl, fsm_output[6]);
  assign mux_2192_nl = MUX_s_1_2_2(mux_2191_nl, mux_2187_nl, fsm_output[0]);
  assign mux_2196_nl = MUX_s_1_2_2(mux_2195_nl, mux_2192_nl, fsm_output[5]);
  assign mux_2181_nl = MUX_s_1_2_2(nand_tmp_134, or_tmp_2223, fsm_output[7]);
  assign mux_2182_nl = MUX_s_1_2_2(mux_2181_nl, mux_tmp_2128, fsm_output[6]);
  assign mux_2173_nl = MUX_s_1_2_2(mux_tmp_1861, or_2336_cse, fsm_output[1]);
  assign mux_2174_nl = MUX_s_1_2_2(or_tmp_2041, mux_2173_nl, fsm_output[7]);
  assign mux_2177_nl = MUX_s_1_2_2(mux_tmp_2124, mux_2174_nl, fsm_output[6]);
  assign mux_2183_nl = MUX_s_1_2_2(mux_2182_nl, mux_2177_nl, fsm_output[0]);
  assign mux_2157_nl = MUX_s_1_2_2(or_tmp_2037, or_1916_cse, fsm_output[1]);
  assign mux_2161_nl = MUX_s_1_2_2(mux_tmp_2108, mux_2157_nl, fsm_output[7]);
  assign mux_2165_nl = MUX_s_1_2_2(mux_tmp_2112, mux_2161_nl, fsm_output[6]);
  assign mux_2172_nl = MUX_s_1_2_2(mux_tmp_2119, mux_2165_nl, fsm_output[0]);
  assign mux_2184_nl = MUX_s_1_2_2(mux_2183_nl, mux_2172_nl, fsm_output[5]);
  assign or_2347_nl = (fsm_output[2]) | (~ (fsm_output[8])) | (fsm_output[9]);
  assign mux_2237_nl = MUX_s_1_2_2(or_2347_nl, mux_tmp_2179, fsm_output[3]);
  assign mux_2238_nl = MUX_s_1_2_2(mux_2237_nl, mux_tmp_2180, fsm_output[0]);
  assign mux_2239_nl = MUX_s_1_2_2(or_212_cse, mux_2238_nl, fsm_output[4]);
  assign mux_2236_nl = MUX_s_1_2_2(mux_1949_cse, or_212_cse, fsm_output[4]);
  assign mux_2240_nl = MUX_s_1_2_2(mux_2239_nl, mux_2236_nl, fsm_output[5]);
  assign mux_2233_nl = MUX_s_1_2_2(mux_tmp_2180, mux_tmp_1861, fsm_output[0]);
  assign mux_2230_nl = MUX_s_1_2_2(mux_1949_cse, mux_tmp_2167, fsm_output[0]);
  assign mux_2234_nl = MUX_s_1_2_2(mux_2233_nl, mux_2230_nl, fsm_output[4]);
  assign mux_2235_nl = MUX_s_1_2_2(mux_2234_nl, mux_tmp_2170, fsm_output[5]);
  assign mux_2241_nl = MUX_s_1_2_2(mux_2240_nl, mux_2235_nl, fsm_output[6]);
  assign mux_2227_nl = MUX_s_1_2_2(mux_tmp_2169, mux_tmp_2165, fsm_output[5]);
  assign mux_2226_nl = MUX_s_1_2_2(mux_tmp_2164, mux_tmp_2159, fsm_output[5]);
  assign mux_2228_nl = MUX_s_1_2_2(mux_2227_nl, mux_2226_nl, fsm_output[6]);
  assign mux_2242_nl = MUX_s_1_2_2(mux_2241_nl, mux_2228_nl, fsm_output[7]);
  assign mux_2223_nl = MUX_s_1_2_2(mux_tmp_2170, mux_tmp_2169, fsm_output[5]);
  assign mux_2218_nl = MUX_s_1_2_2(mux_tmp_2165, mux_tmp_2164, fsm_output[5]);
  assign mux_2224_nl = MUX_s_1_2_2(mux_2223_nl, mux_2218_nl, fsm_output[6]);
  assign mux_2209_nl = MUX_s_1_2_2(mux_tmp_2156, mux_tmp_2150, fsm_output[0]);
  assign mux_2207_nl = MUX_s_1_2_2(mux_tmp_2154, mux_1922_cse, fsm_output[0]);
  assign mux_2210_nl = MUX_s_1_2_2(mux_2209_nl, mux_2207_nl, fsm_output[4]);
  assign mux_2212_nl = MUX_s_1_2_2(mux_tmp_2159, mux_2210_nl, fsm_output[5]);
  assign mux_2203_nl = MUX_s_1_2_2(or_tmp_2037, mux_tmp_2150, fsm_output[4]);
  assign mux_2198_nl = MUX_s_1_2_2(or_tmp_2044, or_212_cse, fsm_output[3]);
  assign mux_2200_nl = MUX_s_1_2_2(mux_1922_cse, mux_2198_nl, fsm_output[0]);
  assign mux_2201_nl = MUX_s_1_2_2(mux_2200_nl, or_tmp_2037, fsm_output[4]);
  assign mux_2204_nl = MUX_s_1_2_2(mux_2203_nl, mux_2201_nl, fsm_output[5]);
  assign mux_2213_nl = MUX_s_1_2_2(mux_2212_nl, mux_2204_nl, fsm_output[6]);
  assign mux_2225_nl = MUX_s_1_2_2(mux_2224_nl, mux_2213_nl, fsm_output[7]);
  assign mux_2243_nl = MUX_s_1_2_2(mux_2242_nl, mux_2225_nl, fsm_output[1]);
  assign nand_396_nl = ~((fsm_output[6]) & (fsm_output[4]) & (fsm_output[0]) & (fsm_output[5])
      & (fsm_output[1]));
  assign mux_2259_nl = MUX_s_1_2_2(mux_tmp_2204, mux_tmp_2199, fsm_output[6]);
  assign mux_2260_nl = MUX_s_1_2_2(nand_396_nl, mux_2259_nl, fsm_output[2]);
  assign nand_397_nl = ~(((fsm_output[0]) | (fsm_output[5])) & (fsm_output[1]));
  assign mux_2257_nl = MUX_s_1_2_2(nand_397_nl, or_tmp_2245, fsm_output[4]);
  assign mux_2258_nl = MUX_s_1_2_2(mux_2257_nl, mux_tmp_2204, fsm_output[6]);
  assign or_2362_nl = (fsm_output[2]) | mux_2258_nl;
  assign mux_2261_nl = MUX_s_1_2_2(mux_2260_nl, or_2362_nl, fsm_output[7]);
  assign nor_797_nl = ~((fsm_output[3]) | mux_2261_nl);
  assign and_700_nl = (fsm_output[7]) & (fsm_output[2]) & (~ mux_2249_itm);
  assign mux_2253_nl = MUX_s_1_2_2(mux_tmp_2196, mux_tmp_2193, fsm_output[6]);
  assign nor_798_nl = ~((fsm_output[2]) | mux_2253_nl);
  assign nor_799_nl = ~((fsm_output[2]) | (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0])
      | (fsm_output[1]));
  assign mux_2254_nl = MUX_s_1_2_2(nor_798_nl, nor_799_nl, fsm_output[7]);
  assign mux_2255_nl = MUX_s_1_2_2(and_700_nl, mux_2254_nl, fsm_output[3]);
  assign mux_2262_nl = MUX_s_1_2_2(nor_797_nl, mux_2255_nl, fsm_output[9]);
  assign or_2356_nl = (fsm_output[7]) | (fsm_output[2]) | (fsm_output[6]) | mux_tmp_2199;
  assign nand_394_nl = ~((fsm_output[2]) & (~ mux_2249_itm));
  assign nand_398_nl = ~((fsm_output[6]) & (fsm_output[0]) & (fsm_output[5]) & (fsm_output[1]));
  assign mux_2246_nl = MUX_s_1_2_2(mux_tmp_2193, or_2348_cse, fsm_output[6]);
  assign mux_2247_nl = MUX_s_1_2_2(nand_398_nl, mux_2246_nl, fsm_output[2]);
  assign mux_2250_nl = MUX_s_1_2_2(nand_394_nl, mux_2247_nl, fsm_output[7]);
  assign mux_2252_nl = MUX_s_1_2_2(or_2356_nl, mux_2250_nl, fsm_output[3]);
  assign nor_800_nl = ~((fsm_output[9]) | mux_2252_nl);
  assign COMP_LOOP_or_27_nl = and_dcpl_52 | and_dcpl_97;
  assign COMP_LOOP_COMP_LOOP_or_3_nl = (VEC_LOOP_j_sva_9_0[9]) | and_dcpl_242 | and_dcpl_246
      | and_dcpl_252 | and_dcpl_255 | and_dcpl_260 | and_dcpl_267 | and_dcpl_272
      | and_dcpl_274 | and_dcpl_279 | and_dcpl_281 | and_dcpl_284;
  assign COMP_LOOP_or_52_nl = and_dcpl_242 | and_dcpl_246 | and_dcpl_252 | and_dcpl_255
      | and_dcpl_260 | and_dcpl_267 | and_dcpl_272 | and_dcpl_274 | and_dcpl_279
      | and_dcpl_281 | and_dcpl_284;
  assign COMP_LOOP_COMP_LOOP_mux_15_nl = MUX_v_9_2_2((VEC_LOOP_j_sva_9_0[8:0]), (~
      (STAGE_LOOP_lshift_psp_sva[9:1])), COMP_LOOP_or_52_nl);
  assign COMP_LOOP_or_53_nl = (~ and_dcpl_238) | and_dcpl_242 | and_dcpl_246 | and_dcpl_252
      | and_dcpl_255 | and_dcpl_260 | and_dcpl_267 | and_dcpl_272 | and_dcpl_274
      | and_dcpl_279 | and_dcpl_281 | and_dcpl_284;
  assign COMP_LOOP_or_54_nl = and_dcpl_238 | and_dcpl_255;
  assign COMP_LOOP_mux1h_271_nl = MUX1HOT_v_4_11_2(4'b0101, 4'b0001, 4'b0010, 4'b0100,
      4'b0110, 4'b1000, 4'b1001, 4'b1010, 4'b1100, 4'b1101, 4'b1110, {COMP_LOOP_or_54_nl
      , and_dcpl_242 , and_dcpl_246 , and_dcpl_252 , and_dcpl_260 , and_dcpl_267
      , and_dcpl_272 , and_dcpl_274 , and_dcpl_279 , and_dcpl_281 , and_dcpl_284});
  assign nl_acc_nl = ({COMP_LOOP_COMP_LOOP_or_3_nl , COMP_LOOP_COMP_LOOP_mux_15_nl
      , COMP_LOOP_or_53_nl}) + conv_u2u_10_11({COMP_LOOP_k_9_4_sva_4_0 , COMP_LOOP_mux1h_271_nl
      , 1'b1});
  assign acc_nl = nl_acc_nl[10:0];
  assign z_out_1 = readslicef_11_10_1(acc_nl);
  assign COMP_LOOP_COMP_LOOP_or_4_nl = (VEC_LOOP_j_sva_9_0[9]) | and_dcpl_300 | and_dcpl_308;
  assign COMP_LOOP_or_55_nl = and_dcpl_300 | and_dcpl_308;
  assign COMP_LOOP_COMP_LOOP_mux_16_nl = MUX_v_7_2_2((VEC_LOOP_j_sva_9_0[8:2]), (~
      (STAGE_LOOP_lshift_psp_sva[9:3])), COMP_LOOP_or_55_nl);
  assign COMP_LOOP_or_56_nl = (~ and_dcpl_293) | and_dcpl_300 | and_dcpl_308;
  assign COMP_LOOP_COMP_LOOP_or_5_nl = (~ and_dcpl_300) | and_dcpl_293;
  assign nl_acc_1_nl = ({COMP_LOOP_COMP_LOOP_or_4_nl , COMP_LOOP_COMP_LOOP_mux_16_nl
      , COMP_LOOP_or_56_nl}) + conv_u2u_8_9({COMP_LOOP_k_9_4_sva_4_0 , COMP_LOOP_COMP_LOOP_or_5_nl
      , and_dcpl_293 , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[8:0];
  assign z_out_2 = readslicef_9_8_1(acc_1_nl);
  assign operator_64_false_1_mux_1_nl = MUX_v_5_2_2((~ COMP_LOOP_k_9_4_sva_4_0),
      COMP_LOOP_k_9_4_sva_4_0, and_551_ssc);
  assign nl_z_out_3 = ({(~ and_551_ssc) , operator_64_false_1_mux_1_nl}) + 6'b000001;
  assign z_out_3 = nl_z_out_3[5:0];
  assign COMP_LOOP_mux_35_nl = MUX_v_6_2_2(({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[9:5]))}),
      (VEC_LOOP_j_sva_9_0[9:4]), and_dcpl_344);
  assign COMP_LOOP_COMP_LOOP_nand_1_nl = ~(and_dcpl_344 & (~((fsm_output==10'b1010110111))));
  assign nl_acc_3_nl = ({COMP_LOOP_mux_35_nl , COMP_LOOP_COMP_LOOP_nand_1_nl}) +
      conv_u2u_6_7({COMP_LOOP_k_9_4_sva_4_0 , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[6:0];
  assign z_out_4 = readslicef_7_6_1(acc_3_nl);
  assign COMP_LOOP_mux_36_nl = MUX_v_7_2_2((VEC_LOOP_j_sva_9_0[9:3]), ({1'b1 , (~
      (STAGE_LOOP_lshift_psp_sva[9:4]))}), and_dcpl_361);
  assign COMP_LOOP_or_57_nl = (~(and_dcpl_236 & and_dcpl_234 & nor_761_cse & (~ (fsm_output[0]))
      & (fsm_output[4]))) | and_dcpl_361;
  assign nl_acc_4_nl = ({COMP_LOOP_mux_36_nl , COMP_LOOP_or_57_nl}) + conv_u2u_7_8({COMP_LOOP_k_9_4_sva_4_0
      , (~ and_dcpl_361) , 1'b1});
  assign acc_4_nl = nl_acc_4_nl[7:0];
  assign z_out_5 = readslicef_8_7_1(acc_4_nl);
  assign and_706_nl = and_dcpl_251 & and_dcpl_376 & (~ (fsm_output[5])) & and_dcpl_32;
  assign and_707_nl = and_dcpl_251 & and_dcpl_382 & and_dcpl_29;
  assign and_708_nl = and_dcpl_70 & (~ (fsm_output[3])) & and_dcpl_256 & and_dcpl_232
      & and_dcpl_29;
  assign and_709_nl = and_dcpl_398 & and_dcpl_396;
  assign and_710_nl = and_dcpl_398 & and_dcpl_403;
  assign and_711_nl = and_dcpl_407 & and_dcpl_232 & and_dcpl_66;
  assign and_712_nl = and_dcpl_407 & and_dcpl_244 & and_dcpl_16;
  assign and_713_nl = and_dcpl_265 & and_dcpl_250 & and_dcpl_402 & and_dcpl_66;
  assign and_714_nl = and_dcpl_417 & and_dcpl_382 & and_dcpl_16;
  assign and_715_nl = and_dcpl_417 & and_dcpl_244 & and_dcpl_66;
  assign and_716_nl = and_dcpl_416 & and_dcpl_250 & and_dcpl_232 & and_dcpl_16;
  assign and_717_nl = and_dcpl_425 & and_dcpl_396;
  assign COMP_LOOP_mux1h_272_nl = MUX1HOT_v_4_14_2(4'b1110, 4'b1101, 4'b1100, 4'b1011,
      4'b1010, 4'b1001, 4'b1000, 4'b0111, 4'b0110, 4'b0101, 4'b0100, 4'b0011, 4'b0010,
      4'b0001, {and_dcpl_246 , and_706_nl , and_707_nl , and_dcpl_255 , and_708_nl
      , and_709_nl , and_710_nl , and_711_nl , and_712_nl , and_713_nl , and_714_nl
      , and_715_nl , and_716_nl , and_717_nl});
  assign COMP_LOOP_COMP_LOOP_nor_63_nl = ~(MUX_v_4_2_2(COMP_LOOP_mux1h_272_nl, 4'b1111,
      and_dcpl_242));
  assign and_718_nl = and_dcpl_425 & and_dcpl_403;
  assign COMP_LOOP_or_58_nl = MUX_v_4_2_2(COMP_LOOP_COMP_LOOP_nor_63_nl, 4'b1111,
      and_718_nl);
  assign nl_acc_5_nl = conv_u2u_9_11({COMP_LOOP_k_9_4_sva_4_0 , COMP_LOOP_or_58_nl})
      + conv_u2u_10_11(VEC_LOOP_j_sva_9_0) + conv_u2u_10_11(STAGE_LOOP_lshift_psp_sva);
  assign acc_5_nl = nl_acc_5_nl[10:0];
  assign z_out_6_10_1 = readslicef_11_10_1(acc_5_nl);
  assign STAGE_LOOP_STAGE_LOOP_or_1_nl = (~((fsm_output[9]) & (fsm_output[8]) & (~
      (fsm_output[3])) & and_dcpl_234 & (fsm_output[1]) & (~ (fsm_output[6])) & (~
      (fsm_output[5])) & (~ (fsm_output[0])) & (~ (fsm_output[4])))) | (~ mux_2066_cse)
      | and_dcpl_444;
  assign STAGE_LOOP_or_2_nl = (~ mux_2066_cse) | and_dcpl_444;
  assign STAGE_LOOP_STAGE_LOOP_mux_2_nl = MUX_v_64_2_2(({60'b000000000000000000000000000000000000000000000000000000000000
      , STAGE_LOOP_i_3_0_sva}), (~ (z_out_9[63:0])), STAGE_LOOP_or_2_nl);
  assign nl_z_out_7 = ({STAGE_LOOP_STAGE_LOOP_or_1_nl , STAGE_LOOP_STAGE_LOOP_mux_2_nl})
      + 65'b00000000000000000000000000000000000000000000000000000000000000001;
  assign z_out_7 = nl_z_out_7[64:0];
  assign operator_64_false_operator_64_false_operator_64_false_nor_1_nl = ~(MUX_v_61_2_2((operator_66_true_div_cmp_z[63:3]),
      61'b1111111111111111111111111111111111111111111111111111111111111, and_dcpl_460));
  assign operator_64_false_mux_1_nl = MUX_v_3_2_2((~ (operator_66_true_div_cmp_z[2:0])),
      (z_out_7[3:1]), and_dcpl_460);
  assign nl_operator_64_false_acc_nl = ({(~ and_dcpl_460) , operator_64_false_operator_64_false_operator_64_false_nor_1_nl
      , operator_64_false_mux_1_nl}) + conv_u2u_2_65({and_dcpl_460 , 1'b1});
  assign operator_64_false_acc_nl = nl_operator_64_false_acc_nl[64:0];
  assign z_out_8_64_2 = readslicef_65_63_2(operator_64_false_acc_nl);
  assign and_719_nl = and_dcpl_236 & and_dcpl_256 & and_dcpl_464;
  assign and_720_nl = and_dcpl_236 & (~ (fsm_output[7])) & (fsm_output[2]) & and_dcpl_464;
  assign operator_64_false_mux1h_1_nl = MUX1HOT_v_64_3_2(p_sva, modExp_dev_exp_sva,
      ({modExp_dev_exp_1_sva_63_9 , COMP_LOOP_acc_10_cse_10_1_1_sva_4_0 , modExp_dev_exp_1_sva_3_0}),
      {and_719_nl , and_720_nl , (~ mux_2066_cse)});
  assign nl_z_out_9 = conv_u2u_64_65(operator_64_false_mux1h_1_nl) + 65'b11111111111111111111111111111111111111111111111111111111111111111;
  assign z_out_9 = nl_z_out_9[64:0];

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_11_2;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [10:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    result = result | ( input_5 & {4{sel[5]}});
    result = result | ( input_6 & {4{sel[6]}});
    result = result | ( input_7 & {4{sel[7]}});
    result = result | ( input_8 & {4{sel[8]}});
    result = result | ( input_9 & {4{sel[9]}});
    result = result | ( input_10 & {4{sel[10]}});
    MUX1HOT_v_4_11_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_14_2;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [13:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    result = result | ( input_5 & {4{sel[5]}});
    result = result | ( input_6 & {4{sel[6]}});
    result = result | ( input_7 & {4{sel[7]}});
    result = result | ( input_8 & {4{sel[8]}});
    result = result | ( input_9 & {4{sel[9]}});
    result = result | ( input_10 & {4{sel[10]}});
    result = result | ( input_11 & {4{sel[11]}});
    result = result | ( input_12 & {4{sel[12]}});
    result = result | ( input_13 & {4{sel[13]}});
    MUX1HOT_v_4_14_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_16_2;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [15:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    result = result | ( input_5 & {4{sel[5]}});
    result = result | ( input_6 & {4{sel[6]}});
    result = result | ( input_7 & {4{sel[7]}});
    result = result | ( input_8 & {4{sel[8]}});
    result = result | ( input_9 & {4{sel[9]}});
    result = result | ( input_10 & {4{sel[10]}});
    result = result | ( input_11 & {4{sel[11]}});
    result = result | ( input_12 & {4{sel[12]}});
    result = result | ( input_13 & {4{sel[13]}});
    result = result | ( input_14 & {4{sel[14]}});
    result = result | ( input_15 & {4{sel[15]}});
    MUX1HOT_v_4_16_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_16_2;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [15:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    MUX1HOT_v_64_16_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_4_2;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [3:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    MUX1HOT_v_64_4_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_17_2;
    input [5:0] input_16;
    input [5:0] input_15;
    input [5:0] input_14;
    input [5:0] input_13;
    input [5:0] input_12;
    input [5:0] input_11;
    input [5:0] input_10;
    input [5:0] input_9;
    input [5:0] input_8;
    input [5:0] input_7;
    input [5:0] input_6;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [16:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    result = result | ( input_3 & {6{sel[3]}});
    result = result | ( input_4 & {6{sel[4]}});
    result = result | ( input_5 & {6{sel[5]}});
    result = result | ( input_6 & {6{sel[6]}});
    result = result | ( input_7 & {6{sel[7]}});
    result = result | ( input_8 & {6{sel[8]}});
    result = result | ( input_9 & {6{sel[9]}});
    result = result | ( input_10 & {6{sel[10]}});
    result = result | ( input_11 & {6{sel[11]}});
    result = result | ( input_12 & {6{sel[12]}});
    result = result | ( input_13 & {6{sel[13]}});
    result = result | ( input_14 & {6{sel[14]}});
    result = result | ( input_15 & {6{sel[15]}});
    result = result | ( input_16 & {6{sel[16]}});
    MUX1HOT_v_6_17_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [54:0] MUX_v_55_2_2;
    input [54:0] input_0;
    input [54:0] input_1;
    input [0:0] sel;
    reg [54:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_55_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [60:0] MUX_v_61_2_2;
    input [60:0] input_0;
    input [60:0] input_1;
    input [0:0] sel;
    reg [60:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_61_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [64:0] MUX_v_65_2_2;
    input [64:0] input_0;
    input [64:0] input_1;
    input [0:0] sel;
    reg [64:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_65_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [9:0] readslicef_11_10_1;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_11_10_1 = tmp[9:0];
  end
  endfunction


  function automatic [62:0] readslicef_65_63_2;
    input [64:0] vector;
    reg [64:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_65_63_2 = tmp[62:0];
  end
  endfunction


  function automatic [5:0] readslicef_7_6_1;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_7_6_1 = tmp[5:0];
  end
  endfunction


  function automatic [6:0] readslicef_8_7_1;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_8_7_1 = tmp[6:0];
  end
  endfunction


  function automatic [7:0] readslicef_9_8_1;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_9_8_1 = tmp[7:0];
  end
  endfunction


  function automatic [64:0] conv_u2s_64_65 ;
    input [63:0]  vector ;
  begin
    conv_u2s_64_65 =  {1'b0, vector};
  end
  endfunction


  function automatic [64:0] conv_u2u_2_65 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_65 = {{63{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_11 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [64:0] conv_u2u_64_65 ;
    input [63:0]  vector ;
  begin
    conv_u2u_64_65 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT
// ------------------------------------------------------------------


module inPlaceNTT_DIT (
  clk, rst, vec_rsc_0_0_wadr, vec_rsc_0_0_d, vec_rsc_0_0_we, vec_rsc_0_0_radr, vec_rsc_0_0_q,
      vec_rsc_triosy_0_0_lz, vec_rsc_0_1_wadr, vec_rsc_0_1_d, vec_rsc_0_1_we, vec_rsc_0_1_radr,
      vec_rsc_0_1_q, vec_rsc_triosy_0_1_lz, vec_rsc_0_2_wadr, vec_rsc_0_2_d, vec_rsc_0_2_we,
      vec_rsc_0_2_radr, vec_rsc_0_2_q, vec_rsc_triosy_0_2_lz, vec_rsc_0_3_wadr, vec_rsc_0_3_d,
      vec_rsc_0_3_we, vec_rsc_0_3_radr, vec_rsc_0_3_q, vec_rsc_triosy_0_3_lz, vec_rsc_0_4_wadr,
      vec_rsc_0_4_d, vec_rsc_0_4_we, vec_rsc_0_4_radr, vec_rsc_0_4_q, vec_rsc_triosy_0_4_lz,
      vec_rsc_0_5_wadr, vec_rsc_0_5_d, vec_rsc_0_5_we, vec_rsc_0_5_radr, vec_rsc_0_5_q,
      vec_rsc_triosy_0_5_lz, vec_rsc_0_6_wadr, vec_rsc_0_6_d, vec_rsc_0_6_we, vec_rsc_0_6_radr,
      vec_rsc_0_6_q, vec_rsc_triosy_0_6_lz, vec_rsc_0_7_wadr, vec_rsc_0_7_d, vec_rsc_0_7_we,
      vec_rsc_0_7_radr, vec_rsc_0_7_q, vec_rsc_triosy_0_7_lz, vec_rsc_0_8_wadr, vec_rsc_0_8_d,
      vec_rsc_0_8_we, vec_rsc_0_8_radr, vec_rsc_0_8_q, vec_rsc_triosy_0_8_lz, vec_rsc_0_9_wadr,
      vec_rsc_0_9_d, vec_rsc_0_9_we, vec_rsc_0_9_radr, vec_rsc_0_9_q, vec_rsc_triosy_0_9_lz,
      vec_rsc_0_10_wadr, vec_rsc_0_10_d, vec_rsc_0_10_we, vec_rsc_0_10_radr, vec_rsc_0_10_q,
      vec_rsc_triosy_0_10_lz, vec_rsc_0_11_wadr, vec_rsc_0_11_d, vec_rsc_0_11_we,
      vec_rsc_0_11_radr, vec_rsc_0_11_q, vec_rsc_triosy_0_11_lz, vec_rsc_0_12_wadr,
      vec_rsc_0_12_d, vec_rsc_0_12_we, vec_rsc_0_12_radr, vec_rsc_0_12_q, vec_rsc_triosy_0_12_lz,
      vec_rsc_0_13_wadr, vec_rsc_0_13_d, vec_rsc_0_13_we, vec_rsc_0_13_radr, vec_rsc_0_13_q,
      vec_rsc_triosy_0_13_lz, vec_rsc_0_14_wadr, vec_rsc_0_14_d, vec_rsc_0_14_we,
      vec_rsc_0_14_radr, vec_rsc_0_14_q, vec_rsc_triosy_0_14_lz, vec_rsc_0_15_wadr,
      vec_rsc_0_15_d, vec_rsc_0_15_we, vec_rsc_0_15_radr, vec_rsc_0_15_q, vec_rsc_triosy_0_15_lz,
      p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz
);
  input clk;
  input rst;
  output [5:0] vec_rsc_0_0_wadr;
  output [63:0] vec_rsc_0_0_d;
  output vec_rsc_0_0_we;
  output [5:0] vec_rsc_0_0_radr;
  input [63:0] vec_rsc_0_0_q;
  output vec_rsc_triosy_0_0_lz;
  output [5:0] vec_rsc_0_1_wadr;
  output [63:0] vec_rsc_0_1_d;
  output vec_rsc_0_1_we;
  output [5:0] vec_rsc_0_1_radr;
  input [63:0] vec_rsc_0_1_q;
  output vec_rsc_triosy_0_1_lz;
  output [5:0] vec_rsc_0_2_wadr;
  output [63:0] vec_rsc_0_2_d;
  output vec_rsc_0_2_we;
  output [5:0] vec_rsc_0_2_radr;
  input [63:0] vec_rsc_0_2_q;
  output vec_rsc_triosy_0_2_lz;
  output [5:0] vec_rsc_0_3_wadr;
  output [63:0] vec_rsc_0_3_d;
  output vec_rsc_0_3_we;
  output [5:0] vec_rsc_0_3_radr;
  input [63:0] vec_rsc_0_3_q;
  output vec_rsc_triosy_0_3_lz;
  output [5:0] vec_rsc_0_4_wadr;
  output [63:0] vec_rsc_0_4_d;
  output vec_rsc_0_4_we;
  output [5:0] vec_rsc_0_4_radr;
  input [63:0] vec_rsc_0_4_q;
  output vec_rsc_triosy_0_4_lz;
  output [5:0] vec_rsc_0_5_wadr;
  output [63:0] vec_rsc_0_5_d;
  output vec_rsc_0_5_we;
  output [5:0] vec_rsc_0_5_radr;
  input [63:0] vec_rsc_0_5_q;
  output vec_rsc_triosy_0_5_lz;
  output [5:0] vec_rsc_0_6_wadr;
  output [63:0] vec_rsc_0_6_d;
  output vec_rsc_0_6_we;
  output [5:0] vec_rsc_0_6_radr;
  input [63:0] vec_rsc_0_6_q;
  output vec_rsc_triosy_0_6_lz;
  output [5:0] vec_rsc_0_7_wadr;
  output [63:0] vec_rsc_0_7_d;
  output vec_rsc_0_7_we;
  output [5:0] vec_rsc_0_7_radr;
  input [63:0] vec_rsc_0_7_q;
  output vec_rsc_triosy_0_7_lz;
  output [5:0] vec_rsc_0_8_wadr;
  output [63:0] vec_rsc_0_8_d;
  output vec_rsc_0_8_we;
  output [5:0] vec_rsc_0_8_radr;
  input [63:0] vec_rsc_0_8_q;
  output vec_rsc_triosy_0_8_lz;
  output [5:0] vec_rsc_0_9_wadr;
  output [63:0] vec_rsc_0_9_d;
  output vec_rsc_0_9_we;
  output [5:0] vec_rsc_0_9_radr;
  input [63:0] vec_rsc_0_9_q;
  output vec_rsc_triosy_0_9_lz;
  output [5:0] vec_rsc_0_10_wadr;
  output [63:0] vec_rsc_0_10_d;
  output vec_rsc_0_10_we;
  output [5:0] vec_rsc_0_10_radr;
  input [63:0] vec_rsc_0_10_q;
  output vec_rsc_triosy_0_10_lz;
  output [5:0] vec_rsc_0_11_wadr;
  output [63:0] vec_rsc_0_11_d;
  output vec_rsc_0_11_we;
  output [5:0] vec_rsc_0_11_radr;
  input [63:0] vec_rsc_0_11_q;
  output vec_rsc_triosy_0_11_lz;
  output [5:0] vec_rsc_0_12_wadr;
  output [63:0] vec_rsc_0_12_d;
  output vec_rsc_0_12_we;
  output [5:0] vec_rsc_0_12_radr;
  input [63:0] vec_rsc_0_12_q;
  output vec_rsc_triosy_0_12_lz;
  output [5:0] vec_rsc_0_13_wadr;
  output [63:0] vec_rsc_0_13_d;
  output vec_rsc_0_13_we;
  output [5:0] vec_rsc_0_13_radr;
  input [63:0] vec_rsc_0_13_q;
  output vec_rsc_triosy_0_13_lz;
  output [5:0] vec_rsc_0_14_wadr;
  output [63:0] vec_rsc_0_14_d;
  output vec_rsc_0_14_we;
  output [5:0] vec_rsc_0_14_radr;
  input [63:0] vec_rsc_0_14_q;
  output vec_rsc_triosy_0_14_lz;
  output [5:0] vec_rsc_0_15_wadr;
  output [63:0] vec_rsc_0_15_d;
  output vec_rsc_0_15_we;
  output [5:0] vec_rsc_0_15_radr;
  input [63:0] vec_rsc_0_15_q;
  output vec_rsc_triosy_0_15_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;


  // Interconnect Declarations
  wire [63:0] vec_rsc_0_0_i_q_d;
  wire vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_1_i_q_d;
  wire vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_2_i_q_d;
  wire vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_3_i_q_d;
  wire vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_4_i_q_d;
  wire vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_5_i_q_d;
  wire vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_6_i_q_d;
  wire vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_7_i_q_d;
  wire vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_8_i_q_d;
  wire vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_9_i_q_d;
  wire vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_10_i_q_d;
  wire vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_11_i_q_d;
  wire vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_12_i_q_d;
  wire vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_13_i_q_d;
  wire vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_14_i_q_d;
  wire vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_15_i_q_d;
  wire vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_0_i_d_d_iff;
  wire [5:0] vec_rsc_0_0_i_radr_d_iff;
  wire [5:0] vec_rsc_0_0_i_wadr_d_iff;
  wire vec_rsc_0_0_i_we_d_iff;
  wire vec_rsc_0_1_i_we_d_iff;
  wire vec_rsc_0_2_i_we_d_iff;
  wire vec_rsc_0_3_i_we_d_iff;
  wire vec_rsc_0_4_i_we_d_iff;
  wire vec_rsc_0_5_i_we_d_iff;
  wire vec_rsc_0_6_i_we_d_iff;
  wire vec_rsc_0_7_i_we_d_iff;
  wire vec_rsc_0_8_i_we_d_iff;
  wire vec_rsc_0_9_i_we_d_iff;
  wire vec_rsc_0_10_i_we_d_iff;
  wire vec_rsc_0_11_i_we_d_iff;
  wire vec_rsc_0_12_i_we_d_iff;
  wire vec_rsc_0_13_i_we_d_iff;
  wire vec_rsc_0_14_i_we_d_iff;
  wire vec_rsc_0_15_i_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_6_64_64_64_64_1_gen vec_rsc_0_0_i
      (
      .q(vec_rsc_0_0_q),
      .radr(vec_rsc_0_0_radr),
      .we(vec_rsc_0_0_we),
      .d(vec_rsc_0_0_d),
      .wadr(vec_rsc_0_0_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_0_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen vec_rsc_0_1_i
      (
      .q(vec_rsc_0_1_q),
      .radr(vec_rsc_0_1_radr),
      .we(vec_rsc_0_1_we),
      .d(vec_rsc_0_1_d),
      .wadr(vec_rsc_0_1_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_1_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_1_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_1_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen vec_rsc_0_2_i
      (
      .q(vec_rsc_0_2_q),
      .radr(vec_rsc_0_2_radr),
      .we(vec_rsc_0_2_we),
      .d(vec_rsc_0_2_d),
      .wadr(vec_rsc_0_2_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_2_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_2_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_2_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen vec_rsc_0_3_i
      (
      .q(vec_rsc_0_3_q),
      .radr(vec_rsc_0_3_radr),
      .we(vec_rsc_0_3_we),
      .d(vec_rsc_0_3_d),
      .wadr(vec_rsc_0_3_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_3_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_3_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_3_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen vec_rsc_0_4_i
      (
      .q(vec_rsc_0_4_q),
      .radr(vec_rsc_0_4_radr),
      .we(vec_rsc_0_4_we),
      .d(vec_rsc_0_4_d),
      .wadr(vec_rsc_0_4_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_4_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_4_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_4_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen vec_rsc_0_5_i
      (
      .q(vec_rsc_0_5_q),
      .radr(vec_rsc_0_5_radr),
      .we(vec_rsc_0_5_we),
      .d(vec_rsc_0_5_d),
      .wadr(vec_rsc_0_5_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_5_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_5_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_5_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen vec_rsc_0_6_i
      (
      .q(vec_rsc_0_6_q),
      .radr(vec_rsc_0_6_radr),
      .we(vec_rsc_0_6_we),
      .d(vec_rsc_0_6_d),
      .wadr(vec_rsc_0_6_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_6_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_6_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_6_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen vec_rsc_0_7_i
      (
      .q(vec_rsc_0_7_q),
      .radr(vec_rsc_0_7_radr),
      .we(vec_rsc_0_7_we),
      .d(vec_rsc_0_7_d),
      .wadr(vec_rsc_0_7_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_7_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_7_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_7_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen vec_rsc_0_8_i
      (
      .q(vec_rsc_0_8_q),
      .radr(vec_rsc_0_8_radr),
      .we(vec_rsc_0_8_we),
      .d(vec_rsc_0_8_d),
      .wadr(vec_rsc_0_8_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_8_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_8_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_8_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen vec_rsc_0_9_i
      (
      .q(vec_rsc_0_9_q),
      .radr(vec_rsc_0_9_radr),
      .we(vec_rsc_0_9_we),
      .d(vec_rsc_0_9_d),
      .wadr(vec_rsc_0_9_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_9_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_9_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_9_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen vec_rsc_0_10_i
      (
      .q(vec_rsc_0_10_q),
      .radr(vec_rsc_0_10_radr),
      .we(vec_rsc_0_10_we),
      .d(vec_rsc_0_10_d),
      .wadr(vec_rsc_0_10_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_10_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_10_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_10_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen vec_rsc_0_11_i
      (
      .q(vec_rsc_0_11_q),
      .radr(vec_rsc_0_11_radr),
      .we(vec_rsc_0_11_we),
      .d(vec_rsc_0_11_d),
      .wadr(vec_rsc_0_11_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_11_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_11_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_11_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen vec_rsc_0_12_i
      (
      .q(vec_rsc_0_12_q),
      .radr(vec_rsc_0_12_radr),
      .we(vec_rsc_0_12_we),
      .d(vec_rsc_0_12_d),
      .wadr(vec_rsc_0_12_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_12_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_12_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_12_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen vec_rsc_0_13_i
      (
      .q(vec_rsc_0_13_q),
      .radr(vec_rsc_0_13_radr),
      .we(vec_rsc_0_13_we),
      .d(vec_rsc_0_13_d),
      .wadr(vec_rsc_0_13_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_13_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_13_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_13_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen vec_rsc_0_14_i
      (
      .q(vec_rsc_0_14_q),
      .radr(vec_rsc_0_14_radr),
      .we(vec_rsc_0_14_we),
      .d(vec_rsc_0_14_d),
      .wadr(vec_rsc_0_14_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_14_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_14_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_14_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen vec_rsc_0_15_i
      (
      .q(vec_rsc_0_15_q),
      .radr(vec_rsc_0_15_radr),
      .we(vec_rsc_0_15_we),
      .d(vec_rsc_0_15_d),
      .wadr(vec_rsc_0_15_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_15_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_15_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_15_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIT_core inPlaceNTT_DIT_core_inst (
      .clk(clk),
      .rst(rst),
      .vec_rsc_triosy_0_0_lz(vec_rsc_triosy_0_0_lz),
      .vec_rsc_triosy_0_1_lz(vec_rsc_triosy_0_1_lz),
      .vec_rsc_triosy_0_2_lz(vec_rsc_triosy_0_2_lz),
      .vec_rsc_triosy_0_3_lz(vec_rsc_triosy_0_3_lz),
      .vec_rsc_triosy_0_4_lz(vec_rsc_triosy_0_4_lz),
      .vec_rsc_triosy_0_5_lz(vec_rsc_triosy_0_5_lz),
      .vec_rsc_triosy_0_6_lz(vec_rsc_triosy_0_6_lz),
      .vec_rsc_triosy_0_7_lz(vec_rsc_triosy_0_7_lz),
      .vec_rsc_triosy_0_8_lz(vec_rsc_triosy_0_8_lz),
      .vec_rsc_triosy_0_9_lz(vec_rsc_triosy_0_9_lz),
      .vec_rsc_triosy_0_10_lz(vec_rsc_triosy_0_10_lz),
      .vec_rsc_triosy_0_11_lz(vec_rsc_triosy_0_11_lz),
      .vec_rsc_triosy_0_12_lz(vec_rsc_triosy_0_12_lz),
      .vec_rsc_triosy_0_13_lz(vec_rsc_triosy_0_13_lz),
      .vec_rsc_triosy_0_14_lz(vec_rsc_triosy_0_14_lz),
      .vec_rsc_triosy_0_15_lz(vec_rsc_triosy_0_15_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_dat(r_rsc_dat),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .vec_rsc_0_0_i_q_d(vec_rsc_0_0_i_q_d),
      .vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_1_i_q_d(vec_rsc_0_1_i_q_d),
      .vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_2_i_q_d(vec_rsc_0_2_i_q_d),
      .vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_3_i_q_d(vec_rsc_0_3_i_q_d),
      .vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_4_i_q_d(vec_rsc_0_4_i_q_d),
      .vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_5_i_q_d(vec_rsc_0_5_i_q_d),
      .vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_6_i_q_d(vec_rsc_0_6_i_q_d),
      .vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_7_i_q_d(vec_rsc_0_7_i_q_d),
      .vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_8_i_q_d(vec_rsc_0_8_i_q_d),
      .vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_9_i_q_d(vec_rsc_0_9_i_q_d),
      .vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_10_i_q_d(vec_rsc_0_10_i_q_d),
      .vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_11_i_q_d(vec_rsc_0_11_i_q_d),
      .vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_12_i_q_d(vec_rsc_0_12_i_q_d),
      .vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_13_i_q_d(vec_rsc_0_13_i_q_d),
      .vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_14_i_q_d(vec_rsc_0_14_i_q_d),
      .vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_15_i_q_d(vec_rsc_0_15_i_q_d),
      .vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_0_i_d_d_pff(vec_rsc_0_0_i_d_d_iff),
      .vec_rsc_0_0_i_radr_d_pff(vec_rsc_0_0_i_radr_d_iff),
      .vec_rsc_0_0_i_wadr_d_pff(vec_rsc_0_0_i_wadr_d_iff),
      .vec_rsc_0_0_i_we_d_pff(vec_rsc_0_0_i_we_d_iff),
      .vec_rsc_0_1_i_we_d_pff(vec_rsc_0_1_i_we_d_iff),
      .vec_rsc_0_2_i_we_d_pff(vec_rsc_0_2_i_we_d_iff),
      .vec_rsc_0_3_i_we_d_pff(vec_rsc_0_3_i_we_d_iff),
      .vec_rsc_0_4_i_we_d_pff(vec_rsc_0_4_i_we_d_iff),
      .vec_rsc_0_5_i_we_d_pff(vec_rsc_0_5_i_we_d_iff),
      .vec_rsc_0_6_i_we_d_pff(vec_rsc_0_6_i_we_d_iff),
      .vec_rsc_0_7_i_we_d_pff(vec_rsc_0_7_i_we_d_iff),
      .vec_rsc_0_8_i_we_d_pff(vec_rsc_0_8_i_we_d_iff),
      .vec_rsc_0_9_i_we_d_pff(vec_rsc_0_9_i_we_d_iff),
      .vec_rsc_0_10_i_we_d_pff(vec_rsc_0_10_i_we_d_iff),
      .vec_rsc_0_11_i_we_d_pff(vec_rsc_0_11_i_we_d_iff),
      .vec_rsc_0_12_i_we_d_pff(vec_rsc_0_12_i_we_d_iff),
      .vec_rsc_0_13_i_we_d_pff(vec_rsc_0_13_i_we_d_iff),
      .vec_rsc_0_14_i_we_d_pff(vec_rsc_0_14_i_we_d_iff),
      .vec_rsc_0_15_i_we_d_pff(vec_rsc_0_15_i_we_d_iff)
    );
endmodule



