
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.v 
module mgc_rem(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_b-1:0] z;  
   reg  [width_b-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  rem_s(a,b,z);
	else
          rem_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> ../td_ccore_solutions/modulo_dev_d3e65941ee7586d7daaa2e36d0d005555a5b_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Thu Aug 26 01:37:26 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    modulo_dev_core
// ------------------------------------------------------------------


module modulo_dev_core (
  base_rsc_dat, m_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [63:0] base_rsc_dat;
  input [63:0] m_rsc_dat;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [63:0] base_rsci_idat;
  wire [63:0] m_rsci_idat;
  reg [63:0] return_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  reg [63:0] result_rem_12_cmp_a;
  reg [63:0] result_rem_12_cmp_b;
  wire [63:0] result_rem_12_cmp_z;
  reg [63:0] result_rem_12_cmp_1_a;
  reg [63:0] result_rem_12_cmp_1_b;
  wire [63:0] result_rem_12_cmp_1_z;
  reg [63:0] result_rem_12_cmp_2_a;
  reg [63:0] result_rem_12_cmp_2_b;
  wire [63:0] result_rem_12_cmp_2_z;
  reg [63:0] result_rem_12_cmp_3_a;
  reg [63:0] result_rem_12_cmp_3_b;
  wire [63:0] result_rem_12_cmp_3_z;
  reg [63:0] result_rem_12_cmp_4_a;
  reg [63:0] result_rem_12_cmp_4_b;
  wire [63:0] result_rem_12_cmp_4_z;
  reg [63:0] result_rem_12_cmp_5_a;
  reg [63:0] result_rem_12_cmp_5_b;
  wire [63:0] result_rem_12_cmp_5_z;
  reg [63:0] result_rem_12_cmp_6_a;
  reg [63:0] result_rem_12_cmp_6_b;
  wire [63:0] result_rem_12_cmp_6_z;
  reg [63:0] result_rem_12_cmp_7_a;
  reg [63:0] result_rem_12_cmp_7_b;
  wire [63:0] result_rem_12_cmp_7_z;
  reg [63:0] result_rem_12_cmp_8_a;
  reg [63:0] result_rem_12_cmp_8_b;
  wire [63:0] result_rem_12_cmp_8_z;
  reg [63:0] result_rem_12_cmp_9_a;
  reg [63:0] result_rem_12_cmp_9_b;
  wire [63:0] result_rem_12_cmp_9_z;
  reg [63:0] result_rem_12_cmp_10_a;
  reg [63:0] result_rem_12_cmp_10_b;
  wire [63:0] result_rem_12_cmp_10_z;
  wire [3:0] result_result_acc_tmp;
  wire [4:0] nl_result_result_acc_tmp;
  wire and_dcpl_1;
  wire and_dcpl_2;
  wire and_dcpl_3;
  wire and_dcpl_4;
  wire and_dcpl_6;
  wire and_dcpl_8;
  wire and_dcpl_9;
  wire and_dcpl_11;
  wire and_dcpl_13;
  wire and_dcpl_18;
  wire and_dcpl_26;
  wire and_dcpl_27;
  wire and_dcpl_28;
  wire and_dcpl_29;
  wire and_dcpl_30;
  wire and_dcpl_31;
  wire and_dcpl_32;
  wire and_dcpl_33;
  wire and_dcpl_34;
  wire and_dcpl_35;
  wire and_dcpl_36;
  wire and_dcpl_37;
  wire and_dcpl_38;
  wire and_dcpl_39;
  wire and_dcpl_40;
  wire and_dcpl_41;
  wire and_dcpl_42;
  wire and_dcpl_43;
  wire and_dcpl_45;
  wire and_dcpl_47;
  wire and_dcpl_50;
  wire and_dcpl_51;
  wire and_dcpl_52;
  wire and_dcpl_53;
  wire and_dcpl_54;
  wire and_dcpl_55;
  wire and_dcpl_56;
  wire and_dcpl_57;
  wire and_dcpl_58;
  wire and_dcpl_59;
  wire and_dcpl_60;
  wire and_dcpl_62;
  wire and_dcpl_63;
  wire and_dcpl_65;
  wire and_dcpl_66;
  wire and_dcpl_68;
  wire and_dcpl_70;
  wire and_dcpl_72;
  wire and_dcpl_73;
  wire and_dcpl_74;
  wire and_dcpl_75;
  wire and_dcpl_76;
  wire and_dcpl_77;
  wire and_dcpl_78;
  wire and_dcpl_79;
  wire and_dcpl_80;
  wire and_dcpl_81;
  wire and_dcpl_82;
  wire and_dcpl_83;
  wire and_dcpl_84;
  wire and_dcpl_85;
  wire and_dcpl_86;
  wire and_dcpl_88;
  wire and_dcpl_89;
  wire and_dcpl_91;
  wire and_dcpl_92;
  wire and_dcpl_94;
  wire and_dcpl_96;
  wire and_dcpl_98;
  wire and_dcpl_99;
  wire and_dcpl_100;
  wire and_dcpl_101;
  wire and_dcpl_102;
  wire and_dcpl_103;
  wire and_dcpl_104;
  wire and_dcpl_105;
  wire and_dcpl_106;
  wire and_dcpl_107;
  wire and_dcpl_108;
  wire and_dcpl_109;
  wire and_dcpl_110;
  wire and_dcpl_111;
  wire and_dcpl_112;
  wire and_dcpl_113;
  wire and_dcpl_114;
  wire and_dcpl_115;
  wire and_dcpl_116;
  wire and_dcpl_117;
  wire and_dcpl_118;
  wire and_dcpl_119;
  wire and_dcpl_120;
  wire and_dcpl_122;
  wire and_dcpl_125;
  wire and_dcpl_127;
  wire and_dcpl_128;
  wire and_dcpl_129;
  wire and_dcpl_130;
  wire and_dcpl_131;
  wire and_dcpl_132;
  wire and_dcpl_133;
  wire and_dcpl_134;
  wire and_dcpl_135;
  wire and_dcpl_136;
  wire and_dcpl_137;
  wire and_dcpl_139;
  wire and_dcpl_140;
  wire and_dcpl_142;
  wire and_dcpl_143;
  wire and_dcpl_145;
  wire and_dcpl_147;
  wire and_dcpl_149;
  wire and_dcpl_150;
  wire and_dcpl_151;
  wire and_dcpl_152;
  wire and_dcpl_153;
  wire and_dcpl_154;
  wire and_dcpl_155;
  wire and_dcpl_156;
  wire and_dcpl_157;
  wire and_dcpl_158;
  wire and_dcpl_159;
  wire and_dcpl_160;
  wire and_dcpl_161;
  wire and_dcpl_162;
  wire and_dcpl_163;
  wire and_dcpl_165;
  wire and_dcpl_166;
  wire and_dcpl_168;
  wire and_dcpl_170;
  wire and_dcpl_171;
  wire and_dcpl_173;
  wire and_dcpl_175;
  wire and_dcpl_176;
  wire and_dcpl_177;
  wire and_dcpl_178;
  wire and_dcpl_179;
  wire and_dcpl_180;
  wire and_dcpl_181;
  wire and_dcpl_182;
  wire and_dcpl_183;
  wire and_dcpl_184;
  wire and_dcpl_185;
  wire and_dcpl_186;
  wire and_dcpl_187;
  wire and_dcpl_188;
  wire and_dcpl_189;
  wire and_dcpl_191;
  wire and_dcpl_192;
  wire and_dcpl_194;
  wire and_dcpl_196;
  wire and_dcpl_197;
  wire and_dcpl_199;
  wire and_dcpl_201;
  wire and_dcpl_202;
  wire and_dcpl_203;
  wire and_dcpl_204;
  wire and_dcpl_205;
  wire and_dcpl_206;
  wire and_dcpl_207;
  wire and_dcpl_208;
  wire and_dcpl_209;
  wire and_dcpl_211;
  wire and_dcpl_212;
  wire and_dcpl_214;
  wire and_dcpl_218;
  wire and_dcpl_221;
  wire and_dcpl_228;
  wire and_dcpl_232;
  wire and_dcpl_233;
  wire and_dcpl_234;
  wire and_dcpl_235;
  wire and_dcpl_237;
  wire and_dcpl_239;
  wire and_dcpl_240;
  wire and_dcpl_244;
  wire and_dcpl_249;
  wire and_dcpl_254;
  wire and_dcpl_260;
  wire and_dcpl_261;
  wire and_dcpl_262;
  wire and_dcpl_263;
  wire or_tmp_2;
  wire and_dcpl_269;
  wire mux_tmp_1;
  wire and_dcpl_275;
  wire mux_tmp_3;
  wire mux_tmp_4;
  wire and_dcpl_281;
  wire mux_tmp_6;
  wire mux_tmp_7;
  wire mux_tmp_8;
  wire and_dcpl_287;
  wire mux_tmp_10;
  wire mux_tmp_11;
  wire mux_tmp_12;
  wire mux_tmp_13;
  wire and_dcpl_293;
  wire mux_tmp_15;
  wire mux_tmp_16;
  wire mux_tmp_17;
  wire mux_tmp_18;
  wire mux_tmp_19;
  wire and_dcpl_299;
  wire mux_tmp_21;
  wire mux_tmp_22;
  wire mux_tmp_23;
  wire mux_tmp_24;
  wire mux_tmp_25;
  wire mux_tmp_26;
  wire and_dcpl_305;
  wire mux_tmp_28;
  wire mux_tmp_29;
  wire mux_tmp_30;
  wire mux_tmp_31;
  wire mux_tmp_32;
  wire mux_tmp_33;
  wire mux_tmp_34;
  wire and_dcpl_311;
  wire and_tmp_6;
  wire mux_tmp_36;
  wire mux_tmp_37;
  wire and_dcpl_318;
  wire and_dcpl_319;
  wire or_tmp_102;
  wire and_dcpl_322;
  wire mux_tmp_39;
  wire and_dcpl_325;
  wire mux_tmp_41;
  wire mux_tmp_42;
  wire and_dcpl_329;
  wire mux_tmp_44;
  wire mux_tmp_45;
  wire mux_tmp_46;
  wire and_dcpl_333;
  wire mux_tmp_48;
  wire mux_tmp_49;
  wire mux_tmp_50;
  wire mux_tmp_51;
  wire and_dcpl_337;
  wire mux_tmp_53;
  wire mux_tmp_54;
  wire mux_tmp_55;
  wire mux_tmp_56;
  wire mux_tmp_57;
  wire and_dcpl_341;
  wire mux_tmp_59;
  wire mux_tmp_60;
  wire mux_tmp_61;
  wire mux_tmp_62;
  wire mux_tmp_63;
  wire mux_tmp_64;
  wire and_dcpl_344;
  wire mux_tmp_66;
  wire mux_tmp_67;
  wire mux_tmp_68;
  wire mux_tmp_69;
  wire mux_tmp_70;
  wire mux_tmp_71;
  wire mux_tmp_72;
  wire and_dcpl_347;
  wire and_tmp_13;
  wire mux_tmp_74;
  wire mux_tmp_75;
  wire and_dcpl_352;
  wire and_dcpl_353;
  wire or_tmp_202;
  wire and_dcpl_357;
  wire mux_tmp_77;
  wire and_dcpl_361;
  wire mux_tmp_79;
  wire mux_tmp_80;
  wire and_dcpl_364;
  wire mux_tmp_82;
  wire mux_tmp_83;
  wire mux_tmp_84;
  wire and_dcpl_367;
  wire mux_tmp_86;
  wire mux_tmp_87;
  wire mux_tmp_88;
  wire mux_tmp_89;
  wire and_dcpl_370;
  wire mux_tmp_91;
  wire mux_tmp_92;
  wire mux_tmp_93;
  wire mux_tmp_94;
  wire mux_tmp_95;
  wire and_dcpl_373;
  wire mux_tmp_97;
  wire mux_tmp_98;
  wire mux_tmp_99;
  wire mux_tmp_100;
  wire mux_tmp_101;
  wire mux_tmp_102;
  wire and_dcpl_377;
  wire mux_tmp_104;
  wire mux_tmp_105;
  wire mux_tmp_106;
  wire mux_tmp_107;
  wire mux_tmp_108;
  wire mux_tmp_109;
  wire mux_tmp_110;
  wire and_dcpl_381;
  wire and_tmp_20;
  wire mux_tmp_112;
  wire mux_tmp_113;
  wire and_dcpl_386;
  wire and_dcpl_387;
  wire or_tmp_302;
  wire and_dcpl_390;
  wire mux_tmp_115;
  wire and_dcpl_393;
  wire mux_tmp_117;
  wire mux_tmp_118;
  wire and_dcpl_396;
  wire mux_tmp_120;
  wire mux_tmp_121;
  wire mux_tmp_122;
  wire and_dcpl_399;
  wire mux_tmp_124;
  wire mux_tmp_125;
  wire mux_tmp_126;
  wire mux_tmp_127;
  wire and_dcpl_402;
  wire mux_tmp_129;
  wire mux_tmp_130;
  wire mux_tmp_131;
  wire mux_tmp_132;
  wire mux_tmp_133;
  wire and_dcpl_405;
  wire mux_tmp_135;
  wire mux_tmp_136;
  wire mux_tmp_137;
  wire mux_tmp_138;
  wire mux_tmp_139;
  wire mux_tmp_140;
  wire and_dcpl_408;
  wire mux_tmp_142;
  wire mux_tmp_143;
  wire mux_tmp_144;
  wire mux_tmp_145;
  wire mux_tmp_146;
  wire mux_tmp_147;
  wire mux_tmp_148;
  wire and_dcpl_411;
  wire and_tmp_27;
  wire mux_tmp_150;
  wire mux_tmp_151;
  wire and_dcpl_417;
  wire and_dcpl_418;
  wire or_tmp_402;
  wire and_dcpl_422;
  wire mux_tmp_153;
  wire and_dcpl_426;
  wire mux_tmp_155;
  wire mux_tmp_156;
  wire and_dcpl_430;
  wire mux_tmp_158;
  wire mux_tmp_159;
  wire mux_tmp_160;
  wire and_dcpl_433;
  wire mux_tmp_162;
  wire mux_tmp_163;
  wire mux_tmp_164;
  wire mux_tmp_165;
  wire and_dcpl_437;
  wire mux_tmp_167;
  wire mux_tmp_168;
  wire mux_tmp_169;
  wire mux_tmp_170;
  wire mux_tmp_171;
  wire and_dcpl_441;
  wire mux_tmp_173;
  wire mux_tmp_174;
  wire mux_tmp_175;
  wire mux_tmp_176;
  wire mux_tmp_177;
  wire mux_tmp_178;
  wire and_dcpl_444;
  wire mux_tmp_180;
  wire mux_tmp_181;
  wire mux_tmp_182;
  wire mux_tmp_183;
  wire mux_tmp_184;
  wire mux_tmp_185;
  wire mux_tmp_186;
  wire and_dcpl_447;
  wire and_tmp_34;
  wire mux_tmp_188;
  wire mux_tmp_189;
  wire and_dcpl_452;
  wire or_tmp_502;
  wire and_dcpl_455;
  wire mux_tmp_191;
  wire and_dcpl_458;
  wire mux_tmp_193;
  wire mux_tmp_194;
  wire and_dcpl_462;
  wire mux_tmp_196;
  wire mux_tmp_197;
  wire mux_tmp_198;
  wire and_dcpl_464;
  wire mux_tmp_200;
  wire mux_tmp_201;
  wire mux_tmp_202;
  wire mux_tmp_203;
  wire and_dcpl_468;
  wire mux_tmp_205;
  wire mux_tmp_206;
  wire mux_tmp_207;
  wire mux_tmp_208;
  wire mux_tmp_209;
  wire and_dcpl_472;
  wire mux_tmp_211;
  wire mux_tmp_212;
  wire mux_tmp_213;
  wire mux_tmp_214;
  wire mux_tmp_215;
  wire mux_tmp_216;
  wire and_dcpl_474;
  wire mux_tmp_218;
  wire mux_tmp_219;
  wire mux_tmp_220;
  wire mux_tmp_221;
  wire mux_tmp_222;
  wire mux_tmp_223;
  wire mux_tmp_224;
  wire and_dcpl_476;
  wire and_tmp_41;
  wire mux_tmp_226;
  wire mux_tmp_227;
  wire and_dcpl_480;
  wire or_tmp_602;
  wire and_dcpl_484;
  wire mux_tmp_229;
  wire and_dcpl_488;
  wire mux_tmp_231;
  wire mux_tmp_232;
  wire and_dcpl_491;
  wire mux_tmp_234;
  wire mux_tmp_235;
  wire mux_tmp_236;
  wire and_dcpl_493;
  wire mux_tmp_238;
  wire mux_tmp_239;
  wire mux_tmp_240;
  wire mux_tmp_241;
  wire and_dcpl_496;
  wire mux_tmp_243;
  wire mux_tmp_244;
  wire mux_tmp_245;
  wire mux_tmp_246;
  wire mux_tmp_247;
  wire and_dcpl_499;
  wire mux_tmp_249;
  wire mux_tmp_250;
  wire mux_tmp_251;
  wire mux_tmp_252;
  wire mux_tmp_253;
  wire mux_tmp_254;
  wire and_dcpl_501;
  wire mux_tmp_256;
  wire mux_tmp_257;
  wire mux_tmp_258;
  wire mux_tmp_259;
  wire mux_tmp_260;
  wire mux_tmp_261;
  wire mux_tmp_262;
  wire and_dcpl_503;
  wire and_tmp_48;
  wire mux_tmp_264;
  wire mux_tmp_265;
  wire and_dcpl_507;
  wire or_tmp_702;
  wire and_dcpl_510;
  wire mux_tmp_267;
  wire and_dcpl_513;
  wire mux_tmp_269;
  wire mux_tmp_270;
  wire and_dcpl_516;
  wire mux_tmp_272;
  wire mux_tmp_273;
  wire mux_tmp_274;
  wire and_dcpl_518;
  wire mux_tmp_276;
  wire mux_tmp_277;
  wire mux_tmp_278;
  wire mux_tmp_279;
  wire and_dcpl_521;
  wire mux_tmp_281;
  wire mux_tmp_282;
  wire mux_tmp_283;
  wire mux_tmp_284;
  wire mux_tmp_285;
  wire and_dcpl_524;
  wire mux_tmp_287;
  wire mux_tmp_288;
  wire mux_tmp_289;
  wire mux_tmp_290;
  wire mux_tmp_291;
  wire mux_tmp_292;
  wire and_dcpl_526;
  wire mux_tmp_294;
  wire mux_tmp_295;
  wire mux_tmp_296;
  wire mux_tmp_297;
  wire mux_tmp_298;
  wire mux_tmp_299;
  wire mux_tmp_300;
  wire and_dcpl_528;
  wire and_tmp_55;
  wire mux_tmp_302;
  wire mux_tmp_303;
  wire and_dcpl_532;
  wire and_dcpl_533;
  wire not_tmp_645;
  wire or_tmp_801;
  wire and_dcpl_536;
  wire mux_tmp_305;
  wire and_dcpl_539;
  wire mux_tmp_307;
  wire mux_tmp_308;
  wire and_dcpl_542;
  wire mux_tmp_310;
  wire mux_tmp_311;
  wire mux_tmp_312;
  wire and_dcpl_546;
  wire mux_tmp_314;
  wire mux_tmp_315;
  wire mux_tmp_316;
  wire mux_tmp_317;
  wire and_dcpl_549;
  wire mux_tmp_319;
  wire mux_tmp_320;
  wire mux_tmp_321;
  wire mux_tmp_322;
  wire mux_tmp_323;
  wire and_dcpl_552;
  wire mux_tmp_325;
  wire mux_tmp_326;
  wire mux_tmp_327;
  wire mux_tmp_328;
  wire mux_tmp_329;
  wire mux_tmp_330;
  wire and_dcpl_556;
  wire mux_tmp_332;
  wire mux_tmp_333;
  wire mux_tmp_334;
  wire mux_tmp_335;
  wire mux_tmp_336;
  wire mux_tmp_337;
  wire mux_tmp_338;
  wire and_dcpl_560;
  wire or_tmp_897;
  wire mux_tmp_340;
  wire mux_tmp_341;
  wire mux_tmp_342;
  wire mux_tmp_343;
  wire mux_tmp_344;
  wire mux_tmp_345;
  wire mux_tmp_346;
  wire mux_tmp_347;
  wire mux_tmp_348;
  wire and_dcpl_566;
  wire or_tmp_909;
  wire and_dcpl_568;
  wire mux_tmp_350;
  wire and_dcpl_570;
  wire mux_tmp_352;
  wire mux_tmp_353;
  wire and_dcpl_572;
  wire mux_tmp_355;
  wire mux_tmp_356;
  wire mux_tmp_357;
  wire and_dcpl_576;
  wire mux_tmp_359;
  wire mux_tmp_360;
  wire mux_tmp_361;
  wire mux_tmp_362;
  wire and_dcpl_578;
  wire mux_tmp_364;
  wire mux_tmp_365;
  wire mux_tmp_366;
  wire mux_tmp_367;
  wire mux_tmp_368;
  wire and_dcpl_580;
  wire mux_tmp_370;
  wire mux_tmp_371;
  wire mux_tmp_372;
  wire mux_tmp_373;
  wire mux_tmp_374;
  wire mux_tmp_375;
  wire and_dcpl_583;
  wire mux_tmp_377;
  wire mux_tmp_378;
  wire mux_tmp_379;
  wire mux_tmp_380;
  wire mux_tmp_381;
  wire mux_tmp_382;
  wire mux_tmp_383;
  wire and_dcpl_586;
  wire or_tmp_1005;
  wire mux_tmp_385;
  wire mux_tmp_386;
  wire mux_tmp_387;
  wire mux_tmp_388;
  wire mux_tmp_389;
  wire mux_tmp_390;
  wire mux_tmp_391;
  wire mux_tmp_392;
  wire mux_tmp_393;
  wire and_dcpl_590;
  wire or_tmp_1017;
  wire and_dcpl_592;
  wire mux_tmp_395;
  wire and_dcpl_594;
  wire mux_tmp_397;
  wire mux_tmp_398;
  wire and_dcpl_596;
  wire mux_tmp_400;
  wire mux_tmp_401;
  wire mux_tmp_402;
  wire and_dcpl_599;
  wire mux_tmp_404;
  wire mux_tmp_405;
  wire mux_tmp_406;
  wire mux_tmp_407;
  wire and_dcpl_601;
  wire mux_tmp_409;
  wire mux_tmp_410;
  wire mux_tmp_411;
  wire mux_tmp_412;
  wire mux_tmp_413;
  wire and_dcpl_603;
  wire mux_tmp_415;
  wire mux_tmp_416;
  wire mux_tmp_417;
  wire mux_tmp_418;
  wire mux_tmp_419;
  wire mux_tmp_420;
  wire and_dcpl_607;
  wire mux_tmp_422;
  wire mux_tmp_423;
  wire mux_tmp_424;
  wire mux_tmp_425;
  wire mux_tmp_426;
  wire mux_tmp_427;
  wire mux_tmp_428;
  wire and_dcpl_611;
  wire or_tmp_1113;
  wire mux_tmp_430;
  wire mux_tmp_431;
  wire mux_tmp_432;
  wire mux_tmp_433;
  wire mux_tmp_434;
  wire mux_tmp_435;
  wire mux_tmp_436;
  wire mux_tmp_437;
  wire mux_tmp_438;
  reg main_stage_0_11;
  reg asn_itm_10;
  reg [3:0] result_rem_11cyc_st_9;
  reg [3:0] result_rem_11cyc_st_8;
  reg [3:0] result_rem_11cyc_st_7;
  reg [3:0] result_rem_11cyc_st_6;
  reg [3:0] result_rem_11cyc_st_5;
  reg [3:0] result_rem_11cyc_st_4;
  reg [3:0] result_rem_11cyc_st_3;
  reg [3:0] result_rem_11cyc_st_2;
  reg [3:0] result_rem_11cyc;
  reg [3:0] result_rem_11cyc_st_11;
  reg asn_itm_11;
  reg main_stage_0_12;
  reg main_stage_0_3;
  reg asn_itm_2;
  reg main_stage_0_4;
  reg asn_itm_3;
  reg main_stage_0_5;
  reg asn_itm_4;
  reg main_stage_0_6;
  reg asn_itm_5;
  reg main_stage_0_7;
  reg asn_itm_6;
  reg main_stage_0_8;
  reg asn_itm_7;
  reg main_stage_0_9;
  reg asn_itm_8;
  reg main_stage_0_10;
  reg asn_itm_9;
  reg main_stage_0_2;
  reg asn_itm_1;
  wire result_and_1_cse;
  wire result_and_3_cse;
  wire result_and_5_cse;
  wire result_and_7_cse;
  wire result_and_9_cse;
  wire result_and_11_cse;
  wire result_and_13_cse;
  wire result_and_15_cse;
  wire result_and_17_cse;
  wire result_and_19_cse;
  wire result_and_21_cse;
  wire or_3_cse;
  wire or_8_cse;
  wire or_15_cse;
  wire or_24_cse;
  wire or_35_cse;
  wire or_48_cse;
  wire or_63_cse;
  wire or_107_cse;
  wire or_112_cse;
  wire or_119_cse;
  wire or_128_cse;
  wire or_139_cse;
  wire or_152_cse;
  wire or_167_cse;
  wire or_209_cse;
  wire or_214_cse;
  wire or_221_cse;
  wire or_230_cse;
  wire or_241_cse;
  wire or_254_cse;
  wire or_269_cse;
  wire or_311_cse;
  wire or_316_cse;
  wire or_323_cse;
  wire or_332_cse;
  wire or_343_cse;
  wire or_356_cse;
  wire or_371_cse;
  wire nand_144_cse;
  wire or_413_cse;
  wire or_418_cse;
  wire or_425_cse;
  wire or_434_cse;
  wire or_445_cse;
  wire or_458_cse;
  wire or_473_cse;
  wire nand_138_cse;
  wire or_516_cse;
  wire or_521_cse;
  wire or_528_cse;
  wire or_537_cse;
  wire and_790_cse;
  wire or_548_cse;
  wire or_561_cse;
  wire or_576_cse;
  wire nand_146_cse;
  wire or_617_cse;
  wire or_622_cse;
  wire or_629_cse;
  wire or_638_cse;
  wire or_649_cse;
  wire or_662_cse;
  wire or_677_cse;
  wire or_718_cse;
  wire nand_112_cse;
  wire nand_108_cse;
  wire nand_103_cse;
  wire nand_97_cse;
  wire or_763_cse;
  wire nand_83_cse;
  wire or_818_cse;
  wire or_823_cse;
  wire or_830_cse;
  wire or_839_cse;
  wire nand_58_cse;
  wire or_850_cse;
  wire nand_55_cse;
  wire or_863_cse;
  wire nand_51_cse;
  wire or_878_cse;
  wire and_749_cse;
  wire or_928_cse;
  wire and_747_cse;
  wire or_933_cse;
  wire and_744_cse;
  wire or_940_cse;
  wire and_740_cse;
  wire or_949_cse;
  wire or_960_cse;
  wire and_731_cse;
  wire or_973_cse;
  wire and_725_cse;
  wire nand_42_cse;
  wire or_988_cse;
  wire or_1037_cse;
  wire or_1042_cse;
  wire or_1049_cse;
  wire or_1058_cse;
  wire or_1069_cse;
  wire or_1082_cse;
  wire or_1097_cse;
  reg [63:0] base_buf_sva_mut_2;
  reg [63:0] base_buf_sva_mut_3;
  reg [63:0] base_buf_sva_mut_4;
  reg [63:0] base_buf_sva_mut_5;
  reg [63:0] base_buf_sva_mut_6;
  reg [63:0] base_buf_sva_mut_7;
  reg [63:0] base_buf_sva_mut_8;
  reg [63:0] base_buf_sva_mut_9;
  reg [63:0] base_buf_sva_mut_10;
  reg [63:0] m_buf_sva_mut_2;
  reg [63:0] m_buf_sva_mut_3;
  reg [63:0] m_buf_sva_mut_4;
  reg [63:0] m_buf_sva_mut_5;
  reg [63:0] m_buf_sva_mut_6;
  reg [63:0] m_buf_sva_mut_7;
  reg [63:0] m_buf_sva_mut_8;
  reg [63:0] m_buf_sva_mut_9;
  reg [63:0] m_buf_sva_mut_10;
  reg [63:0] base_buf_sva_mut_1_2;
  reg [63:0] base_buf_sva_mut_1_3;
  reg [63:0] base_buf_sva_mut_1_4;
  reg [63:0] base_buf_sva_mut_1_5;
  reg [63:0] base_buf_sva_mut_1_6;
  reg [63:0] base_buf_sva_mut_1_7;
  reg [63:0] base_buf_sva_mut_1_8;
  reg [63:0] base_buf_sva_mut_1_9;
  reg [63:0] base_buf_sva_mut_1_10;
  reg [63:0] m_buf_sva_mut_1_2;
  reg [63:0] m_buf_sva_mut_1_3;
  reg [63:0] m_buf_sva_mut_1_4;
  reg [63:0] m_buf_sva_mut_1_5;
  reg [63:0] m_buf_sva_mut_1_6;
  reg [63:0] m_buf_sva_mut_1_7;
  reg [63:0] m_buf_sva_mut_1_8;
  reg [63:0] m_buf_sva_mut_1_9;
  reg [63:0] m_buf_sva_mut_1_10;
  reg [63:0] base_buf_sva_mut_2_2;
  reg [63:0] base_buf_sva_mut_2_3;
  reg [63:0] base_buf_sva_mut_2_4;
  reg [63:0] base_buf_sva_mut_2_5;
  reg [63:0] base_buf_sva_mut_2_6;
  reg [63:0] base_buf_sva_mut_2_7;
  reg [63:0] base_buf_sva_mut_2_8;
  reg [63:0] base_buf_sva_mut_2_9;
  reg [63:0] base_buf_sva_mut_2_10;
  reg [63:0] m_buf_sva_mut_2_2;
  reg [63:0] m_buf_sva_mut_2_3;
  reg [63:0] m_buf_sva_mut_2_4;
  reg [63:0] m_buf_sva_mut_2_5;
  reg [63:0] m_buf_sva_mut_2_6;
  reg [63:0] m_buf_sva_mut_2_7;
  reg [63:0] m_buf_sva_mut_2_8;
  reg [63:0] m_buf_sva_mut_2_9;
  reg [63:0] m_buf_sva_mut_2_10;
  reg [63:0] base_buf_sva_mut_3_2;
  reg [63:0] base_buf_sva_mut_3_3;
  reg [63:0] base_buf_sva_mut_3_4;
  reg [63:0] base_buf_sva_mut_3_5;
  reg [63:0] base_buf_sva_mut_3_6;
  reg [63:0] base_buf_sva_mut_3_7;
  reg [63:0] base_buf_sva_mut_3_8;
  reg [63:0] base_buf_sva_mut_3_9;
  reg [63:0] base_buf_sva_mut_3_10;
  reg [63:0] m_buf_sva_mut_3_2;
  reg [63:0] m_buf_sva_mut_3_3;
  reg [63:0] m_buf_sva_mut_3_4;
  reg [63:0] m_buf_sva_mut_3_5;
  reg [63:0] m_buf_sva_mut_3_6;
  reg [63:0] m_buf_sva_mut_3_7;
  reg [63:0] m_buf_sva_mut_3_8;
  reg [63:0] m_buf_sva_mut_3_9;
  reg [63:0] m_buf_sva_mut_3_10;
  reg [63:0] base_buf_sva_mut_4_2;
  reg [63:0] base_buf_sva_mut_4_3;
  reg [63:0] base_buf_sva_mut_4_4;
  reg [63:0] base_buf_sva_mut_4_5;
  reg [63:0] base_buf_sva_mut_4_6;
  reg [63:0] base_buf_sva_mut_4_7;
  reg [63:0] base_buf_sva_mut_4_8;
  reg [63:0] base_buf_sva_mut_4_9;
  reg [63:0] base_buf_sva_mut_4_10;
  reg [63:0] m_buf_sva_mut_4_2;
  reg [63:0] m_buf_sva_mut_4_3;
  reg [63:0] m_buf_sva_mut_4_4;
  reg [63:0] m_buf_sva_mut_4_5;
  reg [63:0] m_buf_sva_mut_4_6;
  reg [63:0] m_buf_sva_mut_4_7;
  reg [63:0] m_buf_sva_mut_4_8;
  reg [63:0] m_buf_sva_mut_4_9;
  reg [63:0] m_buf_sva_mut_4_10;
  reg [63:0] base_buf_sva_mut_5_2;
  reg [63:0] base_buf_sva_mut_5_3;
  reg [63:0] base_buf_sva_mut_5_4;
  reg [63:0] base_buf_sva_mut_5_5;
  reg [63:0] base_buf_sva_mut_5_6;
  reg [63:0] base_buf_sva_mut_5_7;
  reg [63:0] base_buf_sva_mut_5_8;
  reg [63:0] base_buf_sva_mut_5_9;
  reg [63:0] base_buf_sva_mut_5_10;
  reg [63:0] m_buf_sva_mut_5_2;
  reg [63:0] m_buf_sva_mut_5_3;
  reg [63:0] m_buf_sva_mut_5_4;
  reg [63:0] m_buf_sva_mut_5_5;
  reg [63:0] m_buf_sva_mut_5_6;
  reg [63:0] m_buf_sva_mut_5_7;
  reg [63:0] m_buf_sva_mut_5_8;
  reg [63:0] m_buf_sva_mut_5_9;
  reg [63:0] m_buf_sva_mut_5_10;
  reg [63:0] base_buf_sva_mut_6_2;
  reg [63:0] base_buf_sva_mut_6_3;
  reg [63:0] base_buf_sva_mut_6_4;
  reg [63:0] base_buf_sva_mut_6_5;
  reg [63:0] base_buf_sva_mut_6_6;
  reg [63:0] base_buf_sva_mut_6_7;
  reg [63:0] base_buf_sva_mut_6_8;
  reg [63:0] base_buf_sva_mut_6_9;
  reg [63:0] base_buf_sva_mut_6_10;
  reg [63:0] m_buf_sva_mut_6_2;
  reg [63:0] m_buf_sva_mut_6_3;
  reg [63:0] m_buf_sva_mut_6_4;
  reg [63:0] m_buf_sva_mut_6_5;
  reg [63:0] m_buf_sva_mut_6_6;
  reg [63:0] m_buf_sva_mut_6_7;
  reg [63:0] m_buf_sva_mut_6_8;
  reg [63:0] m_buf_sva_mut_6_9;
  reg [63:0] m_buf_sva_mut_6_10;
  reg [63:0] base_buf_sva_mut_7_2;
  reg [63:0] base_buf_sva_mut_7_3;
  reg [63:0] base_buf_sva_mut_7_4;
  reg [63:0] base_buf_sva_mut_7_5;
  reg [63:0] base_buf_sva_mut_7_6;
  reg [63:0] base_buf_sva_mut_7_7;
  reg [63:0] base_buf_sva_mut_7_8;
  reg [63:0] base_buf_sva_mut_7_9;
  reg [63:0] base_buf_sva_mut_7_10;
  reg [63:0] m_buf_sva_mut_7_2;
  reg [63:0] m_buf_sva_mut_7_3;
  reg [63:0] m_buf_sva_mut_7_4;
  reg [63:0] m_buf_sva_mut_7_5;
  reg [63:0] m_buf_sva_mut_7_6;
  reg [63:0] m_buf_sva_mut_7_7;
  reg [63:0] m_buf_sva_mut_7_8;
  reg [63:0] m_buf_sva_mut_7_9;
  reg [63:0] m_buf_sva_mut_7_10;
  reg [63:0] base_buf_sva_mut_8_2;
  reg [63:0] base_buf_sva_mut_8_3;
  reg [63:0] base_buf_sva_mut_8_4;
  reg [63:0] base_buf_sva_mut_8_5;
  reg [63:0] base_buf_sva_mut_8_6;
  reg [63:0] base_buf_sva_mut_8_7;
  reg [63:0] base_buf_sva_mut_8_8;
  reg [63:0] base_buf_sva_mut_8_9;
  reg [63:0] base_buf_sva_mut_8_10;
  reg [63:0] m_buf_sva_mut_8_2;
  reg [63:0] m_buf_sva_mut_8_3;
  reg [63:0] m_buf_sva_mut_8_4;
  reg [63:0] m_buf_sva_mut_8_5;
  reg [63:0] m_buf_sva_mut_8_6;
  reg [63:0] m_buf_sva_mut_8_7;
  reg [63:0] m_buf_sva_mut_8_8;
  reg [63:0] m_buf_sva_mut_8_9;
  reg [63:0] m_buf_sva_mut_8_10;
  reg [63:0] base_buf_sva_mut_9_2;
  reg [63:0] base_buf_sva_mut_9_3;
  reg [63:0] base_buf_sva_mut_9_4;
  reg [63:0] base_buf_sva_mut_9_5;
  reg [63:0] base_buf_sva_mut_9_6;
  reg [63:0] base_buf_sva_mut_9_7;
  reg [63:0] base_buf_sva_mut_9_8;
  reg [63:0] base_buf_sva_mut_9_9;
  reg [63:0] base_buf_sva_mut_9_10;
  reg [63:0] m_buf_sva_mut_9_2;
  reg [63:0] m_buf_sva_mut_9_3;
  reg [63:0] m_buf_sva_mut_9_4;
  reg [63:0] m_buf_sva_mut_9_5;
  reg [63:0] m_buf_sva_mut_9_6;
  reg [63:0] m_buf_sva_mut_9_7;
  reg [63:0] m_buf_sva_mut_9_8;
  reg [63:0] m_buf_sva_mut_9_9;
  reg [63:0] m_buf_sva_mut_9_10;
  reg [63:0] base_buf_sva_mut_10_2;
  reg [63:0] base_buf_sva_mut_10_3;
  reg [63:0] base_buf_sva_mut_10_4;
  reg [63:0] base_buf_sva_mut_10_5;
  reg [63:0] base_buf_sva_mut_10_6;
  reg [63:0] base_buf_sva_mut_10_7;
  reg [63:0] base_buf_sva_mut_10_8;
  reg [63:0] base_buf_sva_mut_10_9;
  reg [63:0] base_buf_sva_mut_10_10;
  reg [63:0] m_buf_sva_mut_10_2;
  reg [63:0] m_buf_sva_mut_10_3;
  reg [63:0] m_buf_sva_mut_10_4;
  reg [63:0] m_buf_sva_mut_10_5;
  reg [63:0] m_buf_sva_mut_10_6;
  reg [63:0] m_buf_sva_mut_10_7;
  reg [63:0] m_buf_sva_mut_10_8;
  reg [63:0] m_buf_sva_mut_10_9;
  reg [63:0] m_buf_sva_mut_10_10;
  reg [3:0] result_rem_11cyc_st_10;
  wire return_rsci_d_mx0c0;
  wire return_rsci_d_mx0c1;
  wire return_rsci_d_mx0c2;
  wire return_rsci_d_mx0c3;
  wire return_rsci_d_mx0c4;
  wire return_rsci_d_mx0c5;
  wire return_rsci_d_mx0c6;
  wire return_rsci_d_mx0c7;
  wire return_rsci_d_mx0c8;
  wire return_rsci_d_mx0c9;
  wire return_rsci_d_mx0c10;
  wire [3:0] result_acc_imod_1;
  wire [5:0] nl_result_acc_imod_1;
  wire [3:0] result_acc_idiv_1;
  wire [4:0] nl_result_acc_idiv_1;
  wire m_and_cse;
  wire m_and_1_cse;
  wire m_and_2_cse;
  wire m_and_3_cse;
  wire m_and_4_cse;
  wire m_and_5_cse;
  wire m_and_6_cse;
  wire m_and_7_cse;
  wire m_and_8_cse;
  wire m_and_9_cse;
  wire m_and_10_cse;
  wire m_and_11_cse;
  wire m_and_12_cse;
  wire m_and_13_cse;
  wire m_and_14_cse;
  wire m_and_15_cse;
  wire m_and_16_cse;
  wire m_and_17_cse;
  wire m_and_18_cse;
  wire m_and_19_cse;
  wire m_and_20_cse;
  wire m_and_21_cse;
  wire m_and_22_cse;
  wire m_and_23_cse;
  wire m_and_24_cse;
  wire m_and_25_cse;
  wire m_and_26_cse;
  wire m_and_27_cse;
  wire m_and_28_cse;
  wire m_and_29_cse;
  wire m_and_30_cse;
  wire m_and_31_cse;
  wire m_and_32_cse;
  wire m_and_33_cse;
  wire m_and_34_cse;
  wire m_and_35_cse;
  wire m_and_36_cse;
  wire m_and_37_cse;
  wire m_and_38_cse;
  wire m_and_39_cse;
  wire m_and_40_cse;
  wire m_and_41_cse;
  wire m_and_42_cse;
  wire m_and_43_cse;
  wire m_and_44_cse;
  wire m_and_45_cse;
  wire m_and_46_cse;
  wire m_and_47_cse;
  wire m_and_48_cse;
  wire m_and_49_cse;
  wire m_and_50_cse;
  wire m_and_51_cse;
  wire m_and_52_cse;
  wire m_and_53_cse;
  wire m_and_54_cse;
  wire m_and_55_cse;
  wire m_and_56_cse;
  wire m_and_57_cse;
  wire m_and_58_cse;
  wire m_and_59_cse;
  wire m_and_60_cse;
  wire m_and_61_cse;
  wire m_and_62_cse;
  wire m_and_63_cse;
  wire m_and_64_cse;
  wire m_and_65_cse;
  wire m_and_66_cse;
  wire m_and_67_cse;
  wire m_and_68_cse;
  wire m_and_69_cse;
  wire m_and_70_cse;
  wire m_and_71_cse;
  wire m_and_72_cse;
  wire m_and_73_cse;
  wire m_and_74_cse;
  wire m_and_75_cse;
  wire m_and_76_cse;
  wire m_and_77_cse;
  wire m_and_78_cse;
  wire m_and_79_cse;
  wire m_and_80_cse;
  wire m_and_81_cse;
  wire m_and_82_cse;
  wire m_and_83_cse;
  wire m_and_84_cse;
  wire m_and_85_cse;
  wire m_and_86_cse;
  wire m_and_87_cse;
  wire m_and_88_cse;
  wire m_and_89_cse;
  wire m_and_90_cse;
  wire m_and_91_cse;
  wire m_and_92_cse;
  wire m_and_93_cse;
  wire m_and_94_cse;
  wire m_and_95_cse;
  wire m_and_96_cse;
  wire m_and_97_cse;
  wire m_and_98_cse;

  wire[0:0] mux_nl;
  wire[0:0] nor_691_nl;
  wire[0:0] nor_690_nl;
  wire[0:0] or_10_nl;
  wire[0:0] mux_2_nl;
  wire[0:0] nor_689_nl;
  wire[0:0] nor_687_nl;
  wire[0:0] or_17_nl;
  wire[0:0] nor_688_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] nor_686_nl;
  wire[0:0] nor_683_nl;
  wire[0:0] or_26_nl;
  wire[0:0] nor_684_nl;
  wire[0:0] nor_685_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] nor_682_nl;
  wire[0:0] nor_678_nl;
  wire[0:0] or_37_nl;
  wire[0:0] nor_679_nl;
  wire[0:0] nor_680_nl;
  wire[0:0] nor_681_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] nor_677_nl;
  wire[0:0] nor_672_nl;
  wire[0:0] or_50_nl;
  wire[0:0] nor_673_nl;
  wire[0:0] nor_674_nl;
  wire[0:0] nor_675_nl;
  wire[0:0] nor_676_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] nor_671_nl;
  wire[0:0] nor_665_nl;
  wire[0:0] or_65_nl;
  wire[0:0] nor_666_nl;
  wire[0:0] nor_667_nl;
  wire[0:0] nor_668_nl;
  wire[0:0] nor_669_nl;
  wire[0:0] nor_670_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] nor_664_nl;
  wire[0:0] nor_656_nl;
  wire[0:0] or_82_nl;
  wire[0:0] or_80_nl;
  wire[0:0] nor_657_nl;
  wire[0:0] nor_658_nl;
  wire[0:0] nor_659_nl;
  wire[0:0] nor_660_nl;
  wire[0:0] nor_661_nl;
  wire[0:0] nor_662_nl;
  wire[0:0] mux_35_nl;
  wire[0:0] nor_663_nl;
  wire[0:0] nor_654_nl;
  wire[0:0] nor_655_nl;
  wire[0:0] mux_38_nl;
  wire[0:0] nor_653_nl;
  wire[0:0] nor_652_nl;
  wire[0:0] or_114_nl;
  wire[0:0] mux_40_nl;
  wire[0:0] nor_651_nl;
  wire[0:0] nor_649_nl;
  wire[0:0] or_121_nl;
  wire[0:0] nor_650_nl;
  wire[0:0] mux_43_nl;
  wire[0:0] nor_648_nl;
  wire[0:0] nor_645_nl;
  wire[0:0] or_130_nl;
  wire[0:0] nor_646_nl;
  wire[0:0] nor_647_nl;
  wire[0:0] mux_47_nl;
  wire[0:0] nor_644_nl;
  wire[0:0] nor_640_nl;
  wire[0:0] or_141_nl;
  wire[0:0] nor_641_nl;
  wire[0:0] nor_642_nl;
  wire[0:0] nor_643_nl;
  wire[0:0] mux_52_nl;
  wire[0:0] nor_639_nl;
  wire[0:0] nor_634_nl;
  wire[0:0] or_154_nl;
  wire[0:0] nor_635_nl;
  wire[0:0] nor_636_nl;
  wire[0:0] nor_637_nl;
  wire[0:0] nor_638_nl;
  wire[0:0] mux_58_nl;
  wire[0:0] nor_633_nl;
  wire[0:0] nor_627_nl;
  wire[0:0] or_169_nl;
  wire[0:0] nor_628_nl;
  wire[0:0] nor_629_nl;
  wire[0:0] nor_630_nl;
  wire[0:0] nor_631_nl;
  wire[0:0] nor_632_nl;
  wire[0:0] mux_65_nl;
  wire[0:0] nor_626_nl;
  wire[0:0] nor_618_nl;
  wire[0:0] or_186_nl;
  wire[0:0] or_184_nl;
  wire[0:0] nor_619_nl;
  wire[0:0] nor_620_nl;
  wire[0:0] nor_621_nl;
  wire[0:0] nor_622_nl;
  wire[0:0] nor_623_nl;
  wire[0:0] nor_624_nl;
  wire[0:0] mux_73_nl;
  wire[0:0] nor_625_nl;
  wire[0:0] nor_617_nl;
  wire[0:0] and_797_nl;
  wire[0:0] or_195_nl;
  wire[0:0] mux_76_nl;
  wire[0:0] nor_616_nl;
  wire[0:0] nor_615_nl;
  wire[0:0] or_216_nl;
  wire[0:0] mux_78_nl;
  wire[0:0] nor_614_nl;
  wire[0:0] nor_612_nl;
  wire[0:0] or_223_nl;
  wire[0:0] nor_613_nl;
  wire[0:0] mux_81_nl;
  wire[0:0] nor_611_nl;
  wire[0:0] nor_608_nl;
  wire[0:0] or_232_nl;
  wire[0:0] nor_609_nl;
  wire[0:0] nor_610_nl;
  wire[0:0] mux_85_nl;
  wire[0:0] nor_607_nl;
  wire[0:0] nor_603_nl;
  wire[0:0] or_243_nl;
  wire[0:0] nor_604_nl;
  wire[0:0] nor_605_nl;
  wire[0:0] nor_606_nl;
  wire[0:0] mux_90_nl;
  wire[0:0] nor_602_nl;
  wire[0:0] nor_597_nl;
  wire[0:0] or_256_nl;
  wire[0:0] nor_598_nl;
  wire[0:0] nor_599_nl;
  wire[0:0] nor_600_nl;
  wire[0:0] nor_601_nl;
  wire[0:0] mux_96_nl;
  wire[0:0] nor_596_nl;
  wire[0:0] nor_590_nl;
  wire[0:0] or_271_nl;
  wire[0:0] nor_591_nl;
  wire[0:0] nor_592_nl;
  wire[0:0] nor_593_nl;
  wire[0:0] nor_594_nl;
  wire[0:0] nor_595_nl;
  wire[0:0] mux_103_nl;
  wire[0:0] nor_589_nl;
  wire[0:0] nor_581_nl;
  wire[0:0] or_288_nl;
  wire[0:0] or_286_nl;
  wire[0:0] nor_582_nl;
  wire[0:0] nor_583_nl;
  wire[0:0] nor_584_nl;
  wire[0:0] nor_585_nl;
  wire[0:0] nor_586_nl;
  wire[0:0] nor_587_nl;
  wire[0:0] mux_111_nl;
  wire[0:0] nor_588_nl;
  wire[0:0] nor_579_nl;
  wire[0:0] nor_580_nl;
  wire[0:0] mux_114_nl;
  wire[0:0] nor_578_nl;
  wire[0:0] nor_577_nl;
  wire[0:0] or_318_nl;
  wire[0:0] mux_116_nl;
  wire[0:0] nor_576_nl;
  wire[0:0] nor_574_nl;
  wire[0:0] or_325_nl;
  wire[0:0] nor_575_nl;
  wire[0:0] mux_119_nl;
  wire[0:0] nor_573_nl;
  wire[0:0] nor_570_nl;
  wire[0:0] or_334_nl;
  wire[0:0] nor_571_nl;
  wire[0:0] nor_572_nl;
  wire[0:0] mux_123_nl;
  wire[0:0] nor_569_nl;
  wire[0:0] nor_565_nl;
  wire[0:0] or_345_nl;
  wire[0:0] nor_566_nl;
  wire[0:0] nor_567_nl;
  wire[0:0] nor_568_nl;
  wire[0:0] mux_128_nl;
  wire[0:0] nor_564_nl;
  wire[0:0] nor_559_nl;
  wire[0:0] or_358_nl;
  wire[0:0] nor_560_nl;
  wire[0:0] nor_561_nl;
  wire[0:0] nor_562_nl;
  wire[0:0] nor_563_nl;
  wire[0:0] mux_134_nl;
  wire[0:0] nor_558_nl;
  wire[0:0] nor_552_nl;
  wire[0:0] or_373_nl;
  wire[0:0] nor_553_nl;
  wire[0:0] nor_554_nl;
  wire[0:0] nor_555_nl;
  wire[0:0] nor_556_nl;
  wire[0:0] nor_557_nl;
  wire[0:0] mux_141_nl;
  wire[0:0] nor_551_nl;
  wire[0:0] nor_543_nl;
  wire[0:0] or_390_nl;
  wire[0:0] or_388_nl;
  wire[0:0] nor_544_nl;
  wire[0:0] nor_545_nl;
  wire[0:0] nor_546_nl;
  wire[0:0] nor_547_nl;
  wire[0:0] nor_548_nl;
  wire[0:0] nor_549_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] nor_550_nl;
  wire[0:0] nor_542_nl;
  wire[0:0] and_796_nl;
  wire[0:0] or_399_nl;
  wire[0:0] mux_152_nl;
  wire[0:0] and_795_nl;
  wire[0:0] nor_541_nl;
  wire[0:0] or_420_nl;
  wire[0:0] mux_154_nl;
  wire[0:0] and_794_nl;
  wire[0:0] nor_539_nl;
  wire[0:0] or_427_nl;
  wire[0:0] nor_540_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] and_793_nl;
  wire[0:0] nor_536_nl;
  wire[0:0] or_436_nl;
  wire[0:0] nor_537_nl;
  wire[0:0] nor_538_nl;
  wire[0:0] mux_161_nl;
  wire[0:0] and_792_nl;
  wire[0:0] nor_532_nl;
  wire[0:0] or_447_nl;
  wire[0:0] nor_533_nl;
  wire[0:0] nor_534_nl;
  wire[0:0] nor_535_nl;
  wire[0:0] mux_166_nl;
  wire[0:0] and_791_nl;
  wire[0:0] nor_527_nl;
  wire[0:0] or_460_nl;
  wire[0:0] nor_528_nl;
  wire[0:0] nor_529_nl;
  wire[0:0] nor_530_nl;
  wire[0:0] nor_531_nl;
  wire[0:0] mux_172_nl;
  wire[0:0] and_789_nl;
  wire[0:0] nor_522_nl;
  wire[0:0] or_475_nl;
  wire[0:0] and_788_nl;
  wire[0:0] nor_523_nl;
  wire[0:0] nor_524_nl;
  wire[0:0] nor_525_nl;
  wire[0:0] nor_526_nl;
  wire[0:0] mux_179_nl;
  wire[0:0] and_787_nl;
  wire[0:0] nor_516_nl;
  wire[0:0] or_492_nl;
  wire[0:0] or_490_nl;
  wire[0:0] nor_517_nl;
  wire[0:0] and_785_nl;
  wire[0:0] nor_518_nl;
  wire[0:0] nor_519_nl;
  wire[0:0] nor_520_nl;
  wire[0:0] nor_521_nl;
  wire[0:0] mux_187_nl;
  wire[0:0] and_786_nl;
  wire[0:0] nor_514_nl;
  wire[0:0] nor_515_nl;
  wire[0:0] or_501_nl;
  wire[0:0] mux_190_nl;
  wire[0:0] and_784_nl;
  wire[0:0] nor_513_nl;
  wire[0:0] or_523_nl;
  wire[0:0] mux_192_nl;
  wire[0:0] and_783_nl;
  wire[0:0] nor_511_nl;
  wire[0:0] or_530_nl;
  wire[0:0] nor_512_nl;
  wire[0:0] mux_195_nl;
  wire[0:0] and_782_nl;
  wire[0:0] nor_508_nl;
  wire[0:0] or_539_nl;
  wire[0:0] nor_509_nl;
  wire[0:0] nor_510_nl;
  wire[0:0] mux_199_nl;
  wire[0:0] and_781_nl;
  wire[0:0] nor_504_nl;
  wire[0:0] or_550_nl;
  wire[0:0] nor_505_nl;
  wire[0:0] nor_506_nl;
  wire[0:0] nor_507_nl;
  wire[0:0] mux_204_nl;
  wire[0:0] and_780_nl;
  wire[0:0] nor_499_nl;
  wire[0:0] or_563_nl;
  wire[0:0] nor_500_nl;
  wire[0:0] nor_501_nl;
  wire[0:0] nor_502_nl;
  wire[0:0] nor_503_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] and_778_nl;
  wire[0:0] nor_494_nl;
  wire[0:0] or_578_nl;
  wire[0:0] and_777_nl;
  wire[0:0] nor_495_nl;
  wire[0:0] nor_496_nl;
  wire[0:0] nor_497_nl;
  wire[0:0] nor_498_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] and_776_nl;
  wire[0:0] nor_488_nl;
  wire[0:0] or_595_nl;
  wire[0:0] or_593_nl;
  wire[0:0] nor_489_nl;
  wire[0:0] and_774_nl;
  wire[0:0] nor_490_nl;
  wire[0:0] nor_491_nl;
  wire[0:0] nor_492_nl;
  wire[0:0] nor_493_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] and_775_nl;
  wire[0:0] nor_487_nl;
  wire[0:0] and_773_nl;
  wire[0:0] or_604_nl;
  wire[0:0] mux_228_nl;
  wire[0:0] and_772_nl;
  wire[0:0] nor_486_nl;
  wire[0:0] or_624_nl;
  wire[0:0] mux_230_nl;
  wire[0:0] and_771_nl;
  wire[0:0] nor_484_nl;
  wire[0:0] or_631_nl;
  wire[0:0] nor_485_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] and_770_nl;
  wire[0:0] nor_481_nl;
  wire[0:0] or_640_nl;
  wire[0:0] nor_482_nl;
  wire[0:0] nor_483_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] and_769_nl;
  wire[0:0] nor_477_nl;
  wire[0:0] or_651_nl;
  wire[0:0] nor_478_nl;
  wire[0:0] nor_479_nl;
  wire[0:0] nor_480_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] and_768_nl;
  wire[0:0] nor_472_nl;
  wire[0:0] or_664_nl;
  wire[0:0] nor_473_nl;
  wire[0:0] nor_474_nl;
  wire[0:0] nor_475_nl;
  wire[0:0] nor_476_nl;
  wire[0:0] mux_248_nl;
  wire[0:0] and_766_nl;
  wire[0:0] nor_467_nl;
  wire[0:0] or_679_nl;
  wire[0:0] and_765_nl;
  wire[0:0] nor_468_nl;
  wire[0:0] nor_469_nl;
  wire[0:0] nor_470_nl;
  wire[0:0] nor_471_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] and_764_nl;
  wire[0:0] nor_461_nl;
  wire[0:0] or_696_nl;
  wire[0:0] or_694_nl;
  wire[0:0] nor_462_nl;
  wire[0:0] and_762_nl;
  wire[0:0] nor_463_nl;
  wire[0:0] nor_464_nl;
  wire[0:0] nor_465_nl;
  wire[0:0] nor_466_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] and_763_nl;
  wire[0:0] nor_459_nl;
  wire[0:0] nor_460_nl;
  wire[0:0] or_705_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] and_761_nl;
  wire[0:0] nor_458_nl;
  wire[0:0] nand_153_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] and_760_nl;
  wire[0:0] nor_456_nl;
  wire[0:0] nand_152_nl;
  wire[0:0] nor_457_nl;
  wire[0:0] mux_271_nl;
  wire[0:0] and_759_nl;
  wire[0:0] nor_453_nl;
  wire[0:0] nand_151_nl;
  wire[0:0] nor_454_nl;
  wire[0:0] nor_455_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] and_758_nl;
  wire[0:0] nor_449_nl;
  wire[0:0] nand_96_nl;
  wire[0:0] nor_450_nl;
  wire[0:0] nor_451_nl;
  wire[0:0] nor_452_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] and_757_nl;
  wire[0:0] nor_444_nl;
  wire[0:0] nand_150_nl;
  wire[0:0] nor_445_nl;
  wire[0:0] nor_446_nl;
  wire[0:0] nor_447_nl;
  wire[0:0] nor_448_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] and_755_nl;
  wire[0:0] nor_439_nl;
  wire[0:0] nand_149_nl;
  wire[0:0] and_754_nl;
  wire[0:0] nor_440_nl;
  wire[0:0] nor_441_nl;
  wire[0:0] nor_442_nl;
  wire[0:0] nor_443_nl;
  wire[0:0] mux_293_nl;
  wire[0:0] and_753_nl;
  wire[0:0] nor_433_nl;
  wire[0:0] nand_72_nl;
  wire[0:0] nand_73_nl;
  wire[0:0] nor_434_nl;
  wire[0:0] and_751_nl;
  wire[0:0] nor_435_nl;
  wire[0:0] nor_436_nl;
  wire[0:0] nor_437_nl;
  wire[0:0] nor_438_nl;
  wire[0:0] mux_301_nl;
  wire[0:0] and_752_nl;
  wire[0:0] nor_432_nl;
  wire[0:0] and_750_nl;
  wire[0:0] mux_304_nl;
  wire[0:0] nor_431_nl;
  wire[0:0] nor_430_nl;
  wire[0:0] or_825_nl;
  wire[0:0] mux_306_nl;
  wire[0:0] nor_429_nl;
  wire[0:0] nor_428_nl;
  wire[0:0] or_832_nl;
  wire[0:0] and_748_nl;
  wire[0:0] mux_309_nl;
  wire[0:0] nor_427_nl;
  wire[0:0] nor_426_nl;
  wire[0:0] or_841_nl;
  wire[0:0] and_745_nl;
  wire[0:0] and_746_nl;
  wire[0:0] mux_313_nl;
  wire[0:0] nor_425_nl;
  wire[0:0] nor_424_nl;
  wire[0:0] or_852_nl;
  wire[0:0] and_741_nl;
  wire[0:0] and_742_nl;
  wire[0:0] and_743_nl;
  wire[0:0] mux_318_nl;
  wire[0:0] nor_423_nl;
  wire[0:0] nor_422_nl;
  wire[0:0] or_865_nl;
  wire[0:0] and_736_nl;
  wire[0:0] and_737_nl;
  wire[0:0] and_738_nl;
  wire[0:0] and_739_nl;
  wire[0:0] mux_324_nl;
  wire[0:0] nor_421_nl;
  wire[0:0] nor_419_nl;
  wire[0:0] or_880_nl;
  wire[0:0] nor_420_nl;
  wire[0:0] and_732_nl;
  wire[0:0] and_733_nl;
  wire[0:0] and_734_nl;
  wire[0:0] and_735_nl;
  wire[0:0] mux_331_nl;
  wire[0:0] nor_418_nl;
  wire[0:0] nor_415_nl;
  wire[0:0] or_897_nl;
  wire[0:0] or_895_nl;
  wire[0:0] and_726_nl;
  wire[0:0] nor_416_nl;
  wire[0:0] and_727_nl;
  wire[0:0] and_728_nl;
  wire[0:0] and_729_nl;
  wire[0:0] and_730_nl;
  wire[0:0] mux_339_nl;
  wire[0:0] nor_417_nl;
  wire[0:0] nor_407_nl;
  wire[0:0] or_914_nl;
  wire[0:0] nor_408_nl;
  wire[0:0] or_913_nl;
  wire[0:0] nor_409_nl;
  wire[0:0] or_912_nl;
  wire[0:0] nor_410_nl;
  wire[0:0] or_911_nl;
  wire[0:0] nor_411_nl;
  wire[0:0] or_910_nl;
  wire[0:0] nor_412_nl;
  wire[0:0] or_909_nl;
  wire[0:0] nor_413_nl;
  wire[0:0] or_908_nl;
  wire[0:0] and_724_nl;
  wire[0:0] nor_414_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] nor_406_nl;
  wire[0:0] nor_405_nl;
  wire[0:0] or_935_nl;
  wire[0:0] mux_351_nl;
  wire[0:0] nor_404_nl;
  wire[0:0] nor_403_nl;
  wire[0:0] or_942_nl;
  wire[0:0] and_722_nl;
  wire[0:0] mux_354_nl;
  wire[0:0] nor_402_nl;
  wire[0:0] nor_401_nl;
  wire[0:0] or_951_nl;
  wire[0:0] and_719_nl;
  wire[0:0] and_720_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] nor_400_nl;
  wire[0:0] nor_399_nl;
  wire[0:0] or_962_nl;
  wire[0:0] and_715_nl;
  wire[0:0] and_716_nl;
  wire[0:0] and_717_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] nor_398_nl;
  wire[0:0] nor_397_nl;
  wire[0:0] or_975_nl;
  wire[0:0] and_710_nl;
  wire[0:0] and_711_nl;
  wire[0:0] and_712_nl;
  wire[0:0] and_713_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] nor_396_nl;
  wire[0:0] nor_394_nl;
  wire[0:0] or_990_nl;
  wire[0:0] nor_395_nl;
  wire[0:0] and_706_nl;
  wire[0:0] and_707_nl;
  wire[0:0] and_708_nl;
  wire[0:0] and_709_nl;
  wire[0:0] mux_376_nl;
  wire[0:0] nor_393_nl;
  wire[0:0] nor_390_nl;
  wire[0:0] or_1007_nl;
  wire[0:0] or_1005_nl;
  wire[0:0] and_700_nl;
  wire[0:0] nor_391_nl;
  wire[0:0] and_701_nl;
  wire[0:0] and_702_nl;
  wire[0:0] and_703_nl;
  wire[0:0] and_704_nl;
  wire[0:0] mux_384_nl;
  wire[0:0] nor_392_nl;
  wire[0:0] nor_383_nl;
  wire[0:0] or_1024_nl;
  wire[0:0] nor_384_nl;
  wire[0:0] or_1023_nl;
  wire[0:0] nor_385_nl;
  wire[0:0] or_1022_nl;
  wire[0:0] nor_386_nl;
  wire[0:0] or_1021_nl;
  wire[0:0] nor_387_nl;
  wire[0:0] or_1020_nl;
  wire[0:0] nor_388_nl;
  wire[0:0] or_1019_nl;
  wire[0:0] nor_389_nl;
  wire[0:0] or_1018_nl;
  wire[0:0] and_697_nl;
  wire[0:0] and_698_nl;
  wire[0:0] or_1016_nl;
  wire[0:0] mux_394_nl;
  wire[0:0] nor_382_nl;
  wire[0:0] nor_381_nl;
  wire[0:0] or_1044_nl;
  wire[0:0] mux_396_nl;
  wire[0:0] nor_380_nl;
  wire[0:0] nor_379_nl;
  wire[0:0] or_1051_nl;
  wire[0:0] and_695_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] nor_378_nl;
  wire[0:0] nor_377_nl;
  wire[0:0] or_1060_nl;
  wire[0:0] and_692_nl;
  wire[0:0] and_693_nl;
  wire[0:0] mux_403_nl;
  wire[0:0] nor_376_nl;
  wire[0:0] nor_375_nl;
  wire[0:0] or_1071_nl;
  wire[0:0] and_688_nl;
  wire[0:0] and_689_nl;
  wire[0:0] and_690_nl;
  wire[0:0] mux_408_nl;
  wire[0:0] nor_374_nl;
  wire[0:0] nor_373_nl;
  wire[0:0] or_1084_nl;
  wire[0:0] and_683_nl;
  wire[0:0] and_684_nl;
  wire[0:0] and_685_nl;
  wire[0:0] and_686_nl;
  wire[0:0] mux_414_nl;
  wire[0:0] nor_372_nl;
  wire[0:0] nor_370_nl;
  wire[0:0] or_1099_nl;
  wire[0:0] nor_371_nl;
  wire[0:0] and_679_nl;
  wire[0:0] and_680_nl;
  wire[0:0] and_681_nl;
  wire[0:0] and_682_nl;
  wire[0:0] mux_421_nl;
  wire[0:0] nor_369_nl;
  wire[0:0] nor_366_nl;
  wire[0:0] or_1116_nl;
  wire[0:0] or_1114_nl;
  wire[0:0] and_673_nl;
  wire[0:0] nor_367_nl;
  wire[0:0] and_674_nl;
  wire[0:0] and_675_nl;
  wire[0:0] and_676_nl;
  wire[0:0] and_677_nl;
  wire[0:0] mux_429_nl;
  wire[0:0] nor_368_nl;
  wire[0:0] nor_358_nl;
  wire[0:0] or_1133_nl;
  wire[0:0] nor_359_nl;
  wire[0:0] or_1132_nl;
  wire[0:0] nor_360_nl;
  wire[0:0] or_1131_nl;
  wire[0:0] nor_361_nl;
  wire[0:0] or_1130_nl;
  wire[0:0] nor_362_nl;
  wire[0:0] or_1129_nl;
  wire[0:0] nor_363_nl;
  wire[0:0] or_1128_nl;
  wire[0:0] nor_364_nl;
  wire[0:0] or_1127_nl;
  wire[0:0] and_671_nl;
  wire[0:0] nor_365_nl;

  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd64)) base_rsci (
      .dat(base_rsc_dat),
      .idat(base_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd3),
  .width(32'sd64)) return_rsci (
      .d(return_rsci_d),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd8),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp (
      .a(result_rem_12_cmp_a),
      .b(result_rem_12_cmp_b),
      .z(result_rem_12_cmp_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_1 (
      .a(result_rem_12_cmp_1_a),
      .b(result_rem_12_cmp_1_b),
      .z(result_rem_12_cmp_1_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_2 (
      .a(result_rem_12_cmp_2_a),
      .b(result_rem_12_cmp_2_b),
      .z(result_rem_12_cmp_2_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_3 (
      .a(result_rem_12_cmp_3_a),
      .b(result_rem_12_cmp_3_b),
      .z(result_rem_12_cmp_3_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_4 (
      .a(result_rem_12_cmp_4_a),
      .b(result_rem_12_cmp_4_b),
      .z(result_rem_12_cmp_4_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_5 (
      .a(result_rem_12_cmp_5_a),
      .b(result_rem_12_cmp_5_b),
      .z(result_rem_12_cmp_5_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_6 (
      .a(result_rem_12_cmp_6_a),
      .b(result_rem_12_cmp_6_b),
      .z(result_rem_12_cmp_6_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_7 (
      .a(result_rem_12_cmp_7_a),
      .b(result_rem_12_cmp_7_b),
      .z(result_rem_12_cmp_7_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_8 (
      .a(result_rem_12_cmp_8_a),
      .b(result_rem_12_cmp_8_b),
      .z(result_rem_12_cmp_8_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_9 (
      .a(result_rem_12_cmp_9_a),
      .b(result_rem_12_cmp_9_b),
      .z(result_rem_12_cmp_9_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_10 (
      .a(result_rem_12_cmp_10_a),
      .b(result_rem_12_cmp_10_b),
      .z(result_rem_12_cmp_10_z)
    );
  assign result_and_1_cse = ccs_ccore_en & (and_dcpl_263 | and_dcpl_269 | and_dcpl_275
      | and_dcpl_281 | and_dcpl_287 | and_dcpl_293 | and_dcpl_299 | and_dcpl_305
      | and_dcpl_311 | mux_tmp_37);
  assign result_and_3_cse = ccs_ccore_en & (and_dcpl_319 | and_dcpl_322 | and_dcpl_325
      | and_dcpl_329 | and_dcpl_333 | and_dcpl_337 | and_dcpl_341 | and_dcpl_344
      | and_dcpl_347 | mux_tmp_75);
  assign result_and_5_cse = ccs_ccore_en & (and_dcpl_353 | and_dcpl_357 | and_dcpl_361
      | and_dcpl_364 | and_dcpl_367 | and_dcpl_370 | and_dcpl_373 | and_dcpl_377
      | and_dcpl_381 | mux_tmp_113);
  assign result_and_7_cse = ccs_ccore_en & (and_dcpl_387 | and_dcpl_390 | and_dcpl_393
      | and_dcpl_396 | and_dcpl_399 | and_dcpl_402 | and_dcpl_405 | and_dcpl_408
      | and_dcpl_411 | mux_tmp_151);
  assign result_and_9_cse = ccs_ccore_en & (and_dcpl_418 | and_dcpl_422 | and_dcpl_426
      | and_dcpl_430 | and_dcpl_433 | and_dcpl_437 | and_dcpl_441 | and_dcpl_444
      | and_dcpl_447 | mux_tmp_189);
  assign result_and_11_cse = ccs_ccore_en & (and_dcpl_452 | and_dcpl_455 | and_dcpl_458
      | and_dcpl_462 | and_dcpl_464 | and_dcpl_468 | and_dcpl_472 | and_dcpl_474
      | and_dcpl_476 | mux_tmp_227);
  assign result_and_13_cse = ccs_ccore_en & (and_dcpl_480 | and_dcpl_484 | and_dcpl_488
      | and_dcpl_491 | and_dcpl_493 | and_dcpl_496 | and_dcpl_499 | and_dcpl_501
      | and_dcpl_503 | mux_tmp_265);
  assign result_and_15_cse = ccs_ccore_en & (and_dcpl_507 | and_dcpl_510 | and_dcpl_513
      | and_dcpl_516 | and_dcpl_518 | and_dcpl_521 | and_dcpl_524 | and_dcpl_526
      | and_dcpl_528 | mux_tmp_303);
  assign result_and_17_cse = ccs_ccore_en & (and_dcpl_533 | and_dcpl_536 | and_dcpl_539
      | and_dcpl_542 | and_dcpl_546 | and_dcpl_549 | and_dcpl_552 | and_dcpl_556
      | and_dcpl_560 | mux_tmp_348);
  assign result_and_19_cse = ccs_ccore_en & (and_dcpl_566 | and_dcpl_568 | and_dcpl_570
      | and_dcpl_572 | and_dcpl_576 | and_dcpl_578 | and_dcpl_580 | and_dcpl_583
      | and_dcpl_586 | mux_tmp_393);
  assign result_and_21_cse = ccs_ccore_en & (and_dcpl_590 | and_dcpl_592 | and_dcpl_594
      | and_dcpl_596 | and_dcpl_599 | and_dcpl_601 | and_dcpl_603 | and_dcpl_607
      | and_dcpl_611 | mux_tmp_438);
  assign m_and_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_2;
  assign m_and_1_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_6;
  assign m_and_2_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_9;
  assign m_and_3_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_11;
  assign m_and_4_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_2;
  assign m_and_5_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_6;
  assign m_and_6_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_9;
  assign m_and_7_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_11;
  assign m_and_8_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_18 & (~ (result_rem_11cyc_st_9[0]));
  assign m_and_9_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_18 & (result_rem_11cyc_st_9[0]);
  assign m_and_10_cse = ccs_ccore_en & and_dcpl_4 & (result_rem_11cyc_st_9[3]) &
      (result_rem_11cyc_st_9[1]) & (~ (result_rem_11cyc_st_9[0]));
  assign m_and_11_cse = ccs_ccore_en & and_dcpl_30;
  assign m_and_12_cse = ccs_ccore_en & and_dcpl_32;
  assign m_and_13_cse = ccs_ccore_en & and_dcpl_35;
  assign m_and_14_cse = ccs_ccore_en & and_dcpl_37;
  assign m_and_15_cse = ccs_ccore_en & and_dcpl_39;
  assign m_and_16_cse = ccs_ccore_en & and_dcpl_40;
  assign m_and_17_cse = ccs_ccore_en & and_dcpl_41;
  assign m_and_18_cse = ccs_ccore_en & and_dcpl_42;
  assign m_and_19_cse = ccs_ccore_en & and_dcpl_45;
  assign m_and_20_cse = ccs_ccore_en & and_dcpl_47;
  assign m_and_21_cse = ccs_ccore_en & and_dcpl_50;
  assign m_and_22_cse = ccs_ccore_en & and_dcpl_55;
  assign m_and_23_cse = ccs_ccore_en & and_dcpl_58;
  assign m_and_24_cse = ccs_ccore_en & and_dcpl_60;
  assign m_and_25_cse = ccs_ccore_en & and_dcpl_62;
  assign m_and_26_cse = ccs_ccore_en & and_dcpl_65;
  assign m_and_27_cse = ccs_ccore_en & and_dcpl_68;
  assign m_and_28_cse = ccs_ccore_en & and_dcpl_70;
  assign m_and_29_cse = ccs_ccore_en & and_dcpl_72;
  assign m_and_30_cse = ccs_ccore_en & and_dcpl_74;
  assign m_and_31_cse = ccs_ccore_en & and_dcpl_75;
  assign m_and_32_cse = ccs_ccore_en & and_dcpl_76;
  assign m_and_33_cse = ccs_ccore_en & and_dcpl_81;
  assign m_and_34_cse = ccs_ccore_en & and_dcpl_84;
  assign m_and_35_cse = ccs_ccore_en & and_dcpl_86;
  assign m_and_36_cse = ccs_ccore_en & and_dcpl_88;
  assign m_and_37_cse = ccs_ccore_en & and_dcpl_91;
  assign m_and_38_cse = ccs_ccore_en & and_dcpl_94;
  assign m_and_39_cse = ccs_ccore_en & and_dcpl_96;
  assign m_and_40_cse = ccs_ccore_en & and_dcpl_98;
  assign m_and_41_cse = ccs_ccore_en & and_dcpl_100;
  assign m_and_42_cse = ccs_ccore_en & and_dcpl_101;
  assign m_and_43_cse = ccs_ccore_en & and_dcpl_102;
  assign m_and_44_cse = ccs_ccore_en & and_dcpl_107;
  assign m_and_45_cse = ccs_ccore_en & and_dcpl_110;
  assign m_and_46_cse = ccs_ccore_en & and_dcpl_112;
  assign m_and_47_cse = ccs_ccore_en & and_dcpl_114;
  assign m_and_48_cse = ccs_ccore_en & and_dcpl_116;
  assign m_and_49_cse = ccs_ccore_en & and_dcpl_117;
  assign m_and_50_cse = ccs_ccore_en & and_dcpl_118;
  assign m_and_51_cse = ccs_ccore_en & and_dcpl_119;
  assign m_and_52_cse = ccs_ccore_en & and_dcpl_122;
  assign m_and_53_cse = ccs_ccore_en & and_dcpl_125;
  assign m_and_54_cse = ccs_ccore_en & and_dcpl_127;
  assign m_and_55_cse = ccs_ccore_en & and_dcpl_132;
  assign m_and_56_cse = ccs_ccore_en & and_dcpl_135;
  assign m_and_57_cse = ccs_ccore_en & and_dcpl_137;
  assign m_and_58_cse = ccs_ccore_en & and_dcpl_139;
  assign m_and_59_cse = ccs_ccore_en & and_dcpl_142;
  assign m_and_60_cse = ccs_ccore_en & and_dcpl_145;
  assign m_and_61_cse = ccs_ccore_en & and_dcpl_147;
  assign m_and_62_cse = ccs_ccore_en & and_dcpl_149;
  assign m_and_63_cse = ccs_ccore_en & and_dcpl_151;
  assign m_and_64_cse = ccs_ccore_en & and_dcpl_152;
  assign m_and_65_cse = ccs_ccore_en & and_dcpl_153;
  assign m_and_66_cse = ccs_ccore_en & and_dcpl_158;
  assign m_and_67_cse = ccs_ccore_en & and_dcpl_160;
  assign m_and_68_cse = ccs_ccore_en & and_dcpl_163;
  assign m_and_69_cse = ccs_ccore_en & and_dcpl_165;
  assign m_and_70_cse = ccs_ccore_en & and_dcpl_168;
  assign m_and_71_cse = ccs_ccore_en & and_dcpl_170;
  assign m_and_72_cse = ccs_ccore_en & and_dcpl_173;
  assign m_and_73_cse = ccs_ccore_en & and_dcpl_175;
  assign m_and_74_cse = ccs_ccore_en & and_dcpl_177;
  assign m_and_75_cse = ccs_ccore_en & and_dcpl_178;
  assign m_and_76_cse = ccs_ccore_en & and_dcpl_179;
  assign m_and_77_cse = ccs_ccore_en & and_dcpl_184;
  assign m_and_78_cse = ccs_ccore_en & and_dcpl_186;
  assign m_and_79_cse = ccs_ccore_en & and_dcpl_189;
  assign m_and_80_cse = ccs_ccore_en & and_dcpl_191;
  assign m_and_81_cse = ccs_ccore_en & and_dcpl_194;
  assign m_and_82_cse = ccs_ccore_en & and_dcpl_196;
  assign m_and_83_cse = ccs_ccore_en & and_dcpl_199;
  assign m_and_84_cse = ccs_ccore_en & and_dcpl_201;
  assign m_and_85_cse = ccs_ccore_en & and_dcpl_203;
  assign m_and_86_cse = ccs_ccore_en & and_dcpl_204;
  assign m_and_87_cse = ccs_ccore_en & and_dcpl_205;
  assign m_and_88_cse = ccs_ccore_en & and_dcpl_209 & and_dcpl_207;
  assign m_and_89_cse = ccs_ccore_en & and_dcpl_209 & and_dcpl_212;
  assign m_and_90_cse = ccs_ccore_en & and_dcpl_209 & and_dcpl_214;
  assign m_and_91_cse = ccs_ccore_en & and_dcpl_209 & and_dcpl_211 & (result_rem_11cyc[1]);
  assign m_and_92_cse = ccs_ccore_en & and_dcpl_209 & and_dcpl_218 & (~ (result_rem_11cyc[1]));
  assign m_and_93_cse = ccs_ccore_en & and_dcpl_209 & and_dcpl_221 & (~ (result_rem_11cyc[1]));
  assign m_and_94_cse = ccs_ccore_en & and_dcpl_209 & and_dcpl_218 & (result_rem_11cyc[1]);
  assign m_and_95_cse = ccs_ccore_en & and_dcpl_209 & and_dcpl_221 & (result_rem_11cyc[1]);
  assign m_and_96_cse = ccs_ccore_en & and_dcpl_228 & and_dcpl_207;
  assign m_and_97_cse = ccs_ccore_en & and_dcpl_228 & and_dcpl_212;
  assign m_and_98_cse = ccs_ccore_en & and_dcpl_228 & and_dcpl_214;
  assign nl_result_result_acc_tmp = conv_u2u_2_4(signext_2_1(result_acc_imod_1[3]))
      + conv_u2u_3_4(result_acc_imod_1[2:0]);
  assign result_result_acc_tmp = nl_result_result_acc_tmp[3:0];
  assign nl_result_acc_imod_1 = conv_u2s_3_4(result_acc_idiv_1[2:0]) + conv_u2s_3_4({(~
      (result_acc_idiv_1[3])) , 2'b00}) + conv_s2s_3_4({2'b10 , (result_acc_idiv_1[3])});
  assign result_acc_imod_1 = nl_result_acc_imod_1[3:0];
  assign nl_result_acc_idiv_1 = result_rem_11cyc + 4'b0001;
  assign result_acc_idiv_1 = nl_result_acc_idiv_1[3:0];
  assign and_dcpl_1 = ~((result_rem_11cyc_st_9[3]) | (result_rem_11cyc_st_9[1]));
  assign and_dcpl_2 = and_dcpl_1 & (~ (result_rem_11cyc_st_9[0]));
  assign and_dcpl_3 = main_stage_0_10 & asn_itm_9;
  assign and_dcpl_4 = and_dcpl_3 & (~ (result_rem_11cyc_st_9[2]));
  assign and_dcpl_6 = and_dcpl_1 & (result_rem_11cyc_st_9[0]);
  assign and_dcpl_8 = (~ (result_rem_11cyc_st_9[3])) & (result_rem_11cyc_st_9[1]);
  assign and_dcpl_9 = and_dcpl_8 & (~ (result_rem_11cyc_st_9[0]));
  assign and_dcpl_11 = and_dcpl_8 & (result_rem_11cyc_st_9[0]);
  assign and_dcpl_13 = and_dcpl_3 & (result_rem_11cyc_st_9[2]);
  assign and_dcpl_18 = (result_rem_11cyc_st_9[3]) & (~ (result_rem_11cyc_st_9[1]));
  assign and_dcpl_26 = ~((result_rem_11cyc_st_8[3]) | (result_rem_11cyc_st_8[1]));
  assign and_dcpl_27 = and_dcpl_26 & (~ (result_rem_11cyc_st_8[0]));
  assign and_dcpl_28 = main_stage_0_9 & asn_itm_8;
  assign and_dcpl_29 = and_dcpl_28 & (~ (result_rem_11cyc_st_8[2]));
  assign and_dcpl_30 = and_dcpl_29 & and_dcpl_27;
  assign and_dcpl_31 = and_dcpl_26 & (result_rem_11cyc_st_8[0]);
  assign and_dcpl_32 = and_dcpl_29 & and_dcpl_31;
  assign and_dcpl_33 = (~ (result_rem_11cyc_st_8[3])) & (result_rem_11cyc_st_8[1]);
  assign and_dcpl_34 = and_dcpl_33 & (~ (result_rem_11cyc_st_8[0]));
  assign and_dcpl_35 = and_dcpl_29 & and_dcpl_34;
  assign and_dcpl_36 = and_dcpl_33 & (result_rem_11cyc_st_8[0]);
  assign and_dcpl_37 = and_dcpl_29 & and_dcpl_36;
  assign and_dcpl_38 = and_dcpl_28 & (result_rem_11cyc_st_8[2]);
  assign and_dcpl_39 = and_dcpl_38 & and_dcpl_27;
  assign and_dcpl_40 = and_dcpl_38 & and_dcpl_31;
  assign and_dcpl_41 = and_dcpl_38 & and_dcpl_34;
  assign and_dcpl_42 = and_dcpl_38 & and_dcpl_36;
  assign and_dcpl_43 = (result_rem_11cyc_st_8[3]) & (~ (result_rem_11cyc_st_8[1]));
  assign and_dcpl_45 = and_dcpl_29 & and_dcpl_43 & (~ (result_rem_11cyc_st_8[0]));
  assign and_dcpl_47 = and_dcpl_29 & and_dcpl_43 & (result_rem_11cyc_st_8[0]);
  assign and_dcpl_50 = and_dcpl_29 & (result_rem_11cyc_st_8[3]) & (result_rem_11cyc_st_8[1])
      & (~ (result_rem_11cyc_st_8[0]));
  assign and_dcpl_51 = ~((result_rem_11cyc_st_7[2]) | (result_rem_11cyc_st_7[0]));
  assign and_dcpl_52 = and_dcpl_51 & (~ (result_rem_11cyc_st_7[1]));
  assign and_dcpl_53 = main_stage_0_8 & asn_itm_7;
  assign and_dcpl_54 = and_dcpl_53 & (~ (result_rem_11cyc_st_7[3]));
  assign and_dcpl_55 = and_dcpl_54 & and_dcpl_52;
  assign and_dcpl_56 = (~ (result_rem_11cyc_st_7[2])) & (result_rem_11cyc_st_7[0]);
  assign and_dcpl_57 = and_dcpl_56 & (~ (result_rem_11cyc_st_7[1]));
  assign and_dcpl_58 = and_dcpl_54 & and_dcpl_57;
  assign and_dcpl_59 = and_dcpl_51 & (result_rem_11cyc_st_7[1]);
  assign and_dcpl_60 = and_dcpl_54 & and_dcpl_59;
  assign and_dcpl_62 = and_dcpl_54 & and_dcpl_56 & (result_rem_11cyc_st_7[1]);
  assign and_dcpl_63 = (result_rem_11cyc_st_7[2]) & (~ (result_rem_11cyc_st_7[0]));
  assign and_dcpl_65 = and_dcpl_54 & and_dcpl_63 & (~ (result_rem_11cyc_st_7[1]));
  assign and_dcpl_66 = (result_rem_11cyc_st_7[2]) & (result_rem_11cyc_st_7[0]);
  assign and_dcpl_68 = and_dcpl_54 & and_dcpl_66 & (~ (result_rem_11cyc_st_7[1]));
  assign and_dcpl_70 = and_dcpl_54 & and_dcpl_63 & (result_rem_11cyc_st_7[1]);
  assign and_dcpl_72 = and_dcpl_54 & and_dcpl_66 & (result_rem_11cyc_st_7[1]);
  assign and_dcpl_73 = and_dcpl_53 & (result_rem_11cyc_st_7[3]);
  assign and_dcpl_74 = and_dcpl_73 & and_dcpl_52;
  assign and_dcpl_75 = and_dcpl_73 & and_dcpl_57;
  assign and_dcpl_76 = and_dcpl_73 & and_dcpl_59;
  assign and_dcpl_77 = ~((result_rem_11cyc_st_6[2]) | (result_rem_11cyc_st_6[0]));
  assign and_dcpl_78 = and_dcpl_77 & (~ (result_rem_11cyc_st_6[1]));
  assign and_dcpl_79 = main_stage_0_7 & asn_itm_6;
  assign and_dcpl_80 = and_dcpl_79 & (~ (result_rem_11cyc_st_6[3]));
  assign and_dcpl_81 = and_dcpl_80 & and_dcpl_78;
  assign and_dcpl_82 = (~ (result_rem_11cyc_st_6[2])) & (result_rem_11cyc_st_6[0]);
  assign and_dcpl_83 = and_dcpl_82 & (~ (result_rem_11cyc_st_6[1]));
  assign and_dcpl_84 = and_dcpl_80 & and_dcpl_83;
  assign and_dcpl_85 = and_dcpl_77 & (result_rem_11cyc_st_6[1]);
  assign and_dcpl_86 = and_dcpl_80 & and_dcpl_85;
  assign and_dcpl_88 = and_dcpl_80 & and_dcpl_82 & (result_rem_11cyc_st_6[1]);
  assign and_dcpl_89 = (result_rem_11cyc_st_6[2]) & (~ (result_rem_11cyc_st_6[0]));
  assign and_dcpl_91 = and_dcpl_80 & and_dcpl_89 & (~ (result_rem_11cyc_st_6[1]));
  assign and_dcpl_92 = (result_rem_11cyc_st_6[2]) & (result_rem_11cyc_st_6[0]);
  assign and_dcpl_94 = and_dcpl_80 & and_dcpl_92 & (~ (result_rem_11cyc_st_6[1]));
  assign and_dcpl_96 = and_dcpl_80 & and_dcpl_89 & (result_rem_11cyc_st_6[1]);
  assign and_dcpl_98 = and_dcpl_80 & and_dcpl_92 & (result_rem_11cyc_st_6[1]);
  assign and_dcpl_99 = and_dcpl_79 & (result_rem_11cyc_st_6[3]);
  assign and_dcpl_100 = and_dcpl_99 & and_dcpl_78;
  assign and_dcpl_101 = and_dcpl_99 & and_dcpl_83;
  assign and_dcpl_102 = and_dcpl_99 & and_dcpl_85;
  assign and_dcpl_103 = ~((result_rem_11cyc_st_5[3]) | (result_rem_11cyc_st_5[0]));
  assign and_dcpl_104 = and_dcpl_103 & (~ (result_rem_11cyc_st_5[1]));
  assign and_dcpl_105 = main_stage_0_6 & asn_itm_5;
  assign and_dcpl_106 = and_dcpl_105 & (~ (result_rem_11cyc_st_5[2]));
  assign and_dcpl_107 = and_dcpl_106 & and_dcpl_104;
  assign and_dcpl_108 = (~ (result_rem_11cyc_st_5[3])) & (result_rem_11cyc_st_5[0]);
  assign and_dcpl_109 = and_dcpl_108 & (~ (result_rem_11cyc_st_5[1]));
  assign and_dcpl_110 = and_dcpl_106 & and_dcpl_109;
  assign and_dcpl_111 = and_dcpl_103 & (result_rem_11cyc_st_5[1]);
  assign and_dcpl_112 = and_dcpl_106 & and_dcpl_111;
  assign and_dcpl_113 = and_dcpl_108 & (result_rem_11cyc_st_5[1]);
  assign and_dcpl_114 = and_dcpl_106 & and_dcpl_113;
  assign and_dcpl_115 = and_dcpl_105 & (result_rem_11cyc_st_5[2]);
  assign and_dcpl_116 = and_dcpl_115 & and_dcpl_104;
  assign and_dcpl_117 = and_dcpl_115 & and_dcpl_109;
  assign and_dcpl_118 = and_dcpl_115 & and_dcpl_111;
  assign and_dcpl_119 = and_dcpl_115 & and_dcpl_113;
  assign and_dcpl_120 = (result_rem_11cyc_st_5[3]) & (~ (result_rem_11cyc_st_5[0]));
  assign and_dcpl_122 = and_dcpl_106 & and_dcpl_120 & (~ (result_rem_11cyc_st_5[1]));
  assign and_dcpl_125 = and_dcpl_106 & (result_rem_11cyc_st_5[3]) & (result_rem_11cyc_st_5[0])
      & (~ (result_rem_11cyc_st_5[1]));
  assign and_dcpl_127 = and_dcpl_106 & and_dcpl_120 & (result_rem_11cyc_st_5[1]);
  assign and_dcpl_128 = ~((result_rem_11cyc_st_4[2]) | (result_rem_11cyc_st_4[0]));
  assign and_dcpl_129 = and_dcpl_128 & (~ (result_rem_11cyc_st_4[1]));
  assign and_dcpl_130 = main_stage_0_5 & asn_itm_4;
  assign and_dcpl_131 = and_dcpl_130 & (~ (result_rem_11cyc_st_4[3]));
  assign and_dcpl_132 = and_dcpl_131 & and_dcpl_129;
  assign and_dcpl_133 = (~ (result_rem_11cyc_st_4[2])) & (result_rem_11cyc_st_4[0]);
  assign and_dcpl_134 = and_dcpl_133 & (~ (result_rem_11cyc_st_4[1]));
  assign and_dcpl_135 = and_dcpl_131 & and_dcpl_134;
  assign and_dcpl_136 = and_dcpl_128 & (result_rem_11cyc_st_4[1]);
  assign and_dcpl_137 = and_dcpl_131 & and_dcpl_136;
  assign and_dcpl_139 = and_dcpl_131 & and_dcpl_133 & (result_rem_11cyc_st_4[1]);
  assign and_dcpl_140 = (result_rem_11cyc_st_4[2]) & (~ (result_rem_11cyc_st_4[0]));
  assign and_dcpl_142 = and_dcpl_131 & and_dcpl_140 & (~ (result_rem_11cyc_st_4[1]));
  assign and_dcpl_143 = (result_rem_11cyc_st_4[2]) & (result_rem_11cyc_st_4[0]);
  assign and_dcpl_145 = and_dcpl_131 & and_dcpl_143 & (~ (result_rem_11cyc_st_4[1]));
  assign and_dcpl_147 = and_dcpl_131 & and_dcpl_140 & (result_rem_11cyc_st_4[1]);
  assign and_dcpl_149 = and_dcpl_131 & and_dcpl_143 & (result_rem_11cyc_st_4[1]);
  assign and_dcpl_150 = and_dcpl_130 & (result_rem_11cyc_st_4[3]);
  assign and_dcpl_151 = and_dcpl_150 & and_dcpl_129;
  assign and_dcpl_152 = and_dcpl_150 & and_dcpl_134;
  assign and_dcpl_153 = and_dcpl_150 & and_dcpl_136;
  assign and_dcpl_154 = ~((result_rem_11cyc_st_3[2:1]!=2'b00));
  assign and_dcpl_155 = and_dcpl_154 & (~ (result_rem_11cyc_st_3[0]));
  assign and_dcpl_156 = main_stage_0_4 & asn_itm_3;
  assign and_dcpl_157 = and_dcpl_156 & (~ (result_rem_11cyc_st_3[3]));
  assign and_dcpl_158 = and_dcpl_157 & and_dcpl_155;
  assign and_dcpl_159 = and_dcpl_154 & (result_rem_11cyc_st_3[0]);
  assign and_dcpl_160 = and_dcpl_157 & and_dcpl_159;
  assign and_dcpl_161 = (result_rem_11cyc_st_3[2:1]==2'b01);
  assign and_dcpl_162 = and_dcpl_161 & (~ (result_rem_11cyc_st_3[0]));
  assign and_dcpl_163 = and_dcpl_157 & and_dcpl_162;
  assign and_dcpl_165 = and_dcpl_157 & and_dcpl_161 & (result_rem_11cyc_st_3[0]);
  assign and_dcpl_166 = (result_rem_11cyc_st_3[2:1]==2'b10);
  assign and_dcpl_168 = and_dcpl_157 & and_dcpl_166 & (~ (result_rem_11cyc_st_3[0]));
  assign and_dcpl_170 = and_dcpl_157 & and_dcpl_166 & (result_rem_11cyc_st_3[0]);
  assign and_dcpl_171 = (result_rem_11cyc_st_3[2:1]==2'b11);
  assign and_dcpl_173 = and_dcpl_157 & and_dcpl_171 & (~ (result_rem_11cyc_st_3[0]));
  assign and_dcpl_175 = and_dcpl_157 & and_dcpl_171 & (result_rem_11cyc_st_3[0]);
  assign and_dcpl_176 = and_dcpl_156 & (result_rem_11cyc_st_3[3]);
  assign and_dcpl_177 = and_dcpl_176 & and_dcpl_155;
  assign and_dcpl_178 = and_dcpl_176 & and_dcpl_159;
  assign and_dcpl_179 = and_dcpl_176 & and_dcpl_162;
  assign and_dcpl_180 = ~((result_rem_11cyc_st_2[2:1]!=2'b00));
  assign and_dcpl_181 = and_dcpl_180 & (~ (result_rem_11cyc_st_2[0]));
  assign and_dcpl_182 = main_stage_0_3 & asn_itm_2;
  assign and_dcpl_183 = and_dcpl_182 & (~ (result_rem_11cyc_st_2[3]));
  assign and_dcpl_184 = and_dcpl_183 & and_dcpl_181;
  assign and_dcpl_185 = and_dcpl_180 & (result_rem_11cyc_st_2[0]);
  assign and_dcpl_186 = and_dcpl_183 & and_dcpl_185;
  assign and_dcpl_187 = (result_rem_11cyc_st_2[2:1]==2'b01);
  assign and_dcpl_188 = and_dcpl_187 & (~ (result_rem_11cyc_st_2[0]));
  assign and_dcpl_189 = and_dcpl_183 & and_dcpl_188;
  assign and_dcpl_191 = and_dcpl_183 & and_dcpl_187 & (result_rem_11cyc_st_2[0]);
  assign and_dcpl_192 = (result_rem_11cyc_st_2[2:1]==2'b10);
  assign and_dcpl_194 = and_dcpl_183 & and_dcpl_192 & (~ (result_rem_11cyc_st_2[0]));
  assign and_dcpl_196 = and_dcpl_183 & and_dcpl_192 & (result_rem_11cyc_st_2[0]);
  assign and_dcpl_197 = (result_rem_11cyc_st_2[2:1]==2'b11);
  assign and_dcpl_199 = and_dcpl_183 & and_dcpl_197 & (~ (result_rem_11cyc_st_2[0]));
  assign and_dcpl_201 = and_dcpl_183 & and_dcpl_197 & (result_rem_11cyc_st_2[0]);
  assign and_dcpl_202 = and_dcpl_182 & (result_rem_11cyc_st_2[3]);
  assign and_dcpl_203 = and_dcpl_202 & and_dcpl_181;
  assign and_dcpl_204 = and_dcpl_202 & and_dcpl_185;
  assign and_dcpl_205 = and_dcpl_202 & and_dcpl_188;
  assign and_dcpl_206 = ~((result_rem_11cyc[2]) | (result_rem_11cyc[0]));
  assign and_dcpl_207 = and_dcpl_206 & (~ (result_rem_11cyc[1]));
  assign and_dcpl_208 = main_stage_0_2 & asn_itm_1;
  assign and_dcpl_209 = and_dcpl_208 & (~ (result_rem_11cyc[3]));
  assign and_dcpl_211 = (~ (result_rem_11cyc[2])) & (result_rem_11cyc[0]);
  assign and_dcpl_212 = and_dcpl_211 & (~ (result_rem_11cyc[1]));
  assign and_dcpl_214 = and_dcpl_206 & (result_rem_11cyc[1]);
  assign and_dcpl_218 = (result_rem_11cyc[2]) & (~ (result_rem_11cyc[0]));
  assign and_dcpl_221 = (result_rem_11cyc[2]) & (result_rem_11cyc[0]);
  assign and_dcpl_228 = and_dcpl_208 & (result_rem_11cyc[3]);
  assign and_dcpl_232 = ~((result_rem_11cyc_st_11[2:1]!=2'b00));
  assign and_dcpl_233 = and_dcpl_232 & (~ (result_rem_11cyc_st_11[0]));
  assign and_dcpl_234 = main_stage_0_12 & asn_itm_11;
  assign and_dcpl_235 = and_dcpl_234 & (~ (result_rem_11cyc_st_11[3]));
  assign and_dcpl_237 = and_dcpl_232 & (result_rem_11cyc_st_11[0]);
  assign and_dcpl_239 = (result_rem_11cyc_st_11[2:1]==2'b01);
  assign and_dcpl_240 = and_dcpl_239 & (~ (result_rem_11cyc_st_11[0]));
  assign and_dcpl_244 = (result_rem_11cyc_st_11[2:1]==2'b10);
  assign and_dcpl_249 = (result_rem_11cyc_st_11[2:1]==2'b11);
  assign and_dcpl_254 = and_dcpl_234 & (result_rem_11cyc_st_11[3]);
  assign and_dcpl_260 = ~((result_result_acc_tmp[1:0]!=2'b00));
  assign and_dcpl_261 = ccs_ccore_start_rsci_idat & (~ (result_result_acc_tmp[2]));
  assign and_dcpl_262 = and_dcpl_261 & (~ (result_result_acc_tmp[3]));
  assign and_dcpl_263 = and_dcpl_262 & and_dcpl_260;
  assign or_tmp_2 = (result_rem_11cyc!=4'b0000) | (~ and_dcpl_208);
  assign or_3_cse = (result_result_acc_tmp!=4'b0000);
  assign nor_691_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_2));
  assign mux_nl = MUX_s_1_2_2(nor_691_nl, or_tmp_2, or_3_cse);
  assign and_dcpl_269 = mux_nl & and_dcpl_184;
  assign or_8_cse = (result_rem_11cyc!=4'b0000);
  assign nor_690_nl = ~(and_dcpl_208 | and_dcpl_184);
  assign or_10_nl = (result_rem_11cyc_st_2!=4'b0000) | (~ and_dcpl_182);
  assign mux_tmp_1 = MUX_s_1_2_2(nor_690_nl, or_10_nl, or_8_cse);
  assign nor_689_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_1));
  assign mux_2_nl = MUX_s_1_2_2(nor_689_nl, mux_tmp_1, or_3_cse);
  assign and_dcpl_275 = mux_2_nl & and_dcpl_158;
  assign or_15_cse = (result_rem_11cyc_st_2!=4'b0000);
  assign nor_687_nl = ~(and_dcpl_182 | and_dcpl_158);
  assign or_17_nl = (result_rem_11cyc_st_3!=4'b0000) | (~ and_dcpl_156);
  assign mux_tmp_3 = MUX_s_1_2_2(nor_687_nl, or_17_nl, or_15_cse);
  assign nor_688_nl = ~(and_dcpl_208 | (~ mux_tmp_3));
  assign mux_tmp_4 = MUX_s_1_2_2(nor_688_nl, mux_tmp_3, or_8_cse);
  assign nor_686_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_4));
  assign mux_5_nl = MUX_s_1_2_2(nor_686_nl, mux_tmp_4, or_3_cse);
  assign and_dcpl_281 = mux_5_nl & and_dcpl_132;
  assign or_24_cse = (result_rem_11cyc_st_3!=4'b0000);
  assign nor_683_nl = ~(and_dcpl_156 | and_dcpl_132);
  assign or_26_nl = (result_rem_11cyc_st_4!=4'b0000) | (~ and_dcpl_130);
  assign mux_tmp_6 = MUX_s_1_2_2(nor_683_nl, or_26_nl, or_24_cse);
  assign nor_684_nl = ~(and_dcpl_182 | (~ mux_tmp_6));
  assign mux_tmp_7 = MUX_s_1_2_2(nor_684_nl, mux_tmp_6, or_15_cse);
  assign nor_685_nl = ~(and_dcpl_208 | (~ mux_tmp_7));
  assign mux_tmp_8 = MUX_s_1_2_2(nor_685_nl, mux_tmp_7, or_8_cse);
  assign nor_682_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_8));
  assign mux_9_nl = MUX_s_1_2_2(nor_682_nl, mux_tmp_8, or_3_cse);
  assign and_dcpl_287 = mux_9_nl & and_dcpl_107;
  assign or_35_cse = (result_rem_11cyc_st_4!=4'b0000);
  assign nor_678_nl = ~(and_dcpl_130 | and_dcpl_107);
  assign or_37_nl = (result_rem_11cyc_st_5!=4'b0000) | (~ and_dcpl_105);
  assign mux_tmp_10 = MUX_s_1_2_2(nor_678_nl, or_37_nl, or_35_cse);
  assign nor_679_nl = ~(and_dcpl_156 | (~ mux_tmp_10));
  assign mux_tmp_11 = MUX_s_1_2_2(nor_679_nl, mux_tmp_10, or_24_cse);
  assign nor_680_nl = ~(and_dcpl_182 | (~ mux_tmp_11));
  assign mux_tmp_12 = MUX_s_1_2_2(nor_680_nl, mux_tmp_11, or_15_cse);
  assign nor_681_nl = ~(and_dcpl_208 | (~ mux_tmp_12));
  assign mux_tmp_13 = MUX_s_1_2_2(nor_681_nl, mux_tmp_12, or_8_cse);
  assign nor_677_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_13));
  assign mux_14_nl = MUX_s_1_2_2(nor_677_nl, mux_tmp_13, or_3_cse);
  assign and_dcpl_293 = mux_14_nl & and_dcpl_81;
  assign or_48_cse = (result_rem_11cyc_st_5!=4'b0000);
  assign nor_672_nl = ~(and_dcpl_105 | and_dcpl_81);
  assign or_50_nl = (result_rem_11cyc_st_6!=4'b0000) | (~ and_dcpl_79);
  assign mux_tmp_15 = MUX_s_1_2_2(nor_672_nl, or_50_nl, or_48_cse);
  assign nor_673_nl = ~(and_dcpl_130 | (~ mux_tmp_15));
  assign mux_tmp_16 = MUX_s_1_2_2(nor_673_nl, mux_tmp_15, or_35_cse);
  assign nor_674_nl = ~(and_dcpl_156 | (~ mux_tmp_16));
  assign mux_tmp_17 = MUX_s_1_2_2(nor_674_nl, mux_tmp_16, or_24_cse);
  assign nor_675_nl = ~(and_dcpl_182 | (~ mux_tmp_17));
  assign mux_tmp_18 = MUX_s_1_2_2(nor_675_nl, mux_tmp_17, or_15_cse);
  assign nor_676_nl = ~(and_dcpl_208 | (~ mux_tmp_18));
  assign mux_tmp_19 = MUX_s_1_2_2(nor_676_nl, mux_tmp_18, or_8_cse);
  assign nor_671_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_19));
  assign mux_20_nl = MUX_s_1_2_2(nor_671_nl, mux_tmp_19, or_3_cse);
  assign and_dcpl_299 = mux_20_nl & and_dcpl_55;
  assign or_63_cse = (result_rem_11cyc_st_6!=4'b0000);
  assign nor_665_nl = ~(and_dcpl_79 | and_dcpl_55);
  assign or_65_nl = (result_rem_11cyc_st_7!=4'b0000) | (~ and_dcpl_53);
  assign mux_tmp_21 = MUX_s_1_2_2(nor_665_nl, or_65_nl, or_63_cse);
  assign nor_666_nl = ~(and_dcpl_105 | (~ mux_tmp_21));
  assign mux_tmp_22 = MUX_s_1_2_2(nor_666_nl, mux_tmp_21, or_48_cse);
  assign nor_667_nl = ~(and_dcpl_130 | (~ mux_tmp_22));
  assign mux_tmp_23 = MUX_s_1_2_2(nor_667_nl, mux_tmp_22, or_35_cse);
  assign nor_668_nl = ~(and_dcpl_156 | (~ mux_tmp_23));
  assign mux_tmp_24 = MUX_s_1_2_2(nor_668_nl, mux_tmp_23, or_24_cse);
  assign nor_669_nl = ~(and_dcpl_182 | (~ mux_tmp_24));
  assign mux_tmp_25 = MUX_s_1_2_2(nor_669_nl, mux_tmp_24, or_15_cse);
  assign nor_670_nl = ~(and_dcpl_208 | (~ mux_tmp_25));
  assign mux_tmp_26 = MUX_s_1_2_2(nor_670_nl, mux_tmp_25, or_8_cse);
  assign nor_664_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_26));
  assign mux_27_nl = MUX_s_1_2_2(nor_664_nl, mux_tmp_26, or_3_cse);
  assign and_dcpl_305 = mux_27_nl & and_dcpl_30;
  assign nor_656_nl = ~(and_dcpl_53 | and_dcpl_30);
  assign or_82_nl = (result_rem_11cyc_st_8!=4'b0000) | (~ and_dcpl_28);
  assign or_80_nl = (result_rem_11cyc_st_7!=4'b0000);
  assign mux_tmp_28 = MUX_s_1_2_2(nor_656_nl, or_82_nl, or_80_nl);
  assign nor_657_nl = ~(and_dcpl_79 | (~ mux_tmp_28));
  assign mux_tmp_29 = MUX_s_1_2_2(nor_657_nl, mux_tmp_28, or_63_cse);
  assign nor_658_nl = ~(and_dcpl_105 | (~ mux_tmp_29));
  assign mux_tmp_30 = MUX_s_1_2_2(nor_658_nl, mux_tmp_29, or_48_cse);
  assign nor_659_nl = ~(and_dcpl_130 | (~ mux_tmp_30));
  assign mux_tmp_31 = MUX_s_1_2_2(nor_659_nl, mux_tmp_30, or_35_cse);
  assign nor_660_nl = ~(and_dcpl_156 | (~ mux_tmp_31));
  assign mux_tmp_32 = MUX_s_1_2_2(nor_660_nl, mux_tmp_31, or_24_cse);
  assign nor_661_nl = ~(and_dcpl_182 | (~ mux_tmp_32));
  assign mux_tmp_33 = MUX_s_1_2_2(nor_661_nl, mux_tmp_32, or_15_cse);
  assign nor_662_nl = ~(and_dcpl_208 | (~ mux_tmp_33));
  assign mux_tmp_34 = MUX_s_1_2_2(nor_662_nl, mux_tmp_33, or_8_cse);
  assign nor_663_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_34));
  assign mux_35_nl = MUX_s_1_2_2(nor_663_nl, mux_tmp_34, or_3_cse);
  assign and_dcpl_311 = mux_35_nl & and_dcpl_4 & and_dcpl_2;
  assign and_tmp_6 = ((~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2!=4'b0000))
      & ((~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3!=4'b0000)) &
      ((~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4!=4'b0000)) & ((~
      main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5!=4'b0000)) & ((~ main_stage_0_7)
      | (~ asn_itm_6) | (result_rem_11cyc_st_6!=4'b0000)) & ((~ main_stage_0_8) |
      (~ asn_itm_7) | (result_rem_11cyc_st_7!=4'b0000)) & ((~ main_stage_0_9) | (~
      asn_itm_8) | (result_rem_11cyc_st_8!=4'b0000)) & ((~ main_stage_0_10) | (~
      asn_itm_9) | (result_rem_11cyc_st_9!=4'b0000));
  assign nor_654_nl = ~(and_dcpl_208 | (~ and_tmp_6));
  assign mux_tmp_36 = MUX_s_1_2_2(nor_654_nl, and_tmp_6, or_8_cse);
  assign nor_655_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_36));
  assign mux_tmp_37 = MUX_s_1_2_2(nor_655_nl, mux_tmp_36, or_3_cse);
  assign and_dcpl_318 = (result_result_acc_tmp[1:0]==2'b01);
  assign and_dcpl_319 = and_dcpl_262 & and_dcpl_318;
  assign or_tmp_102 = (result_rem_11cyc!=4'b0001) | (~ and_dcpl_208);
  assign or_107_cse = (result_result_acc_tmp!=4'b0001);
  assign nor_653_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_102));
  assign mux_38_nl = MUX_s_1_2_2(nor_653_nl, or_tmp_102, or_107_cse);
  assign and_dcpl_322 = mux_38_nl & and_dcpl_186;
  assign or_112_cse = (result_rem_11cyc!=4'b0001);
  assign nor_652_nl = ~(and_dcpl_208 | and_dcpl_186);
  assign or_114_nl = (result_rem_11cyc_st_2!=4'b0001) | (~ and_dcpl_182);
  assign mux_tmp_39 = MUX_s_1_2_2(nor_652_nl, or_114_nl, or_112_cse);
  assign nor_651_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_39));
  assign mux_40_nl = MUX_s_1_2_2(nor_651_nl, mux_tmp_39, or_107_cse);
  assign and_dcpl_325 = mux_40_nl & and_dcpl_160;
  assign or_119_cse = (result_rem_11cyc_st_2!=4'b0001);
  assign nor_649_nl = ~(and_dcpl_182 | and_dcpl_160);
  assign or_121_nl = (result_rem_11cyc_st_3!=4'b0001) | (~ and_dcpl_156);
  assign mux_tmp_41 = MUX_s_1_2_2(nor_649_nl, or_121_nl, or_119_cse);
  assign nor_650_nl = ~(and_dcpl_208 | (~ mux_tmp_41));
  assign mux_tmp_42 = MUX_s_1_2_2(nor_650_nl, mux_tmp_41, or_112_cse);
  assign nor_648_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_42));
  assign mux_43_nl = MUX_s_1_2_2(nor_648_nl, mux_tmp_42, or_107_cse);
  assign and_dcpl_329 = mux_43_nl & and_dcpl_135;
  assign or_128_cse = (result_rem_11cyc_st_3!=4'b0001);
  assign nor_645_nl = ~(and_dcpl_156 | and_dcpl_135);
  assign or_130_nl = (result_rem_11cyc_st_4!=4'b0001) | (~ and_dcpl_130);
  assign mux_tmp_44 = MUX_s_1_2_2(nor_645_nl, or_130_nl, or_128_cse);
  assign nor_646_nl = ~(and_dcpl_182 | (~ mux_tmp_44));
  assign mux_tmp_45 = MUX_s_1_2_2(nor_646_nl, mux_tmp_44, or_119_cse);
  assign nor_647_nl = ~(and_dcpl_208 | (~ mux_tmp_45));
  assign mux_tmp_46 = MUX_s_1_2_2(nor_647_nl, mux_tmp_45, or_112_cse);
  assign nor_644_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_46));
  assign mux_47_nl = MUX_s_1_2_2(nor_644_nl, mux_tmp_46, or_107_cse);
  assign and_dcpl_333 = mux_47_nl & and_dcpl_110;
  assign or_139_cse = (result_rem_11cyc_st_4!=4'b0001);
  assign nor_640_nl = ~(and_dcpl_130 | and_dcpl_110);
  assign or_141_nl = (result_rem_11cyc_st_5!=4'b0001) | (~ and_dcpl_105);
  assign mux_tmp_48 = MUX_s_1_2_2(nor_640_nl, or_141_nl, or_139_cse);
  assign nor_641_nl = ~(and_dcpl_156 | (~ mux_tmp_48));
  assign mux_tmp_49 = MUX_s_1_2_2(nor_641_nl, mux_tmp_48, or_128_cse);
  assign nor_642_nl = ~(and_dcpl_182 | (~ mux_tmp_49));
  assign mux_tmp_50 = MUX_s_1_2_2(nor_642_nl, mux_tmp_49, or_119_cse);
  assign nor_643_nl = ~(and_dcpl_208 | (~ mux_tmp_50));
  assign mux_tmp_51 = MUX_s_1_2_2(nor_643_nl, mux_tmp_50, or_112_cse);
  assign nor_639_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_51));
  assign mux_52_nl = MUX_s_1_2_2(nor_639_nl, mux_tmp_51, or_107_cse);
  assign and_dcpl_337 = mux_52_nl & and_dcpl_84;
  assign or_152_cse = (result_rem_11cyc_st_5!=4'b0001);
  assign nor_634_nl = ~(and_dcpl_105 | and_dcpl_84);
  assign or_154_nl = (result_rem_11cyc_st_6!=4'b0001) | (~ and_dcpl_79);
  assign mux_tmp_53 = MUX_s_1_2_2(nor_634_nl, or_154_nl, or_152_cse);
  assign nor_635_nl = ~(and_dcpl_130 | (~ mux_tmp_53));
  assign mux_tmp_54 = MUX_s_1_2_2(nor_635_nl, mux_tmp_53, or_139_cse);
  assign nor_636_nl = ~(and_dcpl_156 | (~ mux_tmp_54));
  assign mux_tmp_55 = MUX_s_1_2_2(nor_636_nl, mux_tmp_54, or_128_cse);
  assign nor_637_nl = ~(and_dcpl_182 | (~ mux_tmp_55));
  assign mux_tmp_56 = MUX_s_1_2_2(nor_637_nl, mux_tmp_55, or_119_cse);
  assign nor_638_nl = ~(and_dcpl_208 | (~ mux_tmp_56));
  assign mux_tmp_57 = MUX_s_1_2_2(nor_638_nl, mux_tmp_56, or_112_cse);
  assign nor_633_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_57));
  assign mux_58_nl = MUX_s_1_2_2(nor_633_nl, mux_tmp_57, or_107_cse);
  assign and_dcpl_341 = mux_58_nl & and_dcpl_58;
  assign or_167_cse = (result_rem_11cyc_st_6!=4'b0001);
  assign nor_627_nl = ~(and_dcpl_79 | and_dcpl_58);
  assign or_169_nl = (result_rem_11cyc_st_7!=4'b0001) | (~ and_dcpl_53);
  assign mux_tmp_59 = MUX_s_1_2_2(nor_627_nl, or_169_nl, or_167_cse);
  assign nor_628_nl = ~(and_dcpl_105 | (~ mux_tmp_59));
  assign mux_tmp_60 = MUX_s_1_2_2(nor_628_nl, mux_tmp_59, or_152_cse);
  assign nor_629_nl = ~(and_dcpl_130 | (~ mux_tmp_60));
  assign mux_tmp_61 = MUX_s_1_2_2(nor_629_nl, mux_tmp_60, or_139_cse);
  assign nor_630_nl = ~(and_dcpl_156 | (~ mux_tmp_61));
  assign mux_tmp_62 = MUX_s_1_2_2(nor_630_nl, mux_tmp_61, or_128_cse);
  assign nor_631_nl = ~(and_dcpl_182 | (~ mux_tmp_62));
  assign mux_tmp_63 = MUX_s_1_2_2(nor_631_nl, mux_tmp_62, or_119_cse);
  assign nor_632_nl = ~(and_dcpl_208 | (~ mux_tmp_63));
  assign mux_tmp_64 = MUX_s_1_2_2(nor_632_nl, mux_tmp_63, or_112_cse);
  assign nor_626_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_64));
  assign mux_65_nl = MUX_s_1_2_2(nor_626_nl, mux_tmp_64, or_107_cse);
  assign and_dcpl_344 = mux_65_nl & and_dcpl_32;
  assign nor_618_nl = ~(and_dcpl_53 | and_dcpl_32);
  assign or_186_nl = (result_rem_11cyc_st_8!=4'b0001) | (~ and_dcpl_28);
  assign or_184_nl = (result_rem_11cyc_st_7!=4'b0001);
  assign mux_tmp_66 = MUX_s_1_2_2(nor_618_nl, or_186_nl, or_184_nl);
  assign nor_619_nl = ~(and_dcpl_79 | (~ mux_tmp_66));
  assign mux_tmp_67 = MUX_s_1_2_2(nor_619_nl, mux_tmp_66, or_167_cse);
  assign nor_620_nl = ~(and_dcpl_105 | (~ mux_tmp_67));
  assign mux_tmp_68 = MUX_s_1_2_2(nor_620_nl, mux_tmp_67, or_152_cse);
  assign nor_621_nl = ~(and_dcpl_130 | (~ mux_tmp_68));
  assign mux_tmp_69 = MUX_s_1_2_2(nor_621_nl, mux_tmp_68, or_139_cse);
  assign nor_622_nl = ~(and_dcpl_156 | (~ mux_tmp_69));
  assign mux_tmp_70 = MUX_s_1_2_2(nor_622_nl, mux_tmp_69, or_128_cse);
  assign nor_623_nl = ~(and_dcpl_182 | (~ mux_tmp_70));
  assign mux_tmp_71 = MUX_s_1_2_2(nor_623_nl, mux_tmp_70, or_119_cse);
  assign nor_624_nl = ~(and_dcpl_208 | (~ mux_tmp_71));
  assign mux_tmp_72 = MUX_s_1_2_2(nor_624_nl, mux_tmp_71, or_112_cse);
  assign nor_625_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_72));
  assign mux_73_nl = MUX_s_1_2_2(nor_625_nl, mux_tmp_72, or_107_cse);
  assign and_dcpl_347 = mux_73_nl & and_dcpl_4 & and_dcpl_6;
  assign and_tmp_13 = ((~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2!=4'b0001))
      & ((~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3!=4'b0001)) &
      ((~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4!=4'b0001)) & ((~
      main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5!=4'b0001)) & ((~ main_stage_0_7)
      | (~ asn_itm_6) | (result_rem_11cyc_st_6!=4'b0001)) & ((~ main_stage_0_8) |
      (~ asn_itm_7) | (result_rem_11cyc_st_7!=4'b0001)) & ((~ main_stage_0_9) | (~
      asn_itm_8) | (result_rem_11cyc_st_8!=4'b0001)) & ((~ main_stage_0_10) | (~
      asn_itm_9) | (result_rem_11cyc_st_9!=4'b0001));
  assign nor_617_nl = ~(and_dcpl_208 | (~ and_tmp_13));
  assign mux_tmp_74 = MUX_s_1_2_2(nor_617_nl, and_tmp_13, or_112_cse);
  assign nand_146_cse = ~((result_result_acc_tmp[0]) & ccs_ccore_start_rsci_idat);
  assign and_797_nl = nand_146_cse & mux_tmp_74;
  assign or_195_nl = (result_result_acc_tmp[3:1]!=3'b000);
  assign mux_tmp_75 = MUX_s_1_2_2(and_797_nl, mux_tmp_74, or_195_nl);
  assign and_dcpl_352 = (result_result_acc_tmp[1:0]==2'b10);
  assign and_dcpl_353 = and_dcpl_262 & and_dcpl_352;
  assign or_tmp_202 = (result_rem_11cyc!=4'b0010) | (~ and_dcpl_208);
  assign or_209_cse = (result_result_acc_tmp!=4'b0010);
  assign nor_616_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_202));
  assign mux_76_nl = MUX_s_1_2_2(nor_616_nl, or_tmp_202, or_209_cse);
  assign and_dcpl_357 = mux_76_nl & and_dcpl_189;
  assign or_214_cse = (result_rem_11cyc!=4'b0010);
  assign nor_615_nl = ~(and_dcpl_208 | and_dcpl_189);
  assign or_216_nl = (result_rem_11cyc_st_2!=4'b0010) | (~ and_dcpl_182);
  assign mux_tmp_77 = MUX_s_1_2_2(nor_615_nl, or_216_nl, or_214_cse);
  assign nor_614_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_77));
  assign mux_78_nl = MUX_s_1_2_2(nor_614_nl, mux_tmp_77, or_209_cse);
  assign and_dcpl_361 = mux_78_nl & and_dcpl_163;
  assign or_221_cse = (result_rem_11cyc_st_2!=4'b0010);
  assign nor_612_nl = ~(and_dcpl_182 | and_dcpl_163);
  assign or_223_nl = (result_rem_11cyc_st_3!=4'b0010) | (~ and_dcpl_156);
  assign mux_tmp_79 = MUX_s_1_2_2(nor_612_nl, or_223_nl, or_221_cse);
  assign nor_613_nl = ~(and_dcpl_208 | (~ mux_tmp_79));
  assign mux_tmp_80 = MUX_s_1_2_2(nor_613_nl, mux_tmp_79, or_214_cse);
  assign nor_611_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_80));
  assign mux_81_nl = MUX_s_1_2_2(nor_611_nl, mux_tmp_80, or_209_cse);
  assign and_dcpl_364 = mux_81_nl & and_dcpl_137;
  assign or_230_cse = (result_rem_11cyc_st_3!=4'b0010);
  assign nor_608_nl = ~(and_dcpl_156 | and_dcpl_137);
  assign or_232_nl = (result_rem_11cyc_st_4!=4'b0010) | (~ and_dcpl_130);
  assign mux_tmp_82 = MUX_s_1_2_2(nor_608_nl, or_232_nl, or_230_cse);
  assign nor_609_nl = ~(and_dcpl_182 | (~ mux_tmp_82));
  assign mux_tmp_83 = MUX_s_1_2_2(nor_609_nl, mux_tmp_82, or_221_cse);
  assign nor_610_nl = ~(and_dcpl_208 | (~ mux_tmp_83));
  assign mux_tmp_84 = MUX_s_1_2_2(nor_610_nl, mux_tmp_83, or_214_cse);
  assign nor_607_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_84));
  assign mux_85_nl = MUX_s_1_2_2(nor_607_nl, mux_tmp_84, or_209_cse);
  assign and_dcpl_367 = mux_85_nl & and_dcpl_112;
  assign or_241_cse = (result_rem_11cyc_st_4!=4'b0010);
  assign nor_603_nl = ~(and_dcpl_130 | and_dcpl_112);
  assign or_243_nl = (result_rem_11cyc_st_5!=4'b0010) | (~ and_dcpl_105);
  assign mux_tmp_86 = MUX_s_1_2_2(nor_603_nl, or_243_nl, or_241_cse);
  assign nor_604_nl = ~(and_dcpl_156 | (~ mux_tmp_86));
  assign mux_tmp_87 = MUX_s_1_2_2(nor_604_nl, mux_tmp_86, or_230_cse);
  assign nor_605_nl = ~(and_dcpl_182 | (~ mux_tmp_87));
  assign mux_tmp_88 = MUX_s_1_2_2(nor_605_nl, mux_tmp_87, or_221_cse);
  assign nor_606_nl = ~(and_dcpl_208 | (~ mux_tmp_88));
  assign mux_tmp_89 = MUX_s_1_2_2(nor_606_nl, mux_tmp_88, or_214_cse);
  assign nor_602_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_89));
  assign mux_90_nl = MUX_s_1_2_2(nor_602_nl, mux_tmp_89, or_209_cse);
  assign and_dcpl_370 = mux_90_nl & and_dcpl_86;
  assign or_254_cse = (result_rem_11cyc_st_5!=4'b0010);
  assign nor_597_nl = ~(and_dcpl_105 | and_dcpl_86);
  assign or_256_nl = (result_rem_11cyc_st_6!=4'b0010) | (~ and_dcpl_79);
  assign mux_tmp_91 = MUX_s_1_2_2(nor_597_nl, or_256_nl, or_254_cse);
  assign nor_598_nl = ~(and_dcpl_130 | (~ mux_tmp_91));
  assign mux_tmp_92 = MUX_s_1_2_2(nor_598_nl, mux_tmp_91, or_241_cse);
  assign nor_599_nl = ~(and_dcpl_156 | (~ mux_tmp_92));
  assign mux_tmp_93 = MUX_s_1_2_2(nor_599_nl, mux_tmp_92, or_230_cse);
  assign nor_600_nl = ~(and_dcpl_182 | (~ mux_tmp_93));
  assign mux_tmp_94 = MUX_s_1_2_2(nor_600_nl, mux_tmp_93, or_221_cse);
  assign nor_601_nl = ~(and_dcpl_208 | (~ mux_tmp_94));
  assign mux_tmp_95 = MUX_s_1_2_2(nor_601_nl, mux_tmp_94, or_214_cse);
  assign nor_596_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_95));
  assign mux_96_nl = MUX_s_1_2_2(nor_596_nl, mux_tmp_95, or_209_cse);
  assign and_dcpl_373 = mux_96_nl & and_dcpl_60;
  assign or_269_cse = (result_rem_11cyc_st_6!=4'b0010);
  assign nor_590_nl = ~(and_dcpl_79 | and_dcpl_60);
  assign or_271_nl = (result_rem_11cyc_st_7!=4'b0010) | (~ and_dcpl_53);
  assign mux_tmp_97 = MUX_s_1_2_2(nor_590_nl, or_271_nl, or_269_cse);
  assign nor_591_nl = ~(and_dcpl_105 | (~ mux_tmp_97));
  assign mux_tmp_98 = MUX_s_1_2_2(nor_591_nl, mux_tmp_97, or_254_cse);
  assign nor_592_nl = ~(and_dcpl_130 | (~ mux_tmp_98));
  assign mux_tmp_99 = MUX_s_1_2_2(nor_592_nl, mux_tmp_98, or_241_cse);
  assign nor_593_nl = ~(and_dcpl_156 | (~ mux_tmp_99));
  assign mux_tmp_100 = MUX_s_1_2_2(nor_593_nl, mux_tmp_99, or_230_cse);
  assign nor_594_nl = ~(and_dcpl_182 | (~ mux_tmp_100));
  assign mux_tmp_101 = MUX_s_1_2_2(nor_594_nl, mux_tmp_100, or_221_cse);
  assign nor_595_nl = ~(and_dcpl_208 | (~ mux_tmp_101));
  assign mux_tmp_102 = MUX_s_1_2_2(nor_595_nl, mux_tmp_101, or_214_cse);
  assign nor_589_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_102));
  assign mux_103_nl = MUX_s_1_2_2(nor_589_nl, mux_tmp_102, or_209_cse);
  assign and_dcpl_377 = mux_103_nl & and_dcpl_35;
  assign nor_581_nl = ~(and_dcpl_53 | and_dcpl_35);
  assign or_288_nl = (result_rem_11cyc_st_8!=4'b0010) | (~ and_dcpl_28);
  assign or_286_nl = (result_rem_11cyc_st_7!=4'b0010);
  assign mux_tmp_104 = MUX_s_1_2_2(nor_581_nl, or_288_nl, or_286_nl);
  assign nor_582_nl = ~(and_dcpl_79 | (~ mux_tmp_104));
  assign mux_tmp_105 = MUX_s_1_2_2(nor_582_nl, mux_tmp_104, or_269_cse);
  assign nor_583_nl = ~(and_dcpl_105 | (~ mux_tmp_105));
  assign mux_tmp_106 = MUX_s_1_2_2(nor_583_nl, mux_tmp_105, or_254_cse);
  assign nor_584_nl = ~(and_dcpl_130 | (~ mux_tmp_106));
  assign mux_tmp_107 = MUX_s_1_2_2(nor_584_nl, mux_tmp_106, or_241_cse);
  assign nor_585_nl = ~(and_dcpl_156 | (~ mux_tmp_107));
  assign mux_tmp_108 = MUX_s_1_2_2(nor_585_nl, mux_tmp_107, or_230_cse);
  assign nor_586_nl = ~(and_dcpl_182 | (~ mux_tmp_108));
  assign mux_tmp_109 = MUX_s_1_2_2(nor_586_nl, mux_tmp_108, or_221_cse);
  assign nor_587_nl = ~(and_dcpl_208 | (~ mux_tmp_109));
  assign mux_tmp_110 = MUX_s_1_2_2(nor_587_nl, mux_tmp_109, or_214_cse);
  assign nor_588_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_110));
  assign mux_111_nl = MUX_s_1_2_2(nor_588_nl, mux_tmp_110, or_209_cse);
  assign and_dcpl_381 = mux_111_nl & and_dcpl_4 & and_dcpl_9;
  assign and_tmp_20 = ((~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2!=4'b0010))
      & ((~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3!=4'b0010)) &
      ((~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4!=4'b0010)) & ((~
      main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5!=4'b0010)) & ((~ main_stage_0_7)
      | (~ asn_itm_6) | (result_rem_11cyc_st_6!=4'b0010)) & ((~ main_stage_0_8) |
      (~ asn_itm_7) | (result_rem_11cyc_st_7!=4'b0010)) & ((~ main_stage_0_9) | (~
      asn_itm_8) | (result_rem_11cyc_st_8!=4'b0010)) & ((~ main_stage_0_10) | (~
      asn_itm_9) | (result_rem_11cyc_st_9!=4'b0010));
  assign nor_579_nl = ~(and_dcpl_208 | (~ and_tmp_20));
  assign mux_tmp_112 = MUX_s_1_2_2(nor_579_nl, and_tmp_20, or_214_cse);
  assign nor_580_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_112));
  assign mux_tmp_113 = MUX_s_1_2_2(nor_580_nl, mux_tmp_112, or_209_cse);
  assign and_dcpl_386 = (result_result_acc_tmp[1:0]==2'b11);
  assign and_dcpl_387 = and_dcpl_262 & and_dcpl_386;
  assign or_tmp_302 = (result_rem_11cyc!=4'b0011) | (~ and_dcpl_208);
  assign or_311_cse = (result_result_acc_tmp!=4'b0011);
  assign nor_578_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_302));
  assign mux_114_nl = MUX_s_1_2_2(nor_578_nl, or_tmp_302, or_311_cse);
  assign and_dcpl_390 = mux_114_nl & and_dcpl_191;
  assign or_316_cse = (result_rem_11cyc!=4'b0011);
  assign nor_577_nl = ~(and_dcpl_208 | and_dcpl_191);
  assign or_318_nl = (result_rem_11cyc_st_2!=4'b0011) | (~ and_dcpl_182);
  assign mux_tmp_115 = MUX_s_1_2_2(nor_577_nl, or_318_nl, or_316_cse);
  assign nor_576_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_115));
  assign mux_116_nl = MUX_s_1_2_2(nor_576_nl, mux_tmp_115, or_311_cse);
  assign and_dcpl_393 = mux_116_nl & and_dcpl_165;
  assign or_323_cse = (result_rem_11cyc_st_2!=4'b0011);
  assign nor_574_nl = ~(and_dcpl_182 | and_dcpl_165);
  assign or_325_nl = (result_rem_11cyc_st_3!=4'b0011) | (~ and_dcpl_156);
  assign mux_tmp_117 = MUX_s_1_2_2(nor_574_nl, or_325_nl, or_323_cse);
  assign nor_575_nl = ~(and_dcpl_208 | (~ mux_tmp_117));
  assign mux_tmp_118 = MUX_s_1_2_2(nor_575_nl, mux_tmp_117, or_316_cse);
  assign nor_573_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_118));
  assign mux_119_nl = MUX_s_1_2_2(nor_573_nl, mux_tmp_118, or_311_cse);
  assign and_dcpl_396 = mux_119_nl & and_dcpl_139;
  assign or_332_cse = (result_rem_11cyc_st_3!=4'b0011);
  assign nor_570_nl = ~(and_dcpl_156 | and_dcpl_139);
  assign or_334_nl = (result_rem_11cyc_st_4!=4'b0011) | (~ and_dcpl_130);
  assign mux_tmp_120 = MUX_s_1_2_2(nor_570_nl, or_334_nl, or_332_cse);
  assign nor_571_nl = ~(and_dcpl_182 | (~ mux_tmp_120));
  assign mux_tmp_121 = MUX_s_1_2_2(nor_571_nl, mux_tmp_120, or_323_cse);
  assign nor_572_nl = ~(and_dcpl_208 | (~ mux_tmp_121));
  assign mux_tmp_122 = MUX_s_1_2_2(nor_572_nl, mux_tmp_121, or_316_cse);
  assign nor_569_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_122));
  assign mux_123_nl = MUX_s_1_2_2(nor_569_nl, mux_tmp_122, or_311_cse);
  assign and_dcpl_399 = mux_123_nl & and_dcpl_114;
  assign or_343_cse = (result_rem_11cyc_st_4!=4'b0011);
  assign nor_565_nl = ~(and_dcpl_130 | and_dcpl_114);
  assign or_345_nl = (result_rem_11cyc_st_5!=4'b0011) | (~ and_dcpl_105);
  assign mux_tmp_124 = MUX_s_1_2_2(nor_565_nl, or_345_nl, or_343_cse);
  assign nor_566_nl = ~(and_dcpl_156 | (~ mux_tmp_124));
  assign mux_tmp_125 = MUX_s_1_2_2(nor_566_nl, mux_tmp_124, or_332_cse);
  assign nor_567_nl = ~(and_dcpl_182 | (~ mux_tmp_125));
  assign mux_tmp_126 = MUX_s_1_2_2(nor_567_nl, mux_tmp_125, or_323_cse);
  assign nor_568_nl = ~(and_dcpl_208 | (~ mux_tmp_126));
  assign mux_tmp_127 = MUX_s_1_2_2(nor_568_nl, mux_tmp_126, or_316_cse);
  assign nor_564_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_127));
  assign mux_128_nl = MUX_s_1_2_2(nor_564_nl, mux_tmp_127, or_311_cse);
  assign and_dcpl_402 = mux_128_nl & and_dcpl_88;
  assign or_356_cse = (result_rem_11cyc_st_5!=4'b0011);
  assign nor_559_nl = ~(and_dcpl_105 | and_dcpl_88);
  assign or_358_nl = (result_rem_11cyc_st_6!=4'b0011) | (~ and_dcpl_79);
  assign mux_tmp_129 = MUX_s_1_2_2(nor_559_nl, or_358_nl, or_356_cse);
  assign nor_560_nl = ~(and_dcpl_130 | (~ mux_tmp_129));
  assign mux_tmp_130 = MUX_s_1_2_2(nor_560_nl, mux_tmp_129, or_343_cse);
  assign nor_561_nl = ~(and_dcpl_156 | (~ mux_tmp_130));
  assign mux_tmp_131 = MUX_s_1_2_2(nor_561_nl, mux_tmp_130, or_332_cse);
  assign nor_562_nl = ~(and_dcpl_182 | (~ mux_tmp_131));
  assign mux_tmp_132 = MUX_s_1_2_2(nor_562_nl, mux_tmp_131, or_323_cse);
  assign nor_563_nl = ~(and_dcpl_208 | (~ mux_tmp_132));
  assign mux_tmp_133 = MUX_s_1_2_2(nor_563_nl, mux_tmp_132, or_316_cse);
  assign nor_558_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_133));
  assign mux_134_nl = MUX_s_1_2_2(nor_558_nl, mux_tmp_133, or_311_cse);
  assign and_dcpl_405 = mux_134_nl & and_dcpl_62;
  assign or_371_cse = (result_rem_11cyc_st_6!=4'b0011);
  assign nor_552_nl = ~(and_dcpl_79 | and_dcpl_62);
  assign or_373_nl = (result_rem_11cyc_st_7!=4'b0011) | (~ and_dcpl_53);
  assign mux_tmp_135 = MUX_s_1_2_2(nor_552_nl, or_373_nl, or_371_cse);
  assign nor_553_nl = ~(and_dcpl_105 | (~ mux_tmp_135));
  assign mux_tmp_136 = MUX_s_1_2_2(nor_553_nl, mux_tmp_135, or_356_cse);
  assign nor_554_nl = ~(and_dcpl_130 | (~ mux_tmp_136));
  assign mux_tmp_137 = MUX_s_1_2_2(nor_554_nl, mux_tmp_136, or_343_cse);
  assign nor_555_nl = ~(and_dcpl_156 | (~ mux_tmp_137));
  assign mux_tmp_138 = MUX_s_1_2_2(nor_555_nl, mux_tmp_137, or_332_cse);
  assign nor_556_nl = ~(and_dcpl_182 | (~ mux_tmp_138));
  assign mux_tmp_139 = MUX_s_1_2_2(nor_556_nl, mux_tmp_138, or_323_cse);
  assign nor_557_nl = ~(and_dcpl_208 | (~ mux_tmp_139));
  assign mux_tmp_140 = MUX_s_1_2_2(nor_557_nl, mux_tmp_139, or_316_cse);
  assign nor_551_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_140));
  assign mux_141_nl = MUX_s_1_2_2(nor_551_nl, mux_tmp_140, or_311_cse);
  assign and_dcpl_408 = mux_141_nl & and_dcpl_37;
  assign nor_543_nl = ~(and_dcpl_53 | and_dcpl_37);
  assign or_390_nl = (result_rem_11cyc_st_8!=4'b0011) | (~ and_dcpl_28);
  assign or_388_nl = (result_rem_11cyc_st_7!=4'b0011);
  assign mux_tmp_142 = MUX_s_1_2_2(nor_543_nl, or_390_nl, or_388_nl);
  assign nor_544_nl = ~(and_dcpl_79 | (~ mux_tmp_142));
  assign mux_tmp_143 = MUX_s_1_2_2(nor_544_nl, mux_tmp_142, or_371_cse);
  assign nor_545_nl = ~(and_dcpl_105 | (~ mux_tmp_143));
  assign mux_tmp_144 = MUX_s_1_2_2(nor_545_nl, mux_tmp_143, or_356_cse);
  assign nor_546_nl = ~(and_dcpl_130 | (~ mux_tmp_144));
  assign mux_tmp_145 = MUX_s_1_2_2(nor_546_nl, mux_tmp_144, or_343_cse);
  assign nor_547_nl = ~(and_dcpl_156 | (~ mux_tmp_145));
  assign mux_tmp_146 = MUX_s_1_2_2(nor_547_nl, mux_tmp_145, or_332_cse);
  assign nor_548_nl = ~(and_dcpl_182 | (~ mux_tmp_146));
  assign mux_tmp_147 = MUX_s_1_2_2(nor_548_nl, mux_tmp_146, or_323_cse);
  assign nor_549_nl = ~(and_dcpl_208 | (~ mux_tmp_147));
  assign mux_tmp_148 = MUX_s_1_2_2(nor_549_nl, mux_tmp_147, or_316_cse);
  assign nor_550_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_148));
  assign mux_149_nl = MUX_s_1_2_2(nor_550_nl, mux_tmp_148, or_311_cse);
  assign and_dcpl_411 = mux_149_nl & and_dcpl_4 & and_dcpl_11;
  assign and_tmp_27 = ((~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2!=4'b0011))
      & ((~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3!=4'b0011)) &
      ((~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4!=4'b0011)) & ((~
      main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5!=4'b0011)) & ((~ main_stage_0_7)
      | (~ asn_itm_6) | (result_rem_11cyc_st_6!=4'b0011)) & ((~ main_stage_0_8) |
      (~ asn_itm_7) | (result_rem_11cyc_st_7!=4'b0011)) & ((~ main_stage_0_9) | (~
      asn_itm_8) | (result_rem_11cyc_st_8!=4'b0011)) & ((~ main_stage_0_10) | (~
      asn_itm_9) | (result_rem_11cyc_st_9!=4'b0011));
  assign nor_542_nl = ~(and_dcpl_208 | (~ and_tmp_27));
  assign mux_tmp_150 = MUX_s_1_2_2(nor_542_nl, and_tmp_27, or_316_cse);
  assign and_796_nl = (~((result_result_acc_tmp[1:0]==2'b11) & ccs_ccore_start_rsci_idat))
      & mux_tmp_150;
  assign or_399_nl = (result_result_acc_tmp[3:2]!=2'b00);
  assign mux_tmp_151 = MUX_s_1_2_2(and_796_nl, mux_tmp_150, or_399_nl);
  assign and_dcpl_417 = ccs_ccore_start_rsci_idat & (result_result_acc_tmp[3:2]==2'b01);
  assign and_dcpl_418 = and_dcpl_417 & and_dcpl_260;
  assign or_tmp_402 = (result_rem_11cyc!=4'b0100) | (~ and_dcpl_208);
  assign nand_144_cse = ~((result_result_acc_tmp[2]) & ccs_ccore_start_rsci_idat);
  assign or_413_cse = (result_result_acc_tmp[1]) | (result_result_acc_tmp[0]) | (result_result_acc_tmp[3]);
  assign and_795_nl = nand_144_cse & or_tmp_402;
  assign mux_152_nl = MUX_s_1_2_2(and_795_nl, or_tmp_402, or_413_cse);
  assign and_dcpl_422 = mux_152_nl & and_dcpl_194;
  assign or_418_cse = (result_rem_11cyc!=4'b0100);
  assign nor_541_nl = ~(and_dcpl_208 | and_dcpl_194);
  assign or_420_nl = (result_rem_11cyc_st_2!=4'b0100) | (~ and_dcpl_182);
  assign mux_tmp_153 = MUX_s_1_2_2(nor_541_nl, or_420_nl, or_418_cse);
  assign and_794_nl = nand_144_cse & mux_tmp_153;
  assign mux_154_nl = MUX_s_1_2_2(and_794_nl, mux_tmp_153, or_413_cse);
  assign and_dcpl_426 = mux_154_nl & and_dcpl_168;
  assign or_425_cse = (result_rem_11cyc_st_2!=4'b0100);
  assign nor_539_nl = ~(and_dcpl_182 | and_dcpl_168);
  assign or_427_nl = (result_rem_11cyc_st_3!=4'b0100) | (~ and_dcpl_156);
  assign mux_tmp_155 = MUX_s_1_2_2(nor_539_nl, or_427_nl, or_425_cse);
  assign nor_540_nl = ~(and_dcpl_208 | (~ mux_tmp_155));
  assign mux_tmp_156 = MUX_s_1_2_2(nor_540_nl, mux_tmp_155, or_418_cse);
  assign and_793_nl = nand_144_cse & mux_tmp_156;
  assign mux_157_nl = MUX_s_1_2_2(and_793_nl, mux_tmp_156, or_413_cse);
  assign and_dcpl_430 = mux_157_nl & and_dcpl_142;
  assign or_434_cse = (result_rem_11cyc_st_3!=4'b0100);
  assign nor_536_nl = ~(and_dcpl_156 | and_dcpl_142);
  assign or_436_nl = (result_rem_11cyc_st_4!=4'b0100) | (~ and_dcpl_130);
  assign mux_tmp_158 = MUX_s_1_2_2(nor_536_nl, or_436_nl, or_434_cse);
  assign nor_537_nl = ~(and_dcpl_182 | (~ mux_tmp_158));
  assign mux_tmp_159 = MUX_s_1_2_2(nor_537_nl, mux_tmp_158, or_425_cse);
  assign nor_538_nl = ~(and_dcpl_208 | (~ mux_tmp_159));
  assign mux_tmp_160 = MUX_s_1_2_2(nor_538_nl, mux_tmp_159, or_418_cse);
  assign and_792_nl = nand_144_cse & mux_tmp_160;
  assign mux_161_nl = MUX_s_1_2_2(and_792_nl, mux_tmp_160, or_413_cse);
  assign and_dcpl_433 = mux_161_nl & and_dcpl_116;
  assign or_445_cse = (result_rem_11cyc_st_4!=4'b0100);
  assign nor_532_nl = ~(and_dcpl_130 | and_dcpl_116);
  assign or_447_nl = (result_rem_11cyc_st_5[1]) | (result_rem_11cyc_st_5[0]) | (result_rem_11cyc_st_5[3])
      | (~ and_dcpl_115);
  assign mux_tmp_162 = MUX_s_1_2_2(nor_532_nl, or_447_nl, or_445_cse);
  assign nor_533_nl = ~(and_dcpl_156 | (~ mux_tmp_162));
  assign mux_tmp_163 = MUX_s_1_2_2(nor_533_nl, mux_tmp_162, or_434_cse);
  assign nor_534_nl = ~(and_dcpl_182 | (~ mux_tmp_163));
  assign mux_tmp_164 = MUX_s_1_2_2(nor_534_nl, mux_tmp_163, or_425_cse);
  assign nor_535_nl = ~(and_dcpl_208 | (~ mux_tmp_164));
  assign mux_tmp_165 = MUX_s_1_2_2(nor_535_nl, mux_tmp_164, or_418_cse);
  assign and_791_nl = nand_144_cse & mux_tmp_165;
  assign mux_166_nl = MUX_s_1_2_2(and_791_nl, mux_tmp_165, or_413_cse);
  assign and_dcpl_437 = mux_166_nl & and_dcpl_91;
  assign or_458_cse = (result_rem_11cyc_st_5[1]) | (result_rem_11cyc_st_5[0]) | (result_rem_11cyc_st_5[3]);
  assign and_790_cse = (result_rem_11cyc_st_5[2]) & asn_itm_5 & main_stage_0_6;
  assign nor_527_nl = ~(and_790_cse | and_dcpl_91);
  assign or_460_nl = (result_rem_11cyc_st_6!=4'b0100) | (~ and_dcpl_79);
  assign mux_tmp_167 = MUX_s_1_2_2(nor_527_nl, or_460_nl, or_458_cse);
  assign nor_528_nl = ~(and_dcpl_130 | (~ mux_tmp_167));
  assign mux_tmp_168 = MUX_s_1_2_2(nor_528_nl, mux_tmp_167, or_445_cse);
  assign nor_529_nl = ~(and_dcpl_156 | (~ mux_tmp_168));
  assign mux_tmp_169 = MUX_s_1_2_2(nor_529_nl, mux_tmp_168, or_434_cse);
  assign nor_530_nl = ~(and_dcpl_182 | (~ mux_tmp_169));
  assign mux_tmp_170 = MUX_s_1_2_2(nor_530_nl, mux_tmp_169, or_425_cse);
  assign nor_531_nl = ~(and_dcpl_208 | (~ mux_tmp_170));
  assign mux_tmp_171 = MUX_s_1_2_2(nor_531_nl, mux_tmp_170, or_418_cse);
  assign and_789_nl = nand_144_cse & mux_tmp_171;
  assign mux_172_nl = MUX_s_1_2_2(and_789_nl, mux_tmp_171, or_413_cse);
  assign and_dcpl_441 = mux_172_nl & and_dcpl_65;
  assign or_473_cse = (result_rem_11cyc_st_6!=4'b0100);
  assign nor_522_nl = ~(and_dcpl_79 | and_dcpl_65);
  assign or_475_nl = (result_rem_11cyc_st_7!=4'b0100) | (~ and_dcpl_53);
  assign mux_tmp_173 = MUX_s_1_2_2(nor_522_nl, or_475_nl, or_473_cse);
  assign nand_138_cse = ~((result_rem_11cyc_st_5[2]) & asn_itm_5 & main_stage_0_6);
  assign and_788_nl = nand_138_cse & mux_tmp_173;
  assign mux_tmp_174 = MUX_s_1_2_2(and_788_nl, mux_tmp_173, or_458_cse);
  assign nor_523_nl = ~(and_dcpl_130 | (~ mux_tmp_174));
  assign mux_tmp_175 = MUX_s_1_2_2(nor_523_nl, mux_tmp_174, or_445_cse);
  assign nor_524_nl = ~(and_dcpl_156 | (~ mux_tmp_175));
  assign mux_tmp_176 = MUX_s_1_2_2(nor_524_nl, mux_tmp_175, or_434_cse);
  assign nor_525_nl = ~(and_dcpl_182 | (~ mux_tmp_176));
  assign mux_tmp_177 = MUX_s_1_2_2(nor_525_nl, mux_tmp_176, or_425_cse);
  assign nor_526_nl = ~(and_dcpl_208 | (~ mux_tmp_177));
  assign mux_tmp_178 = MUX_s_1_2_2(nor_526_nl, mux_tmp_177, or_418_cse);
  assign and_787_nl = nand_144_cse & mux_tmp_178;
  assign mux_179_nl = MUX_s_1_2_2(and_787_nl, mux_tmp_178, or_413_cse);
  assign and_dcpl_444 = mux_179_nl & and_dcpl_39;
  assign nor_516_nl = ~(and_dcpl_53 | and_dcpl_39);
  assign or_492_nl = (result_rem_11cyc_st_8[0]) | (result_rem_11cyc_st_8[1]) | (result_rem_11cyc_st_8[3])
      | (~ and_dcpl_38);
  assign or_490_nl = (result_rem_11cyc_st_7!=4'b0100);
  assign mux_tmp_180 = MUX_s_1_2_2(nor_516_nl, or_492_nl, or_490_nl);
  assign nor_517_nl = ~(and_dcpl_79 | (~ mux_tmp_180));
  assign mux_tmp_181 = MUX_s_1_2_2(nor_517_nl, mux_tmp_180, or_473_cse);
  assign and_785_nl = nand_138_cse & mux_tmp_181;
  assign mux_tmp_182 = MUX_s_1_2_2(and_785_nl, mux_tmp_181, or_458_cse);
  assign nor_518_nl = ~(and_dcpl_130 | (~ mux_tmp_182));
  assign mux_tmp_183 = MUX_s_1_2_2(nor_518_nl, mux_tmp_182, or_445_cse);
  assign nor_519_nl = ~(and_dcpl_156 | (~ mux_tmp_183));
  assign mux_tmp_184 = MUX_s_1_2_2(nor_519_nl, mux_tmp_183, or_434_cse);
  assign nor_520_nl = ~(and_dcpl_182 | (~ mux_tmp_184));
  assign mux_tmp_185 = MUX_s_1_2_2(nor_520_nl, mux_tmp_184, or_425_cse);
  assign nor_521_nl = ~(and_dcpl_208 | (~ mux_tmp_185));
  assign mux_tmp_186 = MUX_s_1_2_2(nor_521_nl, mux_tmp_185, or_418_cse);
  assign and_786_nl = nand_144_cse & mux_tmp_186;
  assign mux_187_nl = MUX_s_1_2_2(and_786_nl, mux_tmp_186, or_413_cse);
  assign and_dcpl_447 = mux_187_nl & and_dcpl_13 & and_dcpl_2;
  assign and_tmp_34 = ((~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2!=4'b0100))
      & ((~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3!=4'b0100)) &
      ((~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4!=4'b0100)) & ((~
      main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5!=4'b0100)) & ((~ main_stage_0_7)
      | (~ asn_itm_6) | (result_rem_11cyc_st_6!=4'b0100)) & ((~ main_stage_0_8) |
      (~ asn_itm_7) | (result_rem_11cyc_st_7!=4'b0100)) & ((~ main_stage_0_9) | (~
      asn_itm_8) | (result_rem_11cyc_st_8!=4'b0100)) & ((~ main_stage_0_10) | (~
      asn_itm_9) | (result_rem_11cyc_st_9!=4'b0100));
  assign nor_514_nl = ~(and_dcpl_208 | (~ and_tmp_34));
  assign mux_tmp_188 = MUX_s_1_2_2(nor_514_nl, and_tmp_34, or_418_cse);
  assign nor_515_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_188));
  assign or_501_nl = (result_result_acc_tmp!=4'b0100);
  assign mux_tmp_189 = MUX_s_1_2_2(nor_515_nl, mux_tmp_188, or_501_nl);
  assign and_dcpl_452 = and_dcpl_417 & and_dcpl_318;
  assign or_tmp_502 = (result_rem_11cyc!=4'b0101) | (~ and_dcpl_208);
  assign or_516_cse = (result_result_acc_tmp[1]) | (~ (result_result_acc_tmp[0]))
      | (result_result_acc_tmp[3]);
  assign and_784_nl = nand_144_cse & or_tmp_502;
  assign mux_190_nl = MUX_s_1_2_2(and_784_nl, or_tmp_502, or_516_cse);
  assign and_dcpl_455 = mux_190_nl & and_dcpl_196;
  assign or_521_cse = (result_rem_11cyc!=4'b0101);
  assign nor_513_nl = ~(and_dcpl_208 | and_dcpl_196);
  assign or_523_nl = (result_rem_11cyc_st_2!=4'b0101) | (~ and_dcpl_182);
  assign mux_tmp_191 = MUX_s_1_2_2(nor_513_nl, or_523_nl, or_521_cse);
  assign and_783_nl = nand_144_cse & mux_tmp_191;
  assign mux_192_nl = MUX_s_1_2_2(and_783_nl, mux_tmp_191, or_516_cse);
  assign and_dcpl_458 = mux_192_nl & and_dcpl_170;
  assign or_528_cse = (result_rem_11cyc_st_2!=4'b0101);
  assign nor_511_nl = ~(and_dcpl_182 | and_dcpl_170);
  assign or_530_nl = (result_rem_11cyc_st_3!=4'b0101) | (~ and_dcpl_156);
  assign mux_tmp_193 = MUX_s_1_2_2(nor_511_nl, or_530_nl, or_528_cse);
  assign nor_512_nl = ~(and_dcpl_208 | (~ mux_tmp_193));
  assign mux_tmp_194 = MUX_s_1_2_2(nor_512_nl, mux_tmp_193, or_521_cse);
  assign and_782_nl = nand_144_cse & mux_tmp_194;
  assign mux_195_nl = MUX_s_1_2_2(and_782_nl, mux_tmp_194, or_516_cse);
  assign and_dcpl_462 = mux_195_nl & and_dcpl_145;
  assign or_537_cse = (result_rem_11cyc_st_3!=4'b0101);
  assign nor_508_nl = ~(and_dcpl_156 | and_dcpl_145);
  assign or_539_nl = (result_rem_11cyc_st_4!=4'b0101) | (~ and_dcpl_130);
  assign mux_tmp_196 = MUX_s_1_2_2(nor_508_nl, or_539_nl, or_537_cse);
  assign nor_509_nl = ~(and_dcpl_182 | (~ mux_tmp_196));
  assign mux_tmp_197 = MUX_s_1_2_2(nor_509_nl, mux_tmp_196, or_528_cse);
  assign nor_510_nl = ~(and_dcpl_208 | (~ mux_tmp_197));
  assign mux_tmp_198 = MUX_s_1_2_2(nor_510_nl, mux_tmp_197, or_521_cse);
  assign and_781_nl = nand_144_cse & mux_tmp_198;
  assign mux_199_nl = MUX_s_1_2_2(and_781_nl, mux_tmp_198, or_516_cse);
  assign and_dcpl_464 = mux_199_nl & and_dcpl_117;
  assign or_548_cse = (result_rem_11cyc_st_4!=4'b0101);
  assign nor_504_nl = ~(and_dcpl_130 | and_dcpl_117);
  assign or_550_nl = (result_rem_11cyc_st_5[1]) | (~ (result_rem_11cyc_st_5[0]))
      | (result_rem_11cyc_st_5[3]) | (~ and_dcpl_115);
  assign mux_tmp_200 = MUX_s_1_2_2(nor_504_nl, or_550_nl, or_548_cse);
  assign nor_505_nl = ~(and_dcpl_156 | (~ mux_tmp_200));
  assign mux_tmp_201 = MUX_s_1_2_2(nor_505_nl, mux_tmp_200, or_537_cse);
  assign nor_506_nl = ~(and_dcpl_182 | (~ mux_tmp_201));
  assign mux_tmp_202 = MUX_s_1_2_2(nor_506_nl, mux_tmp_201, or_528_cse);
  assign nor_507_nl = ~(and_dcpl_208 | (~ mux_tmp_202));
  assign mux_tmp_203 = MUX_s_1_2_2(nor_507_nl, mux_tmp_202, or_521_cse);
  assign and_780_nl = nand_144_cse & mux_tmp_203;
  assign mux_204_nl = MUX_s_1_2_2(and_780_nl, mux_tmp_203, or_516_cse);
  assign and_dcpl_468 = mux_204_nl & and_dcpl_94;
  assign or_561_cse = (result_rem_11cyc_st_5[1]) | (~ (result_rem_11cyc_st_5[0]))
      | (result_rem_11cyc_st_5[3]);
  assign nor_499_nl = ~(and_790_cse | and_dcpl_94);
  assign or_563_nl = (result_rem_11cyc_st_6!=4'b0101) | (~ and_dcpl_79);
  assign mux_tmp_205 = MUX_s_1_2_2(nor_499_nl, or_563_nl, or_561_cse);
  assign nor_500_nl = ~(and_dcpl_130 | (~ mux_tmp_205));
  assign mux_tmp_206 = MUX_s_1_2_2(nor_500_nl, mux_tmp_205, or_548_cse);
  assign nor_501_nl = ~(and_dcpl_156 | (~ mux_tmp_206));
  assign mux_tmp_207 = MUX_s_1_2_2(nor_501_nl, mux_tmp_206, or_537_cse);
  assign nor_502_nl = ~(and_dcpl_182 | (~ mux_tmp_207));
  assign mux_tmp_208 = MUX_s_1_2_2(nor_502_nl, mux_tmp_207, or_528_cse);
  assign nor_503_nl = ~(and_dcpl_208 | (~ mux_tmp_208));
  assign mux_tmp_209 = MUX_s_1_2_2(nor_503_nl, mux_tmp_208, or_521_cse);
  assign and_778_nl = nand_144_cse & mux_tmp_209;
  assign mux_210_nl = MUX_s_1_2_2(and_778_nl, mux_tmp_209, or_516_cse);
  assign and_dcpl_472 = mux_210_nl & and_dcpl_68;
  assign or_576_cse = (result_rem_11cyc_st_6!=4'b0101);
  assign nor_494_nl = ~(and_dcpl_79 | and_dcpl_68);
  assign or_578_nl = (result_rem_11cyc_st_7!=4'b0101) | (~ and_dcpl_53);
  assign mux_tmp_211 = MUX_s_1_2_2(nor_494_nl, or_578_nl, or_576_cse);
  assign and_777_nl = nand_138_cse & mux_tmp_211;
  assign mux_tmp_212 = MUX_s_1_2_2(and_777_nl, mux_tmp_211, or_561_cse);
  assign nor_495_nl = ~(and_dcpl_130 | (~ mux_tmp_212));
  assign mux_tmp_213 = MUX_s_1_2_2(nor_495_nl, mux_tmp_212, or_548_cse);
  assign nor_496_nl = ~(and_dcpl_156 | (~ mux_tmp_213));
  assign mux_tmp_214 = MUX_s_1_2_2(nor_496_nl, mux_tmp_213, or_537_cse);
  assign nor_497_nl = ~(and_dcpl_182 | (~ mux_tmp_214));
  assign mux_tmp_215 = MUX_s_1_2_2(nor_497_nl, mux_tmp_214, or_528_cse);
  assign nor_498_nl = ~(and_dcpl_208 | (~ mux_tmp_215));
  assign mux_tmp_216 = MUX_s_1_2_2(nor_498_nl, mux_tmp_215, or_521_cse);
  assign and_776_nl = nand_144_cse & mux_tmp_216;
  assign mux_217_nl = MUX_s_1_2_2(and_776_nl, mux_tmp_216, or_516_cse);
  assign and_dcpl_474 = mux_217_nl & and_dcpl_40;
  assign nor_488_nl = ~(and_dcpl_53 | and_dcpl_40);
  assign or_595_nl = (~ (result_rem_11cyc_st_8[0])) | (result_rem_11cyc_st_8[1])
      | (result_rem_11cyc_st_8[3]) | (~ and_dcpl_38);
  assign or_593_nl = (result_rem_11cyc_st_7!=4'b0101);
  assign mux_tmp_218 = MUX_s_1_2_2(nor_488_nl, or_595_nl, or_593_nl);
  assign nor_489_nl = ~(and_dcpl_79 | (~ mux_tmp_218));
  assign mux_tmp_219 = MUX_s_1_2_2(nor_489_nl, mux_tmp_218, or_576_cse);
  assign and_774_nl = nand_138_cse & mux_tmp_219;
  assign mux_tmp_220 = MUX_s_1_2_2(and_774_nl, mux_tmp_219, or_561_cse);
  assign nor_490_nl = ~(and_dcpl_130 | (~ mux_tmp_220));
  assign mux_tmp_221 = MUX_s_1_2_2(nor_490_nl, mux_tmp_220, or_548_cse);
  assign nor_491_nl = ~(and_dcpl_156 | (~ mux_tmp_221));
  assign mux_tmp_222 = MUX_s_1_2_2(nor_491_nl, mux_tmp_221, or_537_cse);
  assign nor_492_nl = ~(and_dcpl_182 | (~ mux_tmp_222));
  assign mux_tmp_223 = MUX_s_1_2_2(nor_492_nl, mux_tmp_222, or_528_cse);
  assign nor_493_nl = ~(and_dcpl_208 | (~ mux_tmp_223));
  assign mux_tmp_224 = MUX_s_1_2_2(nor_493_nl, mux_tmp_223, or_521_cse);
  assign and_775_nl = nand_144_cse & mux_tmp_224;
  assign mux_225_nl = MUX_s_1_2_2(and_775_nl, mux_tmp_224, or_516_cse);
  assign and_dcpl_476 = mux_225_nl & and_dcpl_13 & and_dcpl_6;
  assign and_tmp_41 = ((~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2!=4'b0101))
      & ((~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3!=4'b0101)) &
      ((~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4!=4'b0101)) & ((~
      main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5!=4'b0101)) & ((~ main_stage_0_7)
      | (~ asn_itm_6) | (result_rem_11cyc_st_6!=4'b0101)) & ((~ main_stage_0_8) |
      (~ asn_itm_7) | (result_rem_11cyc_st_7!=4'b0101)) & ((~ main_stage_0_9) | (~
      asn_itm_8) | (result_rem_11cyc_st_8!=4'b0101)) & ((~ main_stage_0_10) | (~
      asn_itm_9) | (result_rem_11cyc_st_9!=4'b0101));
  assign nor_487_nl = ~(and_dcpl_208 | (~ and_tmp_41));
  assign mux_tmp_226 = MUX_s_1_2_2(nor_487_nl, and_tmp_41, or_521_cse);
  assign and_773_nl = nand_146_cse & mux_tmp_226;
  assign or_604_nl = (result_result_acc_tmp[3:1]!=3'b010);
  assign mux_tmp_227 = MUX_s_1_2_2(and_773_nl, mux_tmp_226, or_604_nl);
  assign and_dcpl_480 = and_dcpl_417 & and_dcpl_352;
  assign or_tmp_602 = (result_rem_11cyc!=4'b0110) | (~ and_dcpl_208);
  assign or_617_cse = (~ (result_result_acc_tmp[1])) | (result_result_acc_tmp[0])
      | (result_result_acc_tmp[3]);
  assign and_772_nl = nand_144_cse & or_tmp_602;
  assign mux_228_nl = MUX_s_1_2_2(and_772_nl, or_tmp_602, or_617_cse);
  assign and_dcpl_484 = mux_228_nl & and_dcpl_199;
  assign or_622_cse = (result_rem_11cyc!=4'b0110);
  assign nor_486_nl = ~(and_dcpl_208 | and_dcpl_199);
  assign or_624_nl = (result_rem_11cyc_st_2!=4'b0110) | (~ and_dcpl_182);
  assign mux_tmp_229 = MUX_s_1_2_2(nor_486_nl, or_624_nl, or_622_cse);
  assign and_771_nl = nand_144_cse & mux_tmp_229;
  assign mux_230_nl = MUX_s_1_2_2(and_771_nl, mux_tmp_229, or_617_cse);
  assign and_dcpl_488 = mux_230_nl & and_dcpl_173;
  assign or_629_cse = (result_rem_11cyc_st_2!=4'b0110);
  assign nor_484_nl = ~(and_dcpl_182 | and_dcpl_173);
  assign or_631_nl = (result_rem_11cyc_st_3!=4'b0110) | (~ and_dcpl_156);
  assign mux_tmp_231 = MUX_s_1_2_2(nor_484_nl, or_631_nl, or_629_cse);
  assign nor_485_nl = ~(and_dcpl_208 | (~ mux_tmp_231));
  assign mux_tmp_232 = MUX_s_1_2_2(nor_485_nl, mux_tmp_231, or_622_cse);
  assign and_770_nl = nand_144_cse & mux_tmp_232;
  assign mux_233_nl = MUX_s_1_2_2(and_770_nl, mux_tmp_232, or_617_cse);
  assign and_dcpl_491 = mux_233_nl & and_dcpl_147;
  assign or_638_cse = (result_rem_11cyc_st_3!=4'b0110);
  assign nor_481_nl = ~(and_dcpl_156 | and_dcpl_147);
  assign or_640_nl = (result_rem_11cyc_st_4!=4'b0110) | (~ and_dcpl_130);
  assign mux_tmp_234 = MUX_s_1_2_2(nor_481_nl, or_640_nl, or_638_cse);
  assign nor_482_nl = ~(and_dcpl_182 | (~ mux_tmp_234));
  assign mux_tmp_235 = MUX_s_1_2_2(nor_482_nl, mux_tmp_234, or_629_cse);
  assign nor_483_nl = ~(and_dcpl_208 | (~ mux_tmp_235));
  assign mux_tmp_236 = MUX_s_1_2_2(nor_483_nl, mux_tmp_235, or_622_cse);
  assign and_769_nl = nand_144_cse & mux_tmp_236;
  assign mux_237_nl = MUX_s_1_2_2(and_769_nl, mux_tmp_236, or_617_cse);
  assign and_dcpl_493 = mux_237_nl & and_dcpl_118;
  assign or_649_cse = (result_rem_11cyc_st_4!=4'b0110);
  assign nor_477_nl = ~(and_dcpl_130 | and_dcpl_118);
  assign or_651_nl = (~ (result_rem_11cyc_st_5[1])) | (result_rem_11cyc_st_5[0])
      | (result_rem_11cyc_st_5[3]) | (~ and_dcpl_115);
  assign mux_tmp_238 = MUX_s_1_2_2(nor_477_nl, or_651_nl, or_649_cse);
  assign nor_478_nl = ~(and_dcpl_156 | (~ mux_tmp_238));
  assign mux_tmp_239 = MUX_s_1_2_2(nor_478_nl, mux_tmp_238, or_638_cse);
  assign nor_479_nl = ~(and_dcpl_182 | (~ mux_tmp_239));
  assign mux_tmp_240 = MUX_s_1_2_2(nor_479_nl, mux_tmp_239, or_629_cse);
  assign nor_480_nl = ~(and_dcpl_208 | (~ mux_tmp_240));
  assign mux_tmp_241 = MUX_s_1_2_2(nor_480_nl, mux_tmp_240, or_622_cse);
  assign and_768_nl = nand_144_cse & mux_tmp_241;
  assign mux_242_nl = MUX_s_1_2_2(and_768_nl, mux_tmp_241, or_617_cse);
  assign and_dcpl_496 = mux_242_nl & and_dcpl_96;
  assign or_662_cse = (~ (result_rem_11cyc_st_5[1])) | (result_rem_11cyc_st_5[0])
      | (result_rem_11cyc_st_5[3]);
  assign nor_472_nl = ~(and_790_cse | and_dcpl_96);
  assign or_664_nl = (result_rem_11cyc_st_6!=4'b0110) | (~ and_dcpl_79);
  assign mux_tmp_243 = MUX_s_1_2_2(nor_472_nl, or_664_nl, or_662_cse);
  assign nor_473_nl = ~(and_dcpl_130 | (~ mux_tmp_243));
  assign mux_tmp_244 = MUX_s_1_2_2(nor_473_nl, mux_tmp_243, or_649_cse);
  assign nor_474_nl = ~(and_dcpl_156 | (~ mux_tmp_244));
  assign mux_tmp_245 = MUX_s_1_2_2(nor_474_nl, mux_tmp_244, or_638_cse);
  assign nor_475_nl = ~(and_dcpl_182 | (~ mux_tmp_245));
  assign mux_tmp_246 = MUX_s_1_2_2(nor_475_nl, mux_tmp_245, or_629_cse);
  assign nor_476_nl = ~(and_dcpl_208 | (~ mux_tmp_246));
  assign mux_tmp_247 = MUX_s_1_2_2(nor_476_nl, mux_tmp_246, or_622_cse);
  assign and_766_nl = nand_144_cse & mux_tmp_247;
  assign mux_248_nl = MUX_s_1_2_2(and_766_nl, mux_tmp_247, or_617_cse);
  assign and_dcpl_499 = mux_248_nl & and_dcpl_70;
  assign or_677_cse = (result_rem_11cyc_st_6!=4'b0110);
  assign nor_467_nl = ~(and_dcpl_79 | and_dcpl_70);
  assign or_679_nl = (result_rem_11cyc_st_7!=4'b0110) | (~ and_dcpl_53);
  assign mux_tmp_249 = MUX_s_1_2_2(nor_467_nl, or_679_nl, or_677_cse);
  assign and_765_nl = nand_138_cse & mux_tmp_249;
  assign mux_tmp_250 = MUX_s_1_2_2(and_765_nl, mux_tmp_249, or_662_cse);
  assign nor_468_nl = ~(and_dcpl_130 | (~ mux_tmp_250));
  assign mux_tmp_251 = MUX_s_1_2_2(nor_468_nl, mux_tmp_250, or_649_cse);
  assign nor_469_nl = ~(and_dcpl_156 | (~ mux_tmp_251));
  assign mux_tmp_252 = MUX_s_1_2_2(nor_469_nl, mux_tmp_251, or_638_cse);
  assign nor_470_nl = ~(and_dcpl_182 | (~ mux_tmp_252));
  assign mux_tmp_253 = MUX_s_1_2_2(nor_470_nl, mux_tmp_252, or_629_cse);
  assign nor_471_nl = ~(and_dcpl_208 | (~ mux_tmp_253));
  assign mux_tmp_254 = MUX_s_1_2_2(nor_471_nl, mux_tmp_253, or_622_cse);
  assign and_764_nl = nand_144_cse & mux_tmp_254;
  assign mux_255_nl = MUX_s_1_2_2(and_764_nl, mux_tmp_254, or_617_cse);
  assign and_dcpl_501 = mux_255_nl & and_dcpl_41;
  assign nor_461_nl = ~(and_dcpl_53 | and_dcpl_41);
  assign or_696_nl = (result_rem_11cyc_st_8[0]) | (~ (result_rem_11cyc_st_8[1]))
      | (result_rem_11cyc_st_8[3]) | (~ and_dcpl_38);
  assign or_694_nl = (result_rem_11cyc_st_7!=4'b0110);
  assign mux_tmp_256 = MUX_s_1_2_2(nor_461_nl, or_696_nl, or_694_nl);
  assign nor_462_nl = ~(and_dcpl_79 | (~ mux_tmp_256));
  assign mux_tmp_257 = MUX_s_1_2_2(nor_462_nl, mux_tmp_256, or_677_cse);
  assign and_762_nl = nand_138_cse & mux_tmp_257;
  assign mux_tmp_258 = MUX_s_1_2_2(and_762_nl, mux_tmp_257, or_662_cse);
  assign nor_463_nl = ~(and_dcpl_130 | (~ mux_tmp_258));
  assign mux_tmp_259 = MUX_s_1_2_2(nor_463_nl, mux_tmp_258, or_649_cse);
  assign nor_464_nl = ~(and_dcpl_156 | (~ mux_tmp_259));
  assign mux_tmp_260 = MUX_s_1_2_2(nor_464_nl, mux_tmp_259, or_638_cse);
  assign nor_465_nl = ~(and_dcpl_182 | (~ mux_tmp_260));
  assign mux_tmp_261 = MUX_s_1_2_2(nor_465_nl, mux_tmp_260, or_629_cse);
  assign nor_466_nl = ~(and_dcpl_208 | (~ mux_tmp_261));
  assign mux_tmp_262 = MUX_s_1_2_2(nor_466_nl, mux_tmp_261, or_622_cse);
  assign and_763_nl = nand_144_cse & mux_tmp_262;
  assign mux_263_nl = MUX_s_1_2_2(and_763_nl, mux_tmp_262, or_617_cse);
  assign and_dcpl_503 = mux_263_nl & and_dcpl_13 & and_dcpl_9;
  assign and_tmp_48 = ((~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2!=4'b0110))
      & ((~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3!=4'b0110)) &
      ((~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4!=4'b0110)) & ((~
      main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5!=4'b0110)) & ((~ main_stage_0_7)
      | (~ asn_itm_6) | (result_rem_11cyc_st_6!=4'b0110)) & ((~ main_stage_0_8) |
      (~ asn_itm_7) | (result_rem_11cyc_st_7!=4'b0110)) & ((~ main_stage_0_9) | (~
      asn_itm_8) | (result_rem_11cyc_st_8!=4'b0110)) & ((~ main_stage_0_10) | (~
      asn_itm_9) | (result_rem_11cyc_st_9!=4'b0110));
  assign nor_459_nl = ~(and_dcpl_208 | (~ and_tmp_48));
  assign mux_tmp_264 = MUX_s_1_2_2(nor_459_nl, and_tmp_48, or_622_cse);
  assign nor_460_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_264));
  assign or_705_nl = (result_result_acc_tmp!=4'b0110);
  assign mux_tmp_265 = MUX_s_1_2_2(nor_460_nl, mux_tmp_264, or_705_nl);
  assign and_dcpl_507 = and_dcpl_417 & and_dcpl_386;
  assign or_tmp_702 = ~((result_rem_11cyc==4'b0111) & and_dcpl_208);
  assign or_718_cse = (~ (result_result_acc_tmp[1])) | (~ (result_result_acc_tmp[0]))
      | (result_result_acc_tmp[3]);
  assign and_761_nl = nand_144_cse & or_tmp_702;
  assign mux_266_nl = MUX_s_1_2_2(and_761_nl, or_tmp_702, or_718_cse);
  assign and_dcpl_510 = mux_266_nl & and_dcpl_201;
  assign nand_112_cse = ~((result_rem_11cyc==4'b0111));
  assign nor_458_nl = ~(and_dcpl_208 | and_dcpl_201);
  assign nand_153_nl = ~((result_rem_11cyc_st_2==4'b0111) & and_dcpl_182);
  assign mux_tmp_267 = MUX_s_1_2_2(nor_458_nl, nand_153_nl, nand_112_cse);
  assign and_760_nl = nand_144_cse & mux_tmp_267;
  assign mux_268_nl = MUX_s_1_2_2(and_760_nl, mux_tmp_267, or_718_cse);
  assign and_dcpl_513 = mux_268_nl & and_dcpl_175;
  assign nand_108_cse = ~((result_rem_11cyc_st_2==4'b0111));
  assign nor_456_nl = ~(and_dcpl_182 | and_dcpl_175);
  assign nand_152_nl = ~((result_rem_11cyc_st_3==4'b0111) & and_dcpl_156);
  assign mux_tmp_269 = MUX_s_1_2_2(nor_456_nl, nand_152_nl, nand_108_cse);
  assign nor_457_nl = ~(and_dcpl_208 | (~ mux_tmp_269));
  assign mux_tmp_270 = MUX_s_1_2_2(nor_457_nl, mux_tmp_269, nand_112_cse);
  assign and_759_nl = nand_144_cse & mux_tmp_270;
  assign mux_271_nl = MUX_s_1_2_2(and_759_nl, mux_tmp_270, or_718_cse);
  assign and_dcpl_516 = mux_271_nl & and_dcpl_149;
  assign nand_103_cse = ~((result_rem_11cyc_st_3==4'b0111));
  assign nor_453_nl = ~(and_dcpl_156 | and_dcpl_149);
  assign nand_151_nl = ~((result_rem_11cyc_st_4==4'b0111) & and_dcpl_130);
  assign mux_tmp_272 = MUX_s_1_2_2(nor_453_nl, nand_151_nl, nand_103_cse);
  assign nor_454_nl = ~(and_dcpl_182 | (~ mux_tmp_272));
  assign mux_tmp_273 = MUX_s_1_2_2(nor_454_nl, mux_tmp_272, nand_108_cse);
  assign nor_455_nl = ~(and_dcpl_208 | (~ mux_tmp_273));
  assign mux_tmp_274 = MUX_s_1_2_2(nor_455_nl, mux_tmp_273, nand_112_cse);
  assign and_758_nl = nand_144_cse & mux_tmp_274;
  assign mux_275_nl = MUX_s_1_2_2(and_758_nl, mux_tmp_274, or_718_cse);
  assign and_dcpl_518 = mux_275_nl & and_dcpl_119;
  assign nand_97_cse = ~((result_rem_11cyc_st_4==4'b0111));
  assign nor_449_nl = ~(and_dcpl_130 | and_dcpl_119);
  assign nand_96_nl = ~((result_rem_11cyc_st_5[1]) & (result_rem_11cyc_st_5[0]) &
      (~ (result_rem_11cyc_st_5[3])) & and_dcpl_115);
  assign mux_tmp_276 = MUX_s_1_2_2(nor_449_nl, nand_96_nl, nand_97_cse);
  assign nor_450_nl = ~(and_dcpl_156 | (~ mux_tmp_276));
  assign mux_tmp_277 = MUX_s_1_2_2(nor_450_nl, mux_tmp_276, nand_103_cse);
  assign nor_451_nl = ~(and_dcpl_182 | (~ mux_tmp_277));
  assign mux_tmp_278 = MUX_s_1_2_2(nor_451_nl, mux_tmp_277, nand_108_cse);
  assign nor_452_nl = ~(and_dcpl_208 | (~ mux_tmp_278));
  assign mux_tmp_279 = MUX_s_1_2_2(nor_452_nl, mux_tmp_278, nand_112_cse);
  assign and_757_nl = nand_144_cse & mux_tmp_279;
  assign mux_280_nl = MUX_s_1_2_2(and_757_nl, mux_tmp_279, or_718_cse);
  assign and_dcpl_521 = mux_280_nl & and_dcpl_98;
  assign or_763_cse = (~ (result_rem_11cyc_st_5[1])) | (~ (result_rem_11cyc_st_5[0]))
      | (result_rem_11cyc_st_5[3]);
  assign nor_444_nl = ~(and_790_cse | and_dcpl_98);
  assign nand_150_nl = ~((result_rem_11cyc_st_6==4'b0111) & and_dcpl_79);
  assign mux_tmp_281 = MUX_s_1_2_2(nor_444_nl, nand_150_nl, or_763_cse);
  assign nor_445_nl = ~(and_dcpl_130 | (~ mux_tmp_281));
  assign mux_tmp_282 = MUX_s_1_2_2(nor_445_nl, mux_tmp_281, nand_97_cse);
  assign nor_446_nl = ~(and_dcpl_156 | (~ mux_tmp_282));
  assign mux_tmp_283 = MUX_s_1_2_2(nor_446_nl, mux_tmp_282, nand_103_cse);
  assign nor_447_nl = ~(and_dcpl_182 | (~ mux_tmp_283));
  assign mux_tmp_284 = MUX_s_1_2_2(nor_447_nl, mux_tmp_283, nand_108_cse);
  assign nor_448_nl = ~(and_dcpl_208 | (~ mux_tmp_284));
  assign mux_tmp_285 = MUX_s_1_2_2(nor_448_nl, mux_tmp_284, nand_112_cse);
  assign and_755_nl = nand_144_cse & mux_tmp_285;
  assign mux_286_nl = MUX_s_1_2_2(and_755_nl, mux_tmp_285, or_718_cse);
  assign and_dcpl_524 = mux_286_nl & and_dcpl_72;
  assign nand_83_cse = ~((result_rem_11cyc_st_6==4'b0111));
  assign nor_439_nl = ~(and_dcpl_79 | and_dcpl_72);
  assign nand_149_nl = ~((result_rem_11cyc_st_7==4'b0111) & and_dcpl_53);
  assign mux_tmp_287 = MUX_s_1_2_2(nor_439_nl, nand_149_nl, nand_83_cse);
  assign and_754_nl = nand_138_cse & mux_tmp_287;
  assign mux_tmp_288 = MUX_s_1_2_2(and_754_nl, mux_tmp_287, or_763_cse);
  assign nor_440_nl = ~(and_dcpl_130 | (~ mux_tmp_288));
  assign mux_tmp_289 = MUX_s_1_2_2(nor_440_nl, mux_tmp_288, nand_97_cse);
  assign nor_441_nl = ~(and_dcpl_156 | (~ mux_tmp_289));
  assign mux_tmp_290 = MUX_s_1_2_2(nor_441_nl, mux_tmp_289, nand_103_cse);
  assign nor_442_nl = ~(and_dcpl_182 | (~ mux_tmp_290));
  assign mux_tmp_291 = MUX_s_1_2_2(nor_442_nl, mux_tmp_290, nand_108_cse);
  assign nor_443_nl = ~(and_dcpl_208 | (~ mux_tmp_291));
  assign mux_tmp_292 = MUX_s_1_2_2(nor_443_nl, mux_tmp_291, nand_112_cse);
  assign and_753_nl = nand_144_cse & mux_tmp_292;
  assign mux_293_nl = MUX_s_1_2_2(and_753_nl, mux_tmp_292, or_718_cse);
  assign and_dcpl_526 = mux_293_nl & and_dcpl_42;
  assign nor_433_nl = ~(and_dcpl_53 | and_dcpl_42);
  assign nand_72_nl = ~((result_rem_11cyc_st_8[0]) & (result_rem_11cyc_st_8[1]) &
      (~ (result_rem_11cyc_st_8[3])) & and_dcpl_38);
  assign nand_73_nl = ~((result_rem_11cyc_st_7==4'b0111));
  assign mux_tmp_294 = MUX_s_1_2_2(nor_433_nl, nand_72_nl, nand_73_nl);
  assign nor_434_nl = ~(and_dcpl_79 | (~ mux_tmp_294));
  assign mux_tmp_295 = MUX_s_1_2_2(nor_434_nl, mux_tmp_294, nand_83_cse);
  assign and_751_nl = nand_138_cse & mux_tmp_295;
  assign mux_tmp_296 = MUX_s_1_2_2(and_751_nl, mux_tmp_295, or_763_cse);
  assign nor_435_nl = ~(and_dcpl_130 | (~ mux_tmp_296));
  assign mux_tmp_297 = MUX_s_1_2_2(nor_435_nl, mux_tmp_296, nand_97_cse);
  assign nor_436_nl = ~(and_dcpl_156 | (~ mux_tmp_297));
  assign mux_tmp_298 = MUX_s_1_2_2(nor_436_nl, mux_tmp_297, nand_103_cse);
  assign nor_437_nl = ~(and_dcpl_182 | (~ mux_tmp_298));
  assign mux_tmp_299 = MUX_s_1_2_2(nor_437_nl, mux_tmp_298, nand_108_cse);
  assign nor_438_nl = ~(and_dcpl_208 | (~ mux_tmp_299));
  assign mux_tmp_300 = MUX_s_1_2_2(nor_438_nl, mux_tmp_299, nand_112_cse);
  assign and_752_nl = nand_144_cse & mux_tmp_300;
  assign mux_301_nl = MUX_s_1_2_2(and_752_nl, mux_tmp_300, or_718_cse);
  assign and_dcpl_528 = mux_301_nl & and_dcpl_13 & and_dcpl_11;
  assign and_tmp_55 = (~(main_stage_0_3 & asn_itm_2 & (result_rem_11cyc_st_2==4'b0111)))
      & (~(main_stage_0_4 & asn_itm_3 & (result_rem_11cyc_st_3==4'b0111))) & (~(main_stage_0_5
      & asn_itm_4 & (result_rem_11cyc_st_4==4'b0111))) & (~(main_stage_0_6 & asn_itm_5
      & (result_rem_11cyc_st_5==4'b0111))) & (~(main_stage_0_7 & asn_itm_6 & (result_rem_11cyc_st_6==4'b0111)))
      & (~(main_stage_0_8 & asn_itm_7 & (result_rem_11cyc_st_7==4'b0111))) & (~(main_stage_0_9
      & asn_itm_8 & (result_rem_11cyc_st_8==4'b0111))) & (~(main_stage_0_10 & asn_itm_9
      & (result_rem_11cyc_st_9==4'b0111)));
  assign nor_432_nl = ~(and_dcpl_208 | (~ and_tmp_55));
  assign mux_tmp_302 = MUX_s_1_2_2(nor_432_nl, and_tmp_55, nand_112_cse);
  assign and_750_nl = (~((result_result_acc_tmp[2:0]==3'b111) & ccs_ccore_start_rsci_idat))
      & mux_tmp_302;
  assign mux_tmp_303 = MUX_s_1_2_2(and_750_nl, mux_tmp_302, result_result_acc_tmp[3]);
  assign and_dcpl_532 = and_dcpl_261 & (result_result_acc_tmp[3]);
  assign and_dcpl_533 = and_dcpl_532 & and_dcpl_260;
  assign not_tmp_645 = ~((result_rem_11cyc[3]) & asn_itm_1 & main_stage_0_2);
  assign or_tmp_801 = (result_rem_11cyc[2:0]!=3'b000) | not_tmp_645;
  assign or_818_cse = (result_result_acc_tmp!=4'b1000);
  assign nor_431_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_801));
  assign mux_304_nl = MUX_s_1_2_2(nor_431_nl, or_tmp_801, or_818_cse);
  assign and_dcpl_536 = mux_304_nl & and_dcpl_203;
  assign or_823_cse = (result_rem_11cyc[2:0]!=3'b000);
  assign and_749_cse = (result_rem_11cyc[3]) & asn_itm_1 & main_stage_0_2;
  assign nor_430_nl = ~(and_749_cse | and_dcpl_203);
  assign or_825_nl = (result_rem_11cyc_st_2[2:0]!=3'b000) | (~ and_dcpl_202);
  assign mux_tmp_305 = MUX_s_1_2_2(nor_430_nl, or_825_nl, or_823_cse);
  assign nor_429_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_305));
  assign mux_306_nl = MUX_s_1_2_2(nor_429_nl, mux_tmp_305, or_818_cse);
  assign and_dcpl_539 = mux_306_nl & and_dcpl_177;
  assign or_830_cse = (result_rem_11cyc_st_2[2:0]!=3'b000);
  assign and_747_cse = (result_rem_11cyc_st_2[3]) & asn_itm_2 & main_stage_0_3;
  assign nor_428_nl = ~(and_747_cse | and_dcpl_177);
  assign or_832_nl = (result_rem_11cyc_st_3[2:0]!=3'b000) | (~ and_dcpl_176);
  assign mux_tmp_307 = MUX_s_1_2_2(nor_428_nl, or_832_nl, or_830_cse);
  assign and_748_nl = not_tmp_645 & mux_tmp_307;
  assign mux_tmp_308 = MUX_s_1_2_2(and_748_nl, mux_tmp_307, or_823_cse);
  assign nor_427_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_308));
  assign mux_309_nl = MUX_s_1_2_2(nor_427_nl, mux_tmp_308, or_818_cse);
  assign and_dcpl_542 = mux_309_nl & and_dcpl_151;
  assign or_839_cse = (result_rem_11cyc_st_3[2:0]!=3'b000);
  assign and_744_cse = (result_rem_11cyc_st_3[3]) & asn_itm_3 & main_stage_0_4;
  assign nor_426_nl = ~(and_744_cse | and_dcpl_151);
  assign or_841_nl = (result_rem_11cyc_st_4[2:0]!=3'b000) | (~ and_dcpl_150);
  assign mux_tmp_310 = MUX_s_1_2_2(nor_426_nl, or_841_nl, or_839_cse);
  assign nand_58_cse = ~((result_rem_11cyc_st_2[3]) & asn_itm_2 & main_stage_0_3);
  assign and_745_nl = nand_58_cse & mux_tmp_310;
  assign mux_tmp_311 = MUX_s_1_2_2(and_745_nl, mux_tmp_310, or_830_cse);
  assign and_746_nl = not_tmp_645 & mux_tmp_311;
  assign mux_tmp_312 = MUX_s_1_2_2(and_746_nl, mux_tmp_311, or_823_cse);
  assign nor_425_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_312));
  assign mux_313_nl = MUX_s_1_2_2(nor_425_nl, mux_tmp_312, or_818_cse);
  assign and_dcpl_546 = mux_313_nl & and_dcpl_122;
  assign or_850_cse = (result_rem_11cyc_st_4[2:0]!=3'b000);
  assign and_740_cse = (result_rem_11cyc_st_4[3]) & asn_itm_4 & main_stage_0_5;
  assign nor_424_nl = ~(and_740_cse | and_dcpl_122);
  assign or_852_nl = (result_rem_11cyc_st_5!=4'b1000) | (~ and_dcpl_105);
  assign mux_tmp_314 = MUX_s_1_2_2(nor_424_nl, or_852_nl, or_850_cse);
  assign nand_55_cse = ~((result_rem_11cyc_st_3[3]) & asn_itm_3 & main_stage_0_4);
  assign and_741_nl = nand_55_cse & mux_tmp_314;
  assign mux_tmp_315 = MUX_s_1_2_2(and_741_nl, mux_tmp_314, or_839_cse);
  assign and_742_nl = nand_58_cse & mux_tmp_315;
  assign mux_tmp_316 = MUX_s_1_2_2(and_742_nl, mux_tmp_315, or_830_cse);
  assign and_743_nl = not_tmp_645 & mux_tmp_316;
  assign mux_tmp_317 = MUX_s_1_2_2(and_743_nl, mux_tmp_316, or_823_cse);
  assign nor_423_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_317));
  assign mux_318_nl = MUX_s_1_2_2(nor_423_nl, mux_tmp_317, or_818_cse);
  assign and_dcpl_549 = mux_318_nl & and_dcpl_100;
  assign or_863_cse = (result_rem_11cyc_st_5!=4'b1000);
  assign nor_422_nl = ~(and_dcpl_105 | and_dcpl_100);
  assign or_865_nl = (result_rem_11cyc_st_6[2:0]!=3'b000) | (~ and_dcpl_99);
  assign mux_tmp_319 = MUX_s_1_2_2(nor_422_nl, or_865_nl, or_863_cse);
  assign nand_51_cse = ~((result_rem_11cyc_st_4[3]) & asn_itm_4 & main_stage_0_5);
  assign and_736_nl = nand_51_cse & mux_tmp_319;
  assign mux_tmp_320 = MUX_s_1_2_2(and_736_nl, mux_tmp_319, or_850_cse);
  assign and_737_nl = nand_55_cse & mux_tmp_320;
  assign mux_tmp_321 = MUX_s_1_2_2(and_737_nl, mux_tmp_320, or_839_cse);
  assign and_738_nl = nand_58_cse & mux_tmp_321;
  assign mux_tmp_322 = MUX_s_1_2_2(and_738_nl, mux_tmp_321, or_830_cse);
  assign and_739_nl = not_tmp_645 & mux_tmp_322;
  assign mux_tmp_323 = MUX_s_1_2_2(and_739_nl, mux_tmp_322, or_823_cse);
  assign nor_421_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_323));
  assign mux_324_nl = MUX_s_1_2_2(nor_421_nl, mux_tmp_323, or_818_cse);
  assign and_dcpl_552 = mux_324_nl & and_dcpl_74;
  assign or_878_cse = (result_rem_11cyc_st_6[2:0]!=3'b000);
  assign and_731_cse = (result_rem_11cyc_st_6[3]) & asn_itm_6 & main_stage_0_7;
  assign nor_419_nl = ~(and_731_cse | and_dcpl_74);
  assign or_880_nl = (result_rem_11cyc_st_7[2:0]!=3'b000) | (~ and_dcpl_73);
  assign mux_tmp_325 = MUX_s_1_2_2(nor_419_nl, or_880_nl, or_878_cse);
  assign nor_420_nl = ~(and_dcpl_105 | (~ mux_tmp_325));
  assign mux_tmp_326 = MUX_s_1_2_2(nor_420_nl, mux_tmp_325, or_863_cse);
  assign and_732_nl = nand_51_cse & mux_tmp_326;
  assign mux_tmp_327 = MUX_s_1_2_2(and_732_nl, mux_tmp_326, or_850_cse);
  assign and_733_nl = nand_55_cse & mux_tmp_327;
  assign mux_tmp_328 = MUX_s_1_2_2(and_733_nl, mux_tmp_327, or_839_cse);
  assign and_734_nl = nand_58_cse & mux_tmp_328;
  assign mux_tmp_329 = MUX_s_1_2_2(and_734_nl, mux_tmp_328, or_830_cse);
  assign and_735_nl = not_tmp_645 & mux_tmp_329;
  assign mux_tmp_330 = MUX_s_1_2_2(and_735_nl, mux_tmp_329, or_823_cse);
  assign nor_418_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_330));
  assign mux_331_nl = MUX_s_1_2_2(nor_418_nl, mux_tmp_330, or_818_cse);
  assign and_dcpl_556 = mux_331_nl & and_dcpl_45;
  assign and_725_cse = (result_rem_11cyc_st_7[3]) & asn_itm_7 & main_stage_0_8;
  assign nor_415_nl = ~(and_725_cse | and_dcpl_45);
  assign or_897_nl = (result_rem_11cyc_st_8!=4'b1000) | (~ and_dcpl_28);
  assign or_895_nl = (result_rem_11cyc_st_7[2:0]!=3'b000);
  assign mux_tmp_332 = MUX_s_1_2_2(nor_415_nl, or_897_nl, or_895_nl);
  assign nand_42_cse = ~((result_rem_11cyc_st_6[3]) & asn_itm_6 & main_stage_0_7);
  assign and_726_nl = nand_42_cse & mux_tmp_332;
  assign mux_tmp_333 = MUX_s_1_2_2(and_726_nl, mux_tmp_332, or_878_cse);
  assign nor_416_nl = ~(and_dcpl_105 | (~ mux_tmp_333));
  assign mux_tmp_334 = MUX_s_1_2_2(nor_416_nl, mux_tmp_333, or_863_cse);
  assign and_727_nl = nand_51_cse & mux_tmp_334;
  assign mux_tmp_335 = MUX_s_1_2_2(and_727_nl, mux_tmp_334, or_850_cse);
  assign and_728_nl = nand_55_cse & mux_tmp_335;
  assign mux_tmp_336 = MUX_s_1_2_2(and_728_nl, mux_tmp_335, or_839_cse);
  assign and_729_nl = nand_58_cse & mux_tmp_336;
  assign mux_tmp_337 = MUX_s_1_2_2(and_729_nl, mux_tmp_336, or_830_cse);
  assign and_730_nl = not_tmp_645 & mux_tmp_337;
  assign mux_tmp_338 = MUX_s_1_2_2(and_730_nl, mux_tmp_337, or_823_cse);
  assign nor_417_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_338));
  assign mux_339_nl = MUX_s_1_2_2(nor_417_nl, mux_tmp_338, or_818_cse);
  assign and_dcpl_560 = mux_339_nl & and_dcpl_4 & and_dcpl_18 & (~ (result_rem_11cyc_st_9[0]));
  assign or_tmp_897 = (~ main_stage_0_10) | (~ asn_itm_9) | (result_rem_11cyc_st_9!=4'b1000);
  assign nor_407_nl = ~((result_rem_11cyc_st_8[3]) | (~ or_tmp_897));
  assign or_914_nl = (~ main_stage_0_9) | (~ asn_itm_8) | (result_rem_11cyc_st_8[2:0]!=3'b000);
  assign mux_tmp_340 = MUX_s_1_2_2(nor_407_nl, or_tmp_897, or_914_nl);
  assign nor_408_nl = ~((result_rem_11cyc_st_7[3]) | (~ mux_tmp_340));
  assign or_913_nl = (~ main_stage_0_8) | (~ asn_itm_7) | (result_rem_11cyc_st_7[2:0]!=3'b000);
  assign mux_tmp_341 = MUX_s_1_2_2(nor_408_nl, mux_tmp_340, or_913_nl);
  assign nor_409_nl = ~((result_rem_11cyc_st_6[3]) | (~ mux_tmp_341));
  assign or_912_nl = (~ main_stage_0_7) | (~ asn_itm_6) | (result_rem_11cyc_st_6[2:0]!=3'b000);
  assign mux_tmp_342 = MUX_s_1_2_2(nor_409_nl, mux_tmp_341, or_912_nl);
  assign nor_410_nl = ~((result_rem_11cyc_st_5[3]) | (~ mux_tmp_342));
  assign or_911_nl = (~ main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5[2:0]!=3'b000);
  assign mux_tmp_343 = MUX_s_1_2_2(nor_410_nl, mux_tmp_342, or_911_nl);
  assign nor_411_nl = ~((result_rem_11cyc_st_4[3]) | (~ mux_tmp_343));
  assign or_910_nl = (~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4[2:0]!=3'b000);
  assign mux_tmp_344 = MUX_s_1_2_2(nor_411_nl, mux_tmp_343, or_910_nl);
  assign nor_412_nl = ~((result_rem_11cyc_st_3[3]) | (~ mux_tmp_344));
  assign or_909_nl = (~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3[2:0]!=3'b000);
  assign mux_tmp_345 = MUX_s_1_2_2(nor_412_nl, mux_tmp_344, or_909_nl);
  assign nor_413_nl = ~((result_rem_11cyc_st_2[3]) | (~ mux_tmp_345));
  assign or_908_nl = (~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2[2:0]!=3'b000);
  assign mux_tmp_346 = MUX_s_1_2_2(nor_413_nl, mux_tmp_345, or_908_nl);
  assign and_724_nl = not_tmp_645 & mux_tmp_346;
  assign mux_tmp_347 = MUX_s_1_2_2(and_724_nl, mux_tmp_346, or_823_cse);
  assign nor_414_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_347));
  assign mux_tmp_348 = MUX_s_1_2_2(nor_414_nl, mux_tmp_347, or_818_cse);
  assign and_dcpl_566 = and_dcpl_532 & and_dcpl_318;
  assign or_tmp_909 = (result_rem_11cyc[2:0]!=3'b001) | not_tmp_645;
  assign or_928_cse = (result_result_acc_tmp!=4'b1001);
  assign nor_406_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_909));
  assign mux_349_nl = MUX_s_1_2_2(nor_406_nl, or_tmp_909, or_928_cse);
  assign and_dcpl_568 = mux_349_nl & and_dcpl_204;
  assign or_933_cse = (result_rem_11cyc[2:0]!=3'b001);
  assign nor_405_nl = ~(and_749_cse | and_dcpl_204);
  assign or_935_nl = (result_rem_11cyc_st_2[2:0]!=3'b001) | (~ and_dcpl_202);
  assign mux_tmp_350 = MUX_s_1_2_2(nor_405_nl, or_935_nl, or_933_cse);
  assign nor_404_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_350));
  assign mux_351_nl = MUX_s_1_2_2(nor_404_nl, mux_tmp_350, or_928_cse);
  assign and_dcpl_570 = mux_351_nl & and_dcpl_178;
  assign or_940_cse = (result_rem_11cyc_st_2[2:0]!=3'b001);
  assign nor_403_nl = ~(and_747_cse | and_dcpl_178);
  assign or_942_nl = (result_rem_11cyc_st_3[2:0]!=3'b001) | (~ and_dcpl_176);
  assign mux_tmp_352 = MUX_s_1_2_2(nor_403_nl, or_942_nl, or_940_cse);
  assign and_722_nl = not_tmp_645 & mux_tmp_352;
  assign mux_tmp_353 = MUX_s_1_2_2(and_722_nl, mux_tmp_352, or_933_cse);
  assign nor_402_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_353));
  assign mux_354_nl = MUX_s_1_2_2(nor_402_nl, mux_tmp_353, or_928_cse);
  assign and_dcpl_572 = mux_354_nl & and_dcpl_152;
  assign or_949_cse = (result_rem_11cyc_st_3[2:0]!=3'b001);
  assign nor_401_nl = ~(and_744_cse | and_dcpl_152);
  assign or_951_nl = (result_rem_11cyc_st_4[2:0]!=3'b001) | (~ and_dcpl_150);
  assign mux_tmp_355 = MUX_s_1_2_2(nor_401_nl, or_951_nl, or_949_cse);
  assign and_719_nl = nand_58_cse & mux_tmp_355;
  assign mux_tmp_356 = MUX_s_1_2_2(and_719_nl, mux_tmp_355, or_940_cse);
  assign and_720_nl = not_tmp_645 & mux_tmp_356;
  assign mux_tmp_357 = MUX_s_1_2_2(and_720_nl, mux_tmp_356, or_933_cse);
  assign nor_400_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_357));
  assign mux_358_nl = MUX_s_1_2_2(nor_400_nl, mux_tmp_357, or_928_cse);
  assign and_dcpl_576 = mux_358_nl & and_dcpl_125;
  assign or_960_cse = (result_rem_11cyc_st_4[2:0]!=3'b001);
  assign nor_399_nl = ~(and_740_cse | and_dcpl_125);
  assign or_962_nl = (result_rem_11cyc_st_5!=4'b1001) | (~ and_dcpl_105);
  assign mux_tmp_359 = MUX_s_1_2_2(nor_399_nl, or_962_nl, or_960_cse);
  assign and_715_nl = nand_55_cse & mux_tmp_359;
  assign mux_tmp_360 = MUX_s_1_2_2(and_715_nl, mux_tmp_359, or_949_cse);
  assign and_716_nl = nand_58_cse & mux_tmp_360;
  assign mux_tmp_361 = MUX_s_1_2_2(and_716_nl, mux_tmp_360, or_940_cse);
  assign and_717_nl = not_tmp_645 & mux_tmp_361;
  assign mux_tmp_362 = MUX_s_1_2_2(and_717_nl, mux_tmp_361, or_933_cse);
  assign nor_398_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_362));
  assign mux_363_nl = MUX_s_1_2_2(nor_398_nl, mux_tmp_362, or_928_cse);
  assign and_dcpl_578 = mux_363_nl & and_dcpl_101;
  assign or_973_cse = (result_rem_11cyc_st_5!=4'b1001);
  assign nor_397_nl = ~(and_dcpl_105 | and_dcpl_101);
  assign or_975_nl = (result_rem_11cyc_st_6[2:0]!=3'b001) | (~ and_dcpl_99);
  assign mux_tmp_364 = MUX_s_1_2_2(nor_397_nl, or_975_nl, or_973_cse);
  assign and_710_nl = nand_51_cse & mux_tmp_364;
  assign mux_tmp_365 = MUX_s_1_2_2(and_710_nl, mux_tmp_364, or_960_cse);
  assign and_711_nl = nand_55_cse & mux_tmp_365;
  assign mux_tmp_366 = MUX_s_1_2_2(and_711_nl, mux_tmp_365, or_949_cse);
  assign and_712_nl = nand_58_cse & mux_tmp_366;
  assign mux_tmp_367 = MUX_s_1_2_2(and_712_nl, mux_tmp_366, or_940_cse);
  assign and_713_nl = not_tmp_645 & mux_tmp_367;
  assign mux_tmp_368 = MUX_s_1_2_2(and_713_nl, mux_tmp_367, or_933_cse);
  assign nor_396_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_368));
  assign mux_369_nl = MUX_s_1_2_2(nor_396_nl, mux_tmp_368, or_928_cse);
  assign and_dcpl_580 = mux_369_nl & and_dcpl_75;
  assign or_988_cse = (result_rem_11cyc_st_6[2:0]!=3'b001);
  assign nor_394_nl = ~(and_731_cse | and_dcpl_75);
  assign or_990_nl = (result_rem_11cyc_st_7[2:0]!=3'b001) | (~ and_dcpl_73);
  assign mux_tmp_370 = MUX_s_1_2_2(nor_394_nl, or_990_nl, or_988_cse);
  assign nor_395_nl = ~(and_dcpl_105 | (~ mux_tmp_370));
  assign mux_tmp_371 = MUX_s_1_2_2(nor_395_nl, mux_tmp_370, or_973_cse);
  assign and_706_nl = nand_51_cse & mux_tmp_371;
  assign mux_tmp_372 = MUX_s_1_2_2(and_706_nl, mux_tmp_371, or_960_cse);
  assign and_707_nl = nand_55_cse & mux_tmp_372;
  assign mux_tmp_373 = MUX_s_1_2_2(and_707_nl, mux_tmp_372, or_949_cse);
  assign and_708_nl = nand_58_cse & mux_tmp_373;
  assign mux_tmp_374 = MUX_s_1_2_2(and_708_nl, mux_tmp_373, or_940_cse);
  assign and_709_nl = not_tmp_645 & mux_tmp_374;
  assign mux_tmp_375 = MUX_s_1_2_2(and_709_nl, mux_tmp_374, or_933_cse);
  assign nor_393_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_375));
  assign mux_376_nl = MUX_s_1_2_2(nor_393_nl, mux_tmp_375, or_928_cse);
  assign and_dcpl_583 = mux_376_nl & and_dcpl_47;
  assign nor_390_nl = ~(and_725_cse | and_dcpl_47);
  assign or_1007_nl = (result_rem_11cyc_st_8!=4'b1001) | (~ and_dcpl_28);
  assign or_1005_nl = (result_rem_11cyc_st_7[2:0]!=3'b001);
  assign mux_tmp_377 = MUX_s_1_2_2(nor_390_nl, or_1007_nl, or_1005_nl);
  assign and_700_nl = nand_42_cse & mux_tmp_377;
  assign mux_tmp_378 = MUX_s_1_2_2(and_700_nl, mux_tmp_377, or_988_cse);
  assign nor_391_nl = ~(and_dcpl_105 | (~ mux_tmp_378));
  assign mux_tmp_379 = MUX_s_1_2_2(nor_391_nl, mux_tmp_378, or_973_cse);
  assign and_701_nl = nand_51_cse & mux_tmp_379;
  assign mux_tmp_380 = MUX_s_1_2_2(and_701_nl, mux_tmp_379, or_960_cse);
  assign and_702_nl = nand_55_cse & mux_tmp_380;
  assign mux_tmp_381 = MUX_s_1_2_2(and_702_nl, mux_tmp_380, or_949_cse);
  assign and_703_nl = nand_58_cse & mux_tmp_381;
  assign mux_tmp_382 = MUX_s_1_2_2(and_703_nl, mux_tmp_381, or_940_cse);
  assign and_704_nl = not_tmp_645 & mux_tmp_382;
  assign mux_tmp_383 = MUX_s_1_2_2(and_704_nl, mux_tmp_382, or_933_cse);
  assign nor_392_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_383));
  assign mux_384_nl = MUX_s_1_2_2(nor_392_nl, mux_tmp_383, or_928_cse);
  assign and_dcpl_586 = mux_384_nl & and_dcpl_4 & and_dcpl_18 & (result_rem_11cyc_st_9[0]);
  assign or_tmp_1005 = (~ main_stage_0_10) | (~ asn_itm_9) | (result_rem_11cyc_st_9!=4'b1001);
  assign nor_383_nl = ~((result_rem_11cyc_st_8[3]) | (~ or_tmp_1005));
  assign or_1024_nl = (~ main_stage_0_9) | (~ asn_itm_8) | (result_rem_11cyc_st_8[2:0]!=3'b001);
  assign mux_tmp_385 = MUX_s_1_2_2(nor_383_nl, or_tmp_1005, or_1024_nl);
  assign nor_384_nl = ~((result_rem_11cyc_st_7[3]) | (~ mux_tmp_385));
  assign or_1023_nl = (~ main_stage_0_8) | (~ asn_itm_7) | (result_rem_11cyc_st_7[2:0]!=3'b001);
  assign mux_tmp_386 = MUX_s_1_2_2(nor_384_nl, mux_tmp_385, or_1023_nl);
  assign nor_385_nl = ~((result_rem_11cyc_st_6[3]) | (~ mux_tmp_386));
  assign or_1022_nl = (~ main_stage_0_7) | (~ asn_itm_6) | (result_rem_11cyc_st_6[2:0]!=3'b001);
  assign mux_tmp_387 = MUX_s_1_2_2(nor_385_nl, mux_tmp_386, or_1022_nl);
  assign nor_386_nl = ~((result_rem_11cyc_st_5[3]) | (~ mux_tmp_387));
  assign or_1021_nl = (~ main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5[2:0]!=3'b001);
  assign mux_tmp_388 = MUX_s_1_2_2(nor_386_nl, mux_tmp_387, or_1021_nl);
  assign nor_387_nl = ~((result_rem_11cyc_st_4[3]) | (~ mux_tmp_388));
  assign or_1020_nl = (~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4[2:0]!=3'b001);
  assign mux_tmp_389 = MUX_s_1_2_2(nor_387_nl, mux_tmp_388, or_1020_nl);
  assign nor_388_nl = ~((result_rem_11cyc_st_3[3]) | (~ mux_tmp_389));
  assign or_1019_nl = (~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3[2:0]!=3'b001);
  assign mux_tmp_390 = MUX_s_1_2_2(nor_388_nl, mux_tmp_389, or_1019_nl);
  assign nor_389_nl = ~((result_rem_11cyc_st_2[3]) | (~ mux_tmp_390));
  assign or_1018_nl = (~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2[2:0]!=3'b001);
  assign mux_tmp_391 = MUX_s_1_2_2(nor_389_nl, mux_tmp_390, or_1018_nl);
  assign and_697_nl = not_tmp_645 & mux_tmp_391;
  assign mux_tmp_392 = MUX_s_1_2_2(and_697_nl, mux_tmp_391, or_933_cse);
  assign and_698_nl = nand_146_cse & mux_tmp_392;
  assign or_1016_nl = (result_result_acc_tmp[3:1]!=3'b100);
  assign mux_tmp_393 = MUX_s_1_2_2(and_698_nl, mux_tmp_392, or_1016_nl);
  assign and_dcpl_590 = and_dcpl_532 & and_dcpl_352;
  assign or_tmp_1017 = (result_rem_11cyc[2:0]!=3'b010) | not_tmp_645;
  assign or_1037_cse = (result_result_acc_tmp!=4'b1010);
  assign nor_382_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_1017));
  assign mux_394_nl = MUX_s_1_2_2(nor_382_nl, or_tmp_1017, or_1037_cse);
  assign and_dcpl_592 = mux_394_nl & and_dcpl_205;
  assign or_1042_cse = (result_rem_11cyc[2:0]!=3'b010);
  assign nor_381_nl = ~(and_749_cse | and_dcpl_205);
  assign or_1044_nl = (result_rem_11cyc_st_2[2:0]!=3'b010) | (~ and_dcpl_202);
  assign mux_tmp_395 = MUX_s_1_2_2(nor_381_nl, or_1044_nl, or_1042_cse);
  assign nor_380_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_395));
  assign mux_396_nl = MUX_s_1_2_2(nor_380_nl, mux_tmp_395, or_1037_cse);
  assign and_dcpl_594 = mux_396_nl & and_dcpl_179;
  assign or_1049_cse = (result_rem_11cyc_st_2[2:0]!=3'b010);
  assign nor_379_nl = ~(and_747_cse | and_dcpl_179);
  assign or_1051_nl = (result_rem_11cyc_st_3[2:0]!=3'b010) | (~ and_dcpl_176);
  assign mux_tmp_397 = MUX_s_1_2_2(nor_379_nl, or_1051_nl, or_1049_cse);
  assign and_695_nl = not_tmp_645 & mux_tmp_397;
  assign mux_tmp_398 = MUX_s_1_2_2(and_695_nl, mux_tmp_397, or_1042_cse);
  assign nor_378_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_398));
  assign mux_399_nl = MUX_s_1_2_2(nor_378_nl, mux_tmp_398, or_1037_cse);
  assign and_dcpl_596 = mux_399_nl & and_dcpl_153;
  assign or_1058_cse = (result_rem_11cyc_st_3[2:0]!=3'b010);
  assign nor_377_nl = ~(and_744_cse | and_dcpl_153);
  assign or_1060_nl = (result_rem_11cyc_st_4[2:0]!=3'b010) | (~ and_dcpl_150);
  assign mux_tmp_400 = MUX_s_1_2_2(nor_377_nl, or_1060_nl, or_1058_cse);
  assign and_692_nl = nand_58_cse & mux_tmp_400;
  assign mux_tmp_401 = MUX_s_1_2_2(and_692_nl, mux_tmp_400, or_1049_cse);
  assign and_693_nl = not_tmp_645 & mux_tmp_401;
  assign mux_tmp_402 = MUX_s_1_2_2(and_693_nl, mux_tmp_401, or_1042_cse);
  assign nor_376_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_402));
  assign mux_403_nl = MUX_s_1_2_2(nor_376_nl, mux_tmp_402, or_1037_cse);
  assign and_dcpl_599 = mux_403_nl & and_dcpl_127;
  assign or_1069_cse = (result_rem_11cyc_st_4[2:0]!=3'b010);
  assign nor_375_nl = ~(and_740_cse | and_dcpl_127);
  assign or_1071_nl = (result_rem_11cyc_st_5!=4'b1010) | (~ and_dcpl_105);
  assign mux_tmp_404 = MUX_s_1_2_2(nor_375_nl, or_1071_nl, or_1069_cse);
  assign and_688_nl = nand_55_cse & mux_tmp_404;
  assign mux_tmp_405 = MUX_s_1_2_2(and_688_nl, mux_tmp_404, or_1058_cse);
  assign and_689_nl = nand_58_cse & mux_tmp_405;
  assign mux_tmp_406 = MUX_s_1_2_2(and_689_nl, mux_tmp_405, or_1049_cse);
  assign and_690_nl = not_tmp_645 & mux_tmp_406;
  assign mux_tmp_407 = MUX_s_1_2_2(and_690_nl, mux_tmp_406, or_1042_cse);
  assign nor_374_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_407));
  assign mux_408_nl = MUX_s_1_2_2(nor_374_nl, mux_tmp_407, or_1037_cse);
  assign and_dcpl_601 = mux_408_nl & and_dcpl_102;
  assign or_1082_cse = (result_rem_11cyc_st_5!=4'b1010);
  assign nor_373_nl = ~(and_dcpl_105 | and_dcpl_102);
  assign or_1084_nl = (result_rem_11cyc_st_6[2:0]!=3'b010) | (~ and_dcpl_99);
  assign mux_tmp_409 = MUX_s_1_2_2(nor_373_nl, or_1084_nl, or_1082_cse);
  assign and_683_nl = nand_51_cse & mux_tmp_409;
  assign mux_tmp_410 = MUX_s_1_2_2(and_683_nl, mux_tmp_409, or_1069_cse);
  assign and_684_nl = nand_55_cse & mux_tmp_410;
  assign mux_tmp_411 = MUX_s_1_2_2(and_684_nl, mux_tmp_410, or_1058_cse);
  assign and_685_nl = nand_58_cse & mux_tmp_411;
  assign mux_tmp_412 = MUX_s_1_2_2(and_685_nl, mux_tmp_411, or_1049_cse);
  assign and_686_nl = not_tmp_645 & mux_tmp_412;
  assign mux_tmp_413 = MUX_s_1_2_2(and_686_nl, mux_tmp_412, or_1042_cse);
  assign nor_372_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_413));
  assign mux_414_nl = MUX_s_1_2_2(nor_372_nl, mux_tmp_413, or_1037_cse);
  assign and_dcpl_603 = mux_414_nl & and_dcpl_76;
  assign or_1097_cse = (result_rem_11cyc_st_6[2:0]!=3'b010);
  assign nor_370_nl = ~(and_731_cse | and_dcpl_76);
  assign or_1099_nl = (result_rem_11cyc_st_7[2:0]!=3'b010) | (~ and_dcpl_73);
  assign mux_tmp_415 = MUX_s_1_2_2(nor_370_nl, or_1099_nl, or_1097_cse);
  assign nor_371_nl = ~(and_dcpl_105 | (~ mux_tmp_415));
  assign mux_tmp_416 = MUX_s_1_2_2(nor_371_nl, mux_tmp_415, or_1082_cse);
  assign and_679_nl = nand_51_cse & mux_tmp_416;
  assign mux_tmp_417 = MUX_s_1_2_2(and_679_nl, mux_tmp_416, or_1069_cse);
  assign and_680_nl = nand_55_cse & mux_tmp_417;
  assign mux_tmp_418 = MUX_s_1_2_2(and_680_nl, mux_tmp_417, or_1058_cse);
  assign and_681_nl = nand_58_cse & mux_tmp_418;
  assign mux_tmp_419 = MUX_s_1_2_2(and_681_nl, mux_tmp_418, or_1049_cse);
  assign and_682_nl = not_tmp_645 & mux_tmp_419;
  assign mux_tmp_420 = MUX_s_1_2_2(and_682_nl, mux_tmp_419, or_1042_cse);
  assign nor_369_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_420));
  assign mux_421_nl = MUX_s_1_2_2(nor_369_nl, mux_tmp_420, or_1037_cse);
  assign and_dcpl_607 = mux_421_nl & and_dcpl_50;
  assign nor_366_nl = ~(and_725_cse | and_dcpl_50);
  assign or_1116_nl = (result_rem_11cyc_st_8!=4'b1010) | (~ and_dcpl_28);
  assign or_1114_nl = (result_rem_11cyc_st_7[2:0]!=3'b010);
  assign mux_tmp_422 = MUX_s_1_2_2(nor_366_nl, or_1116_nl, or_1114_nl);
  assign and_673_nl = nand_42_cse & mux_tmp_422;
  assign mux_tmp_423 = MUX_s_1_2_2(and_673_nl, mux_tmp_422, or_1097_cse);
  assign nor_367_nl = ~(and_dcpl_105 | (~ mux_tmp_423));
  assign mux_tmp_424 = MUX_s_1_2_2(nor_367_nl, mux_tmp_423, or_1082_cse);
  assign and_674_nl = nand_51_cse & mux_tmp_424;
  assign mux_tmp_425 = MUX_s_1_2_2(and_674_nl, mux_tmp_424, or_1069_cse);
  assign and_675_nl = nand_55_cse & mux_tmp_425;
  assign mux_tmp_426 = MUX_s_1_2_2(and_675_nl, mux_tmp_425, or_1058_cse);
  assign and_676_nl = nand_58_cse & mux_tmp_426;
  assign mux_tmp_427 = MUX_s_1_2_2(and_676_nl, mux_tmp_426, or_1049_cse);
  assign and_677_nl = not_tmp_645 & mux_tmp_427;
  assign mux_tmp_428 = MUX_s_1_2_2(and_677_nl, mux_tmp_427, or_1042_cse);
  assign nor_368_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_428));
  assign mux_429_nl = MUX_s_1_2_2(nor_368_nl, mux_tmp_428, or_1037_cse);
  assign and_dcpl_611 = mux_429_nl & and_dcpl_4 & (result_rem_11cyc_st_9[3]) & (result_rem_11cyc_st_9[1])
      & (~ (result_rem_11cyc_st_9[0]));
  assign or_tmp_1113 = (~ main_stage_0_10) | (~ asn_itm_9) | (result_rem_11cyc_st_9!=4'b1010);
  assign nor_358_nl = ~((result_rem_11cyc_st_8[3]) | (~ or_tmp_1113));
  assign or_1133_nl = (~ main_stage_0_9) | (~ asn_itm_8) | (result_rem_11cyc_st_8[2:0]!=3'b010);
  assign mux_tmp_430 = MUX_s_1_2_2(nor_358_nl, or_tmp_1113, or_1133_nl);
  assign nor_359_nl = ~((result_rem_11cyc_st_7[3]) | (~ mux_tmp_430));
  assign or_1132_nl = (~ main_stage_0_8) | (~ asn_itm_7) | (result_rem_11cyc_st_7[2:0]!=3'b010);
  assign mux_tmp_431 = MUX_s_1_2_2(nor_359_nl, mux_tmp_430, or_1132_nl);
  assign nor_360_nl = ~((result_rem_11cyc_st_6[3]) | (~ mux_tmp_431));
  assign or_1131_nl = (~ main_stage_0_7) | (~ asn_itm_6) | (result_rem_11cyc_st_6[2:0]!=3'b010);
  assign mux_tmp_432 = MUX_s_1_2_2(nor_360_nl, mux_tmp_431, or_1131_nl);
  assign nor_361_nl = ~((result_rem_11cyc_st_5[3]) | (~ mux_tmp_432));
  assign or_1130_nl = (~ main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5[2:0]!=3'b010);
  assign mux_tmp_433 = MUX_s_1_2_2(nor_361_nl, mux_tmp_432, or_1130_nl);
  assign nor_362_nl = ~((result_rem_11cyc_st_4[3]) | (~ mux_tmp_433));
  assign or_1129_nl = (~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4[2:0]!=3'b010);
  assign mux_tmp_434 = MUX_s_1_2_2(nor_362_nl, mux_tmp_433, or_1129_nl);
  assign nor_363_nl = ~((result_rem_11cyc_st_3[3]) | (~ mux_tmp_434));
  assign or_1128_nl = (~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3[2:0]!=3'b010);
  assign mux_tmp_435 = MUX_s_1_2_2(nor_363_nl, mux_tmp_434, or_1128_nl);
  assign nor_364_nl = ~((result_rem_11cyc_st_2[3]) | (~ mux_tmp_435));
  assign or_1127_nl = (~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2[2:0]!=3'b010);
  assign mux_tmp_436 = MUX_s_1_2_2(nor_364_nl, mux_tmp_435, or_1127_nl);
  assign and_671_nl = not_tmp_645 & mux_tmp_436;
  assign mux_tmp_437 = MUX_s_1_2_2(and_671_nl, mux_tmp_436, or_1042_cse);
  assign nor_365_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_437));
  assign mux_tmp_438 = MUX_s_1_2_2(nor_365_nl, mux_tmp_437, or_1037_cse);
  assign return_rsci_d_mx0c0 = and_dcpl_235 & and_dcpl_233;
  assign return_rsci_d_mx0c1 = and_dcpl_235 & and_dcpl_237;
  assign return_rsci_d_mx0c2 = and_dcpl_235 & and_dcpl_240;
  assign return_rsci_d_mx0c3 = and_dcpl_235 & and_dcpl_239 & (result_rem_11cyc_st_11[0]);
  assign return_rsci_d_mx0c4 = and_dcpl_235 & and_dcpl_244 & (~ (result_rem_11cyc_st_11[0]));
  assign return_rsci_d_mx0c5 = and_dcpl_235 & and_dcpl_244 & (result_rem_11cyc_st_11[0]);
  assign return_rsci_d_mx0c6 = and_dcpl_235 & and_dcpl_249 & (~ (result_rem_11cyc_st_11[0]));
  assign return_rsci_d_mx0c7 = and_dcpl_235 & and_dcpl_249 & (result_rem_11cyc_st_11[0]);
  assign return_rsci_d_mx0c8 = and_dcpl_254 & and_dcpl_233;
  assign return_rsci_d_mx0c9 = and_dcpl_254 & and_dcpl_237;
  assign return_rsci_d_mx0c10 = and_dcpl_254 & and_dcpl_240;
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_en & (return_rsci_d_mx0c0 | return_rsci_d_mx0c1 | return_rsci_d_mx0c2
        | return_rsci_d_mx0c3 | return_rsci_d_mx0c4 | return_rsci_d_mx0c5 | return_rsci_d_mx0c6
        | return_rsci_d_mx0c7 | return_rsci_d_mx0c8 | return_rsci_d_mx0c9 | return_rsci_d_mx0c10)
        ) begin
      return_rsci_d <= MUX1HOT_v_64_11_2(result_rem_12_cmp_1_z, result_rem_12_cmp_2_z,
          result_rem_12_cmp_3_z, result_rem_12_cmp_4_z, result_rem_12_cmp_5_z, result_rem_12_cmp_6_z,
          result_rem_12_cmp_7_z, result_rem_12_cmp_8_z, result_rem_12_cmp_9_z, result_rem_12_cmp_10_z,
          result_rem_12_cmp_z, {return_rsci_d_mx0c0 , return_rsci_d_mx0c1 , return_rsci_d_mx0c2
          , return_rsci_d_mx0c3 , return_rsci_d_mx0c4 , return_rsci_d_mx0c5 , return_rsci_d_mx0c6
          , return_rsci_d_mx0c7 , return_rsci_d_mx0c8 , return_rsci_d_mx0c9 , return_rsci_d_mx0c10});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_11 <= 4'b0000;
    end
    else if ( ccs_ccore_en & main_stage_0_11 & asn_itm_10 ) begin
      result_rem_11cyc_st_11 <= result_rem_11cyc_st_10;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      asn_itm_11 <= 1'b0;
      asn_itm_10 <= 1'b0;
      asn_itm_9 <= 1'b0;
      asn_itm_8 <= 1'b0;
      asn_itm_7 <= 1'b0;
      asn_itm_6 <= 1'b0;
      asn_itm_5 <= 1'b0;
      asn_itm_4 <= 1'b0;
      asn_itm_3 <= 1'b0;
      asn_itm_2 <= 1'b0;
      asn_itm_1 <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
      main_stage_0_5 <= 1'b0;
      main_stage_0_6 <= 1'b0;
      main_stage_0_7 <= 1'b0;
      main_stage_0_8 <= 1'b0;
      main_stage_0_9 <= 1'b0;
      main_stage_0_10 <= 1'b0;
      main_stage_0_11 <= 1'b0;
      main_stage_0_12 <= 1'b0;
    end
    else if ( ccs_ccore_en ) begin
      asn_itm_11 <= asn_itm_10;
      asn_itm_10 <= asn_itm_9;
      asn_itm_9 <= asn_itm_8;
      asn_itm_8 <= asn_itm_7;
      asn_itm_7 <= asn_itm_6;
      asn_itm_6 <= asn_itm_5;
      asn_itm_5 <= asn_itm_4;
      asn_itm_4 <= asn_itm_3;
      asn_itm_3 <= asn_itm_2;
      asn_itm_2 <= asn_itm_1;
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
      main_stage_0_4 <= main_stage_0_3;
      main_stage_0_5 <= main_stage_0_4;
      main_stage_0_6 <= main_stage_0_5;
      main_stage_0_7 <= main_stage_0_6;
      main_stage_0_8 <= main_stage_0_7;
      main_stage_0_9 <= main_stage_0_8;
      main_stage_0_10 <= main_stage_0_9;
      main_stage_0_11 <= main_stage_0_10;
      main_stage_0_12 <= main_stage_0_11;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_1_cse ) begin
      result_rem_12_cmp_1_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_1_2,
          m_buf_sva_mut_1_3, m_buf_sva_mut_1_4, m_buf_sva_mut_1_5, m_buf_sva_mut_1_6,
          m_buf_sva_mut_1_7, m_buf_sva_mut_1_8, m_buf_sva_mut_1_9, m_buf_sva_mut_1_10,
          {and_dcpl_263 , and_dcpl_269 , and_dcpl_275 , and_dcpl_281 , and_dcpl_287
          , and_dcpl_293 , and_dcpl_299 , and_dcpl_305 , and_dcpl_311 , mux_tmp_37});
      result_rem_12_cmp_1_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_1_2,
          base_buf_sva_mut_1_3, base_buf_sva_mut_1_4, base_buf_sva_mut_1_5, base_buf_sva_mut_1_6,
          base_buf_sva_mut_1_7, base_buf_sva_mut_1_8, base_buf_sva_mut_1_9, base_buf_sva_mut_1_10,
          {and_dcpl_263 , and_dcpl_269 , and_dcpl_275 , and_dcpl_281 , and_dcpl_287
          , and_dcpl_293 , and_dcpl_299 , and_dcpl_305 , and_dcpl_311 , mux_tmp_37});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_3_cse ) begin
      result_rem_12_cmp_2_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_2_2,
          m_buf_sva_mut_2_3, m_buf_sva_mut_2_4, m_buf_sva_mut_2_5, m_buf_sva_mut_2_6,
          m_buf_sva_mut_2_7, m_buf_sva_mut_2_8, m_buf_sva_mut_2_9, m_buf_sva_mut_2_10,
          {and_dcpl_319 , and_dcpl_322 , and_dcpl_325 , and_dcpl_329 , and_dcpl_333
          , and_dcpl_337 , and_dcpl_341 , and_dcpl_344 , and_dcpl_347 , mux_tmp_75});
      result_rem_12_cmp_2_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_2_2,
          base_buf_sva_mut_2_3, base_buf_sva_mut_2_4, base_buf_sva_mut_2_5, base_buf_sva_mut_2_6,
          base_buf_sva_mut_2_7, base_buf_sva_mut_2_8, base_buf_sva_mut_2_9, base_buf_sva_mut_2_10,
          {and_dcpl_319 , and_dcpl_322 , and_dcpl_325 , and_dcpl_329 , and_dcpl_333
          , and_dcpl_337 , and_dcpl_341 , and_dcpl_344 , and_dcpl_347 , mux_tmp_75});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_5_cse ) begin
      result_rem_12_cmp_3_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_3_2,
          m_buf_sva_mut_3_3, m_buf_sva_mut_3_4, m_buf_sva_mut_3_5, m_buf_sva_mut_3_6,
          m_buf_sva_mut_3_7, m_buf_sva_mut_3_8, m_buf_sva_mut_3_9, m_buf_sva_mut_3_10,
          {and_dcpl_353 , and_dcpl_357 , and_dcpl_361 , and_dcpl_364 , and_dcpl_367
          , and_dcpl_370 , and_dcpl_373 , and_dcpl_377 , and_dcpl_381 , mux_tmp_113});
      result_rem_12_cmp_3_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_3_2,
          base_buf_sva_mut_3_3, base_buf_sva_mut_3_4, base_buf_sva_mut_3_5, base_buf_sva_mut_3_6,
          base_buf_sva_mut_3_7, base_buf_sva_mut_3_8, base_buf_sva_mut_3_9, base_buf_sva_mut_3_10,
          {and_dcpl_353 , and_dcpl_357 , and_dcpl_361 , and_dcpl_364 , and_dcpl_367
          , and_dcpl_370 , and_dcpl_373 , and_dcpl_377 , and_dcpl_381 , mux_tmp_113});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_7_cse ) begin
      result_rem_12_cmp_4_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_4_2,
          m_buf_sva_mut_4_3, m_buf_sva_mut_4_4, m_buf_sva_mut_4_5, m_buf_sva_mut_4_6,
          m_buf_sva_mut_4_7, m_buf_sva_mut_4_8, m_buf_sva_mut_4_9, m_buf_sva_mut_4_10,
          {and_dcpl_387 , and_dcpl_390 , and_dcpl_393 , and_dcpl_396 , and_dcpl_399
          , and_dcpl_402 , and_dcpl_405 , and_dcpl_408 , and_dcpl_411 , mux_tmp_151});
      result_rem_12_cmp_4_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_4_2,
          base_buf_sva_mut_4_3, base_buf_sva_mut_4_4, base_buf_sva_mut_4_5, base_buf_sva_mut_4_6,
          base_buf_sva_mut_4_7, base_buf_sva_mut_4_8, base_buf_sva_mut_4_9, base_buf_sva_mut_4_10,
          {and_dcpl_387 , and_dcpl_390 , and_dcpl_393 , and_dcpl_396 , and_dcpl_399
          , and_dcpl_402 , and_dcpl_405 , and_dcpl_408 , and_dcpl_411 , mux_tmp_151});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_9_cse ) begin
      result_rem_12_cmp_5_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_5_2,
          m_buf_sva_mut_5_3, m_buf_sva_mut_5_4, m_buf_sva_mut_5_5, m_buf_sva_mut_5_6,
          m_buf_sva_mut_5_7, m_buf_sva_mut_5_8, m_buf_sva_mut_5_9, m_buf_sva_mut_5_10,
          {and_dcpl_418 , and_dcpl_422 , and_dcpl_426 , and_dcpl_430 , and_dcpl_433
          , and_dcpl_437 , and_dcpl_441 , and_dcpl_444 , and_dcpl_447 , mux_tmp_189});
      result_rem_12_cmp_5_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_5_2,
          base_buf_sva_mut_5_3, base_buf_sva_mut_5_4, base_buf_sva_mut_5_5, base_buf_sva_mut_5_6,
          base_buf_sva_mut_5_7, base_buf_sva_mut_5_8, base_buf_sva_mut_5_9, base_buf_sva_mut_5_10,
          {and_dcpl_418 , and_dcpl_422 , and_dcpl_426 , and_dcpl_430 , and_dcpl_433
          , and_dcpl_437 , and_dcpl_441 , and_dcpl_444 , and_dcpl_447 , mux_tmp_189});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_11_cse ) begin
      result_rem_12_cmp_6_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_6_2,
          m_buf_sva_mut_6_3, m_buf_sva_mut_6_4, m_buf_sva_mut_6_5, m_buf_sva_mut_6_6,
          m_buf_sva_mut_6_7, m_buf_sva_mut_6_8, m_buf_sva_mut_6_9, m_buf_sva_mut_6_10,
          {and_dcpl_452 , and_dcpl_455 , and_dcpl_458 , and_dcpl_462 , and_dcpl_464
          , and_dcpl_468 , and_dcpl_472 , and_dcpl_474 , and_dcpl_476 , mux_tmp_227});
      result_rem_12_cmp_6_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_6_2,
          base_buf_sva_mut_6_3, base_buf_sva_mut_6_4, base_buf_sva_mut_6_5, base_buf_sva_mut_6_6,
          base_buf_sva_mut_6_7, base_buf_sva_mut_6_8, base_buf_sva_mut_6_9, base_buf_sva_mut_6_10,
          {and_dcpl_452 , and_dcpl_455 , and_dcpl_458 , and_dcpl_462 , and_dcpl_464
          , and_dcpl_468 , and_dcpl_472 , and_dcpl_474 , and_dcpl_476 , mux_tmp_227});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_13_cse ) begin
      result_rem_12_cmp_7_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_7_2,
          m_buf_sva_mut_7_3, m_buf_sva_mut_7_4, m_buf_sva_mut_7_5, m_buf_sva_mut_7_6,
          m_buf_sva_mut_7_7, m_buf_sva_mut_7_8, m_buf_sva_mut_7_9, m_buf_sva_mut_7_10,
          {and_dcpl_480 , and_dcpl_484 , and_dcpl_488 , and_dcpl_491 , and_dcpl_493
          , and_dcpl_496 , and_dcpl_499 , and_dcpl_501 , and_dcpl_503 , mux_tmp_265});
      result_rem_12_cmp_7_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_7_2,
          base_buf_sva_mut_7_3, base_buf_sva_mut_7_4, base_buf_sva_mut_7_5, base_buf_sva_mut_7_6,
          base_buf_sva_mut_7_7, base_buf_sva_mut_7_8, base_buf_sva_mut_7_9, base_buf_sva_mut_7_10,
          {and_dcpl_480 , and_dcpl_484 , and_dcpl_488 , and_dcpl_491 , and_dcpl_493
          , and_dcpl_496 , and_dcpl_499 , and_dcpl_501 , and_dcpl_503 , mux_tmp_265});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_15_cse ) begin
      result_rem_12_cmp_8_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_8_2,
          m_buf_sva_mut_8_3, m_buf_sva_mut_8_4, m_buf_sva_mut_8_5, m_buf_sva_mut_8_6,
          m_buf_sva_mut_8_7, m_buf_sva_mut_8_8, m_buf_sva_mut_8_9, m_buf_sva_mut_8_10,
          {and_dcpl_507 , and_dcpl_510 , and_dcpl_513 , and_dcpl_516 , and_dcpl_518
          , and_dcpl_521 , and_dcpl_524 , and_dcpl_526 , and_dcpl_528 , mux_tmp_303});
      result_rem_12_cmp_8_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_8_2,
          base_buf_sva_mut_8_3, base_buf_sva_mut_8_4, base_buf_sva_mut_8_5, base_buf_sva_mut_8_6,
          base_buf_sva_mut_8_7, base_buf_sva_mut_8_8, base_buf_sva_mut_8_9, base_buf_sva_mut_8_10,
          {and_dcpl_507 , and_dcpl_510 , and_dcpl_513 , and_dcpl_516 , and_dcpl_518
          , and_dcpl_521 , and_dcpl_524 , and_dcpl_526 , and_dcpl_528 , mux_tmp_303});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_17_cse ) begin
      result_rem_12_cmp_9_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_9_2,
          m_buf_sva_mut_9_3, m_buf_sva_mut_9_4, m_buf_sva_mut_9_5, m_buf_sva_mut_9_6,
          m_buf_sva_mut_9_7, m_buf_sva_mut_9_8, m_buf_sva_mut_9_9, m_buf_sva_mut_9_10,
          {and_dcpl_533 , and_dcpl_536 , and_dcpl_539 , and_dcpl_542 , and_dcpl_546
          , and_dcpl_549 , and_dcpl_552 , and_dcpl_556 , and_dcpl_560 , mux_tmp_348});
      result_rem_12_cmp_9_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_9_2,
          base_buf_sva_mut_9_3, base_buf_sva_mut_9_4, base_buf_sva_mut_9_5, base_buf_sva_mut_9_6,
          base_buf_sva_mut_9_7, base_buf_sva_mut_9_8, base_buf_sva_mut_9_9, base_buf_sva_mut_9_10,
          {and_dcpl_533 , and_dcpl_536 , and_dcpl_539 , and_dcpl_542 , and_dcpl_546
          , and_dcpl_549 , and_dcpl_552 , and_dcpl_556 , and_dcpl_560 , mux_tmp_348});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_19_cse ) begin
      result_rem_12_cmp_10_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_10_2,
          m_buf_sva_mut_10_3, m_buf_sva_mut_10_4, m_buf_sva_mut_10_5, m_buf_sva_mut_10_6,
          m_buf_sva_mut_10_7, m_buf_sva_mut_10_8, m_buf_sva_mut_10_9, m_buf_sva_mut_10_10,
          {and_dcpl_566 , and_dcpl_568 , and_dcpl_570 , and_dcpl_572 , and_dcpl_576
          , and_dcpl_578 , and_dcpl_580 , and_dcpl_583 , and_dcpl_586 , mux_tmp_393});
      result_rem_12_cmp_10_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_10_2,
          base_buf_sva_mut_10_3, base_buf_sva_mut_10_4, base_buf_sva_mut_10_5, base_buf_sva_mut_10_6,
          base_buf_sva_mut_10_7, base_buf_sva_mut_10_8, base_buf_sva_mut_10_9, base_buf_sva_mut_10_10,
          {and_dcpl_566 , and_dcpl_568 , and_dcpl_570 , and_dcpl_572 , and_dcpl_576
          , and_dcpl_578 , and_dcpl_580 , and_dcpl_583 , and_dcpl_586 , mux_tmp_393});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_21_cse ) begin
      result_rem_12_cmp_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_2, m_buf_sva_mut_3,
          m_buf_sva_mut_4, m_buf_sva_mut_5, m_buf_sva_mut_6, m_buf_sva_mut_7, m_buf_sva_mut_8,
          m_buf_sva_mut_9, m_buf_sva_mut_10, {and_dcpl_590 , and_dcpl_592 , and_dcpl_594
          , and_dcpl_596 , and_dcpl_599 , and_dcpl_601 , and_dcpl_603 , and_dcpl_607
          , and_dcpl_611 , mux_tmp_438});
      result_rem_12_cmp_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_2,
          base_buf_sva_mut_3, base_buf_sva_mut_4, base_buf_sva_mut_5, base_buf_sva_mut_6,
          base_buf_sva_mut_7, base_buf_sva_mut_8, base_buf_sva_mut_9, base_buf_sva_mut_10,
          {and_dcpl_590 , and_dcpl_592 , and_dcpl_594 , and_dcpl_596 , and_dcpl_599
          , and_dcpl_601 , and_dcpl_603 , and_dcpl_607 , and_dcpl_611 , mux_tmp_438});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_cse ) begin
      m_buf_sva_mut_1_10 <= m_buf_sva_mut_1_9;
      base_buf_sva_mut_1_10 <= base_buf_sva_mut_1_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_1_cse ) begin
      m_buf_sva_mut_2_10 <= m_buf_sva_mut_2_9;
      base_buf_sva_mut_2_10 <= base_buf_sva_mut_2_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_2_cse ) begin
      m_buf_sva_mut_3_10 <= m_buf_sva_mut_3_9;
      base_buf_sva_mut_3_10 <= base_buf_sva_mut_3_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_3_cse ) begin
      m_buf_sva_mut_4_10 <= m_buf_sva_mut_4_9;
      base_buf_sva_mut_4_10 <= base_buf_sva_mut_4_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_4_cse ) begin
      m_buf_sva_mut_5_10 <= m_buf_sva_mut_5_9;
      base_buf_sva_mut_5_10 <= base_buf_sva_mut_5_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_5_cse ) begin
      m_buf_sva_mut_6_10 <= m_buf_sva_mut_6_9;
      base_buf_sva_mut_6_10 <= base_buf_sva_mut_6_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_6_cse ) begin
      m_buf_sva_mut_7_10 <= m_buf_sva_mut_7_9;
      base_buf_sva_mut_7_10 <= base_buf_sva_mut_7_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_7_cse ) begin
      m_buf_sva_mut_8_10 <= m_buf_sva_mut_8_9;
      base_buf_sva_mut_8_10 <= base_buf_sva_mut_8_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_8_cse ) begin
      m_buf_sva_mut_9_10 <= m_buf_sva_mut_9_9;
      base_buf_sva_mut_9_10 <= base_buf_sva_mut_9_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_9_cse ) begin
      m_buf_sva_mut_10_10 <= m_buf_sva_mut_10_9;
      base_buf_sva_mut_10_10 <= base_buf_sva_mut_10_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_10_cse ) begin
      m_buf_sva_mut_10 <= m_buf_sva_mut_9;
      base_buf_sva_mut_10 <= base_buf_sva_mut_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_10 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_3 ) begin
      result_rem_11cyc_st_10 <= result_rem_11cyc_st_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_11_cse ) begin
      m_buf_sva_mut_1_9 <= m_buf_sva_mut_1_8;
      base_buf_sva_mut_1_9 <= base_buf_sva_mut_1_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_12_cse ) begin
      m_buf_sva_mut_2_9 <= m_buf_sva_mut_2_8;
      base_buf_sva_mut_2_9 <= base_buf_sva_mut_2_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_13_cse ) begin
      m_buf_sva_mut_3_9 <= m_buf_sva_mut_3_8;
      base_buf_sva_mut_3_9 <= base_buf_sva_mut_3_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_14_cse ) begin
      m_buf_sva_mut_4_9 <= m_buf_sva_mut_4_8;
      base_buf_sva_mut_4_9 <= base_buf_sva_mut_4_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_15_cse ) begin
      m_buf_sva_mut_5_9 <= m_buf_sva_mut_5_8;
      base_buf_sva_mut_5_9 <= base_buf_sva_mut_5_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_16_cse ) begin
      m_buf_sva_mut_6_9 <= m_buf_sva_mut_6_8;
      base_buf_sva_mut_6_9 <= base_buf_sva_mut_6_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_17_cse ) begin
      m_buf_sva_mut_7_9 <= m_buf_sva_mut_7_8;
      base_buf_sva_mut_7_9 <= base_buf_sva_mut_7_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_18_cse ) begin
      m_buf_sva_mut_8_9 <= m_buf_sva_mut_8_8;
      base_buf_sva_mut_8_9 <= base_buf_sva_mut_8_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_19_cse ) begin
      m_buf_sva_mut_9_9 <= m_buf_sva_mut_9_8;
      base_buf_sva_mut_9_9 <= base_buf_sva_mut_9_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_20_cse ) begin
      m_buf_sva_mut_10_9 <= m_buf_sva_mut_10_8;
      base_buf_sva_mut_10_9 <= base_buf_sva_mut_10_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_21_cse ) begin
      m_buf_sva_mut_9 <= m_buf_sva_mut_8;
      base_buf_sva_mut_9 <= base_buf_sva_mut_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_9 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_28 ) begin
      result_rem_11cyc_st_9 <= result_rem_11cyc_st_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_22_cse ) begin
      m_buf_sva_mut_1_8 <= m_buf_sva_mut_1_7;
      base_buf_sva_mut_1_8 <= base_buf_sva_mut_1_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_23_cse ) begin
      m_buf_sva_mut_2_8 <= m_buf_sva_mut_2_7;
      base_buf_sva_mut_2_8 <= base_buf_sva_mut_2_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_24_cse ) begin
      m_buf_sva_mut_3_8 <= m_buf_sva_mut_3_7;
      base_buf_sva_mut_3_8 <= base_buf_sva_mut_3_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_25_cse ) begin
      m_buf_sva_mut_4_8 <= m_buf_sva_mut_4_7;
      base_buf_sva_mut_4_8 <= base_buf_sva_mut_4_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_26_cse ) begin
      m_buf_sva_mut_5_8 <= m_buf_sva_mut_5_7;
      base_buf_sva_mut_5_8 <= base_buf_sva_mut_5_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_27_cse ) begin
      m_buf_sva_mut_6_8 <= m_buf_sva_mut_6_7;
      base_buf_sva_mut_6_8 <= base_buf_sva_mut_6_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_28_cse ) begin
      m_buf_sva_mut_7_8 <= m_buf_sva_mut_7_7;
      base_buf_sva_mut_7_8 <= base_buf_sva_mut_7_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_29_cse ) begin
      m_buf_sva_mut_8_8 <= m_buf_sva_mut_8_7;
      base_buf_sva_mut_8_8 <= base_buf_sva_mut_8_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_30_cse ) begin
      m_buf_sva_mut_9_8 <= m_buf_sva_mut_9_7;
      base_buf_sva_mut_9_8 <= base_buf_sva_mut_9_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_31_cse ) begin
      m_buf_sva_mut_10_8 <= m_buf_sva_mut_10_7;
      base_buf_sva_mut_10_8 <= base_buf_sva_mut_10_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_32_cse ) begin
      m_buf_sva_mut_8 <= m_buf_sva_mut_7;
      base_buf_sva_mut_8 <= base_buf_sva_mut_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_8 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_53 ) begin
      result_rem_11cyc_st_8 <= result_rem_11cyc_st_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_33_cse ) begin
      m_buf_sva_mut_1_7 <= m_buf_sva_mut_1_6;
      base_buf_sva_mut_1_7 <= base_buf_sva_mut_1_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_34_cse ) begin
      m_buf_sva_mut_2_7 <= m_buf_sva_mut_2_6;
      base_buf_sva_mut_2_7 <= base_buf_sva_mut_2_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_35_cse ) begin
      m_buf_sva_mut_3_7 <= m_buf_sva_mut_3_6;
      base_buf_sva_mut_3_7 <= base_buf_sva_mut_3_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_36_cse ) begin
      m_buf_sva_mut_4_7 <= m_buf_sva_mut_4_6;
      base_buf_sva_mut_4_7 <= base_buf_sva_mut_4_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_37_cse ) begin
      m_buf_sva_mut_5_7 <= m_buf_sva_mut_5_6;
      base_buf_sva_mut_5_7 <= base_buf_sva_mut_5_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_38_cse ) begin
      m_buf_sva_mut_6_7 <= m_buf_sva_mut_6_6;
      base_buf_sva_mut_6_7 <= base_buf_sva_mut_6_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_39_cse ) begin
      m_buf_sva_mut_7_7 <= m_buf_sva_mut_7_6;
      base_buf_sva_mut_7_7 <= base_buf_sva_mut_7_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_40_cse ) begin
      m_buf_sva_mut_8_7 <= m_buf_sva_mut_8_6;
      base_buf_sva_mut_8_7 <= base_buf_sva_mut_8_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_41_cse ) begin
      m_buf_sva_mut_9_7 <= m_buf_sva_mut_9_6;
      base_buf_sva_mut_9_7 <= base_buf_sva_mut_9_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_42_cse ) begin
      m_buf_sva_mut_10_7 <= m_buf_sva_mut_10_6;
      base_buf_sva_mut_10_7 <= base_buf_sva_mut_10_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_43_cse ) begin
      m_buf_sva_mut_7 <= m_buf_sva_mut_6;
      base_buf_sva_mut_7 <= base_buf_sva_mut_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_7 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_79 ) begin
      result_rem_11cyc_st_7 <= result_rem_11cyc_st_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_44_cse ) begin
      m_buf_sva_mut_1_6 <= m_buf_sva_mut_1_5;
      base_buf_sva_mut_1_6 <= base_buf_sva_mut_1_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_45_cse ) begin
      m_buf_sva_mut_2_6 <= m_buf_sva_mut_2_5;
      base_buf_sva_mut_2_6 <= base_buf_sva_mut_2_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_46_cse ) begin
      m_buf_sva_mut_3_6 <= m_buf_sva_mut_3_5;
      base_buf_sva_mut_3_6 <= base_buf_sva_mut_3_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_47_cse ) begin
      m_buf_sva_mut_4_6 <= m_buf_sva_mut_4_5;
      base_buf_sva_mut_4_6 <= base_buf_sva_mut_4_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_48_cse ) begin
      m_buf_sva_mut_5_6 <= m_buf_sva_mut_5_5;
      base_buf_sva_mut_5_6 <= base_buf_sva_mut_5_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_49_cse ) begin
      m_buf_sva_mut_6_6 <= m_buf_sva_mut_6_5;
      base_buf_sva_mut_6_6 <= base_buf_sva_mut_6_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_50_cse ) begin
      m_buf_sva_mut_7_6 <= m_buf_sva_mut_7_5;
      base_buf_sva_mut_7_6 <= base_buf_sva_mut_7_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_51_cse ) begin
      m_buf_sva_mut_8_6 <= m_buf_sva_mut_8_5;
      base_buf_sva_mut_8_6 <= base_buf_sva_mut_8_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_52_cse ) begin
      m_buf_sva_mut_9_6 <= m_buf_sva_mut_9_5;
      base_buf_sva_mut_9_6 <= base_buf_sva_mut_9_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_53_cse ) begin
      m_buf_sva_mut_10_6 <= m_buf_sva_mut_10_5;
      base_buf_sva_mut_10_6 <= base_buf_sva_mut_10_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_54_cse ) begin
      m_buf_sva_mut_6 <= m_buf_sva_mut_5;
      base_buf_sva_mut_6 <= base_buf_sva_mut_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_6 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_105 ) begin
      result_rem_11cyc_st_6 <= result_rem_11cyc_st_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_55_cse ) begin
      m_buf_sva_mut_1_5 <= m_buf_sva_mut_1_4;
      base_buf_sva_mut_1_5 <= base_buf_sva_mut_1_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_56_cse ) begin
      m_buf_sva_mut_2_5 <= m_buf_sva_mut_2_4;
      base_buf_sva_mut_2_5 <= base_buf_sva_mut_2_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_57_cse ) begin
      m_buf_sva_mut_3_5 <= m_buf_sva_mut_3_4;
      base_buf_sva_mut_3_5 <= base_buf_sva_mut_3_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_58_cse ) begin
      m_buf_sva_mut_4_5 <= m_buf_sva_mut_4_4;
      base_buf_sva_mut_4_5 <= base_buf_sva_mut_4_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_59_cse ) begin
      m_buf_sva_mut_5_5 <= m_buf_sva_mut_5_4;
      base_buf_sva_mut_5_5 <= base_buf_sva_mut_5_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_60_cse ) begin
      m_buf_sva_mut_6_5 <= m_buf_sva_mut_6_4;
      base_buf_sva_mut_6_5 <= base_buf_sva_mut_6_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_61_cse ) begin
      m_buf_sva_mut_7_5 <= m_buf_sva_mut_7_4;
      base_buf_sva_mut_7_5 <= base_buf_sva_mut_7_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_62_cse ) begin
      m_buf_sva_mut_8_5 <= m_buf_sva_mut_8_4;
      base_buf_sva_mut_8_5 <= base_buf_sva_mut_8_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_63_cse ) begin
      m_buf_sva_mut_9_5 <= m_buf_sva_mut_9_4;
      base_buf_sva_mut_9_5 <= base_buf_sva_mut_9_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_64_cse ) begin
      m_buf_sva_mut_10_5 <= m_buf_sva_mut_10_4;
      base_buf_sva_mut_10_5 <= base_buf_sva_mut_10_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_65_cse ) begin
      m_buf_sva_mut_5 <= m_buf_sva_mut_4;
      base_buf_sva_mut_5 <= base_buf_sva_mut_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_5 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_130 ) begin
      result_rem_11cyc_st_5 <= result_rem_11cyc_st_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_66_cse ) begin
      m_buf_sva_mut_1_4 <= m_buf_sva_mut_1_3;
      base_buf_sva_mut_1_4 <= base_buf_sva_mut_1_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_67_cse ) begin
      m_buf_sva_mut_2_4 <= m_buf_sva_mut_2_3;
      base_buf_sva_mut_2_4 <= base_buf_sva_mut_2_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_68_cse ) begin
      m_buf_sva_mut_3_4 <= m_buf_sva_mut_3_3;
      base_buf_sva_mut_3_4 <= base_buf_sva_mut_3_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_69_cse ) begin
      m_buf_sva_mut_4_4 <= m_buf_sva_mut_4_3;
      base_buf_sva_mut_4_4 <= base_buf_sva_mut_4_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_70_cse ) begin
      m_buf_sva_mut_5_4 <= m_buf_sva_mut_5_3;
      base_buf_sva_mut_5_4 <= base_buf_sva_mut_5_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_71_cse ) begin
      m_buf_sva_mut_6_4 <= m_buf_sva_mut_6_3;
      base_buf_sva_mut_6_4 <= base_buf_sva_mut_6_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_72_cse ) begin
      m_buf_sva_mut_7_4 <= m_buf_sva_mut_7_3;
      base_buf_sva_mut_7_4 <= base_buf_sva_mut_7_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_73_cse ) begin
      m_buf_sva_mut_8_4 <= m_buf_sva_mut_8_3;
      base_buf_sva_mut_8_4 <= base_buf_sva_mut_8_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_74_cse ) begin
      m_buf_sva_mut_9_4 <= m_buf_sva_mut_9_3;
      base_buf_sva_mut_9_4 <= base_buf_sva_mut_9_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_75_cse ) begin
      m_buf_sva_mut_10_4 <= m_buf_sva_mut_10_3;
      base_buf_sva_mut_10_4 <= base_buf_sva_mut_10_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_76_cse ) begin
      m_buf_sva_mut_4 <= m_buf_sva_mut_3;
      base_buf_sva_mut_4 <= base_buf_sva_mut_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_4 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_156 ) begin
      result_rem_11cyc_st_4 <= result_rem_11cyc_st_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_77_cse ) begin
      m_buf_sva_mut_1_3 <= m_buf_sva_mut_1_2;
      base_buf_sva_mut_1_3 <= base_buf_sva_mut_1_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_78_cse ) begin
      m_buf_sva_mut_2_3 <= m_buf_sva_mut_2_2;
      base_buf_sva_mut_2_3 <= base_buf_sva_mut_2_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_79_cse ) begin
      m_buf_sva_mut_3_3 <= m_buf_sva_mut_3_2;
      base_buf_sva_mut_3_3 <= base_buf_sva_mut_3_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_80_cse ) begin
      m_buf_sva_mut_4_3 <= m_buf_sva_mut_4_2;
      base_buf_sva_mut_4_3 <= base_buf_sva_mut_4_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_81_cse ) begin
      m_buf_sva_mut_5_3 <= m_buf_sva_mut_5_2;
      base_buf_sva_mut_5_3 <= base_buf_sva_mut_5_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_82_cse ) begin
      m_buf_sva_mut_6_3 <= m_buf_sva_mut_6_2;
      base_buf_sva_mut_6_3 <= base_buf_sva_mut_6_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_83_cse ) begin
      m_buf_sva_mut_7_3 <= m_buf_sva_mut_7_2;
      base_buf_sva_mut_7_3 <= base_buf_sva_mut_7_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_84_cse ) begin
      m_buf_sva_mut_8_3 <= m_buf_sva_mut_8_2;
      base_buf_sva_mut_8_3 <= base_buf_sva_mut_8_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_85_cse ) begin
      m_buf_sva_mut_9_3 <= m_buf_sva_mut_9_2;
      base_buf_sva_mut_9_3 <= base_buf_sva_mut_9_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_86_cse ) begin
      m_buf_sva_mut_10_3 <= m_buf_sva_mut_10_2;
      base_buf_sva_mut_10_3 <= base_buf_sva_mut_10_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_87_cse ) begin
      m_buf_sva_mut_3 <= m_buf_sva_mut_2;
      base_buf_sva_mut_3 <= base_buf_sva_mut_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_3 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_182 ) begin
      result_rem_11cyc_st_3 <= result_rem_11cyc_st_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_88_cse ) begin
      m_buf_sva_mut_1_2 <= result_rem_12_cmp_1_b;
      base_buf_sva_mut_1_2 <= result_rem_12_cmp_1_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_89_cse ) begin
      m_buf_sva_mut_2_2 <= result_rem_12_cmp_2_b;
      base_buf_sva_mut_2_2 <= result_rem_12_cmp_2_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_90_cse ) begin
      m_buf_sva_mut_3_2 <= result_rem_12_cmp_3_b;
      base_buf_sva_mut_3_2 <= result_rem_12_cmp_3_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_91_cse ) begin
      m_buf_sva_mut_4_2 <= result_rem_12_cmp_4_b;
      base_buf_sva_mut_4_2 <= result_rem_12_cmp_4_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_92_cse ) begin
      m_buf_sva_mut_5_2 <= result_rem_12_cmp_5_b;
      base_buf_sva_mut_5_2 <= result_rem_12_cmp_5_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_93_cse ) begin
      m_buf_sva_mut_6_2 <= result_rem_12_cmp_6_b;
      base_buf_sva_mut_6_2 <= result_rem_12_cmp_6_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_94_cse ) begin
      m_buf_sva_mut_7_2 <= result_rem_12_cmp_7_b;
      base_buf_sva_mut_7_2 <= result_rem_12_cmp_7_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_95_cse ) begin
      m_buf_sva_mut_8_2 <= result_rem_12_cmp_8_b;
      base_buf_sva_mut_8_2 <= result_rem_12_cmp_8_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_96_cse ) begin
      m_buf_sva_mut_9_2 <= result_rem_12_cmp_9_b;
      base_buf_sva_mut_9_2 <= result_rem_12_cmp_9_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_97_cse ) begin
      m_buf_sva_mut_10_2 <= result_rem_12_cmp_10_b;
      base_buf_sva_mut_10_2 <= result_rem_12_cmp_10_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_98_cse ) begin
      m_buf_sva_mut_2 <= result_rem_12_cmp_b;
      base_buf_sva_mut_2 <= result_rem_12_cmp_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_2 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_208 ) begin
      result_rem_11cyc_st_2 <= result_rem_11cyc;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc <= 4'b0000;
    end
    else if ( ccs_ccore_en & ccs_ccore_start_rsci_idat ) begin
      result_rem_11cyc <= result_result_acc_tmp;
    end
  end

  function automatic [63:0] MUX1HOT_v_64_10_2;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [9:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    MUX1HOT_v_64_10_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_11_2;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [10:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    MUX1HOT_v_64_11_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function automatic [3:0] conv_s2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_s2s_3_4 = {vector[2], vector};
  end
  endfunction


  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_2_4 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_4 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    modulo_dev
// ------------------------------------------------------------------


module modulo_dev (
  base_rsc_dat, m_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [63:0] base_rsc_dat;
  input [63:0] m_rsc_dat;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  modulo_dev_core modulo_dev_core_inst (
      .base_rsc_dat(base_rsc_dat),
      .m_rsc_dat(m_rsc_dat),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Thu Aug 26 04:29:45 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_72_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_72_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_71_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_71_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_70_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_70_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_69_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_69_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_68_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_68_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_67_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_67_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_66_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_66_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_65_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_65_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_64_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_64_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_63_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_63_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_62_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_62_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_61_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_61_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_60_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_60_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_59_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_59_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_58_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_58_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_57_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_57_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_56_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_56_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_55_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_55_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_54_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_54_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_53_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_53_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_52_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_52_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_51_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_51_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_50_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_50_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_49_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_49_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_48_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_48_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_47_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_47_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_46_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_46_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_45_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_45_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_44_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_44_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_43_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_43_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_42_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_42_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_41_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_41_5_64_32_32_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output [63:0] q_d;
  input [4:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_5_64_32_32_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_5_64_32_32_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [4:0] radr;
  output we;
  output [63:0] d;
  output [4:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [4:0] radr_d;
  input [4:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module inPlaceNTT_DIF_core_core_fsm (
  clk, rst, fsm_output, COMP_LOOP_C_28_tr0, COMP_LOOP_C_56_tr0, COMP_LOOP_C_84_tr0,
      COMP_LOOP_C_112_tr0, COMP_LOOP_C_140_tr0, COMP_LOOP_C_168_tr0, COMP_LOOP_C_196_tr0,
      COMP_LOOP_C_224_tr0, VEC_LOOP_C_0_tr0, STAGE_LOOP_C_1_tr0
);
  input clk;
  input rst;
  output [7:0] fsm_output;
  reg [7:0] fsm_output;
  input COMP_LOOP_C_28_tr0;
  input COMP_LOOP_C_56_tr0;
  input COMP_LOOP_C_84_tr0;
  input COMP_LOOP_C_112_tr0;
  input COMP_LOOP_C_140_tr0;
  input COMP_LOOP_C_168_tr0;
  input COMP_LOOP_C_196_tr0;
  input COMP_LOOP_C_224_tr0;
  input VEC_LOOP_C_0_tr0;
  input STAGE_LOOP_C_1_tr0;


  // FSM State Type Declaration for inPlaceNTT_DIF_core_core_fsm_1
  parameter
    main_C_0 = 8'd0,
    STAGE_LOOP_C_0 = 8'd1,
    COMP_LOOP_C_0 = 8'd2,
    COMP_LOOP_C_1 = 8'd3,
    COMP_LOOP_C_2 = 8'd4,
    COMP_LOOP_C_3 = 8'd5,
    COMP_LOOP_C_4 = 8'd6,
    COMP_LOOP_C_5 = 8'd7,
    COMP_LOOP_C_6 = 8'd8,
    COMP_LOOP_C_7 = 8'd9,
    COMP_LOOP_C_8 = 8'd10,
    COMP_LOOP_C_9 = 8'd11,
    COMP_LOOP_C_10 = 8'd12,
    COMP_LOOP_C_11 = 8'd13,
    COMP_LOOP_C_12 = 8'd14,
    COMP_LOOP_C_13 = 8'd15,
    COMP_LOOP_C_14 = 8'd16,
    COMP_LOOP_C_15 = 8'd17,
    COMP_LOOP_C_16 = 8'd18,
    COMP_LOOP_C_17 = 8'd19,
    COMP_LOOP_C_18 = 8'd20,
    COMP_LOOP_C_19 = 8'd21,
    COMP_LOOP_C_20 = 8'd22,
    COMP_LOOP_C_21 = 8'd23,
    COMP_LOOP_C_22 = 8'd24,
    COMP_LOOP_C_23 = 8'd25,
    COMP_LOOP_C_24 = 8'd26,
    COMP_LOOP_C_25 = 8'd27,
    COMP_LOOP_C_26 = 8'd28,
    COMP_LOOP_C_27 = 8'd29,
    COMP_LOOP_C_28 = 8'd30,
    COMP_LOOP_C_29 = 8'd31,
    COMP_LOOP_C_30 = 8'd32,
    COMP_LOOP_C_31 = 8'd33,
    COMP_LOOP_C_32 = 8'd34,
    COMP_LOOP_C_33 = 8'd35,
    COMP_LOOP_C_34 = 8'd36,
    COMP_LOOP_C_35 = 8'd37,
    COMP_LOOP_C_36 = 8'd38,
    COMP_LOOP_C_37 = 8'd39,
    COMP_LOOP_C_38 = 8'd40,
    COMP_LOOP_C_39 = 8'd41,
    COMP_LOOP_C_40 = 8'd42,
    COMP_LOOP_C_41 = 8'd43,
    COMP_LOOP_C_42 = 8'd44,
    COMP_LOOP_C_43 = 8'd45,
    COMP_LOOP_C_44 = 8'd46,
    COMP_LOOP_C_45 = 8'd47,
    COMP_LOOP_C_46 = 8'd48,
    COMP_LOOP_C_47 = 8'd49,
    COMP_LOOP_C_48 = 8'd50,
    COMP_LOOP_C_49 = 8'd51,
    COMP_LOOP_C_50 = 8'd52,
    COMP_LOOP_C_51 = 8'd53,
    COMP_LOOP_C_52 = 8'd54,
    COMP_LOOP_C_53 = 8'd55,
    COMP_LOOP_C_54 = 8'd56,
    COMP_LOOP_C_55 = 8'd57,
    COMP_LOOP_C_56 = 8'd58,
    COMP_LOOP_C_57 = 8'd59,
    COMP_LOOP_C_58 = 8'd60,
    COMP_LOOP_C_59 = 8'd61,
    COMP_LOOP_C_60 = 8'd62,
    COMP_LOOP_C_61 = 8'd63,
    COMP_LOOP_C_62 = 8'd64,
    COMP_LOOP_C_63 = 8'd65,
    COMP_LOOP_C_64 = 8'd66,
    COMP_LOOP_C_65 = 8'd67,
    COMP_LOOP_C_66 = 8'd68,
    COMP_LOOP_C_67 = 8'd69,
    COMP_LOOP_C_68 = 8'd70,
    COMP_LOOP_C_69 = 8'd71,
    COMP_LOOP_C_70 = 8'd72,
    COMP_LOOP_C_71 = 8'd73,
    COMP_LOOP_C_72 = 8'd74,
    COMP_LOOP_C_73 = 8'd75,
    COMP_LOOP_C_74 = 8'd76,
    COMP_LOOP_C_75 = 8'd77,
    COMP_LOOP_C_76 = 8'd78,
    COMP_LOOP_C_77 = 8'd79,
    COMP_LOOP_C_78 = 8'd80,
    COMP_LOOP_C_79 = 8'd81,
    COMP_LOOP_C_80 = 8'd82,
    COMP_LOOP_C_81 = 8'd83,
    COMP_LOOP_C_82 = 8'd84,
    COMP_LOOP_C_83 = 8'd85,
    COMP_LOOP_C_84 = 8'd86,
    COMP_LOOP_C_85 = 8'd87,
    COMP_LOOP_C_86 = 8'd88,
    COMP_LOOP_C_87 = 8'd89,
    COMP_LOOP_C_88 = 8'd90,
    COMP_LOOP_C_89 = 8'd91,
    COMP_LOOP_C_90 = 8'd92,
    COMP_LOOP_C_91 = 8'd93,
    COMP_LOOP_C_92 = 8'd94,
    COMP_LOOP_C_93 = 8'd95,
    COMP_LOOP_C_94 = 8'd96,
    COMP_LOOP_C_95 = 8'd97,
    COMP_LOOP_C_96 = 8'd98,
    COMP_LOOP_C_97 = 8'd99,
    COMP_LOOP_C_98 = 8'd100,
    COMP_LOOP_C_99 = 8'd101,
    COMP_LOOP_C_100 = 8'd102,
    COMP_LOOP_C_101 = 8'd103,
    COMP_LOOP_C_102 = 8'd104,
    COMP_LOOP_C_103 = 8'd105,
    COMP_LOOP_C_104 = 8'd106,
    COMP_LOOP_C_105 = 8'd107,
    COMP_LOOP_C_106 = 8'd108,
    COMP_LOOP_C_107 = 8'd109,
    COMP_LOOP_C_108 = 8'd110,
    COMP_LOOP_C_109 = 8'd111,
    COMP_LOOP_C_110 = 8'd112,
    COMP_LOOP_C_111 = 8'd113,
    COMP_LOOP_C_112 = 8'd114,
    COMP_LOOP_C_113 = 8'd115,
    COMP_LOOP_C_114 = 8'd116,
    COMP_LOOP_C_115 = 8'd117,
    COMP_LOOP_C_116 = 8'd118,
    COMP_LOOP_C_117 = 8'd119,
    COMP_LOOP_C_118 = 8'd120,
    COMP_LOOP_C_119 = 8'd121,
    COMP_LOOP_C_120 = 8'd122,
    COMP_LOOP_C_121 = 8'd123,
    COMP_LOOP_C_122 = 8'd124,
    COMP_LOOP_C_123 = 8'd125,
    COMP_LOOP_C_124 = 8'd126,
    COMP_LOOP_C_125 = 8'd127,
    COMP_LOOP_C_126 = 8'd128,
    COMP_LOOP_C_127 = 8'd129,
    COMP_LOOP_C_128 = 8'd130,
    COMP_LOOP_C_129 = 8'd131,
    COMP_LOOP_C_130 = 8'd132,
    COMP_LOOP_C_131 = 8'd133,
    COMP_LOOP_C_132 = 8'd134,
    COMP_LOOP_C_133 = 8'd135,
    COMP_LOOP_C_134 = 8'd136,
    COMP_LOOP_C_135 = 8'd137,
    COMP_LOOP_C_136 = 8'd138,
    COMP_LOOP_C_137 = 8'd139,
    COMP_LOOP_C_138 = 8'd140,
    COMP_LOOP_C_139 = 8'd141,
    COMP_LOOP_C_140 = 8'd142,
    COMP_LOOP_C_141 = 8'd143,
    COMP_LOOP_C_142 = 8'd144,
    COMP_LOOP_C_143 = 8'd145,
    COMP_LOOP_C_144 = 8'd146,
    COMP_LOOP_C_145 = 8'd147,
    COMP_LOOP_C_146 = 8'd148,
    COMP_LOOP_C_147 = 8'd149,
    COMP_LOOP_C_148 = 8'd150,
    COMP_LOOP_C_149 = 8'd151,
    COMP_LOOP_C_150 = 8'd152,
    COMP_LOOP_C_151 = 8'd153,
    COMP_LOOP_C_152 = 8'd154,
    COMP_LOOP_C_153 = 8'd155,
    COMP_LOOP_C_154 = 8'd156,
    COMP_LOOP_C_155 = 8'd157,
    COMP_LOOP_C_156 = 8'd158,
    COMP_LOOP_C_157 = 8'd159,
    COMP_LOOP_C_158 = 8'd160,
    COMP_LOOP_C_159 = 8'd161,
    COMP_LOOP_C_160 = 8'd162,
    COMP_LOOP_C_161 = 8'd163,
    COMP_LOOP_C_162 = 8'd164,
    COMP_LOOP_C_163 = 8'd165,
    COMP_LOOP_C_164 = 8'd166,
    COMP_LOOP_C_165 = 8'd167,
    COMP_LOOP_C_166 = 8'd168,
    COMP_LOOP_C_167 = 8'd169,
    COMP_LOOP_C_168 = 8'd170,
    COMP_LOOP_C_169 = 8'd171,
    COMP_LOOP_C_170 = 8'd172,
    COMP_LOOP_C_171 = 8'd173,
    COMP_LOOP_C_172 = 8'd174,
    COMP_LOOP_C_173 = 8'd175,
    COMP_LOOP_C_174 = 8'd176,
    COMP_LOOP_C_175 = 8'd177,
    COMP_LOOP_C_176 = 8'd178,
    COMP_LOOP_C_177 = 8'd179,
    COMP_LOOP_C_178 = 8'd180,
    COMP_LOOP_C_179 = 8'd181,
    COMP_LOOP_C_180 = 8'd182,
    COMP_LOOP_C_181 = 8'd183,
    COMP_LOOP_C_182 = 8'd184,
    COMP_LOOP_C_183 = 8'd185,
    COMP_LOOP_C_184 = 8'd186,
    COMP_LOOP_C_185 = 8'd187,
    COMP_LOOP_C_186 = 8'd188,
    COMP_LOOP_C_187 = 8'd189,
    COMP_LOOP_C_188 = 8'd190,
    COMP_LOOP_C_189 = 8'd191,
    COMP_LOOP_C_190 = 8'd192,
    COMP_LOOP_C_191 = 8'd193,
    COMP_LOOP_C_192 = 8'd194,
    COMP_LOOP_C_193 = 8'd195,
    COMP_LOOP_C_194 = 8'd196,
    COMP_LOOP_C_195 = 8'd197,
    COMP_LOOP_C_196 = 8'd198,
    COMP_LOOP_C_197 = 8'd199,
    COMP_LOOP_C_198 = 8'd200,
    COMP_LOOP_C_199 = 8'd201,
    COMP_LOOP_C_200 = 8'd202,
    COMP_LOOP_C_201 = 8'd203,
    COMP_LOOP_C_202 = 8'd204,
    COMP_LOOP_C_203 = 8'd205,
    COMP_LOOP_C_204 = 8'd206,
    COMP_LOOP_C_205 = 8'd207,
    COMP_LOOP_C_206 = 8'd208,
    COMP_LOOP_C_207 = 8'd209,
    COMP_LOOP_C_208 = 8'd210,
    COMP_LOOP_C_209 = 8'd211,
    COMP_LOOP_C_210 = 8'd212,
    COMP_LOOP_C_211 = 8'd213,
    COMP_LOOP_C_212 = 8'd214,
    COMP_LOOP_C_213 = 8'd215,
    COMP_LOOP_C_214 = 8'd216,
    COMP_LOOP_C_215 = 8'd217,
    COMP_LOOP_C_216 = 8'd218,
    COMP_LOOP_C_217 = 8'd219,
    COMP_LOOP_C_218 = 8'd220,
    COMP_LOOP_C_219 = 8'd221,
    COMP_LOOP_C_220 = 8'd222,
    COMP_LOOP_C_221 = 8'd223,
    COMP_LOOP_C_222 = 8'd224,
    COMP_LOOP_C_223 = 8'd225,
    COMP_LOOP_C_224 = 8'd226,
    VEC_LOOP_C_0 = 8'd227,
    STAGE_LOOP_C_1 = 8'd228,
    main_C_1 = 8'd229;

  reg [7:0] state_var;
  reg [7:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : inPlaceNTT_DIF_core_core_fsm_1
    case (state_var)
      STAGE_LOOP_C_0 : begin
        fsm_output = 8'b00000001;
        state_var_NS = COMP_LOOP_C_0;
      end
      COMP_LOOP_C_0 : begin
        fsm_output = 8'b00000010;
        state_var_NS = COMP_LOOP_C_1;
      end
      COMP_LOOP_C_1 : begin
        fsm_output = 8'b00000011;
        state_var_NS = COMP_LOOP_C_2;
      end
      COMP_LOOP_C_2 : begin
        fsm_output = 8'b00000100;
        state_var_NS = COMP_LOOP_C_3;
      end
      COMP_LOOP_C_3 : begin
        fsm_output = 8'b00000101;
        state_var_NS = COMP_LOOP_C_4;
      end
      COMP_LOOP_C_4 : begin
        fsm_output = 8'b00000110;
        state_var_NS = COMP_LOOP_C_5;
      end
      COMP_LOOP_C_5 : begin
        fsm_output = 8'b00000111;
        state_var_NS = COMP_LOOP_C_6;
      end
      COMP_LOOP_C_6 : begin
        fsm_output = 8'b00001000;
        state_var_NS = COMP_LOOP_C_7;
      end
      COMP_LOOP_C_7 : begin
        fsm_output = 8'b00001001;
        state_var_NS = COMP_LOOP_C_8;
      end
      COMP_LOOP_C_8 : begin
        fsm_output = 8'b00001010;
        state_var_NS = COMP_LOOP_C_9;
      end
      COMP_LOOP_C_9 : begin
        fsm_output = 8'b00001011;
        state_var_NS = COMP_LOOP_C_10;
      end
      COMP_LOOP_C_10 : begin
        fsm_output = 8'b00001100;
        state_var_NS = COMP_LOOP_C_11;
      end
      COMP_LOOP_C_11 : begin
        fsm_output = 8'b00001101;
        state_var_NS = COMP_LOOP_C_12;
      end
      COMP_LOOP_C_12 : begin
        fsm_output = 8'b00001110;
        state_var_NS = COMP_LOOP_C_13;
      end
      COMP_LOOP_C_13 : begin
        fsm_output = 8'b00001111;
        state_var_NS = COMP_LOOP_C_14;
      end
      COMP_LOOP_C_14 : begin
        fsm_output = 8'b00010000;
        state_var_NS = COMP_LOOP_C_15;
      end
      COMP_LOOP_C_15 : begin
        fsm_output = 8'b00010001;
        state_var_NS = COMP_LOOP_C_16;
      end
      COMP_LOOP_C_16 : begin
        fsm_output = 8'b00010010;
        state_var_NS = COMP_LOOP_C_17;
      end
      COMP_LOOP_C_17 : begin
        fsm_output = 8'b00010011;
        state_var_NS = COMP_LOOP_C_18;
      end
      COMP_LOOP_C_18 : begin
        fsm_output = 8'b00010100;
        state_var_NS = COMP_LOOP_C_19;
      end
      COMP_LOOP_C_19 : begin
        fsm_output = 8'b00010101;
        state_var_NS = COMP_LOOP_C_20;
      end
      COMP_LOOP_C_20 : begin
        fsm_output = 8'b00010110;
        state_var_NS = COMP_LOOP_C_21;
      end
      COMP_LOOP_C_21 : begin
        fsm_output = 8'b00010111;
        state_var_NS = COMP_LOOP_C_22;
      end
      COMP_LOOP_C_22 : begin
        fsm_output = 8'b00011000;
        state_var_NS = COMP_LOOP_C_23;
      end
      COMP_LOOP_C_23 : begin
        fsm_output = 8'b00011001;
        state_var_NS = COMP_LOOP_C_24;
      end
      COMP_LOOP_C_24 : begin
        fsm_output = 8'b00011010;
        state_var_NS = COMP_LOOP_C_25;
      end
      COMP_LOOP_C_25 : begin
        fsm_output = 8'b00011011;
        state_var_NS = COMP_LOOP_C_26;
      end
      COMP_LOOP_C_26 : begin
        fsm_output = 8'b00011100;
        state_var_NS = COMP_LOOP_C_27;
      end
      COMP_LOOP_C_27 : begin
        fsm_output = 8'b00011101;
        state_var_NS = COMP_LOOP_C_28;
      end
      COMP_LOOP_C_28 : begin
        fsm_output = 8'b00011110;
        if ( COMP_LOOP_C_28_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_29;
        end
      end
      COMP_LOOP_C_29 : begin
        fsm_output = 8'b00011111;
        state_var_NS = COMP_LOOP_C_30;
      end
      COMP_LOOP_C_30 : begin
        fsm_output = 8'b00100000;
        state_var_NS = COMP_LOOP_C_31;
      end
      COMP_LOOP_C_31 : begin
        fsm_output = 8'b00100001;
        state_var_NS = COMP_LOOP_C_32;
      end
      COMP_LOOP_C_32 : begin
        fsm_output = 8'b00100010;
        state_var_NS = COMP_LOOP_C_33;
      end
      COMP_LOOP_C_33 : begin
        fsm_output = 8'b00100011;
        state_var_NS = COMP_LOOP_C_34;
      end
      COMP_LOOP_C_34 : begin
        fsm_output = 8'b00100100;
        state_var_NS = COMP_LOOP_C_35;
      end
      COMP_LOOP_C_35 : begin
        fsm_output = 8'b00100101;
        state_var_NS = COMP_LOOP_C_36;
      end
      COMP_LOOP_C_36 : begin
        fsm_output = 8'b00100110;
        state_var_NS = COMP_LOOP_C_37;
      end
      COMP_LOOP_C_37 : begin
        fsm_output = 8'b00100111;
        state_var_NS = COMP_LOOP_C_38;
      end
      COMP_LOOP_C_38 : begin
        fsm_output = 8'b00101000;
        state_var_NS = COMP_LOOP_C_39;
      end
      COMP_LOOP_C_39 : begin
        fsm_output = 8'b00101001;
        state_var_NS = COMP_LOOP_C_40;
      end
      COMP_LOOP_C_40 : begin
        fsm_output = 8'b00101010;
        state_var_NS = COMP_LOOP_C_41;
      end
      COMP_LOOP_C_41 : begin
        fsm_output = 8'b00101011;
        state_var_NS = COMP_LOOP_C_42;
      end
      COMP_LOOP_C_42 : begin
        fsm_output = 8'b00101100;
        state_var_NS = COMP_LOOP_C_43;
      end
      COMP_LOOP_C_43 : begin
        fsm_output = 8'b00101101;
        state_var_NS = COMP_LOOP_C_44;
      end
      COMP_LOOP_C_44 : begin
        fsm_output = 8'b00101110;
        state_var_NS = COMP_LOOP_C_45;
      end
      COMP_LOOP_C_45 : begin
        fsm_output = 8'b00101111;
        state_var_NS = COMP_LOOP_C_46;
      end
      COMP_LOOP_C_46 : begin
        fsm_output = 8'b00110000;
        state_var_NS = COMP_LOOP_C_47;
      end
      COMP_LOOP_C_47 : begin
        fsm_output = 8'b00110001;
        state_var_NS = COMP_LOOP_C_48;
      end
      COMP_LOOP_C_48 : begin
        fsm_output = 8'b00110010;
        state_var_NS = COMP_LOOP_C_49;
      end
      COMP_LOOP_C_49 : begin
        fsm_output = 8'b00110011;
        state_var_NS = COMP_LOOP_C_50;
      end
      COMP_LOOP_C_50 : begin
        fsm_output = 8'b00110100;
        state_var_NS = COMP_LOOP_C_51;
      end
      COMP_LOOP_C_51 : begin
        fsm_output = 8'b00110101;
        state_var_NS = COMP_LOOP_C_52;
      end
      COMP_LOOP_C_52 : begin
        fsm_output = 8'b00110110;
        state_var_NS = COMP_LOOP_C_53;
      end
      COMP_LOOP_C_53 : begin
        fsm_output = 8'b00110111;
        state_var_NS = COMP_LOOP_C_54;
      end
      COMP_LOOP_C_54 : begin
        fsm_output = 8'b00111000;
        state_var_NS = COMP_LOOP_C_55;
      end
      COMP_LOOP_C_55 : begin
        fsm_output = 8'b00111001;
        state_var_NS = COMP_LOOP_C_56;
      end
      COMP_LOOP_C_56 : begin
        fsm_output = 8'b00111010;
        if ( COMP_LOOP_C_56_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_57;
        end
      end
      COMP_LOOP_C_57 : begin
        fsm_output = 8'b00111011;
        state_var_NS = COMP_LOOP_C_58;
      end
      COMP_LOOP_C_58 : begin
        fsm_output = 8'b00111100;
        state_var_NS = COMP_LOOP_C_59;
      end
      COMP_LOOP_C_59 : begin
        fsm_output = 8'b00111101;
        state_var_NS = COMP_LOOP_C_60;
      end
      COMP_LOOP_C_60 : begin
        fsm_output = 8'b00111110;
        state_var_NS = COMP_LOOP_C_61;
      end
      COMP_LOOP_C_61 : begin
        fsm_output = 8'b00111111;
        state_var_NS = COMP_LOOP_C_62;
      end
      COMP_LOOP_C_62 : begin
        fsm_output = 8'b01000000;
        state_var_NS = COMP_LOOP_C_63;
      end
      COMP_LOOP_C_63 : begin
        fsm_output = 8'b01000001;
        state_var_NS = COMP_LOOP_C_64;
      end
      COMP_LOOP_C_64 : begin
        fsm_output = 8'b01000010;
        state_var_NS = COMP_LOOP_C_65;
      end
      COMP_LOOP_C_65 : begin
        fsm_output = 8'b01000011;
        state_var_NS = COMP_LOOP_C_66;
      end
      COMP_LOOP_C_66 : begin
        fsm_output = 8'b01000100;
        state_var_NS = COMP_LOOP_C_67;
      end
      COMP_LOOP_C_67 : begin
        fsm_output = 8'b01000101;
        state_var_NS = COMP_LOOP_C_68;
      end
      COMP_LOOP_C_68 : begin
        fsm_output = 8'b01000110;
        state_var_NS = COMP_LOOP_C_69;
      end
      COMP_LOOP_C_69 : begin
        fsm_output = 8'b01000111;
        state_var_NS = COMP_LOOP_C_70;
      end
      COMP_LOOP_C_70 : begin
        fsm_output = 8'b01001000;
        state_var_NS = COMP_LOOP_C_71;
      end
      COMP_LOOP_C_71 : begin
        fsm_output = 8'b01001001;
        state_var_NS = COMP_LOOP_C_72;
      end
      COMP_LOOP_C_72 : begin
        fsm_output = 8'b01001010;
        state_var_NS = COMP_LOOP_C_73;
      end
      COMP_LOOP_C_73 : begin
        fsm_output = 8'b01001011;
        state_var_NS = COMP_LOOP_C_74;
      end
      COMP_LOOP_C_74 : begin
        fsm_output = 8'b01001100;
        state_var_NS = COMP_LOOP_C_75;
      end
      COMP_LOOP_C_75 : begin
        fsm_output = 8'b01001101;
        state_var_NS = COMP_LOOP_C_76;
      end
      COMP_LOOP_C_76 : begin
        fsm_output = 8'b01001110;
        state_var_NS = COMP_LOOP_C_77;
      end
      COMP_LOOP_C_77 : begin
        fsm_output = 8'b01001111;
        state_var_NS = COMP_LOOP_C_78;
      end
      COMP_LOOP_C_78 : begin
        fsm_output = 8'b01010000;
        state_var_NS = COMP_LOOP_C_79;
      end
      COMP_LOOP_C_79 : begin
        fsm_output = 8'b01010001;
        state_var_NS = COMP_LOOP_C_80;
      end
      COMP_LOOP_C_80 : begin
        fsm_output = 8'b01010010;
        state_var_NS = COMP_LOOP_C_81;
      end
      COMP_LOOP_C_81 : begin
        fsm_output = 8'b01010011;
        state_var_NS = COMP_LOOP_C_82;
      end
      COMP_LOOP_C_82 : begin
        fsm_output = 8'b01010100;
        state_var_NS = COMP_LOOP_C_83;
      end
      COMP_LOOP_C_83 : begin
        fsm_output = 8'b01010101;
        state_var_NS = COMP_LOOP_C_84;
      end
      COMP_LOOP_C_84 : begin
        fsm_output = 8'b01010110;
        if ( COMP_LOOP_C_84_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_85;
        end
      end
      COMP_LOOP_C_85 : begin
        fsm_output = 8'b01010111;
        state_var_NS = COMP_LOOP_C_86;
      end
      COMP_LOOP_C_86 : begin
        fsm_output = 8'b01011000;
        state_var_NS = COMP_LOOP_C_87;
      end
      COMP_LOOP_C_87 : begin
        fsm_output = 8'b01011001;
        state_var_NS = COMP_LOOP_C_88;
      end
      COMP_LOOP_C_88 : begin
        fsm_output = 8'b01011010;
        state_var_NS = COMP_LOOP_C_89;
      end
      COMP_LOOP_C_89 : begin
        fsm_output = 8'b01011011;
        state_var_NS = COMP_LOOP_C_90;
      end
      COMP_LOOP_C_90 : begin
        fsm_output = 8'b01011100;
        state_var_NS = COMP_LOOP_C_91;
      end
      COMP_LOOP_C_91 : begin
        fsm_output = 8'b01011101;
        state_var_NS = COMP_LOOP_C_92;
      end
      COMP_LOOP_C_92 : begin
        fsm_output = 8'b01011110;
        state_var_NS = COMP_LOOP_C_93;
      end
      COMP_LOOP_C_93 : begin
        fsm_output = 8'b01011111;
        state_var_NS = COMP_LOOP_C_94;
      end
      COMP_LOOP_C_94 : begin
        fsm_output = 8'b01100000;
        state_var_NS = COMP_LOOP_C_95;
      end
      COMP_LOOP_C_95 : begin
        fsm_output = 8'b01100001;
        state_var_NS = COMP_LOOP_C_96;
      end
      COMP_LOOP_C_96 : begin
        fsm_output = 8'b01100010;
        state_var_NS = COMP_LOOP_C_97;
      end
      COMP_LOOP_C_97 : begin
        fsm_output = 8'b01100011;
        state_var_NS = COMP_LOOP_C_98;
      end
      COMP_LOOP_C_98 : begin
        fsm_output = 8'b01100100;
        state_var_NS = COMP_LOOP_C_99;
      end
      COMP_LOOP_C_99 : begin
        fsm_output = 8'b01100101;
        state_var_NS = COMP_LOOP_C_100;
      end
      COMP_LOOP_C_100 : begin
        fsm_output = 8'b01100110;
        state_var_NS = COMP_LOOP_C_101;
      end
      COMP_LOOP_C_101 : begin
        fsm_output = 8'b01100111;
        state_var_NS = COMP_LOOP_C_102;
      end
      COMP_LOOP_C_102 : begin
        fsm_output = 8'b01101000;
        state_var_NS = COMP_LOOP_C_103;
      end
      COMP_LOOP_C_103 : begin
        fsm_output = 8'b01101001;
        state_var_NS = COMP_LOOP_C_104;
      end
      COMP_LOOP_C_104 : begin
        fsm_output = 8'b01101010;
        state_var_NS = COMP_LOOP_C_105;
      end
      COMP_LOOP_C_105 : begin
        fsm_output = 8'b01101011;
        state_var_NS = COMP_LOOP_C_106;
      end
      COMP_LOOP_C_106 : begin
        fsm_output = 8'b01101100;
        state_var_NS = COMP_LOOP_C_107;
      end
      COMP_LOOP_C_107 : begin
        fsm_output = 8'b01101101;
        state_var_NS = COMP_LOOP_C_108;
      end
      COMP_LOOP_C_108 : begin
        fsm_output = 8'b01101110;
        state_var_NS = COMP_LOOP_C_109;
      end
      COMP_LOOP_C_109 : begin
        fsm_output = 8'b01101111;
        state_var_NS = COMP_LOOP_C_110;
      end
      COMP_LOOP_C_110 : begin
        fsm_output = 8'b01110000;
        state_var_NS = COMP_LOOP_C_111;
      end
      COMP_LOOP_C_111 : begin
        fsm_output = 8'b01110001;
        state_var_NS = COMP_LOOP_C_112;
      end
      COMP_LOOP_C_112 : begin
        fsm_output = 8'b01110010;
        if ( COMP_LOOP_C_112_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_113;
        end
      end
      COMP_LOOP_C_113 : begin
        fsm_output = 8'b01110011;
        state_var_NS = COMP_LOOP_C_114;
      end
      COMP_LOOP_C_114 : begin
        fsm_output = 8'b01110100;
        state_var_NS = COMP_LOOP_C_115;
      end
      COMP_LOOP_C_115 : begin
        fsm_output = 8'b01110101;
        state_var_NS = COMP_LOOP_C_116;
      end
      COMP_LOOP_C_116 : begin
        fsm_output = 8'b01110110;
        state_var_NS = COMP_LOOP_C_117;
      end
      COMP_LOOP_C_117 : begin
        fsm_output = 8'b01110111;
        state_var_NS = COMP_LOOP_C_118;
      end
      COMP_LOOP_C_118 : begin
        fsm_output = 8'b01111000;
        state_var_NS = COMP_LOOP_C_119;
      end
      COMP_LOOP_C_119 : begin
        fsm_output = 8'b01111001;
        state_var_NS = COMP_LOOP_C_120;
      end
      COMP_LOOP_C_120 : begin
        fsm_output = 8'b01111010;
        state_var_NS = COMP_LOOP_C_121;
      end
      COMP_LOOP_C_121 : begin
        fsm_output = 8'b01111011;
        state_var_NS = COMP_LOOP_C_122;
      end
      COMP_LOOP_C_122 : begin
        fsm_output = 8'b01111100;
        state_var_NS = COMP_LOOP_C_123;
      end
      COMP_LOOP_C_123 : begin
        fsm_output = 8'b01111101;
        state_var_NS = COMP_LOOP_C_124;
      end
      COMP_LOOP_C_124 : begin
        fsm_output = 8'b01111110;
        state_var_NS = COMP_LOOP_C_125;
      end
      COMP_LOOP_C_125 : begin
        fsm_output = 8'b01111111;
        state_var_NS = COMP_LOOP_C_126;
      end
      COMP_LOOP_C_126 : begin
        fsm_output = 8'b10000000;
        state_var_NS = COMP_LOOP_C_127;
      end
      COMP_LOOP_C_127 : begin
        fsm_output = 8'b10000001;
        state_var_NS = COMP_LOOP_C_128;
      end
      COMP_LOOP_C_128 : begin
        fsm_output = 8'b10000010;
        state_var_NS = COMP_LOOP_C_129;
      end
      COMP_LOOP_C_129 : begin
        fsm_output = 8'b10000011;
        state_var_NS = COMP_LOOP_C_130;
      end
      COMP_LOOP_C_130 : begin
        fsm_output = 8'b10000100;
        state_var_NS = COMP_LOOP_C_131;
      end
      COMP_LOOP_C_131 : begin
        fsm_output = 8'b10000101;
        state_var_NS = COMP_LOOP_C_132;
      end
      COMP_LOOP_C_132 : begin
        fsm_output = 8'b10000110;
        state_var_NS = COMP_LOOP_C_133;
      end
      COMP_LOOP_C_133 : begin
        fsm_output = 8'b10000111;
        state_var_NS = COMP_LOOP_C_134;
      end
      COMP_LOOP_C_134 : begin
        fsm_output = 8'b10001000;
        state_var_NS = COMP_LOOP_C_135;
      end
      COMP_LOOP_C_135 : begin
        fsm_output = 8'b10001001;
        state_var_NS = COMP_LOOP_C_136;
      end
      COMP_LOOP_C_136 : begin
        fsm_output = 8'b10001010;
        state_var_NS = COMP_LOOP_C_137;
      end
      COMP_LOOP_C_137 : begin
        fsm_output = 8'b10001011;
        state_var_NS = COMP_LOOP_C_138;
      end
      COMP_LOOP_C_138 : begin
        fsm_output = 8'b10001100;
        state_var_NS = COMP_LOOP_C_139;
      end
      COMP_LOOP_C_139 : begin
        fsm_output = 8'b10001101;
        state_var_NS = COMP_LOOP_C_140;
      end
      COMP_LOOP_C_140 : begin
        fsm_output = 8'b10001110;
        if ( COMP_LOOP_C_140_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_141;
        end
      end
      COMP_LOOP_C_141 : begin
        fsm_output = 8'b10001111;
        state_var_NS = COMP_LOOP_C_142;
      end
      COMP_LOOP_C_142 : begin
        fsm_output = 8'b10010000;
        state_var_NS = COMP_LOOP_C_143;
      end
      COMP_LOOP_C_143 : begin
        fsm_output = 8'b10010001;
        state_var_NS = COMP_LOOP_C_144;
      end
      COMP_LOOP_C_144 : begin
        fsm_output = 8'b10010010;
        state_var_NS = COMP_LOOP_C_145;
      end
      COMP_LOOP_C_145 : begin
        fsm_output = 8'b10010011;
        state_var_NS = COMP_LOOP_C_146;
      end
      COMP_LOOP_C_146 : begin
        fsm_output = 8'b10010100;
        state_var_NS = COMP_LOOP_C_147;
      end
      COMP_LOOP_C_147 : begin
        fsm_output = 8'b10010101;
        state_var_NS = COMP_LOOP_C_148;
      end
      COMP_LOOP_C_148 : begin
        fsm_output = 8'b10010110;
        state_var_NS = COMP_LOOP_C_149;
      end
      COMP_LOOP_C_149 : begin
        fsm_output = 8'b10010111;
        state_var_NS = COMP_LOOP_C_150;
      end
      COMP_LOOP_C_150 : begin
        fsm_output = 8'b10011000;
        state_var_NS = COMP_LOOP_C_151;
      end
      COMP_LOOP_C_151 : begin
        fsm_output = 8'b10011001;
        state_var_NS = COMP_LOOP_C_152;
      end
      COMP_LOOP_C_152 : begin
        fsm_output = 8'b10011010;
        state_var_NS = COMP_LOOP_C_153;
      end
      COMP_LOOP_C_153 : begin
        fsm_output = 8'b10011011;
        state_var_NS = COMP_LOOP_C_154;
      end
      COMP_LOOP_C_154 : begin
        fsm_output = 8'b10011100;
        state_var_NS = COMP_LOOP_C_155;
      end
      COMP_LOOP_C_155 : begin
        fsm_output = 8'b10011101;
        state_var_NS = COMP_LOOP_C_156;
      end
      COMP_LOOP_C_156 : begin
        fsm_output = 8'b10011110;
        state_var_NS = COMP_LOOP_C_157;
      end
      COMP_LOOP_C_157 : begin
        fsm_output = 8'b10011111;
        state_var_NS = COMP_LOOP_C_158;
      end
      COMP_LOOP_C_158 : begin
        fsm_output = 8'b10100000;
        state_var_NS = COMP_LOOP_C_159;
      end
      COMP_LOOP_C_159 : begin
        fsm_output = 8'b10100001;
        state_var_NS = COMP_LOOP_C_160;
      end
      COMP_LOOP_C_160 : begin
        fsm_output = 8'b10100010;
        state_var_NS = COMP_LOOP_C_161;
      end
      COMP_LOOP_C_161 : begin
        fsm_output = 8'b10100011;
        state_var_NS = COMP_LOOP_C_162;
      end
      COMP_LOOP_C_162 : begin
        fsm_output = 8'b10100100;
        state_var_NS = COMP_LOOP_C_163;
      end
      COMP_LOOP_C_163 : begin
        fsm_output = 8'b10100101;
        state_var_NS = COMP_LOOP_C_164;
      end
      COMP_LOOP_C_164 : begin
        fsm_output = 8'b10100110;
        state_var_NS = COMP_LOOP_C_165;
      end
      COMP_LOOP_C_165 : begin
        fsm_output = 8'b10100111;
        state_var_NS = COMP_LOOP_C_166;
      end
      COMP_LOOP_C_166 : begin
        fsm_output = 8'b10101000;
        state_var_NS = COMP_LOOP_C_167;
      end
      COMP_LOOP_C_167 : begin
        fsm_output = 8'b10101001;
        state_var_NS = COMP_LOOP_C_168;
      end
      COMP_LOOP_C_168 : begin
        fsm_output = 8'b10101010;
        if ( COMP_LOOP_C_168_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_169;
        end
      end
      COMP_LOOP_C_169 : begin
        fsm_output = 8'b10101011;
        state_var_NS = COMP_LOOP_C_170;
      end
      COMP_LOOP_C_170 : begin
        fsm_output = 8'b10101100;
        state_var_NS = COMP_LOOP_C_171;
      end
      COMP_LOOP_C_171 : begin
        fsm_output = 8'b10101101;
        state_var_NS = COMP_LOOP_C_172;
      end
      COMP_LOOP_C_172 : begin
        fsm_output = 8'b10101110;
        state_var_NS = COMP_LOOP_C_173;
      end
      COMP_LOOP_C_173 : begin
        fsm_output = 8'b10101111;
        state_var_NS = COMP_LOOP_C_174;
      end
      COMP_LOOP_C_174 : begin
        fsm_output = 8'b10110000;
        state_var_NS = COMP_LOOP_C_175;
      end
      COMP_LOOP_C_175 : begin
        fsm_output = 8'b10110001;
        state_var_NS = COMP_LOOP_C_176;
      end
      COMP_LOOP_C_176 : begin
        fsm_output = 8'b10110010;
        state_var_NS = COMP_LOOP_C_177;
      end
      COMP_LOOP_C_177 : begin
        fsm_output = 8'b10110011;
        state_var_NS = COMP_LOOP_C_178;
      end
      COMP_LOOP_C_178 : begin
        fsm_output = 8'b10110100;
        state_var_NS = COMP_LOOP_C_179;
      end
      COMP_LOOP_C_179 : begin
        fsm_output = 8'b10110101;
        state_var_NS = COMP_LOOP_C_180;
      end
      COMP_LOOP_C_180 : begin
        fsm_output = 8'b10110110;
        state_var_NS = COMP_LOOP_C_181;
      end
      COMP_LOOP_C_181 : begin
        fsm_output = 8'b10110111;
        state_var_NS = COMP_LOOP_C_182;
      end
      COMP_LOOP_C_182 : begin
        fsm_output = 8'b10111000;
        state_var_NS = COMP_LOOP_C_183;
      end
      COMP_LOOP_C_183 : begin
        fsm_output = 8'b10111001;
        state_var_NS = COMP_LOOP_C_184;
      end
      COMP_LOOP_C_184 : begin
        fsm_output = 8'b10111010;
        state_var_NS = COMP_LOOP_C_185;
      end
      COMP_LOOP_C_185 : begin
        fsm_output = 8'b10111011;
        state_var_NS = COMP_LOOP_C_186;
      end
      COMP_LOOP_C_186 : begin
        fsm_output = 8'b10111100;
        state_var_NS = COMP_LOOP_C_187;
      end
      COMP_LOOP_C_187 : begin
        fsm_output = 8'b10111101;
        state_var_NS = COMP_LOOP_C_188;
      end
      COMP_LOOP_C_188 : begin
        fsm_output = 8'b10111110;
        state_var_NS = COMP_LOOP_C_189;
      end
      COMP_LOOP_C_189 : begin
        fsm_output = 8'b10111111;
        state_var_NS = COMP_LOOP_C_190;
      end
      COMP_LOOP_C_190 : begin
        fsm_output = 8'b11000000;
        state_var_NS = COMP_LOOP_C_191;
      end
      COMP_LOOP_C_191 : begin
        fsm_output = 8'b11000001;
        state_var_NS = COMP_LOOP_C_192;
      end
      COMP_LOOP_C_192 : begin
        fsm_output = 8'b11000010;
        state_var_NS = COMP_LOOP_C_193;
      end
      COMP_LOOP_C_193 : begin
        fsm_output = 8'b11000011;
        state_var_NS = COMP_LOOP_C_194;
      end
      COMP_LOOP_C_194 : begin
        fsm_output = 8'b11000100;
        state_var_NS = COMP_LOOP_C_195;
      end
      COMP_LOOP_C_195 : begin
        fsm_output = 8'b11000101;
        state_var_NS = COMP_LOOP_C_196;
      end
      COMP_LOOP_C_196 : begin
        fsm_output = 8'b11000110;
        if ( COMP_LOOP_C_196_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_197;
        end
      end
      COMP_LOOP_C_197 : begin
        fsm_output = 8'b11000111;
        state_var_NS = COMP_LOOP_C_198;
      end
      COMP_LOOP_C_198 : begin
        fsm_output = 8'b11001000;
        state_var_NS = COMP_LOOP_C_199;
      end
      COMP_LOOP_C_199 : begin
        fsm_output = 8'b11001001;
        state_var_NS = COMP_LOOP_C_200;
      end
      COMP_LOOP_C_200 : begin
        fsm_output = 8'b11001010;
        state_var_NS = COMP_LOOP_C_201;
      end
      COMP_LOOP_C_201 : begin
        fsm_output = 8'b11001011;
        state_var_NS = COMP_LOOP_C_202;
      end
      COMP_LOOP_C_202 : begin
        fsm_output = 8'b11001100;
        state_var_NS = COMP_LOOP_C_203;
      end
      COMP_LOOP_C_203 : begin
        fsm_output = 8'b11001101;
        state_var_NS = COMP_LOOP_C_204;
      end
      COMP_LOOP_C_204 : begin
        fsm_output = 8'b11001110;
        state_var_NS = COMP_LOOP_C_205;
      end
      COMP_LOOP_C_205 : begin
        fsm_output = 8'b11001111;
        state_var_NS = COMP_LOOP_C_206;
      end
      COMP_LOOP_C_206 : begin
        fsm_output = 8'b11010000;
        state_var_NS = COMP_LOOP_C_207;
      end
      COMP_LOOP_C_207 : begin
        fsm_output = 8'b11010001;
        state_var_NS = COMP_LOOP_C_208;
      end
      COMP_LOOP_C_208 : begin
        fsm_output = 8'b11010010;
        state_var_NS = COMP_LOOP_C_209;
      end
      COMP_LOOP_C_209 : begin
        fsm_output = 8'b11010011;
        state_var_NS = COMP_LOOP_C_210;
      end
      COMP_LOOP_C_210 : begin
        fsm_output = 8'b11010100;
        state_var_NS = COMP_LOOP_C_211;
      end
      COMP_LOOP_C_211 : begin
        fsm_output = 8'b11010101;
        state_var_NS = COMP_LOOP_C_212;
      end
      COMP_LOOP_C_212 : begin
        fsm_output = 8'b11010110;
        state_var_NS = COMP_LOOP_C_213;
      end
      COMP_LOOP_C_213 : begin
        fsm_output = 8'b11010111;
        state_var_NS = COMP_LOOP_C_214;
      end
      COMP_LOOP_C_214 : begin
        fsm_output = 8'b11011000;
        state_var_NS = COMP_LOOP_C_215;
      end
      COMP_LOOP_C_215 : begin
        fsm_output = 8'b11011001;
        state_var_NS = COMP_LOOP_C_216;
      end
      COMP_LOOP_C_216 : begin
        fsm_output = 8'b11011010;
        state_var_NS = COMP_LOOP_C_217;
      end
      COMP_LOOP_C_217 : begin
        fsm_output = 8'b11011011;
        state_var_NS = COMP_LOOP_C_218;
      end
      COMP_LOOP_C_218 : begin
        fsm_output = 8'b11011100;
        state_var_NS = COMP_LOOP_C_219;
      end
      COMP_LOOP_C_219 : begin
        fsm_output = 8'b11011101;
        state_var_NS = COMP_LOOP_C_220;
      end
      COMP_LOOP_C_220 : begin
        fsm_output = 8'b11011110;
        state_var_NS = COMP_LOOP_C_221;
      end
      COMP_LOOP_C_221 : begin
        fsm_output = 8'b11011111;
        state_var_NS = COMP_LOOP_C_222;
      end
      COMP_LOOP_C_222 : begin
        fsm_output = 8'b11100000;
        state_var_NS = COMP_LOOP_C_223;
      end
      COMP_LOOP_C_223 : begin
        fsm_output = 8'b11100001;
        state_var_NS = COMP_LOOP_C_224;
      end
      COMP_LOOP_C_224 : begin
        fsm_output = 8'b11100010;
        if ( COMP_LOOP_C_224_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_C_0 : begin
        fsm_output = 8'b11100011;
        if ( VEC_LOOP_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      STAGE_LOOP_C_1 : begin
        fsm_output = 8'b11100100;
        if ( STAGE_LOOP_C_1_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = STAGE_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 8'b11100101;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 8'b00000000;
        state_var_NS = STAGE_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_core_wait_dp
// ------------------------------------------------------------------


module inPlaceNTT_DIF_core_wait_dp (
  ensig_cgo_iro, ensig_cgo, COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en
);
  input ensig_cgo_iro;
  input ensig_cgo;
  output COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  assign COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en = ensig_cgo | ensig_cgo_iro;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_core
// ------------------------------------------------------------------


module inPlaceNTT_DIF_core (
  clk, rst, vec_rsc_triosy_0_0_lz, vec_rsc_triosy_0_1_lz, vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz, vec_rsc_triosy_0_4_lz, vec_rsc_triosy_0_5_lz, vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz, vec_rsc_triosy_0_8_lz, vec_rsc_triosy_0_9_lz, vec_rsc_triosy_0_10_lz,
      vec_rsc_triosy_0_11_lz, vec_rsc_triosy_0_12_lz, vec_rsc_triosy_0_13_lz, vec_rsc_triosy_0_14_lz,
      vec_rsc_triosy_0_15_lz, vec_rsc_triosy_0_16_lz, vec_rsc_triosy_0_17_lz, vec_rsc_triosy_0_18_lz,
      vec_rsc_triosy_0_19_lz, vec_rsc_triosy_0_20_lz, vec_rsc_triosy_0_21_lz, vec_rsc_triosy_0_22_lz,
      vec_rsc_triosy_0_23_lz, vec_rsc_triosy_0_24_lz, vec_rsc_triosy_0_25_lz, vec_rsc_triosy_0_26_lz,
      vec_rsc_triosy_0_27_lz, vec_rsc_triosy_0_28_lz, vec_rsc_triosy_0_29_lz, vec_rsc_triosy_0_30_lz,
      vec_rsc_triosy_0_31_lz, p_rsc_dat, p_rsc_triosy_lz, r_rsc_triosy_lz, twiddle_rsc_triosy_0_0_lz,
      twiddle_rsc_triosy_0_1_lz, twiddle_rsc_triosy_0_2_lz, twiddle_rsc_triosy_0_3_lz,
      twiddle_rsc_triosy_0_4_lz, twiddle_rsc_triosy_0_5_lz, twiddle_rsc_triosy_0_6_lz,
      twiddle_rsc_triosy_0_7_lz, twiddle_rsc_triosy_0_8_lz, twiddle_rsc_triosy_0_9_lz,
      twiddle_rsc_triosy_0_10_lz, twiddle_rsc_triosy_0_11_lz, twiddle_rsc_triosy_0_12_lz,
      twiddle_rsc_triosy_0_13_lz, twiddle_rsc_triosy_0_14_lz, twiddle_rsc_triosy_0_15_lz,
      twiddle_rsc_triosy_0_16_lz, twiddle_rsc_triosy_0_17_lz, twiddle_rsc_triosy_0_18_lz,
      twiddle_rsc_triosy_0_19_lz, twiddle_rsc_triosy_0_20_lz, twiddle_rsc_triosy_0_21_lz,
      twiddle_rsc_triosy_0_22_lz, twiddle_rsc_triosy_0_23_lz, twiddle_rsc_triosy_0_24_lz,
      twiddle_rsc_triosy_0_25_lz, twiddle_rsc_triosy_0_26_lz, twiddle_rsc_triosy_0_27_lz,
      twiddle_rsc_triosy_0_28_lz, twiddle_rsc_triosy_0_29_lz, twiddle_rsc_triosy_0_30_lz,
      twiddle_rsc_triosy_0_31_lz, vec_rsc_0_0_i_q_d, vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_1_i_q_d, vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_2_i_q_d,
      vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_3_i_q_d, vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_4_i_q_d, vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_5_i_q_d,
      vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_6_i_q_d, vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_7_i_q_d, vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_8_i_q_d,
      vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_9_i_q_d, vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_10_i_q_d, vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_11_i_q_d,
      vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_12_i_q_d, vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_13_i_q_d, vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_14_i_q_d,
      vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_15_i_q_d, vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_16_i_q_d, vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_17_i_q_d,
      vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_18_i_q_d, vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_19_i_q_d, vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_20_i_q_d,
      vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_21_i_q_d, vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_22_i_q_d, vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_23_i_q_d,
      vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_24_i_q_d, vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_25_i_q_d, vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_26_i_q_d,
      vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_27_i_q_d, vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_28_i_q_d, vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_29_i_q_d,
      vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_30_i_q_d, vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_31_i_q_d, vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_0_i_q_d,
      twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_1_i_q_d,
      twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_2_i_q_d,
      twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_3_i_q_d,
      twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_4_i_q_d,
      twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_5_i_q_d,
      twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_6_i_q_d,
      twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_7_i_q_d,
      twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_8_i_q_d,
      twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_9_i_q_d,
      twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_10_i_q_d,
      twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_11_i_q_d,
      twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_12_i_q_d,
      twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_13_i_q_d,
      twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_14_i_q_d,
      twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_15_i_q_d,
      twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_16_i_q_d,
      twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_17_i_q_d,
      twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_18_i_q_d,
      twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_19_i_q_d,
      twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_20_i_q_d,
      twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_21_i_q_d,
      twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_22_i_q_d,
      twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_23_i_q_d,
      twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_24_i_q_d,
      twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_25_i_q_d,
      twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_26_i_q_d,
      twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_27_i_q_d,
      twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_28_i_q_d,
      twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_29_i_q_d,
      twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_30_i_q_d,
      twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_31_i_q_d,
      twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_0_i_d_d_pff,
      vec_rsc_0_0_i_radr_d_pff, vec_rsc_0_0_i_wadr_d_pff, vec_rsc_0_0_i_we_d_pff,
      vec_rsc_0_1_i_we_d_pff, vec_rsc_0_2_i_we_d_pff, vec_rsc_0_3_i_we_d_pff, vec_rsc_0_4_i_we_d_pff,
      vec_rsc_0_5_i_we_d_pff, vec_rsc_0_6_i_we_d_pff, vec_rsc_0_7_i_we_d_pff, vec_rsc_0_8_i_we_d_pff,
      vec_rsc_0_9_i_we_d_pff, vec_rsc_0_10_i_we_d_pff, vec_rsc_0_11_i_we_d_pff, vec_rsc_0_12_i_we_d_pff,
      vec_rsc_0_13_i_we_d_pff, vec_rsc_0_14_i_we_d_pff, vec_rsc_0_15_i_we_d_pff,
      vec_rsc_0_16_i_we_d_pff, vec_rsc_0_17_i_we_d_pff, vec_rsc_0_18_i_we_d_pff,
      vec_rsc_0_19_i_we_d_pff, vec_rsc_0_20_i_we_d_pff, vec_rsc_0_21_i_we_d_pff,
      vec_rsc_0_22_i_we_d_pff, vec_rsc_0_23_i_we_d_pff, vec_rsc_0_24_i_we_d_pff,
      vec_rsc_0_25_i_we_d_pff, vec_rsc_0_26_i_we_d_pff, vec_rsc_0_27_i_we_d_pff,
      vec_rsc_0_28_i_we_d_pff, vec_rsc_0_29_i_we_d_pff, vec_rsc_0_30_i_we_d_pff,
      vec_rsc_0_31_i_we_d_pff, twiddle_rsc_0_0_i_radr_d_pff, twiddle_rsc_0_1_i_radr_d_pff,
      twiddle_rsc_0_2_i_radr_d_pff, twiddle_rsc_0_4_i_radr_d_pff
);
  input clk;
  input rst;
  output vec_rsc_triosy_0_0_lz;
  output vec_rsc_triosy_0_1_lz;
  output vec_rsc_triosy_0_2_lz;
  output vec_rsc_triosy_0_3_lz;
  output vec_rsc_triosy_0_4_lz;
  output vec_rsc_triosy_0_5_lz;
  output vec_rsc_triosy_0_6_lz;
  output vec_rsc_triosy_0_7_lz;
  output vec_rsc_triosy_0_8_lz;
  output vec_rsc_triosy_0_9_lz;
  output vec_rsc_triosy_0_10_lz;
  output vec_rsc_triosy_0_11_lz;
  output vec_rsc_triosy_0_12_lz;
  output vec_rsc_triosy_0_13_lz;
  output vec_rsc_triosy_0_14_lz;
  output vec_rsc_triosy_0_15_lz;
  output vec_rsc_triosy_0_16_lz;
  output vec_rsc_triosy_0_17_lz;
  output vec_rsc_triosy_0_18_lz;
  output vec_rsc_triosy_0_19_lz;
  output vec_rsc_triosy_0_20_lz;
  output vec_rsc_triosy_0_21_lz;
  output vec_rsc_triosy_0_22_lz;
  output vec_rsc_triosy_0_23_lz;
  output vec_rsc_triosy_0_24_lz;
  output vec_rsc_triosy_0_25_lz;
  output vec_rsc_triosy_0_26_lz;
  output vec_rsc_triosy_0_27_lz;
  output vec_rsc_triosy_0_28_lz;
  output vec_rsc_triosy_0_29_lz;
  output vec_rsc_triosy_0_30_lz;
  output vec_rsc_triosy_0_31_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  output r_rsc_triosy_lz;
  output twiddle_rsc_triosy_0_0_lz;
  output twiddle_rsc_triosy_0_1_lz;
  output twiddle_rsc_triosy_0_2_lz;
  output twiddle_rsc_triosy_0_3_lz;
  output twiddle_rsc_triosy_0_4_lz;
  output twiddle_rsc_triosy_0_5_lz;
  output twiddle_rsc_triosy_0_6_lz;
  output twiddle_rsc_triosy_0_7_lz;
  output twiddle_rsc_triosy_0_8_lz;
  output twiddle_rsc_triosy_0_9_lz;
  output twiddle_rsc_triosy_0_10_lz;
  output twiddle_rsc_triosy_0_11_lz;
  output twiddle_rsc_triosy_0_12_lz;
  output twiddle_rsc_triosy_0_13_lz;
  output twiddle_rsc_triosy_0_14_lz;
  output twiddle_rsc_triosy_0_15_lz;
  output twiddle_rsc_triosy_0_16_lz;
  output twiddle_rsc_triosy_0_17_lz;
  output twiddle_rsc_triosy_0_18_lz;
  output twiddle_rsc_triosy_0_19_lz;
  output twiddle_rsc_triosy_0_20_lz;
  output twiddle_rsc_triosy_0_21_lz;
  output twiddle_rsc_triosy_0_22_lz;
  output twiddle_rsc_triosy_0_23_lz;
  output twiddle_rsc_triosy_0_24_lz;
  output twiddle_rsc_triosy_0_25_lz;
  output twiddle_rsc_triosy_0_26_lz;
  output twiddle_rsc_triosy_0_27_lz;
  output twiddle_rsc_triosy_0_28_lz;
  output twiddle_rsc_triosy_0_29_lz;
  output twiddle_rsc_triosy_0_30_lz;
  output twiddle_rsc_triosy_0_31_lz;
  input [63:0] vec_rsc_0_0_i_q_d;
  output vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_1_i_q_d;
  output vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_2_i_q_d;
  output vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_3_i_q_d;
  output vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_4_i_q_d;
  output vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_5_i_q_d;
  output vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_6_i_q_d;
  output vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_7_i_q_d;
  output vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_8_i_q_d;
  output vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_9_i_q_d;
  output vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_10_i_q_d;
  output vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_11_i_q_d;
  output vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_12_i_q_d;
  output vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_13_i_q_d;
  output vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_14_i_q_d;
  output vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_15_i_q_d;
  output vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_16_i_q_d;
  output vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_17_i_q_d;
  output vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_18_i_q_d;
  output vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_19_i_q_d;
  output vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_20_i_q_d;
  output vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_21_i_q_d;
  output vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_22_i_q_d;
  output vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_23_i_q_d;
  output vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_24_i_q_d;
  output vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_25_i_q_d;
  output vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_26_i_q_d;
  output vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_27_i_q_d;
  output vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_28_i_q_d;
  output vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_29_i_q_d;
  output vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_30_i_q_d;
  output vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_31_i_q_d;
  output vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_0_i_q_d;
  output twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_1_i_q_d;
  output twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_2_i_q_d;
  output twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_3_i_q_d;
  output twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_4_i_q_d;
  output twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_5_i_q_d;
  output twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_6_i_q_d;
  output twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_7_i_q_d;
  output twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_8_i_q_d;
  output twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_9_i_q_d;
  output twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_10_i_q_d;
  output twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_11_i_q_d;
  output twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_12_i_q_d;
  output twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_13_i_q_d;
  output twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_14_i_q_d;
  output twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_15_i_q_d;
  output twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_16_i_q_d;
  output twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_17_i_q_d;
  output twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_18_i_q_d;
  output twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_19_i_q_d;
  output twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_20_i_q_d;
  output twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_21_i_q_d;
  output twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_22_i_q_d;
  output twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_23_i_q_d;
  output twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_24_i_q_d;
  output twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_25_i_q_d;
  output twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_26_i_q_d;
  output twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_27_i_q_d;
  output twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_28_i_q_d;
  output twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_29_i_q_d;
  output twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_30_i_q_d;
  output twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_31_i_q_d;
  output twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d;
  output [63:0] vec_rsc_0_0_i_d_d_pff;
  output [4:0] vec_rsc_0_0_i_radr_d_pff;
  output [4:0] vec_rsc_0_0_i_wadr_d_pff;
  output vec_rsc_0_0_i_we_d_pff;
  output vec_rsc_0_1_i_we_d_pff;
  output vec_rsc_0_2_i_we_d_pff;
  output vec_rsc_0_3_i_we_d_pff;
  output vec_rsc_0_4_i_we_d_pff;
  output vec_rsc_0_5_i_we_d_pff;
  output vec_rsc_0_6_i_we_d_pff;
  output vec_rsc_0_7_i_we_d_pff;
  output vec_rsc_0_8_i_we_d_pff;
  output vec_rsc_0_9_i_we_d_pff;
  output vec_rsc_0_10_i_we_d_pff;
  output vec_rsc_0_11_i_we_d_pff;
  output vec_rsc_0_12_i_we_d_pff;
  output vec_rsc_0_13_i_we_d_pff;
  output vec_rsc_0_14_i_we_d_pff;
  output vec_rsc_0_15_i_we_d_pff;
  output vec_rsc_0_16_i_we_d_pff;
  output vec_rsc_0_17_i_we_d_pff;
  output vec_rsc_0_18_i_we_d_pff;
  output vec_rsc_0_19_i_we_d_pff;
  output vec_rsc_0_20_i_we_d_pff;
  output vec_rsc_0_21_i_we_d_pff;
  output vec_rsc_0_22_i_we_d_pff;
  output vec_rsc_0_23_i_we_d_pff;
  output vec_rsc_0_24_i_we_d_pff;
  output vec_rsc_0_25_i_we_d_pff;
  output vec_rsc_0_26_i_we_d_pff;
  output vec_rsc_0_27_i_we_d_pff;
  output vec_rsc_0_28_i_we_d_pff;
  output vec_rsc_0_29_i_we_d_pff;
  output vec_rsc_0_30_i_we_d_pff;
  output vec_rsc_0_31_i_we_d_pff;
  output [4:0] twiddle_rsc_0_0_i_radr_d_pff;
  output [4:0] twiddle_rsc_0_1_i_radr_d_pff;
  output [4:0] twiddle_rsc_0_2_i_radr_d_pff;
  output [4:0] twiddle_rsc_0_4_i_radr_d_pff;


  // Interconnect Declarations
  wire [63:0] p_rsci_idat;
  wire [63:0] COMP_LOOP_1_modulo_dev_cmp_return_rsc_z;
  wire COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en;
  wire [7:0] fsm_output;
  wire nor_tmp_53;
  wire or_tmp_142;
  wire and_dcpl_28;
  wire and_dcpl_29;
  wire and_dcpl_30;
  wire and_dcpl_31;
  wire and_dcpl_33;
  wire and_dcpl_35;
  wire and_dcpl_36;
  wire and_dcpl_38;
  wire nor_tmp_95;
  wire and_dcpl_40;
  wire and_dcpl_44;
  wire and_dcpl_45;
  wire and_dcpl_46;
  wire and_dcpl_48;
  wire and_dcpl_49;
  wire and_dcpl_50;
  wire and_dcpl_52;
  wire and_dcpl_54;
  wire and_dcpl_55;
  wire and_dcpl_56;
  wire and_dcpl_58;
  wire and_dcpl_59;
  wire and_dcpl_60;
  wire and_dcpl_61;
  wire and_dcpl_62;
  wire and_dcpl_64;
  wire and_dcpl_65;
  wire and_dcpl_66;
  wire and_dcpl_68;
  wire and_dcpl_69;
  wire and_dcpl_70;
  wire and_dcpl_71;
  wire and_dcpl_72;
  wire and_dcpl_74;
  wire and_dcpl_75;
  wire and_dcpl_76;
  wire and_dcpl_78;
  wire and_dcpl_79;
  wire and_dcpl_82;
  wire and_dcpl_83;
  wire and_dcpl_85;
  wire and_dcpl_89;
  wire and_dcpl_91;
  wire and_dcpl_95;
  wire and_dcpl_97;
  wire and_dcpl_102;
  wire and_dcpl_104;
  wire mux_tmp_311;
  wire mux_tmp_373;
  wire mux_tmp_435;
  wire mux_tmp_497;
  wire mux_tmp_559;
  wire mux_tmp_621;
  wire mux_tmp_683;
  wire mux_tmp_745;
  wire mux_tmp_807;
  wire mux_tmp_869;
  wire mux_tmp_931;
  wire mux_tmp_993;
  wire mux_tmp_1055;
  wire mux_tmp_1117;
  wire mux_tmp_1179;
  wire mux_tmp_1241;
  wire and_dcpl_171;
  wire and_dcpl_172;
  wire and_dcpl_173;
  wire and_dcpl_174;
  wire and_dcpl_175;
  wire and_dcpl_176;
  wire and_dcpl_177;
  wire and_dcpl_178;
  wire and_dcpl_179;
  wire not_tmp_617;
  wire not_tmp_618;
  wire not_tmp_625;
  wire not_tmp_632;
  wire mux_tmp_1423;
  wire or_tmp_2024;
  wire mux_tmp_1424;
  wire or_tmp_2025;
  wire mux_tmp_1430;
  wire and_dcpl_220;
  wire and_dcpl_222;
  wire and_dcpl_223;
  wire and_dcpl_226;
  wire and_dcpl_229;
  wire and_dcpl_232;
  wire and_dcpl_234;
  wire and_dcpl_236;
  wire and_dcpl_238;
  wire nand_tmp_184;
  wire mux_tmp_1437;
  wire and_dcpl_244;
  wire or_dcpl_84;
  wire or_tmp_2048;
  wire mux_tmp_1452;
  wire mux_tmp_1456;
  wire mux_tmp_1459;
  wire and_tmp_11;
  wire or_tmp_2054;
  wire not_tmp_692;
  wire or_tmp_2057;
  wire and_dcpl_252;
  wire mux_tmp_1468;
  wire and_tmp_13;
  wire and_dcpl_256;
  wire nor_tmp_324;
  wire and_dcpl_259;
  wire mux_tmp_1482;
  wire mux_tmp_1487;
  wire and_dcpl_260;
  wire not_tmp_717;
  wire and_dcpl_262;
  wire and_dcpl_264;
  wire and_dcpl_278;
  wire or_tmp_2075;
  wire or_dcpl_109;
  reg COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm;
  wire [9:0] COMP_LOOP_acc_1_cse_6_sva_1;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_6_sva_1;
  reg [9:0] VEC_LOOP_j_10_0_sva_9_0;
  wire [9:0] COMP_LOOP_acc_1_cse_4_sva_1;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_4_sva_1;
  reg [6:0] COMP_LOOP_k_10_3_sva_6_0;
  reg COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm;
  reg COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm;
  reg COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm;
  reg [9:0] COMP_LOOP_2_tmp_lshift_ncse_sva;
  reg COMP_LOOP_tmp_nor_42_itm;
  reg [9:0] COMP_LOOP_2_tmp_mul_idiv_sva;
  reg COMP_LOOP_tmp_nor_1_itm;
  reg [8:0] COMP_LOOP_3_tmp_lshift_ncse_sva;
  reg COMP_LOOP_tmp_nor_25_itm;
  reg COMP_LOOP_tmp_nor_49_itm;
  reg COMP_LOOP_tmp_nor_14_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_124_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_122_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_128_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_132_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_126_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_130_itm;
  reg [6:0] COMP_LOOP_acc_psp_sva;
  reg [7:0] COMP_LOOP_acc_13_psp_sva;
  wire [8:0] nl_COMP_LOOP_acc_13_psp_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_1_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_5_sva;
  reg [8:0] COMP_LOOP_acc_11_psp_sva;
  wire [9:0] nl_COMP_LOOP_acc_11_psp_sva;
  reg [8:0] COMP_LOOP_acc_14_psp_sva;
  wire [9:0] nl_COMP_LOOP_acc_14_psp_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_3_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_7_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_2_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_6_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_2_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_6_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_4_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_sva;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_4_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_sva;
  reg [7:0] COMP_LOOP_5_tmp_mul_idiv_sva;
  reg [1:0] COMP_LOOP_1_tmp_mul_idiv_sva_1_0;
  reg [10:0] STAGE_LOOP_lshift_psp_sva;
  wire [9:0] COMP_LOOP_acc_1_cse_2_sva_1;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_2_sva_1;
  wire [6:0] COMP_LOOP_acc_psp_sva_mx0w0;
  wire [7:0] nl_COMP_LOOP_acc_psp_sva_mx0w0;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_rgt;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_rgt;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_rgt;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_rgt;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_119_rgt;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_121_rgt;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_125_rgt;
  wire mux_1592_tmp;
  wire and_298_m1c;
  wire nor_1117_tmp;
  wire nor_tmp;
  wire nor_1119_tmp;
  wire and_294_tmp;
  reg [6:0] reg_COMP_LOOP_k_10_3_ftd;
  wire or_285_cse;
  wire nand_443_cse;
  wire nand_444_cse;
  wire or_493_cse;
  wire or_701_cse;
  wire nand_394_cse;
  wire or_1113_cse;
  wire nand_356_cse;
  wire nand_336_cse;
  wire nand_300_cse;
  wire nand_293_cse;
  wire nand_264_cse;
  wire nand_204_cse;
  wire nand_205_cse;
  reg reg_vec_rsc_triosy_0_31_obj_ld_cse;
  reg reg_ensig_cgo_cse;
  wire or_220_cse;
  wire or_212_cse;
  wire and_496_cse;
  wire and_316_cse;
  wire or_32_cse;
  wire mux_189_cse;
  wire COMP_LOOP_tmp_or_cse;
  wire COMP_LOOP_tmp_or_12_cse;
  wire COMP_LOOP_tmp_or_17_cse;
  wire COMP_LOOP_tmp_or_35_cse;
  wire COMP_LOOP_tmp_or_40_cse;
  wire and_4_cse;
  wire and_1_cse;
  wire nor_1025_cse;
  wire and_464_cse;
  wire and_490_cse;
  wire and_449_cse;
  wire and_479_cse;
  wire mux_322_cse;
  wire nand_445_cse;
  wire nand_447_cse;
  wire nand_441_cse;
  wire nand_442_cse;
  wire mux_353_cse;
  wire nand_446_cse;
  wire nand_448_cse;
  wire nor_98_cse;
  wire mux_446_cse;
  wire nand_423_cse;
  wire mux_477_cse;
  wire mux_570_cse;
  wire nand_435_cse;
  wire nand_411_cse;
  wire nand_437_cse;
  wire mux_601_cse;
  wire mux_694_cse;
  wire nand_371_cse;
  wire nand_385_cse;
  wire mux_725_cse;
  wire nand_364_cse;
  wire nand_365_cse;
  wire nand_357_cse;
  wire nand_353_cse;
  wire nand_417_cse;
  wire nand_419_cse;
  wire nand_302_cse;
  wire nand_303_cse;
  wire nand_294_cse;
  wire nand_289_cse;
  wire nand_266_cse;
  wire nand_297_cse;
  wire mux_1190_cse;
  wire mux_1221_cse;
  wire or_167_cse;
  wire or_145_cse;
  wire nor_1023_cse;
  wire and_491_cse;
  wire and_485_cse;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm;
  wire mux_348_cse;
  wire mux_410_cse;
  wire mux_472_cse;
  wire mux_534_cse;
  wire mux_596_cse;
  wire mux_658_cse;
  wire mux_720_cse;
  wire mux_782_cse;
  wire mux_844_cse;
  wire mux_818_cse;
  wire mux_849_cse;
  wire mux_906_cse;
  wire mux_968_cse;
  wire mux_942_cse;
  wire mux_973_cse;
  wire mux_1030_cse;
  wire mux_1092_cse;
  wire mux_1066_cse;
  wire mux_1097_cse;
  wire mux_1154_cse;
  wire mux_1216_cse;
  wire mux_1278_cse;
  wire and_33_cse;
  wire and_456_cse;
  wire mux_1462_rmff;
  reg [63:0] COMP_LOOP_1_acc_8_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_1_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_2_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_3_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_4_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_5_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_6_itm;
  reg [63:0] tmp_21_sva_1;
  reg [63:0] p_sva;
  wire mux_1489_itm;
  wire mux_1531_itm;
  wire mux_1536_itm;
  wire mux_1538_itm;
  wire mux_1543_itm;
  wire [10:0] z_out;
  wire [9:0] z_out_1;
  wire [7:0] z_out_2;
  wire [8:0] nl_z_out_2;
  wire and_dcpl_334;
  wire [10:0] z_out_3;
  wire and_dcpl_347;
  wire [3:0] z_out_4;
  wire [4:0] nl_z_out_4;
  wire and_dcpl_353;
  wire and_dcpl_365;
  wire and_dcpl_372;
  wire and_dcpl_419;
  wire and_dcpl_420;
  wire and_dcpl_422;
  wire and_dcpl_423;
  wire and_dcpl_425;
  wire and_dcpl_428;
  wire and_dcpl_429;
  wire and_dcpl_433;
  wire and_dcpl_434;
  wire and_dcpl_435;
  wire and_dcpl_436;
  wire [9:0] z_out_7;
  wire [19:0] nl_z_out_7;
  wire and_dcpl_448;
  wire and_dcpl_452;
  wire and_dcpl_456;
  wire and_dcpl_458;
  wire and_dcpl_461;
  wire and_dcpl_465;
  wire and_dcpl_468;
  wire and_dcpl_472;
  wire [63:0] z_out_8;
  wire [127:0] nl_z_out_8;
  wire and_dcpl_479;
  wire [63:0] z_out_9;
  reg [3:0] STAGE_LOOP_i_3_0_sva;
  reg [3:0] COMP_LOOP_1_tmp_acc_cse_sva;
  reg [63:0] tmp_21_sva_2;
  reg [63:0] tmp_21_sva_3;
  reg [63:0] tmp_21_sva_5;
  reg [63:0] tmp_21_sva_6;
  reg [63:0] tmp_21_sva_7;
  reg [63:0] tmp_21_sva_9;
  reg [63:0] tmp_21_sva_11;
  reg [63:0] tmp_21_sva_13;
  reg [63:0] tmp_21_sva_14;
  reg [63:0] tmp_21_sva_15;
  reg [63:0] tmp_21_sva_17;
  reg [63:0] tmp_21_sva_18;
  reg [63:0] tmp_21_sva_19;
  reg [63:0] tmp_21_sva_21;
  reg [63:0] tmp_21_sva_22;
  reg [63:0] tmp_21_sva_23;
  reg [63:0] tmp_21_sva_25;
  reg [63:0] tmp_21_sva_26;
  reg [63:0] tmp_21_sva_27;
  reg [63:0] tmp_21_sva_29;
  reg [63:0] tmp_21_sva_30;
  reg [63:0] tmp_21_sva_31;
  reg COMP_LOOP_COMP_LOOP_nor_itm;
  reg COMP_LOOP_COMP_LOOP_and_6_itm;
  reg COMP_LOOP_COMP_LOOP_and_10_itm;
  reg COMP_LOOP_COMP_LOOP_and_12_itm;
  reg COMP_LOOP_COMP_LOOP_and_13_itm;
  reg COMP_LOOP_COMP_LOOP_and_14_itm;
  reg COMP_LOOP_COMP_LOOP_and_18_itm;
  reg COMP_LOOP_COMP_LOOP_and_20_itm;
  reg COMP_LOOP_COMP_LOOP_and_21_itm;
  reg COMP_LOOP_COMP_LOOP_and_22_itm;
  reg COMP_LOOP_COMP_LOOP_and_23_itm;
  reg COMP_LOOP_COMP_LOOP_and_24_itm;
  reg COMP_LOOP_COMP_LOOP_and_25_itm;
  reg COMP_LOOP_COMP_LOOP_and_26_itm;
  reg COMP_LOOP_COMP_LOOP_and_27_itm;
  reg COMP_LOOP_COMP_LOOP_and_28_itm;
  reg COMP_LOOP_COMP_LOOP_and_29_itm;
  reg COMP_LOOP_COMP_LOOP_and_30_itm;
  reg COMP_LOOP_COMP_LOOP_and_126_itm;
  reg COMP_LOOP_COMP_LOOP_and_128_itm;
  reg COMP_LOOP_COMP_LOOP_and_129_itm;
  reg COMP_LOOP_COMP_LOOP_and_130_itm;
  reg COMP_LOOP_COMP_LOOP_and_132_itm;
  reg COMP_LOOP_COMP_LOOP_and_133_itm;
  reg COMP_LOOP_COMP_LOOP_and_134_itm;
  reg COMP_LOOP_COMP_LOOP_and_136_itm;
  reg COMP_LOOP_COMP_LOOP_and_140_itm;
  reg COMP_LOOP_COMP_LOOP_and_141_itm;
  reg COMP_LOOP_COMP_LOOP_and_142_itm;
  reg COMP_LOOP_COMP_LOOP_and_144_itm;
  reg COMP_LOOP_COMP_LOOP_nor_5_itm;
  reg COMP_LOOP_nor_126_itm;
  reg COMP_LOOP_nor_127_itm;
  reg COMP_LOOP_COMP_LOOP_and_157_itm;
  reg COMP_LOOP_nor_129_itm;
  reg COMP_LOOP_COMP_LOOP_and_159_itm;
  reg COMP_LOOP_COMP_LOOP_and_160_itm;
  reg COMP_LOOP_COMP_LOOP_and_161_itm;
  reg COMP_LOOP_nor_133_itm;
  reg COMP_LOOP_COMP_LOOP_and_163_itm;
  reg COMP_LOOP_COMP_LOOP_and_164_itm;
  reg COMP_LOOP_COMP_LOOP_and_165_itm;
  reg COMP_LOOP_COMP_LOOP_and_166_itm;
  reg COMP_LOOP_COMP_LOOP_and_167_itm;
  reg COMP_LOOP_COMP_LOOP_and_168_itm;
  reg COMP_LOOP_COMP_LOOP_and_169_itm;
  reg COMP_LOOP_nor_140_itm;
  reg COMP_LOOP_COMP_LOOP_and_171_itm;
  reg COMP_LOOP_COMP_LOOP_and_172_itm;
  reg COMP_LOOP_COMP_LOOP_and_173_itm;
  reg COMP_LOOP_COMP_LOOP_and_174_itm;
  reg COMP_LOOP_COMP_LOOP_and_175_itm;
  reg COMP_LOOP_COMP_LOOP_and_176_itm;
  reg COMP_LOOP_COMP_LOOP_and_177_itm;
  reg COMP_LOOP_COMP_LOOP_and_178_itm;
  reg COMP_LOOP_COMP_LOOP_and_179_itm;
  reg COMP_LOOP_COMP_LOOP_and_180_itm;
  reg COMP_LOOP_COMP_LOOP_and_181_itm;
  reg COMP_LOOP_COMP_LOOP_and_182_itm;
  reg COMP_LOOP_COMP_LOOP_and_183_itm;
  reg COMP_LOOP_COMP_LOOP_and_184_itm;
  reg COMP_LOOP_COMP_LOOP_and_185_itm;
  reg COMP_LOOP_tmp_nor_3_itm;
  reg COMP_LOOP_COMP_LOOP_nor_9_itm;
  reg COMP_LOOP_nor_226_itm;
  reg COMP_LOOP_nor_227_itm;
  reg COMP_LOOP_COMP_LOOP_and_281_itm;
  reg COMP_LOOP_nor_229_itm;
  reg COMP_LOOP_COMP_LOOP_and_283_itm;
  reg COMP_LOOP_COMP_LOOP_and_284_itm;
  reg COMP_LOOP_COMP_LOOP_and_285_itm;
  reg COMP_LOOP_nor_233_itm;
  reg COMP_LOOP_COMP_LOOP_and_287_itm;
  reg COMP_LOOP_COMP_LOOP_and_288_itm;
  reg COMP_LOOP_COMP_LOOP_and_289_itm;
  reg COMP_LOOP_COMP_LOOP_and_290_itm;
  reg COMP_LOOP_COMP_LOOP_and_291_itm;
  reg COMP_LOOP_COMP_LOOP_and_292_itm;
  reg COMP_LOOP_COMP_LOOP_and_293_itm;
  reg COMP_LOOP_nor_240_itm;
  reg COMP_LOOP_COMP_LOOP_and_295_itm;
  reg COMP_LOOP_COMP_LOOP_and_296_itm;
  reg COMP_LOOP_COMP_LOOP_and_297_itm;
  reg COMP_LOOP_COMP_LOOP_and_298_itm;
  reg COMP_LOOP_COMP_LOOP_and_299_itm;
  reg COMP_LOOP_COMP_LOOP_and_300_itm;
  reg COMP_LOOP_COMP_LOOP_and_301_itm;
  reg COMP_LOOP_COMP_LOOP_and_302_itm;
  reg COMP_LOOP_COMP_LOOP_and_303_itm;
  reg COMP_LOOP_COMP_LOOP_and_304_itm;
  reg COMP_LOOP_COMP_LOOP_and_305_itm;
  reg COMP_LOOP_COMP_LOOP_and_306_itm;
  reg COMP_LOOP_COMP_LOOP_and_307_itm;
  reg COMP_LOOP_COMP_LOOP_and_308_itm;
  reg COMP_LOOP_COMP_LOOP_and_309_itm;
  reg COMP_LOOP_tmp_nor_26_itm;
  reg COMP_LOOP_tmp_nor_28_itm;
  reg COMP_LOOP_tmp_nor_31_itm;
  reg COMP_LOOP_COMP_LOOP_and_377_itm;
  reg COMP_LOOP_COMP_LOOP_nor_13_itm;
  reg COMP_LOOP_nor_326_itm;
  reg COMP_LOOP_nor_327_itm;
  reg COMP_LOOP_COMP_LOOP_and_405_itm;
  reg COMP_LOOP_nor_329_itm;
  reg COMP_LOOP_COMP_LOOP_and_407_itm;
  reg COMP_LOOP_COMP_LOOP_and_408_itm;
  reg COMP_LOOP_COMP_LOOP_and_409_itm;
  reg COMP_LOOP_nor_333_itm;
  reg COMP_LOOP_COMP_LOOP_and_411_itm;
  reg COMP_LOOP_COMP_LOOP_and_412_itm;
  reg COMP_LOOP_COMP_LOOP_and_413_itm;
  reg COMP_LOOP_COMP_LOOP_and_414_itm;
  reg COMP_LOOP_COMP_LOOP_and_415_itm;
  reg COMP_LOOP_COMP_LOOP_and_416_itm;
  reg COMP_LOOP_COMP_LOOP_and_417_itm;
  reg COMP_LOOP_nor_340_itm;
  reg COMP_LOOP_COMP_LOOP_and_419_itm;
  reg COMP_LOOP_COMP_LOOP_and_420_itm;
  reg COMP_LOOP_COMP_LOOP_and_421_itm;
  reg COMP_LOOP_COMP_LOOP_and_422_itm;
  reg COMP_LOOP_COMP_LOOP_and_423_itm;
  reg COMP_LOOP_COMP_LOOP_and_424_itm;
  reg COMP_LOOP_COMP_LOOP_and_425_itm;
  reg COMP_LOOP_COMP_LOOP_and_426_itm;
  reg COMP_LOOP_COMP_LOOP_and_427_itm;
  reg COMP_LOOP_COMP_LOOP_and_428_itm;
  reg COMP_LOOP_COMP_LOOP_and_429_itm;
  reg COMP_LOOP_COMP_LOOP_and_430_itm;
  reg COMP_LOOP_COMP_LOOP_and_431_itm;
  reg COMP_LOOP_COMP_LOOP_and_432_itm;
  reg COMP_LOOP_COMP_LOOP_and_433_itm;
  reg COMP_LOOP_COMP_LOOP_nor_17_itm;
  reg COMP_LOOP_nor_426_itm;
  reg COMP_LOOP_nor_427_itm;
  reg COMP_LOOP_COMP_LOOP_and_529_itm;
  reg COMP_LOOP_nor_429_itm;
  reg COMP_LOOP_COMP_LOOP_and_531_itm;
  reg COMP_LOOP_COMP_LOOP_and_532_itm;
  reg COMP_LOOP_COMP_LOOP_and_533_itm;
  reg COMP_LOOP_nor_433_itm;
  reg COMP_LOOP_COMP_LOOP_and_535_itm;
  reg COMP_LOOP_COMP_LOOP_and_536_itm;
  reg COMP_LOOP_COMP_LOOP_and_537_itm;
  reg COMP_LOOP_COMP_LOOP_and_538_itm;
  reg COMP_LOOP_COMP_LOOP_and_539_itm;
  reg COMP_LOOP_COMP_LOOP_and_540_itm;
  reg COMP_LOOP_COMP_LOOP_and_541_itm;
  reg COMP_LOOP_nor_440_itm;
  reg COMP_LOOP_COMP_LOOP_and_543_itm;
  reg COMP_LOOP_COMP_LOOP_and_544_itm;
  reg COMP_LOOP_COMP_LOOP_and_545_itm;
  reg COMP_LOOP_COMP_LOOP_and_546_itm;
  reg COMP_LOOP_COMP_LOOP_and_547_itm;
  reg COMP_LOOP_COMP_LOOP_and_548_itm;
  reg COMP_LOOP_COMP_LOOP_and_549_itm;
  reg COMP_LOOP_COMP_LOOP_and_550_itm;
  reg COMP_LOOP_COMP_LOOP_and_551_itm;
  reg COMP_LOOP_COMP_LOOP_and_552_itm;
  reg COMP_LOOP_COMP_LOOP_and_553_itm;
  reg COMP_LOOP_COMP_LOOP_and_554_itm;
  reg COMP_LOOP_COMP_LOOP_and_555_itm;
  reg COMP_LOOP_COMP_LOOP_and_556_itm;
  reg COMP_LOOP_COMP_LOOP_and_557_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_82_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_84_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_85_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_86_itm;
  reg COMP_LOOP_COMP_LOOP_and_625_itm;
  reg COMP_LOOP_COMP_LOOP_nor_21_itm;
  reg COMP_LOOP_nor_526_itm;
  reg COMP_LOOP_nor_527_itm;
  reg COMP_LOOP_COMP_LOOP_and_653_itm;
  reg COMP_LOOP_nor_529_itm;
  reg COMP_LOOP_COMP_LOOP_and_655_itm;
  reg COMP_LOOP_COMP_LOOP_and_656_itm;
  reg COMP_LOOP_COMP_LOOP_and_657_itm;
  reg COMP_LOOP_nor_533_itm;
  reg COMP_LOOP_COMP_LOOP_and_659_itm;
  reg COMP_LOOP_COMP_LOOP_and_660_itm;
  reg COMP_LOOP_COMP_LOOP_and_661_itm;
  reg COMP_LOOP_COMP_LOOP_and_662_itm;
  reg COMP_LOOP_COMP_LOOP_and_663_itm;
  reg COMP_LOOP_COMP_LOOP_and_664_itm;
  reg COMP_LOOP_COMP_LOOP_and_665_itm;
  reg COMP_LOOP_nor_540_itm;
  reg COMP_LOOP_COMP_LOOP_and_667_itm;
  reg COMP_LOOP_COMP_LOOP_and_668_itm;
  reg COMP_LOOP_COMP_LOOP_and_669_itm;
  reg COMP_LOOP_COMP_LOOP_and_670_itm;
  reg COMP_LOOP_COMP_LOOP_and_671_itm;
  reg COMP_LOOP_COMP_LOOP_and_672_itm;
  reg COMP_LOOP_COMP_LOOP_and_673_itm;
  reg COMP_LOOP_COMP_LOOP_and_674_itm;
  reg COMP_LOOP_COMP_LOOP_and_675_itm;
  reg COMP_LOOP_COMP_LOOP_and_676_itm;
  reg COMP_LOOP_COMP_LOOP_and_677_itm;
  reg COMP_LOOP_COMP_LOOP_and_678_itm;
  reg COMP_LOOP_COMP_LOOP_and_679_itm;
  reg COMP_LOOP_COMP_LOOP_and_680_itm;
  reg COMP_LOOP_COMP_LOOP_and_681_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm;
  reg COMP_LOOP_COMP_LOOP_nor_25_itm;
  reg COMP_LOOP_nor_626_itm;
  reg COMP_LOOP_nor_627_itm;
  reg COMP_LOOP_COMP_LOOP_and_777_itm;
  reg COMP_LOOP_nor_629_itm;
  reg COMP_LOOP_COMP_LOOP_and_779_itm;
  reg COMP_LOOP_COMP_LOOP_and_780_itm;
  reg COMP_LOOP_COMP_LOOP_and_781_itm;
  reg COMP_LOOP_nor_633_itm;
  reg COMP_LOOP_COMP_LOOP_and_783_itm;
  reg COMP_LOOP_COMP_LOOP_and_784_itm;
  reg COMP_LOOP_COMP_LOOP_and_785_itm;
  reg COMP_LOOP_COMP_LOOP_and_786_itm;
  reg COMP_LOOP_COMP_LOOP_and_787_itm;
  reg COMP_LOOP_COMP_LOOP_and_788_itm;
  reg COMP_LOOP_COMP_LOOP_and_789_itm;
  reg COMP_LOOP_nor_640_itm;
  reg COMP_LOOP_COMP_LOOP_and_791_itm;
  reg COMP_LOOP_COMP_LOOP_and_792_itm;
  reg COMP_LOOP_COMP_LOOP_and_793_itm;
  reg COMP_LOOP_COMP_LOOP_and_794_itm;
  reg COMP_LOOP_COMP_LOOP_and_795_itm;
  reg COMP_LOOP_COMP_LOOP_and_796_itm;
  reg COMP_LOOP_COMP_LOOP_and_797_itm;
  reg COMP_LOOP_COMP_LOOP_and_798_itm;
  reg COMP_LOOP_COMP_LOOP_and_799_itm;
  reg COMP_LOOP_COMP_LOOP_and_800_itm;
  reg COMP_LOOP_COMP_LOOP_and_801_itm;
  reg COMP_LOOP_COMP_LOOP_and_802_itm;
  reg COMP_LOOP_COMP_LOOP_and_803_itm;
  reg COMP_LOOP_COMP_LOOP_and_804_itm;
  reg COMP_LOOP_COMP_LOOP_and_805_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_123_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_127_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_129_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_131_itm;
  reg COMP_LOOP_COMP_LOOP_nor_29_itm;
  reg COMP_LOOP_nor_726_itm;
  reg COMP_LOOP_nor_727_itm;
  reg COMP_LOOP_COMP_LOOP_and_901_itm;
  reg COMP_LOOP_nor_729_itm;
  reg COMP_LOOP_COMP_LOOP_and_903_itm;
  reg COMP_LOOP_COMP_LOOP_and_904_itm;
  reg COMP_LOOP_COMP_LOOP_and_905_itm;
  reg COMP_LOOP_nor_733_itm;
  reg COMP_LOOP_COMP_LOOP_and_907_itm;
  reg COMP_LOOP_COMP_LOOP_and_908_itm;
  reg COMP_LOOP_COMP_LOOP_and_909_itm;
  reg COMP_LOOP_COMP_LOOP_and_910_itm;
  reg COMP_LOOP_COMP_LOOP_and_911_itm;
  reg COMP_LOOP_COMP_LOOP_and_912_itm;
  reg COMP_LOOP_COMP_LOOP_and_913_itm;
  reg COMP_LOOP_nor_740_itm;
  reg COMP_LOOP_COMP_LOOP_and_915_itm;
  reg COMP_LOOP_COMP_LOOP_and_916_itm;
  reg COMP_LOOP_COMP_LOOP_and_917_itm;
  reg COMP_LOOP_COMP_LOOP_and_918_itm;
  reg COMP_LOOP_COMP_LOOP_and_919_itm;
  reg COMP_LOOP_COMP_LOOP_and_920_itm;
  reg COMP_LOOP_COMP_LOOP_and_921_itm;
  reg COMP_LOOP_COMP_LOOP_and_922_itm;
  reg COMP_LOOP_COMP_LOOP_and_923_itm;
  reg COMP_LOOP_COMP_LOOP_and_924_itm;
  reg COMP_LOOP_COMP_LOOP_and_925_itm;
  reg COMP_LOOP_COMP_LOOP_and_926_itm;
  reg COMP_LOOP_COMP_LOOP_and_927_itm;
  reg COMP_LOOP_COMP_LOOP_and_928_itm;
  reg COMP_LOOP_COMP_LOOP_and_929_itm;
  wire STAGE_LOOP_i_3_0_sva_mx0c1;
  wire VEC_LOOP_j_10_0_sva_9_0_mx0c0;
  wire COMP_LOOP_tmp_mux1h_itm_mx0c0;
  wire COMP_LOOP_tmp_mux1h_itm_mx0c1;
  wire COMP_LOOP_tmp_mux1h_itm_mx0c2;
  wire COMP_LOOP_tmp_mux1h_itm_mx0c3;
  wire COMP_LOOP_1_acc_8_itm_mx0c4;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_165;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_167;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_169;
  reg [3:0] COMP_LOOP_3_tmp_mul_idiv_sva_3_0;
  wire COMP_LOOP_or_59_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse;
  wire COMP_LOOP_tmp_nor_27_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse;
  wire COMP_LOOP_tmp_nor_29_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse;
  wire COMP_LOOP_tmp_nor_30_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_cse;
  wire COMP_LOOP_tmp_nor_32_cse;
  wire COMP_LOOP_tmp_nor_33_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_cse;
  wire COMP_LOOP_tmp_nor_34_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_40_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_44_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_46_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_47_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse;
  wire COMP_LOOP_tmp_nor_1_cse;
  wire COMP_LOOP_or_41_cse;
  wire COMP_LOOP_tmp_nor_101_cse;
  wire COMP_LOOP_tmp_nor_105_cse;
  wire COMP_LOOP_tmp_nor_35_cse;
  wire COMP_LOOP_or_39_cse;
  wire COMP_LOOP_tmp_nor_78_cse;
  wire COMP_LOOP_tmp_nor_79_cse;
  wire COMP_LOOP_tmp_nor_81_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_48_cse;
  wire COMP_LOOP_or_42_cse;
  wire nor_489_cse;
  wire nor_480_cse;
  wire nor_479_cse;
  wire nor_461_cse;
  wire nor_460_cse;
  wire nor_450_cse;
  wire nor_441_cse;
  wire nor_440_cse;
  wire nor_422_cse;
  wire nor_421_cse;
  wire nor_411_cse;
  wire nor_402_cse;
  wire nor_401_cse;
  wire nor_383_cse;
  wire nor_382_cse;
  wire nor_372_cse;
  wire nor_363_cse;
  wire nor_362_cse;
  wire nor_347_cse;
  wire and_325_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_36_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_38_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_39_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_42_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_43_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_45_cse;
  wire and_628_cse;
  wire and_605_cse;
  wire and_609_cse;
  wire and_614_cse;
  wire and_617_cse;
  wire and_621_cse;
  wire and_624_cse;
  wire or_tmp_2098;
  wire mux_tmp_1564;
  wire COMP_LOOP_or_36_itm;
  wire COMP_LOOP_or_33_itm;
  wire COMP_LOOP_tmp_or_71_itm;
  wire [9:0] COMP_LOOP_1_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_2_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_3_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_4_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_5_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_6_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_7_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_8_acc_10_itm_10_1_1;
  wire COMP_LOOP_tmp_or_54_ssc;
  wire [63:0] COMP_LOOP_mux_385_cse;
  wire COMP_LOOP_tmp_nor_135_cse;

  wire[0:0] nor_1019_nl;
  wire[0:0] mux_320_nl;
  wire[0:0] mux_347_nl;
  wire[0:0] nand_11_nl;
  wire[0:0] nand_22_nl;
  wire[0:0] mux_409_nl;
  wire[0:0] mux_471_nl;
  wire[0:0] nand_33_nl;
  wire[0:0] nand_44_nl;
  wire[0:0] mux_533_nl;
  wire[0:0] mux_595_nl;
  wire[0:0] nand_55_nl;
  wire[0:0] nand_66_nl;
  wire[0:0] mux_657_nl;
  wire[0:0] mux_719_nl;
  wire[0:0] nand_77_nl;
  wire[0:0] nand_88_nl;
  wire[0:0] mux_781_nl;
  wire[0:0] or_1066_nl;
  wire[0:0] or_1064_nl;
  wire[0:0] mux_843_nl;
  wire[0:0] nand_99_nl;
  wire[0:0] nor_730_nl;
  wire[0:0] nor_731_nl;
  wire[0:0] nand_110_nl;
  wire[0:0] mux_905_nl;
  wire[0:0] or_1274_nl;
  wire[0:0] or_1272_nl;
  wire[0:0] mux_967_nl;
  wire[0:0] nand_121_nl;
  wire[0:0] nor_662_nl;
  wire[0:0] nor_663_nl;
  wire[0:0] nand_132_nl;
  wire[0:0] mux_1029_nl;
  wire[0:0] or_1481_nl;
  wire[0:0] or_1480_nl;
  wire[0:0] mux_1091_nl;
  wire[0:0] nand_143_nl;
  wire[0:0] nor_595_nl;
  wire[0:0] nor_596_nl;
  wire[0:0] nand_154_nl;
  wire[0:0] mux_1153_nl;
  wire[0:0] mux_1215_nl;
  wire[0:0] nand_165_nl;
  wire[0:0] nand_176_nl;
  wire[0:0] mux_1277_nl;
  wire[0:0] mux_1461_nl;
  wire[0:0] mux_1460_nl;
  wire[0:0] mux_1457_nl;
  wire[0:0] mux_1456_nl;
  wire[0:0] mux_1455_nl;
  wire[0:0] VEC_LOOP_j_not_1_nl;
  wire[0:0] nor_1160_nl;
  wire[0:0] and_nl;
  wire[0:0] nand_nl;
  wire[0:0] mux_312_nl;
  wire[0:0] nor_1021_nl;
  wire[0:0] and_451_nl;
  wire[0:0] mux_1604_nl;
  wire[0:0] or_2285_nl;
  wire[0:0] mux_1603_nl;
  wire[0:0] or_2284_nl;
  wire[0:0] mux_1602_nl;
  wire[0:0] mux_nl;
  wire[0:0] or_nl;
  wire[0:0] mux_1492_nl;
  wire[0:0] mux_1497_nl;
  wire[0:0] mux_1496_nl;
  wire[0:0] mux_1499_nl;
  wire[0:0] mux_1498_nl;
  wire[0:0] and_260_nl;
  wire[0:0] mux_1500_nl;
  wire[10:0] COMP_LOOP_3_acc_nl;
  wire[11:0] nl_COMP_LOOP_3_acc_nl;
  wire[0:0] mux_1502_nl;
  wire[0:0] mux_1501_nl;
  wire[0:0] and_310_nl;
  wire[0:0] mux_1505_nl;
  wire[0:0] mux_1504_nl;
  wire[0:0] mux_1507_nl;
  wire[0:0] mux_1506_nl;
  wire[8:0] COMP_LOOP_acc_12_nl;
  wire[9:0] nl_COMP_LOOP_acc_12_nl;
  wire[0:0] mux_1509_nl;
  wire[0:0] mux_1508_nl;
  wire[0:0] mux_1511_nl;
  wire[10:0] COMP_LOOP_5_acc_nl;
  wire[11:0] nl_COMP_LOOP_5_acc_nl;
  wire[0:0] mux_1513_nl;
  wire[0:0] mux_1512_nl;
  wire[0:0] mux_1518_nl;
  wire[0:0] mux_1520_nl;
  wire[10:0] COMP_LOOP_6_acc_nl;
  wire[11:0] nl_COMP_LOOP_6_acc_nl;
  wire[0:0] mux_1523_nl;
  wire[10:0] COMP_LOOP_7_acc_nl;
  wire[11:0] nl_COMP_LOOP_7_acc_nl;
  wire[0:0] mux_1528_nl;
  wire[0:0] mux_1532_nl;
  wire[0:0] or_162_nl;
  wire[7:0] COMP_LOOP_acc_15_nl;
  wire[8:0] nl_COMP_LOOP_acc_15_nl;
  wire[0:0] and_305_nl;
  wire[10:0] COMP_LOOP_1_acc_nl;
  wire[11:0] nl_COMP_LOOP_1_acc_nl;
  wire[0:0] and_304_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_33_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_35_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_36_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_37_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_39_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_40_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_41_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_42_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_43_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_44_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_45_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_47_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_48_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_49_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_50_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_51_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_52_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_53_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_54_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_55_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_56_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_57_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_58_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_59_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_60_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_61_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_nor_1_nl;
  wire[0:0] COMP_LOOP_nor_26_nl;
  wire[0:0] COMP_LOOP_nor_27_nl;
  wire[0:0] COMP_LOOP_nor_29_nl;
  wire[0:0] COMP_LOOP_nor_33_nl;
  wire[0:0] COMP_LOOP_nor_40_nl;
  wire[63:0] COMP_LOOP_acc_17_nl;
  wire[64:0] nl_COMP_LOOP_acc_17_nl;
  wire[63:0] COMP_LOOP_COMP_LOOP_mux_2_nl;
  wire[0:0] COMP_LOOP_or_nl;
  wire[0:0] COMP_LOOP_or_1_nl;
  wire[0:0] COMP_LOOP_or_2_nl;
  wire[0:0] COMP_LOOP_or_3_nl;
  wire[0:0] COMP_LOOP_or_4_nl;
  wire[0:0] COMP_LOOP_or_5_nl;
  wire[0:0] COMP_LOOP_or_6_nl;
  wire[0:0] COMP_LOOP_or_7_nl;
  wire[0:0] COMP_LOOP_or_8_nl;
  wire[0:0] COMP_LOOP_or_9_nl;
  wire[0:0] COMP_LOOP_or_10_nl;
  wire[0:0] COMP_LOOP_or_11_nl;
  wire[0:0] COMP_LOOP_or_12_nl;
  wire[0:0] COMP_LOOP_or_13_nl;
  wire[0:0] COMP_LOOP_or_14_nl;
  wire[0:0] COMP_LOOP_or_15_nl;
  wire[0:0] COMP_LOOP_or_16_nl;
  wire[0:0] COMP_LOOP_or_17_nl;
  wire[0:0] COMP_LOOP_or_18_nl;
  wire[0:0] COMP_LOOP_or_19_nl;
  wire[0:0] COMP_LOOP_or_20_nl;
  wire[0:0] COMP_LOOP_or_21_nl;
  wire[0:0] COMP_LOOP_or_22_nl;
  wire[0:0] COMP_LOOP_or_23_nl;
  wire[0:0] COMP_LOOP_or_24_nl;
  wire[0:0] COMP_LOOP_or_25_nl;
  wire[0:0] COMP_LOOP_or_26_nl;
  wire[0:0] COMP_LOOP_or_27_nl;
  wire[0:0] COMP_LOOP_or_28_nl;
  wire[0:0] COMP_LOOP_or_29_nl;
  wire[0:0] COMP_LOOP_or_30_nl;
  wire[0:0] COMP_LOOP_or_31_nl;
  wire[0:0] COMP_LOOP_tmp_and_127_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_nl;
  wire[0:0] COMP_LOOP_tmp_and_128_nl;
  wire[0:0] COMP_LOOP_tmp_and_129_nl;
  wire[0:0] COMP_LOOP_tmp_and_130_nl;
  wire[0:0] COMP_LOOP_tmp_and_131_nl;
  wire[0:0] COMP_LOOP_tmp_and_132_nl;
  wire[0:0] COMP_LOOP_tmp_and_133_nl;
  wire[0:0] COMP_LOOP_tmp_and_134_nl;
  wire[0:0] COMP_LOOP_tmp_and_135_nl;
  wire[0:0] COMP_LOOP_tmp_and_136_nl;
  wire[0:0] COMP_LOOP_tmp_and_137_nl;
  wire[0:0] COMP_LOOP_tmp_and_138_nl;
  wire[0:0] COMP_LOOP_tmp_and_139_nl;
  wire[0:0] COMP_LOOP_tmp_and_140_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_18_nl;
  wire[0:0] COMP_LOOP_tmp_and_141_nl;
  wire[0:0] COMP_LOOP_tmp_and_142_nl;
  wire[0:0] COMP_LOOP_tmp_and_143_nl;
  wire[0:0] COMP_LOOP_tmp_and_144_nl;
  wire[0:0] COMP_LOOP_tmp_and_145_nl;
  wire[0:0] COMP_LOOP_tmp_and_146_nl;
  wire[0:0] COMP_LOOP_tmp_and_147_nl;
  wire[0:0] COMP_LOOP_tmp_and_148_nl;
  wire[0:0] COMP_LOOP_tmp_and_149_nl;
  wire[0:0] COMP_LOOP_tmp_and_150_nl;
  wire[0:0] COMP_LOOP_tmp_and_151_nl;
  wire[0:0] COMP_LOOP_tmp_and_152_nl;
  wire[0:0] COMP_LOOP_tmp_and_153_nl;
  wire[0:0] COMP_LOOP_tmp_and_154_nl;
  wire[0:0] COMP_LOOP_tmp_and_155_nl;
  wire[0:0] COMP_LOOP_tmp_and_115_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_34_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_35_nl;
  wire[0:0] COMP_LOOP_tmp_and_116_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_37_nl;
  wire[0:0] COMP_LOOP_tmp_and_117_nl;
  wire[0:0] COMP_LOOP_tmp_and_118_nl;
  wire[0:0] COMP_LOOP_tmp_and_119_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_41_nl;
  wire[0:0] COMP_LOOP_tmp_and_120_nl;
  wire[0:0] COMP_LOOP_tmp_and_121_nl;
  wire[0:0] COMP_LOOP_tmp_and_122_nl;
  wire[0:0] COMP_LOOP_tmp_and_123_nl;
  wire[0:0] COMP_LOOP_tmp_and_124_nl;
  wire[0:0] COMP_LOOP_tmp_and_125_nl;
  wire[0:0] COMP_LOOP_tmp_and_126_nl;
  wire[0:0] COMP_LOOP_tmp_and_83_nl;
  wire[0:0] COMP_LOOP_tmp_and_84_nl;
  wire[0:0] COMP_LOOP_tmp_and_85_nl;
  wire[0:0] COMP_LOOP_tmp_and_86_nl;
  wire[0:0] COMP_LOOP_tmp_and_87_nl;
  wire[0:0] COMP_LOOP_tmp_and_88_nl;
  wire[0:0] COMP_LOOP_tmp_and_89_nl;
  wire[0:0] COMP_LOOP_tmp_and_90_nl;
  wire[0:0] COMP_LOOP_tmp_and_91_nl;
  wire[0:0] COMP_LOOP_tmp_and_92_nl;
  wire[0:0] COMP_LOOP_tmp_and_93_nl;
  wire[0:0] COMP_LOOP_tmp_and_94_nl;
  wire[0:0] COMP_LOOP_tmp_and_95_nl;
  wire[0:0] COMP_LOOP_tmp_and_96_nl;
  wire[0:0] COMP_LOOP_tmp_and_97_nl;
  wire[0:0] COMP_LOOP_tmp_and_98_nl;
  wire[0:0] COMP_LOOP_tmp_and_99_nl;
  wire[0:0] COMP_LOOP_tmp_and_100_nl;
  wire[0:0] COMP_LOOP_tmp_and_101_nl;
  wire[0:0] COMP_LOOP_tmp_and_102_nl;
  wire[0:0] COMP_LOOP_tmp_and_103_nl;
  wire[0:0] COMP_LOOP_tmp_and_104_nl;
  wire[0:0] COMP_LOOP_tmp_and_105_nl;
  wire[0:0] COMP_LOOP_tmp_and_106_nl;
  wire[0:0] COMP_LOOP_tmp_and_107_nl;
  wire[0:0] COMP_LOOP_tmp_and_108_nl;
  wire[0:0] COMP_LOOP_tmp_and_109_nl;
  wire[0:0] COMP_LOOP_tmp_and_110_nl;
  wire[0:0] COMP_LOOP_tmp_and_111_nl;
  wire[0:0] COMP_LOOP_tmp_and_112_nl;
  wire[0:0] COMP_LOOP_tmp_and_113_nl;
  wire[0:0] COMP_LOOP_tmp_and_114_nl;
  wire[0:0] COMP_LOOP_tmp_and_78_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_80_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_81_nl;
  wire[0:0] COMP_LOOP_tmp_and_79_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_83_nl;
  wire[0:0] COMP_LOOP_tmp_and_80_nl;
  wire[0:0] COMP_LOOP_tmp_and_81_nl;
  wire[0:0] COMP_LOOP_tmp_and_82_nl;
  wire[0:0] COMP_LOOP_tmp_and_47_nl;
  wire[0:0] COMP_LOOP_tmp_and_48_nl;
  wire[0:0] COMP_LOOP_tmp_and_49_nl;
  wire[0:0] COMP_LOOP_tmp_and_50_nl;
  wire[0:0] COMP_LOOP_tmp_and_51_nl;
  wire[0:0] COMP_LOOP_tmp_and_52_nl;
  wire[0:0] COMP_LOOP_tmp_and_53_nl;
  wire[0:0] COMP_LOOP_tmp_and_54_nl;
  wire[0:0] COMP_LOOP_tmp_and_55_nl;
  wire[0:0] COMP_LOOP_tmp_and_56_nl;
  wire[0:0] COMP_LOOP_tmp_and_57_nl;
  wire[0:0] COMP_LOOP_tmp_and_58_nl;
  wire[0:0] COMP_LOOP_tmp_and_59_nl;
  wire[0:0] COMP_LOOP_tmp_and_60_nl;
  wire[0:0] COMP_LOOP_tmp_and_61_nl;
  wire[0:0] COMP_LOOP_tmp_and_62_nl;
  wire[0:0] COMP_LOOP_tmp_and_63_nl;
  wire[0:0] COMP_LOOP_tmp_and_64_nl;
  wire[0:0] COMP_LOOP_tmp_and_65_nl;
  wire[0:0] COMP_LOOP_tmp_and_66_nl;
  wire[0:0] COMP_LOOP_tmp_and_67_nl;
  wire[0:0] COMP_LOOP_tmp_and_68_nl;
  wire[0:0] COMP_LOOP_tmp_and_69_nl;
  wire[0:0] COMP_LOOP_tmp_and_70_nl;
  wire[0:0] COMP_LOOP_tmp_and_71_nl;
  wire[0:0] COMP_LOOP_tmp_and_72_nl;
  wire[0:0] COMP_LOOP_tmp_and_73_nl;
  wire[0:0] COMP_LOOP_tmp_and_74_nl;
  wire[0:0] COMP_LOOP_tmp_and_75_nl;
  wire[0:0] COMP_LOOP_tmp_and_76_nl;
  wire[0:0] COMP_LOOP_tmp_and_77_nl;
  wire[0:0] mux_1585_nl;
  wire[0:0] mux_1584_nl;
  wire[0:0] mux_1583_nl;
  wire[0:0] nor_337_nl;
  wire[0:0] mux_1582_nl;
  wire[0:0] mux_1591_nl;
  wire[0:0] mux_1590_nl;
  wire[0:0] mux_1589_nl;
  wire[0:0] mux_1588_nl;
  wire[0:0] mux_1587_nl;
  wire[0:0] mux_1586_nl;
  wire[0:0] COMP_LOOP_tmp_and_15_nl;
  wire[0:0] COMP_LOOP_tmp_and_16_nl;
  wire[0:0] COMP_LOOP_tmp_and_17_nl;
  wire[0:0] COMP_LOOP_tmp_and_18_nl;
  wire[0:0] COMP_LOOP_tmp_and_19_nl;
  wire[0:0] COMP_LOOP_tmp_and_20_nl;
  wire[0:0] COMP_LOOP_tmp_and_21_nl;
  wire[0:0] COMP_LOOP_tmp_and_22_nl;
  wire[0:0] COMP_LOOP_tmp_and_23_nl;
  wire[0:0] COMP_LOOP_tmp_and_24_nl;
  wire[0:0] COMP_LOOP_tmp_and_25_nl;
  wire[0:0] COMP_LOOP_tmp_and_26_nl;
  wire[0:0] COMP_LOOP_tmp_and_27_nl;
  wire[0:0] COMP_LOOP_tmp_and_28_nl;
  wire[0:0] COMP_LOOP_tmp_and_29_nl;
  wire[0:0] COMP_LOOP_tmp_and_30_nl;
  wire[0:0] COMP_LOOP_tmp_and_31_nl;
  wire[0:0] COMP_LOOP_tmp_and_32_nl;
  wire[0:0] COMP_LOOP_tmp_and_33_nl;
  wire[0:0] COMP_LOOP_tmp_and_34_nl;
  wire[0:0] COMP_LOOP_tmp_and_35_nl;
  wire[0:0] COMP_LOOP_tmp_and_36_nl;
  wire[0:0] COMP_LOOP_tmp_and_37_nl;
  wire[0:0] COMP_LOOP_tmp_and_38_nl;
  wire[0:0] COMP_LOOP_tmp_and_39_nl;
  wire[0:0] COMP_LOOP_tmp_and_40_nl;
  wire[0:0] COMP_LOOP_tmp_and_41_nl;
  wire[0:0] COMP_LOOP_tmp_and_42_nl;
  wire[0:0] COMP_LOOP_tmp_and_43_nl;
  wire[0:0] COMP_LOOP_tmp_and_44_nl;
  wire[0:0] COMP_LOOP_tmp_and_45_nl;
  wire[0:0] COMP_LOOP_tmp_and_46_nl;
  wire[0:0] COMP_LOOP_tmp_and_nl;
  wire[0:0] COMP_LOOP_tmp_and_1_nl;
  wire[0:0] COMP_LOOP_tmp_and_2_nl;
  wire[0:0] COMP_LOOP_tmp_and_3_nl;
  wire[0:0] COMP_LOOP_tmp_and_4_nl;
  wire[0:0] COMP_LOOP_tmp_and_5_nl;
  wire[0:0] COMP_LOOP_tmp_and_6_nl;
  wire[0:0] COMP_LOOP_tmp_and_7_nl;
  wire[0:0] COMP_LOOP_tmp_and_8_nl;
  wire[0:0] COMP_LOOP_tmp_and_9_nl;
  wire[0:0] COMP_LOOP_tmp_and_10_nl;
  wire[0:0] COMP_LOOP_tmp_and_11_nl;
  wire[0:0] COMP_LOOP_tmp_and_12_nl;
  wire[0:0] COMP_LOOP_tmp_and_13_nl;
  wire[0:0] COMP_LOOP_tmp_and_14_nl;
  wire[0:0] mux_1597_nl;
  wire[0:0] mux_1596_nl;
  wire[0:0] mux_1595_nl;
  wire[0:0] mux_1594_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] and_478_nl;
  wire[10:0] COMP_LOOP_1_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_1_acc_10_nl;
  wire[10:0] COMP_LOOP_2_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_2_acc_10_nl;
  wire[10:0] COMP_LOOP_3_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_3_acc_10_nl;
  wire[10:0] COMP_LOOP_4_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_4_acc_10_nl;
  wire[10:0] COMP_LOOP_5_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_5_acc_10_nl;
  wire[10:0] COMP_LOOP_6_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_6_acc_10_nl;
  wire[10:0] COMP_LOOP_7_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_7_acc_10_nl;
  wire[10:0] COMP_LOOP_8_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_8_acc_10_nl;
  wire[0:0] or_238_nl;
  wire[0:0] or_236_nl;
  wire[0:0] or_284_nl;
  wire[0:0] or_282_nl;
  wire[0:0] nor_1001_nl;
  wire[0:0] nor_1002_nl;
  wire[0:0] or_388_nl;
  wire[0:0] or_386_nl;
  wire[0:0] or_446_nl;
  wire[0:0] or_444_nl;
  wire[0:0] or_492_nl;
  wire[0:0] or_490_nl;
  wire[0:0] nor_933_nl;
  wire[0:0] nor_934_nl;
  wire[0:0] or_596_nl;
  wire[0:0] or_594_nl;
  wire[0:0] or_654_nl;
  wire[0:0] or_652_nl;
  wire[0:0] or_700_nl;
  wire[0:0] or_698_nl;
  wire[0:0] nor_865_nl;
  wire[0:0] nor_866_nl;
  wire[0:0] or_804_nl;
  wire[0:0] or_802_nl;
  wire[0:0] nand_518_nl;
  wire[0:0] or_860_nl;
  wire[0:0] or_908_nl;
  wire[0:0] or_906_nl;
  wire[0:0] and_532_nl;
  wire[0:0] nor_798_nl;
  wire[0:0] nand_472_nl;
  wire[0:0] or_1009_nl;
  wire[0:0] or_1112_nl;
  wire[0:0] or_1110_nl;
  wire[0:0] or_1216_nl;
  wire[0:0] or_1214_nl;
  wire[0:0] or_1320_nl;
  wire[0:0] or_1318_nl;
  wire[0:0] nand_469_nl;
  wire[0:0] or_1422_nl;
  wire[0:0] or_1527_nl;
  wire[0:0] or_1525_nl;
  wire[0:0] nand_466_nl;
  wire[0:0] or_1627_nl;
  wire[0:0] nand_268_nl;
  wire[0:0] nand_269_nl;
  wire[0:0] nand_463_nl;
  wire[0:0] or_1727_nl;
  wire[0:0] and_353_nl;
  wire[0:0] and_354_nl;
  wire[0:0] nand_459_nl;
  wire[0:0] nand_236_nl;
  wire[0:0] mux_1470_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] or_2109_nl;
  wire[0:0] mux_1488_nl;
  wire[0:0] mux_1486_nl;
  wire[0:0] mux_1490_nl;
  wire[0:0] and_448_nl;
  wire[0:0] mux_1606_nl;
  wire[0:0] nor_340_nl;
  wire[0:0] and_511_nl;
  wire[0:0] mux_1510_nl;
  wire[0:0] nand_188_nl;
  wire[0:0] mux_1515_nl;
  wire[0:0] mux_1514_nl;
  wire[0:0] mux_1516_nl;
  wire[0:0] mux_1599_nl;
  wire[0:0] and_446_nl;
  wire[0:0] mux_1526_nl;
  wire[0:0] mux_1525_nl;
  wire[0:0] mux_1530_nl;
  wire[0:0] mux_1535_nl;
  wire[0:0] and_306_nl;
  wire[0:0] mux_1537_nl;
  wire[0:0] mux_1542_nl;
  wire[0:0] mux_1551_nl;
  wire[0:0] nor_1128_nl;
  wire[0:0] nor_1129_nl;
  wire[0:0] mux_1555_nl;
  wire[0:0] mux_1554_nl;
  wire[0:0] mux_1553_nl;
  wire[0:0] nand_185_nl;
  wire[0:0] mux_1552_nl;
  wire[0:0] nand_473_nl;
  wire[0:0] or_2171_nl;
  wire[0:0] mux_1575_nl;
  wire[0:0] mux_1574_nl;
  wire[0:0] or_229_nl;
  wire[0:0] mux_1573_nl;
  wire[0:0] mux_1579_nl;
  wire[0:0] mux_1578_nl;
  wire[0:0] mux_1577_nl;
  wire[0:0] mux_1576_nl;
  wire[0:0] nor_1059_nl;
  wire[0:0] mux_1581_nl;
  wire[0:0] mux_1580_nl;
  wire[0:0] nor_1062_nl;
  wire[0:0] nor_1063_nl;
  wire[0:0] and_520_nl;
  wire[0:0] and_54_nl;
  wire[0:0] and_64_nl;
  wire[0:0] and_68_nl;
  wire[0:0] and_74_nl;
  wire[0:0] and_78_nl;
  wire[0:0] and_84_nl;
  wire[0:0] and_88_nl;
  wire[0:0] and_92_nl;
  wire[0:0] and_95_nl;
  wire[0:0] and_97_nl;
  wire[0:0] and_98_nl;
  wire[0:0] and_99_nl;
  wire[0:0] and_101_nl;
  wire[0:0] and_103_nl;
  wire[0:0] and_104_nl;
  wire[0:0] and_105_nl;
  wire[0:0] and_107_nl;
  wire[0:0] and_109_nl;
  wire[0:0] and_110_nl;
  wire[0:0] and_111_nl;
  wire[0:0] and_112_nl;
  wire[0:0] and_114_nl;
  wire[0:0] and_116_nl;
  wire[0:0] and_117_nl;
  wire[0:0] mux_336_nl;
  wire[0:0] nand_506_nl;
  wire[0:0] mux_335_nl;
  wire[0:0] and_443_nl;
  wire[0:0] mux_334_nl;
  wire[0:0] mux_333_nl;
  wire[0:0] nor_1010_nl;
  wire[0:0] nor_1011_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] nor_1012_nl;
  wire[0:0] nor_1013_nl;
  wire[0:0] nor_1014_nl;
  wire[0:0] mux_331_nl;
  wire[0:0] mux_330_nl;
  wire[0:0] or_257_nl;
  wire[0:0] or_255_nl;
  wire[0:0] mux_329_nl;
  wire[0:0] or_254_nl;
  wire[0:0] or_252_nl;
  wire[0:0] or_2280_nl;
  wire[0:0] mux_328_nl;
  wire[0:0] nand_8_nl;
  wire[0:0] mux_327_nl;
  wire[0:0] mux_326_nl;
  wire[0:0] nor_1016_nl;
  wire[0:0] nor_1017_nl;
  wire[0:0] nor_1018_nl;
  wire[0:0] mux_325_nl;
  wire[0:0] or_246_nl;
  wire[0:0] or_244_nl;
  wire[0:0] or_243_nl;
  wire[0:0] mux_324_nl;
  wire[0:0] mux_323_nl;
  wire[0:0] or_242_nl;
  wire[0:0] or_240_nl;
  wire[0:0] or_239_nl;
  wire[0:0] mux_352_nl;
  wire[0:0] mux_351_nl;
  wire[0:0] mux_350_nl;
  wire[0:0] nor_1003_nl;
  wire[0:0] nor_1004_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] nor_1005_nl;
  wire[0:0] mux_345_nl;
  wire[0:0] nor_1006_nl;
  wire[0:0] mux_344_nl;
  wire[0:0] nor_1007_nl;
  wire[0:0] nor_1008_nl;
  wire[0:0] nor_1009_nl;
  wire[0:0] mux_343_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] mux_341_nl;
  wire[0:0] or_276_nl;
  wire[0:0] or_274_nl;
  wire[0:0] mux_340_nl;
  wire[0:0] or_273_nl;
  wire[0:0] or_271_nl;
  wire[0:0] mux_339_nl;
  wire[0:0] mux_338_nl;
  wire[0:0] or_270_nl;
  wire[0:0] or_268_nl;
  wire[0:0] mux_337_nl;
  wire[0:0] or_267_nl;
  wire[0:0] or_265_nl;
  wire[0:0] mux_367_nl;
  wire[0:0] nand_505_nl;
  wire[0:0] mux_366_nl;
  wire[0:0] and_440_nl;
  wire[0:0] mux_365_nl;
  wire[0:0] mux_364_nl;
  wire[0:0] nor_991_nl;
  wire[0:0] nor_992_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] nor_993_nl;
  wire[0:0] nor_994_nl;
  wire[0:0] nor_995_nl;
  wire[0:0] mux_362_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] or_308_nl;
  wire[0:0] or_306_nl;
  wire[0:0] mux_360_nl;
  wire[0:0] or_305_nl;
  wire[0:0] or_303_nl;
  wire[0:0] or_2279_nl;
  wire[0:0] mux_359_nl;
  wire[0:0] nand_14_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] mux_357_nl;
  wire[0:0] nor_997_nl;
  wire[0:0] nor_998_nl;
  wire[0:0] and_441_nl;
  wire[0:0] mux_356_nl;
  wire[0:0] nor_999_nl;
  wire[0:0] nor_1000_nl;
  wire[0:0] or_295_nl;
  wire[0:0] mux_355_nl;
  wire[0:0] mux_354_nl;
  wire[0:0] or_294_nl;
  wire[0:0] or_292_nl;
  wire[0:0] nand_12_nl;
  wire[0:0] mux_383_nl;
  wire[0:0] mux_382_nl;
  wire[0:0] mux_381_nl;
  wire[0:0] nor_985_nl;
  wire[0:0] nor_986_nl;
  wire[0:0] mux_380_nl;
  wire[0:0] and_438_nl;
  wire[0:0] mux_376_nl;
  wire[0:0] nor_987_nl;
  wire[0:0] mux_375_nl;
  wire[0:0] nor_988_nl;
  wire[0:0] nor_989_nl;
  wire[0:0] nor_990_nl;
  wire[0:0] mux_374_nl;
  wire[0:0] mux_373_nl;
  wire[0:0] mux_372_nl;
  wire[0:0] or_327_nl;
  wire[0:0] or_325_nl;
  wire[0:0] mux_371_nl;
  wire[0:0] or_324_nl;
  wire[0:0] or_322_nl;
  wire[0:0] mux_370_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] or_321_nl;
  wire[0:0] or_319_nl;
  wire[0:0] mux_368_nl;
  wire[0:0] or_318_nl;
  wire[0:0] or_316_nl;
  wire[0:0] mux_398_nl;
  wire[0:0] nand_504_nl;
  wire[0:0] mux_397_nl;
  wire[0:0] and_437_nl;
  wire[0:0] mux_396_nl;
  wire[0:0] mux_395_nl;
  wire[0:0] nor_976_nl;
  wire[0:0] nor_977_nl;
  wire[0:0] mux_394_nl;
  wire[0:0] nor_978_nl;
  wire[0:0] nor_979_nl;
  wire[0:0] nor_980_nl;
  wire[0:0] mux_393_nl;
  wire[0:0] mux_392_nl;
  wire[0:0] or_361_nl;
  wire[0:0] or_359_nl;
  wire[0:0] mux_391_nl;
  wire[0:0] or_358_nl;
  wire[0:0] or_356_nl;
  wire[0:0] or_2278_nl;
  wire[0:0] mux_390_nl;
  wire[0:0] nand_19_nl;
  wire[0:0] mux_389_nl;
  wire[0:0] mux_388_nl;
  wire[0:0] nor_982_nl;
  wire[0:0] nor_983_nl;
  wire[0:0] nor_984_nl;
  wire[0:0] mux_387_nl;
  wire[0:0] or_350_nl;
  wire[0:0] or_348_nl;
  wire[0:0] or_347_nl;
  wire[0:0] mux_386_nl;
  wire[0:0] mux_385_nl;
  wire[0:0] or_346_nl;
  wire[0:0] or_344_nl;
  wire[0:0] or_343_nl;
  wire[0:0] mux_414_nl;
  wire[0:0] mux_413_nl;
  wire[0:0] mux_412_nl;
  wire[0:0] nor_969_nl;
  wire[0:0] nor_970_nl;
  wire[0:0] mux_411_nl;
  wire[0:0] nor_971_nl;
  wire[0:0] mux_407_nl;
  wire[0:0] nor_972_nl;
  wire[0:0] mux_406_nl;
  wire[0:0] nor_973_nl;
  wire[0:0] nor_974_nl;
  wire[0:0] nor_975_nl;
  wire[0:0] mux_405_nl;
  wire[0:0] mux_404_nl;
  wire[0:0] mux_403_nl;
  wire[0:0] or_380_nl;
  wire[0:0] or_378_nl;
  wire[0:0] mux_402_nl;
  wire[0:0] or_377_nl;
  wire[0:0] or_375_nl;
  wire[0:0] mux_401_nl;
  wire[0:0] mux_400_nl;
  wire[0:0] or_374_nl;
  wire[0:0] or_372_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] or_371_nl;
  wire[0:0] or_369_nl;
  wire[0:0] mux_429_nl;
  wire[0:0] nand_503_nl;
  wire[0:0] mux_428_nl;
  wire[0:0] and_434_nl;
  wire[0:0] mux_427_nl;
  wire[0:0] mux_426_nl;
  wire[0:0] nor_957_nl;
  wire[0:0] nor_958_nl;
  wire[0:0] mux_425_nl;
  wire[0:0] nor_959_nl;
  wire[0:0] nor_960_nl;
  wire[0:0] nor_961_nl;
  wire[0:0] mux_424_nl;
  wire[0:0] mux_423_nl;
  wire[0:0] or_412_nl;
  wire[0:0] or_410_nl;
  wire[0:0] mux_422_nl;
  wire[0:0] or_409_nl;
  wire[0:0] or_407_nl;
  wire[0:0] or_2277_nl;
  wire[0:0] mux_421_nl;
  wire[0:0] nand_25_nl;
  wire[0:0] mux_420_nl;
  wire[0:0] mux_419_nl;
  wire[0:0] nor_963_nl;
  wire[0:0] nor_964_nl;
  wire[0:0] and_435_nl;
  wire[0:0] mux_418_nl;
  wire[0:0] nor_965_nl;
  wire[0:0] nor_966_nl;
  wire[0:0] or_399_nl;
  wire[0:0] mux_417_nl;
  wire[0:0] mux_416_nl;
  wire[0:0] or_398_nl;
  wire[0:0] or_396_nl;
  wire[0:0] nand_23_nl;
  wire[0:0] mux_445_nl;
  wire[0:0] mux_444_nl;
  wire[0:0] mux_443_nl;
  wire[0:0] nor_951_nl;
  wire[0:0] nor_952_nl;
  wire[0:0] mux_442_nl;
  wire[0:0] and_432_nl;
  wire[0:0] mux_438_nl;
  wire[0:0] nor_953_nl;
  wire[0:0] mux_437_nl;
  wire[0:0] nor_954_nl;
  wire[0:0] nor_955_nl;
  wire[0:0] nor_956_nl;
  wire[0:0] mux_436_nl;
  wire[0:0] mux_435_nl;
  wire[0:0] mux_434_nl;
  wire[0:0] or_431_nl;
  wire[0:0] or_429_nl;
  wire[0:0] mux_433_nl;
  wire[0:0] or_428_nl;
  wire[0:0] or_426_nl;
  wire[0:0] mux_432_nl;
  wire[0:0] mux_431_nl;
  wire[0:0] or_425_nl;
  wire[0:0] or_423_nl;
  wire[0:0] mux_430_nl;
  wire[0:0] or_422_nl;
  wire[0:0] or_420_nl;
  wire[0:0] mux_460_nl;
  wire[0:0] nand_502_nl;
  wire[0:0] mux_459_nl;
  wire[0:0] and_431_nl;
  wire[0:0] mux_458_nl;
  wire[0:0] mux_457_nl;
  wire[0:0] nor_942_nl;
  wire[0:0] nor_943_nl;
  wire[0:0] mux_456_nl;
  wire[0:0] nor_944_nl;
  wire[0:0] nor_945_nl;
  wire[0:0] nor_946_nl;
  wire[0:0] mux_455_nl;
  wire[0:0] mux_454_nl;
  wire[0:0] or_465_nl;
  wire[0:0] or_463_nl;
  wire[0:0] mux_453_nl;
  wire[0:0] or_462_nl;
  wire[0:0] or_460_nl;
  wire[0:0] or_2276_nl;
  wire[0:0] mux_452_nl;
  wire[0:0] nand_30_nl;
  wire[0:0] mux_451_nl;
  wire[0:0] mux_450_nl;
  wire[0:0] nor_948_nl;
  wire[0:0] nor_949_nl;
  wire[0:0] nor_950_nl;
  wire[0:0] mux_449_nl;
  wire[0:0] or_454_nl;
  wire[0:0] or_452_nl;
  wire[0:0] or_451_nl;
  wire[0:0] mux_448_nl;
  wire[0:0] mux_447_nl;
  wire[0:0] or_450_nl;
  wire[0:0] or_448_nl;
  wire[0:0] or_447_nl;
  wire[0:0] mux_476_nl;
  wire[0:0] mux_475_nl;
  wire[0:0] mux_474_nl;
  wire[0:0] nor_935_nl;
  wire[0:0] nor_936_nl;
  wire[0:0] mux_473_nl;
  wire[0:0] nor_937_nl;
  wire[0:0] mux_469_nl;
  wire[0:0] nor_938_nl;
  wire[0:0] mux_468_nl;
  wire[0:0] nor_939_nl;
  wire[0:0] nor_940_nl;
  wire[0:0] nor_941_nl;
  wire[0:0] mux_467_nl;
  wire[0:0] mux_466_nl;
  wire[0:0] mux_465_nl;
  wire[0:0] or_484_nl;
  wire[0:0] or_482_nl;
  wire[0:0] mux_464_nl;
  wire[0:0] or_481_nl;
  wire[0:0] or_479_nl;
  wire[0:0] mux_463_nl;
  wire[0:0] mux_462_nl;
  wire[0:0] or_478_nl;
  wire[0:0] or_476_nl;
  wire[0:0] mux_461_nl;
  wire[0:0] or_475_nl;
  wire[0:0] or_473_nl;
  wire[0:0] mux_491_nl;
  wire[0:0] nand_501_nl;
  wire[0:0] mux_490_nl;
  wire[0:0] and_428_nl;
  wire[0:0] mux_489_nl;
  wire[0:0] mux_488_nl;
  wire[0:0] nor_923_nl;
  wire[0:0] nor_924_nl;
  wire[0:0] mux_487_nl;
  wire[0:0] nor_925_nl;
  wire[0:0] nor_926_nl;
  wire[0:0] nor_927_nl;
  wire[0:0] mux_486_nl;
  wire[0:0] mux_485_nl;
  wire[0:0] or_516_nl;
  wire[0:0] or_514_nl;
  wire[0:0] mux_484_nl;
  wire[0:0] or_513_nl;
  wire[0:0] or_511_nl;
  wire[0:0] or_2275_nl;
  wire[0:0] mux_483_nl;
  wire[0:0] nand_36_nl;
  wire[0:0] mux_482_nl;
  wire[0:0] mux_481_nl;
  wire[0:0] nor_929_nl;
  wire[0:0] nor_930_nl;
  wire[0:0] and_429_nl;
  wire[0:0] mux_480_nl;
  wire[0:0] nor_931_nl;
  wire[0:0] nor_932_nl;
  wire[0:0] or_503_nl;
  wire[0:0] mux_479_nl;
  wire[0:0] mux_478_nl;
  wire[0:0] or_502_nl;
  wire[0:0] or_500_nl;
  wire[0:0] nand_34_nl;
  wire[0:0] mux_507_nl;
  wire[0:0] mux_506_nl;
  wire[0:0] mux_505_nl;
  wire[0:0] nor_917_nl;
  wire[0:0] nor_918_nl;
  wire[0:0] mux_504_nl;
  wire[0:0] and_426_nl;
  wire[0:0] mux_500_nl;
  wire[0:0] nor_919_nl;
  wire[0:0] mux_499_nl;
  wire[0:0] nor_920_nl;
  wire[0:0] nor_921_nl;
  wire[0:0] nor_922_nl;
  wire[0:0] mux_498_nl;
  wire[0:0] mux_497_nl;
  wire[0:0] mux_496_nl;
  wire[0:0] or_535_nl;
  wire[0:0] or_533_nl;
  wire[0:0] mux_495_nl;
  wire[0:0] or_532_nl;
  wire[0:0] or_530_nl;
  wire[0:0] mux_494_nl;
  wire[0:0] mux_493_nl;
  wire[0:0] or_529_nl;
  wire[0:0] or_527_nl;
  wire[0:0] mux_492_nl;
  wire[0:0] or_526_nl;
  wire[0:0] or_524_nl;
  wire[0:0] mux_522_nl;
  wire[0:0] nand_500_nl;
  wire[0:0] mux_521_nl;
  wire[0:0] and_425_nl;
  wire[0:0] mux_520_nl;
  wire[0:0] mux_519_nl;
  wire[0:0] nor_908_nl;
  wire[0:0] nor_909_nl;
  wire[0:0] mux_518_nl;
  wire[0:0] nor_910_nl;
  wire[0:0] nor_911_nl;
  wire[0:0] nor_912_nl;
  wire[0:0] mux_517_nl;
  wire[0:0] mux_516_nl;
  wire[0:0] or_569_nl;
  wire[0:0] or_567_nl;
  wire[0:0] mux_515_nl;
  wire[0:0] or_566_nl;
  wire[0:0] or_564_nl;
  wire[0:0] or_2274_nl;
  wire[0:0] mux_514_nl;
  wire[0:0] nand_41_nl;
  wire[0:0] mux_513_nl;
  wire[0:0] mux_512_nl;
  wire[0:0] nor_914_nl;
  wire[0:0] nor_915_nl;
  wire[0:0] nor_916_nl;
  wire[0:0] mux_511_nl;
  wire[0:0] or_558_nl;
  wire[0:0] or_556_nl;
  wire[0:0] or_555_nl;
  wire[0:0] mux_510_nl;
  wire[0:0] mux_509_nl;
  wire[0:0] or_554_nl;
  wire[0:0] or_552_nl;
  wire[0:0] or_551_nl;
  wire[0:0] mux_538_nl;
  wire[0:0] mux_537_nl;
  wire[0:0] mux_536_nl;
  wire[0:0] nor_901_nl;
  wire[0:0] nor_902_nl;
  wire[0:0] mux_535_nl;
  wire[0:0] nor_903_nl;
  wire[0:0] mux_531_nl;
  wire[0:0] nor_904_nl;
  wire[0:0] mux_530_nl;
  wire[0:0] nor_905_nl;
  wire[0:0] nor_906_nl;
  wire[0:0] nor_907_nl;
  wire[0:0] mux_529_nl;
  wire[0:0] mux_528_nl;
  wire[0:0] mux_527_nl;
  wire[0:0] or_588_nl;
  wire[0:0] or_586_nl;
  wire[0:0] mux_526_nl;
  wire[0:0] or_585_nl;
  wire[0:0] or_583_nl;
  wire[0:0] mux_525_nl;
  wire[0:0] mux_524_nl;
  wire[0:0] or_582_nl;
  wire[0:0] or_580_nl;
  wire[0:0] mux_523_nl;
  wire[0:0] or_579_nl;
  wire[0:0] or_577_nl;
  wire[0:0] mux_553_nl;
  wire[0:0] nand_499_nl;
  wire[0:0] mux_552_nl;
  wire[0:0] and_422_nl;
  wire[0:0] mux_551_nl;
  wire[0:0] mux_550_nl;
  wire[0:0] nor_889_nl;
  wire[0:0] nor_890_nl;
  wire[0:0] mux_549_nl;
  wire[0:0] nor_891_nl;
  wire[0:0] nor_892_nl;
  wire[0:0] nor_893_nl;
  wire[0:0] mux_548_nl;
  wire[0:0] mux_547_nl;
  wire[0:0] or_620_nl;
  wire[0:0] or_618_nl;
  wire[0:0] mux_546_nl;
  wire[0:0] or_617_nl;
  wire[0:0] or_615_nl;
  wire[0:0] or_2273_nl;
  wire[0:0] mux_545_nl;
  wire[0:0] nand_47_nl;
  wire[0:0] mux_544_nl;
  wire[0:0] mux_543_nl;
  wire[0:0] nor_895_nl;
  wire[0:0] nor_896_nl;
  wire[0:0] and_423_nl;
  wire[0:0] mux_542_nl;
  wire[0:0] nor_897_nl;
  wire[0:0] nor_898_nl;
  wire[0:0] or_607_nl;
  wire[0:0] mux_541_nl;
  wire[0:0] mux_540_nl;
  wire[0:0] or_606_nl;
  wire[0:0] or_604_nl;
  wire[0:0] nand_45_nl;
  wire[0:0] mux_569_nl;
  wire[0:0] mux_568_nl;
  wire[0:0] mux_567_nl;
  wire[0:0] nor_883_nl;
  wire[0:0] nor_884_nl;
  wire[0:0] mux_566_nl;
  wire[0:0] and_420_nl;
  wire[0:0] mux_562_nl;
  wire[0:0] nor_885_nl;
  wire[0:0] mux_561_nl;
  wire[0:0] nor_886_nl;
  wire[0:0] nor_887_nl;
  wire[0:0] nor_888_nl;
  wire[0:0] mux_560_nl;
  wire[0:0] mux_559_nl;
  wire[0:0] mux_558_nl;
  wire[0:0] or_639_nl;
  wire[0:0] or_637_nl;
  wire[0:0] mux_557_nl;
  wire[0:0] or_636_nl;
  wire[0:0] or_634_nl;
  wire[0:0] mux_556_nl;
  wire[0:0] mux_555_nl;
  wire[0:0] or_633_nl;
  wire[0:0] or_631_nl;
  wire[0:0] mux_554_nl;
  wire[0:0] or_630_nl;
  wire[0:0] or_628_nl;
  wire[0:0] mux_584_nl;
  wire[0:0] nand_498_nl;
  wire[0:0] mux_583_nl;
  wire[0:0] and_419_nl;
  wire[0:0] mux_582_nl;
  wire[0:0] mux_581_nl;
  wire[0:0] nor_874_nl;
  wire[0:0] nor_875_nl;
  wire[0:0] mux_580_nl;
  wire[0:0] nor_876_nl;
  wire[0:0] nor_877_nl;
  wire[0:0] nor_878_nl;
  wire[0:0] mux_579_nl;
  wire[0:0] mux_578_nl;
  wire[0:0] or_673_nl;
  wire[0:0] or_671_nl;
  wire[0:0] mux_577_nl;
  wire[0:0] or_670_nl;
  wire[0:0] or_668_nl;
  wire[0:0] or_2272_nl;
  wire[0:0] mux_576_nl;
  wire[0:0] nand_52_nl;
  wire[0:0] mux_575_nl;
  wire[0:0] mux_574_nl;
  wire[0:0] nor_880_nl;
  wire[0:0] nor_881_nl;
  wire[0:0] nor_882_nl;
  wire[0:0] mux_573_nl;
  wire[0:0] or_662_nl;
  wire[0:0] or_660_nl;
  wire[0:0] or_659_nl;
  wire[0:0] mux_572_nl;
  wire[0:0] mux_571_nl;
  wire[0:0] or_658_nl;
  wire[0:0] or_656_nl;
  wire[0:0] or_655_nl;
  wire[0:0] mux_600_nl;
  wire[0:0] mux_599_nl;
  wire[0:0] mux_598_nl;
  wire[0:0] nor_867_nl;
  wire[0:0] nor_868_nl;
  wire[0:0] mux_597_nl;
  wire[0:0] nor_869_nl;
  wire[0:0] mux_593_nl;
  wire[0:0] nor_870_nl;
  wire[0:0] mux_592_nl;
  wire[0:0] nor_871_nl;
  wire[0:0] nor_872_nl;
  wire[0:0] nor_873_nl;
  wire[0:0] mux_591_nl;
  wire[0:0] mux_590_nl;
  wire[0:0] mux_589_nl;
  wire[0:0] or_692_nl;
  wire[0:0] or_690_nl;
  wire[0:0] mux_588_nl;
  wire[0:0] or_689_nl;
  wire[0:0] or_687_nl;
  wire[0:0] mux_587_nl;
  wire[0:0] mux_586_nl;
  wire[0:0] or_686_nl;
  wire[0:0] or_684_nl;
  wire[0:0] mux_585_nl;
  wire[0:0] or_683_nl;
  wire[0:0] or_681_nl;
  wire[0:0] mux_615_nl;
  wire[0:0] nand_497_nl;
  wire[0:0] mux_614_nl;
  wire[0:0] and_416_nl;
  wire[0:0] mux_613_nl;
  wire[0:0] mux_612_nl;
  wire[0:0] nor_855_nl;
  wire[0:0] nor_856_nl;
  wire[0:0] mux_611_nl;
  wire[0:0] nor_857_nl;
  wire[0:0] nor_858_nl;
  wire[0:0] nor_859_nl;
  wire[0:0] mux_610_nl;
  wire[0:0] mux_609_nl;
  wire[0:0] or_724_nl;
  wire[0:0] or_722_nl;
  wire[0:0] mux_608_nl;
  wire[0:0] or_721_nl;
  wire[0:0] or_719_nl;
  wire[0:0] or_2271_nl;
  wire[0:0] mux_607_nl;
  wire[0:0] nand_58_nl;
  wire[0:0] mux_606_nl;
  wire[0:0] mux_605_nl;
  wire[0:0] nor_861_nl;
  wire[0:0] nor_862_nl;
  wire[0:0] and_417_nl;
  wire[0:0] mux_604_nl;
  wire[0:0] nor_863_nl;
  wire[0:0] nor_864_nl;
  wire[0:0] or_711_nl;
  wire[0:0] mux_603_nl;
  wire[0:0] mux_602_nl;
  wire[0:0] or_710_nl;
  wire[0:0] or_708_nl;
  wire[0:0] nand_56_nl;
  wire[0:0] mux_631_nl;
  wire[0:0] mux_630_nl;
  wire[0:0] mux_629_nl;
  wire[0:0] nor_849_nl;
  wire[0:0] nor_850_nl;
  wire[0:0] mux_628_nl;
  wire[0:0] and_414_nl;
  wire[0:0] mux_624_nl;
  wire[0:0] nor_851_nl;
  wire[0:0] mux_623_nl;
  wire[0:0] nor_852_nl;
  wire[0:0] nor_853_nl;
  wire[0:0] nor_854_nl;
  wire[0:0] mux_622_nl;
  wire[0:0] mux_621_nl;
  wire[0:0] mux_620_nl;
  wire[0:0] or_743_nl;
  wire[0:0] or_741_nl;
  wire[0:0] mux_619_nl;
  wire[0:0] or_740_nl;
  wire[0:0] or_738_nl;
  wire[0:0] mux_618_nl;
  wire[0:0] mux_617_nl;
  wire[0:0] or_737_nl;
  wire[0:0] or_735_nl;
  wire[0:0] mux_616_nl;
  wire[0:0] or_734_nl;
  wire[0:0] or_732_nl;
  wire[0:0] mux_646_nl;
  wire[0:0] nand_496_nl;
  wire[0:0] mux_645_nl;
  wire[0:0] and_413_nl;
  wire[0:0] mux_644_nl;
  wire[0:0] mux_643_nl;
  wire[0:0] nor_840_nl;
  wire[0:0] nor_841_nl;
  wire[0:0] mux_642_nl;
  wire[0:0] nor_842_nl;
  wire[0:0] nor_843_nl;
  wire[0:0] nor_844_nl;
  wire[0:0] mux_641_nl;
  wire[0:0] mux_640_nl;
  wire[0:0] or_777_nl;
  wire[0:0] or_775_nl;
  wire[0:0] mux_639_nl;
  wire[0:0] or_774_nl;
  wire[0:0] or_772_nl;
  wire[0:0] or_2270_nl;
  wire[0:0] mux_638_nl;
  wire[0:0] nand_63_nl;
  wire[0:0] mux_637_nl;
  wire[0:0] mux_636_nl;
  wire[0:0] nor_846_nl;
  wire[0:0] nor_847_nl;
  wire[0:0] nor_848_nl;
  wire[0:0] mux_635_nl;
  wire[0:0] or_766_nl;
  wire[0:0] or_764_nl;
  wire[0:0] or_763_nl;
  wire[0:0] mux_634_nl;
  wire[0:0] mux_633_nl;
  wire[0:0] or_762_nl;
  wire[0:0] or_760_nl;
  wire[0:0] or_759_nl;
  wire[0:0] mux_662_nl;
  wire[0:0] mux_661_nl;
  wire[0:0] mux_660_nl;
  wire[0:0] nor_833_nl;
  wire[0:0] nor_834_nl;
  wire[0:0] mux_659_nl;
  wire[0:0] nor_835_nl;
  wire[0:0] mux_655_nl;
  wire[0:0] nor_836_nl;
  wire[0:0] mux_654_nl;
  wire[0:0] nor_837_nl;
  wire[0:0] nor_838_nl;
  wire[0:0] nor_839_nl;
  wire[0:0] mux_653_nl;
  wire[0:0] mux_652_nl;
  wire[0:0] mux_651_nl;
  wire[0:0] or_796_nl;
  wire[0:0] or_794_nl;
  wire[0:0] mux_650_nl;
  wire[0:0] or_793_nl;
  wire[0:0] or_791_nl;
  wire[0:0] mux_649_nl;
  wire[0:0] mux_648_nl;
  wire[0:0] or_790_nl;
  wire[0:0] or_788_nl;
  wire[0:0] mux_647_nl;
  wire[0:0] or_787_nl;
  wire[0:0] or_785_nl;
  wire[0:0] mux_677_nl;
  wire[0:0] nand_495_nl;
  wire[0:0] mux_676_nl;
  wire[0:0] and_410_nl;
  wire[0:0] mux_675_nl;
  wire[0:0] mux_674_nl;
  wire[0:0] nor_821_nl;
  wire[0:0] nor_822_nl;
  wire[0:0] mux_673_nl;
  wire[0:0] nor_823_nl;
  wire[0:0] nor_824_nl;
  wire[0:0] nor_825_nl;
  wire[0:0] mux_672_nl;
  wire[0:0] mux_671_nl;
  wire[0:0] or_828_nl;
  wire[0:0] or_826_nl;
  wire[0:0] mux_670_nl;
  wire[0:0] or_825_nl;
  wire[0:0] or_823_nl;
  wire[0:0] or_2269_nl;
  wire[0:0] mux_669_nl;
  wire[0:0] nand_69_nl;
  wire[0:0] mux_668_nl;
  wire[0:0] mux_667_nl;
  wire[0:0] nor_827_nl;
  wire[0:0] nor_828_nl;
  wire[0:0] and_411_nl;
  wire[0:0] mux_666_nl;
  wire[0:0] nor_829_nl;
  wire[0:0] nor_830_nl;
  wire[0:0] or_815_nl;
  wire[0:0] mux_665_nl;
  wire[0:0] mux_664_nl;
  wire[0:0] or_814_nl;
  wire[0:0] or_812_nl;
  wire[0:0] nand_67_nl;
  wire[0:0] mux_693_nl;
  wire[0:0] mux_692_nl;
  wire[0:0] mux_691_nl;
  wire[0:0] nor_815_nl;
  wire[0:0] nor_816_nl;
  wire[0:0] mux_690_nl;
  wire[0:0] and_408_nl;
  wire[0:0] mux_686_nl;
  wire[0:0] nor_817_nl;
  wire[0:0] mux_685_nl;
  wire[0:0] nor_818_nl;
  wire[0:0] nor_819_nl;
  wire[0:0] nor_820_nl;
  wire[0:0] mux_684_nl;
  wire[0:0] mux_683_nl;
  wire[0:0] mux_682_nl;
  wire[0:0] or_847_nl;
  wire[0:0] or_845_nl;
  wire[0:0] mux_681_nl;
  wire[0:0] or_844_nl;
  wire[0:0] or_842_nl;
  wire[0:0] mux_680_nl;
  wire[0:0] mux_679_nl;
  wire[0:0] or_841_nl;
  wire[0:0] or_839_nl;
  wire[0:0] mux_678_nl;
  wire[0:0] or_838_nl;
  wire[0:0] or_836_nl;
  wire[0:0] mux_708_nl;
  wire[0:0] nand_494_nl;
  wire[0:0] mux_707_nl;
  wire[0:0] and_407_nl;
  wire[0:0] mux_706_nl;
  wire[0:0] mux_705_nl;
  wire[0:0] nor_806_nl;
  wire[0:0] nor_807_nl;
  wire[0:0] mux_704_nl;
  wire[0:0] nor_808_nl;
  wire[0:0] nor_809_nl;
  wire[0:0] nor_810_nl;
  wire[0:0] mux_703_nl;
  wire[0:0] mux_702_nl;
  wire[0:0] or_881_nl;
  wire[0:0] or_879_nl;
  wire[0:0] mux_701_nl;
  wire[0:0] or_878_nl;
  wire[0:0] or_876_nl;
  wire[0:0] or_2268_nl;
  wire[0:0] mux_700_nl;
  wire[0:0] nand_74_nl;
  wire[0:0] mux_699_nl;
  wire[0:0] mux_698_nl;
  wire[0:0] nor_812_nl;
  wire[0:0] nor_813_nl;
  wire[0:0] nor_814_nl;
  wire[0:0] mux_697_nl;
  wire[0:0] or_870_nl;
  wire[0:0] or_868_nl;
  wire[0:0] or_867_nl;
  wire[0:0] mux_696_nl;
  wire[0:0] mux_695_nl;
  wire[0:0] or_866_nl;
  wire[0:0] or_864_nl;
  wire[0:0] or_863_nl;
  wire[0:0] mux_724_nl;
  wire[0:0] mux_723_nl;
  wire[0:0] mux_722_nl;
  wire[0:0] nor_799_nl;
  wire[0:0] nor_800_nl;
  wire[0:0] mux_721_nl;
  wire[0:0] nor_801_nl;
  wire[0:0] mux_717_nl;
  wire[0:0] nor_802_nl;
  wire[0:0] mux_716_nl;
  wire[0:0] nor_803_nl;
  wire[0:0] nor_804_nl;
  wire[0:0] nor_805_nl;
  wire[0:0] mux_715_nl;
  wire[0:0] mux_714_nl;
  wire[0:0] mux_713_nl;
  wire[0:0] or_900_nl;
  wire[0:0] or_898_nl;
  wire[0:0] mux_712_nl;
  wire[0:0] or_897_nl;
  wire[0:0] or_895_nl;
  wire[0:0] mux_711_nl;
  wire[0:0] mux_710_nl;
  wire[0:0] or_894_nl;
  wire[0:0] or_892_nl;
  wire[0:0] mux_709_nl;
  wire[0:0] or_891_nl;
  wire[0:0] or_889_nl;
  wire[0:0] mux_739_nl;
  wire[0:0] nand_493_nl;
  wire[0:0] mux_738_nl;
  wire[0:0] and_404_nl;
  wire[0:0] mux_737_nl;
  wire[0:0] mux_736_nl;
  wire[0:0] nor_787_nl;
  wire[0:0] nor_788_nl;
  wire[0:0] mux_735_nl;
  wire[0:0] nor_789_nl;
  wire[0:0] nor_790_nl;
  wire[0:0] nor_791_nl;
  wire[0:0] mux_734_nl;
  wire[0:0] mux_733_nl;
  wire[0:0] or_932_nl;
  wire[0:0] or_930_nl;
  wire[0:0] mux_732_nl;
  wire[0:0] or_929_nl;
  wire[0:0] or_927_nl;
  wire[0:0] or_2267_nl;
  wire[0:0] mux_731_nl;
  wire[0:0] nand_80_nl;
  wire[0:0] mux_730_nl;
  wire[0:0] mux_729_nl;
  wire[0:0] nor_793_nl;
  wire[0:0] nor_794_nl;
  wire[0:0] and_405_nl;
  wire[0:0] mux_728_nl;
  wire[0:0] nor_795_nl;
  wire[0:0] nor_796_nl;
  wire[0:0] or_919_nl;
  wire[0:0] mux_727_nl;
  wire[0:0] mux_726_nl;
  wire[0:0] or_918_nl;
  wire[0:0] or_916_nl;
  wire[0:0] nand_78_nl;
  wire[0:0] mux_755_nl;
  wire[0:0] mux_754_nl;
  wire[0:0] mux_753_nl;
  wire[0:0] nor_781_nl;
  wire[0:0] nor_782_nl;
  wire[0:0] mux_752_nl;
  wire[0:0] and_402_nl;
  wire[0:0] mux_748_nl;
  wire[0:0] nor_783_nl;
  wire[0:0] mux_747_nl;
  wire[0:0] nor_784_nl;
  wire[0:0] nor_785_nl;
  wire[0:0] nor_786_nl;
  wire[0:0] mux_746_nl;
  wire[0:0] mux_745_nl;
  wire[0:0] mux_744_nl;
  wire[0:0] or_951_nl;
  wire[0:0] or_949_nl;
  wire[0:0] mux_743_nl;
  wire[0:0] or_948_nl;
  wire[0:0] or_946_nl;
  wire[0:0] mux_742_nl;
  wire[0:0] mux_741_nl;
  wire[0:0] or_945_nl;
  wire[0:0] or_943_nl;
  wire[0:0] mux_740_nl;
  wire[0:0] or_942_nl;
  wire[0:0] or_940_nl;
  wire[0:0] mux_770_nl;
  wire[0:0] nand_492_nl;
  wire[0:0] mux_769_nl;
  wire[0:0] and_401_nl;
  wire[0:0] mux_768_nl;
  wire[0:0] mux_767_nl;
  wire[0:0] nor_772_nl;
  wire[0:0] nor_773_nl;
  wire[0:0] mux_766_nl;
  wire[0:0] nor_774_nl;
  wire[0:0] nor_775_nl;
  wire[0:0] nor_776_nl;
  wire[0:0] mux_765_nl;
  wire[0:0] mux_764_nl;
  wire[0:0] or_984_nl;
  wire[0:0] or_982_nl;
  wire[0:0] mux_763_nl;
  wire[0:0] or_981_nl;
  wire[0:0] or_979_nl;
  wire[0:0] or_2266_nl;
  wire[0:0] mux_762_nl;
  wire[0:0] nand_85_nl;
  wire[0:0] mux_761_nl;
  wire[0:0] mux_760_nl;
  wire[0:0] nor_778_nl;
  wire[0:0] nor_779_nl;
  wire[0:0] nor_780_nl;
  wire[0:0] mux_759_nl;
  wire[0:0] or_973_nl;
  wire[0:0] or_972_nl;
  wire[0:0] or_971_nl;
  wire[0:0] mux_758_nl;
  wire[0:0] mux_757_nl;
  wire[0:0] or_970_nl;
  wire[0:0] or_968_nl;
  wire[0:0] or_967_nl;
  wire[0:0] mux_786_nl;
  wire[0:0] mux_785_nl;
  wire[0:0] mux_784_nl;
  wire[0:0] nor_765_nl;
  wire[0:0] nor_766_nl;
  wire[0:0] mux_783_nl;
  wire[0:0] nor_767_nl;
  wire[0:0] mux_779_nl;
  wire[0:0] nor_768_nl;
  wire[0:0] mux_778_nl;
  wire[0:0] nor_769_nl;
  wire[0:0] nor_770_nl;
  wire[0:0] nor_771_nl;
  wire[0:0] mux_777_nl;
  wire[0:0] mux_776_nl;
  wire[0:0] mux_775_nl;
  wire[0:0] or_1003_nl;
  wire[0:0] or_1001_nl;
  wire[0:0] mux_774_nl;
  wire[0:0] or_1000_nl;
  wire[0:0] or_998_nl;
  wire[0:0] mux_773_nl;
  wire[0:0] mux_772_nl;
  wire[0:0] or_997_nl;
  wire[0:0] or_995_nl;
  wire[0:0] mux_771_nl;
  wire[0:0] or_994_nl;
  wire[0:0] or_992_nl;
  wire[0:0] mux_801_nl;
  wire[0:0] nand_491_nl;
  wire[0:0] mux_800_nl;
  wire[0:0] and_398_nl;
  wire[0:0] mux_799_nl;
  wire[0:0] mux_798_nl;
  wire[0:0] nor_753_nl;
  wire[0:0] nor_754_nl;
  wire[0:0] mux_797_nl;
  wire[0:0] nor_755_nl;
  wire[0:0] nor_756_nl;
  wire[0:0] nor_757_nl;
  wire[0:0] mux_796_nl;
  wire[0:0] mux_795_nl;
  wire[0:0] nand_516_nl;
  wire[0:0] or_1031_nl;
  wire[0:0] mux_794_nl;
  wire[0:0] or_1030_nl;
  wire[0:0] or_1028_nl;
  wire[0:0] or_2265_nl;
  wire[0:0] mux_793_nl;
  wire[0:0] nand_91_nl;
  wire[0:0] mux_792_nl;
  wire[0:0] mux_791_nl;
  wire[0:0] nor_759_nl;
  wire[0:0] nor_760_nl;
  wire[0:0] and_399_nl;
  wire[0:0] mux_790_nl;
  wire[0:0] nor_761_nl;
  wire[0:0] nor_762_nl;
  wire[0:0] or_1022_nl;
  wire[0:0] mux_789_nl;
  wire[0:0] mux_788_nl;
  wire[0:0] or_1021_nl;
  wire[0:0] or_1019_nl;
  wire[0:0] nand_89_nl;
  wire[0:0] mux_817_nl;
  wire[0:0] mux_816_nl;
  wire[0:0] mux_815_nl;
  wire[0:0] nor_748_nl;
  wire[0:0] nor_749_nl;
  wire[0:0] mux_814_nl;
  wire[0:0] and_395_nl;
  wire[0:0] mux_810_nl;
  wire[0:0] and_396_nl;
  wire[0:0] mux_809_nl;
  wire[0:0] and_527_nl;
  wire[0:0] nor_751_nl;
  wire[0:0] nor_752_nl;
  wire[0:0] mux_808_nl;
  wire[0:0] mux_807_nl;
  wire[0:0] mux_806_nl;
  wire[0:0] or_1051_nl;
  wire[0:0] nand_369_nl;
  wire[0:0] mux_805_nl;
  wire[0:0] nand_515_nl;
  wire[0:0] or_1046_nl;
  wire[0:0] mux_804_nl;
  wire[0:0] mux_803_nl;
  wire[0:0] or_1045_nl;
  wire[0:0] nand_373_nl;
  wire[0:0] mux_802_nl;
  wire[0:0] nand_471_nl;
  wire[0:0] or_1040_nl;
  wire[0:0] mux_832_nl;
  wire[0:0] nand_490_nl;
  wire[0:0] mux_831_nl;
  wire[0:0] and_394_nl;
  wire[0:0] mux_830_nl;
  wire[0:0] mux_829_nl;
  wire[0:0] nor_739_nl;
  wire[0:0] nor_740_nl;
  wire[0:0] mux_828_nl;
  wire[0:0] nor_741_nl;
  wire[0:0] nor_742_nl;
  wire[0:0] nor_743_nl;
  wire[0:0] mux_827_nl;
  wire[0:0] mux_826_nl;
  wire[0:0] or_1085_nl;
  wire[0:0] or_1083_nl;
  wire[0:0] mux_825_nl;
  wire[0:0] or_1082_nl;
  wire[0:0] or_1080_nl;
  wire[0:0] or_2264_nl;
  wire[0:0] mux_824_nl;
  wire[0:0] nand_96_nl;
  wire[0:0] mux_823_nl;
  wire[0:0] mux_822_nl;
  wire[0:0] nor_745_nl;
  wire[0:0] nor_746_nl;
  wire[0:0] nor_747_nl;
  wire[0:0] mux_821_nl;
  wire[0:0] or_1074_nl;
  wire[0:0] or_1072_nl;
  wire[0:0] or_1071_nl;
  wire[0:0] mux_820_nl;
  wire[0:0] mux_819_nl;
  wire[0:0] or_1070_nl;
  wire[0:0] or_1068_nl;
  wire[0:0] or_1067_nl;
  wire[0:0] mux_848_nl;
  wire[0:0] mux_847_nl;
  wire[0:0] mux_846_nl;
  wire[0:0] nor_732_nl;
  wire[0:0] nor_733_nl;
  wire[0:0] mux_845_nl;
  wire[0:0] nor_734_nl;
  wire[0:0] mux_841_nl;
  wire[0:0] nor_735_nl;
  wire[0:0] mux_840_nl;
  wire[0:0] nor_736_nl;
  wire[0:0] nor_737_nl;
  wire[0:0] nor_738_nl;
  wire[0:0] mux_839_nl;
  wire[0:0] mux_838_nl;
  wire[0:0] mux_837_nl;
  wire[0:0] or_1104_nl;
  wire[0:0] or_1102_nl;
  wire[0:0] mux_836_nl;
  wire[0:0] or_1101_nl;
  wire[0:0] or_1099_nl;
  wire[0:0] mux_835_nl;
  wire[0:0] mux_834_nl;
  wire[0:0] or_1098_nl;
  wire[0:0] or_1096_nl;
  wire[0:0] mux_833_nl;
  wire[0:0] or_1095_nl;
  wire[0:0] or_1093_nl;
  wire[0:0] mux_863_nl;
  wire[0:0] nand_489_nl;
  wire[0:0] mux_862_nl;
  wire[0:0] and_391_nl;
  wire[0:0] mux_861_nl;
  wire[0:0] mux_860_nl;
  wire[0:0] nor_720_nl;
  wire[0:0] nor_721_nl;
  wire[0:0] mux_859_nl;
  wire[0:0] nor_722_nl;
  wire[0:0] nor_723_nl;
  wire[0:0] nor_724_nl;
  wire[0:0] mux_858_nl;
  wire[0:0] mux_857_nl;
  wire[0:0] or_1136_nl;
  wire[0:0] or_1134_nl;
  wire[0:0] mux_856_nl;
  wire[0:0] or_1133_nl;
  wire[0:0] or_1131_nl;
  wire[0:0] or_2263_nl;
  wire[0:0] mux_855_nl;
  wire[0:0] nand_102_nl;
  wire[0:0] mux_854_nl;
  wire[0:0] mux_853_nl;
  wire[0:0] nor_726_nl;
  wire[0:0] nor_727_nl;
  wire[0:0] and_392_nl;
  wire[0:0] mux_852_nl;
  wire[0:0] nor_728_nl;
  wire[0:0] nor_729_nl;
  wire[0:0] or_1123_nl;
  wire[0:0] mux_851_nl;
  wire[0:0] mux_850_nl;
  wire[0:0] or_1122_nl;
  wire[0:0] or_1120_nl;
  wire[0:0] nand_100_nl;
  wire[0:0] mux_879_nl;
  wire[0:0] mux_878_nl;
  wire[0:0] mux_877_nl;
  wire[0:0] nor_714_nl;
  wire[0:0] nor_715_nl;
  wire[0:0] mux_876_nl;
  wire[0:0] and_389_nl;
  wire[0:0] mux_872_nl;
  wire[0:0] nor_716_nl;
  wire[0:0] mux_871_nl;
  wire[0:0] nor_717_nl;
  wire[0:0] nor_718_nl;
  wire[0:0] nor_719_nl;
  wire[0:0] mux_870_nl;
  wire[0:0] mux_869_nl;
  wire[0:0] mux_868_nl;
  wire[0:0] or_1155_nl;
  wire[0:0] or_1153_nl;
  wire[0:0] mux_867_nl;
  wire[0:0] or_1152_nl;
  wire[0:0] or_1150_nl;
  wire[0:0] mux_866_nl;
  wire[0:0] mux_865_nl;
  wire[0:0] or_1149_nl;
  wire[0:0] or_1147_nl;
  wire[0:0] mux_864_nl;
  wire[0:0] or_1146_nl;
  wire[0:0] or_1144_nl;
  wire[0:0] mux_894_nl;
  wire[0:0] nand_488_nl;
  wire[0:0] mux_893_nl;
  wire[0:0] and_388_nl;
  wire[0:0] mux_892_nl;
  wire[0:0] mux_891_nl;
  wire[0:0] nor_705_nl;
  wire[0:0] nor_706_nl;
  wire[0:0] mux_890_nl;
  wire[0:0] nor_707_nl;
  wire[0:0] nor_708_nl;
  wire[0:0] nor_709_nl;
  wire[0:0] mux_889_nl;
  wire[0:0] mux_888_nl;
  wire[0:0] or_1189_nl;
  wire[0:0] or_1187_nl;
  wire[0:0] mux_887_nl;
  wire[0:0] or_1186_nl;
  wire[0:0] or_1184_nl;
  wire[0:0] or_2262_nl;
  wire[0:0] mux_886_nl;
  wire[0:0] nand_107_nl;
  wire[0:0] mux_885_nl;
  wire[0:0] mux_884_nl;
  wire[0:0] nor_711_nl;
  wire[0:0] nor_712_nl;
  wire[0:0] nor_713_nl;
  wire[0:0] mux_883_nl;
  wire[0:0] or_1178_nl;
  wire[0:0] or_1176_nl;
  wire[0:0] or_1175_nl;
  wire[0:0] mux_882_nl;
  wire[0:0] mux_881_nl;
  wire[0:0] or_1174_nl;
  wire[0:0] or_1172_nl;
  wire[0:0] or_1171_nl;
  wire[0:0] mux_910_nl;
  wire[0:0] mux_909_nl;
  wire[0:0] mux_908_nl;
  wire[0:0] nor_698_nl;
  wire[0:0] nor_699_nl;
  wire[0:0] mux_907_nl;
  wire[0:0] nor_700_nl;
  wire[0:0] mux_903_nl;
  wire[0:0] nor_701_nl;
  wire[0:0] mux_902_nl;
  wire[0:0] nor_702_nl;
  wire[0:0] nor_703_nl;
  wire[0:0] nor_704_nl;
  wire[0:0] mux_901_nl;
  wire[0:0] mux_900_nl;
  wire[0:0] mux_899_nl;
  wire[0:0] or_1208_nl;
  wire[0:0] or_1206_nl;
  wire[0:0] mux_898_nl;
  wire[0:0] or_1205_nl;
  wire[0:0] or_1203_nl;
  wire[0:0] mux_897_nl;
  wire[0:0] mux_896_nl;
  wire[0:0] or_1202_nl;
  wire[0:0] or_1200_nl;
  wire[0:0] mux_895_nl;
  wire[0:0] or_1199_nl;
  wire[0:0] or_1197_nl;
  wire[0:0] mux_925_nl;
  wire[0:0] nand_487_nl;
  wire[0:0] mux_924_nl;
  wire[0:0] and_385_nl;
  wire[0:0] mux_923_nl;
  wire[0:0] mux_922_nl;
  wire[0:0] nor_686_nl;
  wire[0:0] nor_687_nl;
  wire[0:0] mux_921_nl;
  wire[0:0] nor_688_nl;
  wire[0:0] nor_689_nl;
  wire[0:0] nor_690_nl;
  wire[0:0] mux_920_nl;
  wire[0:0] mux_919_nl;
  wire[0:0] or_1240_nl;
  wire[0:0] or_1238_nl;
  wire[0:0] mux_918_nl;
  wire[0:0] or_1237_nl;
  wire[0:0] or_1235_nl;
  wire[0:0] or_2261_nl;
  wire[0:0] mux_917_nl;
  wire[0:0] nand_113_nl;
  wire[0:0] mux_916_nl;
  wire[0:0] mux_915_nl;
  wire[0:0] nor_692_nl;
  wire[0:0] nor_693_nl;
  wire[0:0] and_386_nl;
  wire[0:0] mux_914_nl;
  wire[0:0] nor_694_nl;
  wire[0:0] nor_695_nl;
  wire[0:0] or_1227_nl;
  wire[0:0] mux_913_nl;
  wire[0:0] mux_912_nl;
  wire[0:0] or_1226_nl;
  wire[0:0] or_1224_nl;
  wire[0:0] nand_111_nl;
  wire[0:0] mux_941_nl;
  wire[0:0] mux_940_nl;
  wire[0:0] mux_939_nl;
  wire[0:0] nor_680_nl;
  wire[0:0] nor_681_nl;
  wire[0:0] mux_938_nl;
  wire[0:0] and_383_nl;
  wire[0:0] mux_934_nl;
  wire[0:0] nor_682_nl;
  wire[0:0] mux_933_nl;
  wire[0:0] nor_683_nl;
  wire[0:0] nor_684_nl;
  wire[0:0] nor_685_nl;
  wire[0:0] mux_932_nl;
  wire[0:0] mux_931_nl;
  wire[0:0] mux_930_nl;
  wire[0:0] or_1259_nl;
  wire[0:0] or_1257_nl;
  wire[0:0] mux_929_nl;
  wire[0:0] or_1256_nl;
  wire[0:0] or_1254_nl;
  wire[0:0] mux_928_nl;
  wire[0:0] mux_927_nl;
  wire[0:0] or_1253_nl;
  wire[0:0] or_1251_nl;
  wire[0:0] mux_926_nl;
  wire[0:0] or_1250_nl;
  wire[0:0] or_1248_nl;
  wire[0:0] mux_956_nl;
  wire[0:0] nand_486_nl;
  wire[0:0] mux_955_nl;
  wire[0:0] and_382_nl;
  wire[0:0] mux_954_nl;
  wire[0:0] mux_953_nl;
  wire[0:0] nor_671_nl;
  wire[0:0] nor_672_nl;
  wire[0:0] mux_952_nl;
  wire[0:0] nor_673_nl;
  wire[0:0] nor_674_nl;
  wire[0:0] nor_675_nl;
  wire[0:0] mux_951_nl;
  wire[0:0] mux_950_nl;
  wire[0:0] or_1293_nl;
  wire[0:0] or_1291_nl;
  wire[0:0] mux_949_nl;
  wire[0:0] or_1290_nl;
  wire[0:0] or_1288_nl;
  wire[0:0] or_2260_nl;
  wire[0:0] mux_948_nl;
  wire[0:0] nand_118_nl;
  wire[0:0] mux_947_nl;
  wire[0:0] mux_946_nl;
  wire[0:0] nor_677_nl;
  wire[0:0] nor_678_nl;
  wire[0:0] nor_679_nl;
  wire[0:0] mux_945_nl;
  wire[0:0] or_1282_nl;
  wire[0:0] or_1280_nl;
  wire[0:0] or_1279_nl;
  wire[0:0] mux_944_nl;
  wire[0:0] mux_943_nl;
  wire[0:0] or_1278_nl;
  wire[0:0] or_1276_nl;
  wire[0:0] or_1275_nl;
  wire[0:0] mux_972_nl;
  wire[0:0] mux_971_nl;
  wire[0:0] mux_970_nl;
  wire[0:0] nor_664_nl;
  wire[0:0] nor_665_nl;
  wire[0:0] mux_969_nl;
  wire[0:0] nor_666_nl;
  wire[0:0] mux_965_nl;
  wire[0:0] nor_667_nl;
  wire[0:0] mux_964_nl;
  wire[0:0] nor_668_nl;
  wire[0:0] nor_669_nl;
  wire[0:0] nor_670_nl;
  wire[0:0] mux_963_nl;
  wire[0:0] mux_962_nl;
  wire[0:0] mux_961_nl;
  wire[0:0] or_1312_nl;
  wire[0:0] or_1310_nl;
  wire[0:0] mux_960_nl;
  wire[0:0] or_1309_nl;
  wire[0:0] or_1307_nl;
  wire[0:0] mux_959_nl;
  wire[0:0] mux_958_nl;
  wire[0:0] or_1306_nl;
  wire[0:0] or_1304_nl;
  wire[0:0] mux_957_nl;
  wire[0:0] or_1303_nl;
  wire[0:0] or_1301_nl;
  wire[0:0] mux_987_nl;
  wire[0:0] nand_485_nl;
  wire[0:0] mux_986_nl;
  wire[0:0] and_379_nl;
  wire[0:0] mux_985_nl;
  wire[0:0] mux_984_nl;
  wire[0:0] nor_652_nl;
  wire[0:0] nor_653_nl;
  wire[0:0] mux_983_nl;
  wire[0:0] nor_654_nl;
  wire[0:0] nor_655_nl;
  wire[0:0] nor_656_nl;
  wire[0:0] mux_982_nl;
  wire[0:0] mux_981_nl;
  wire[0:0] or_1344_nl;
  wire[0:0] or_1342_nl;
  wire[0:0] mux_980_nl;
  wire[0:0] or_1341_nl;
  wire[0:0] or_1339_nl;
  wire[0:0] or_2259_nl;
  wire[0:0] mux_979_nl;
  wire[0:0] nand_124_nl;
  wire[0:0] mux_978_nl;
  wire[0:0] mux_977_nl;
  wire[0:0] nor_658_nl;
  wire[0:0] nor_659_nl;
  wire[0:0] and_380_nl;
  wire[0:0] mux_976_nl;
  wire[0:0] nor_660_nl;
  wire[0:0] nor_661_nl;
  wire[0:0] or_1331_nl;
  wire[0:0] mux_975_nl;
  wire[0:0] mux_974_nl;
  wire[0:0] or_1330_nl;
  wire[0:0] or_1328_nl;
  wire[0:0] nand_122_nl;
  wire[0:0] mux_1003_nl;
  wire[0:0] mux_1002_nl;
  wire[0:0] mux_1001_nl;
  wire[0:0] nor_646_nl;
  wire[0:0] nor_647_nl;
  wire[0:0] mux_1000_nl;
  wire[0:0] and_377_nl;
  wire[0:0] mux_996_nl;
  wire[0:0] nor_648_nl;
  wire[0:0] mux_995_nl;
  wire[0:0] nor_649_nl;
  wire[0:0] nor_650_nl;
  wire[0:0] nor_651_nl;
  wire[0:0] mux_994_nl;
  wire[0:0] mux_993_nl;
  wire[0:0] mux_992_nl;
  wire[0:0] or_1363_nl;
  wire[0:0] or_1361_nl;
  wire[0:0] mux_991_nl;
  wire[0:0] or_1360_nl;
  wire[0:0] or_1358_nl;
  wire[0:0] mux_990_nl;
  wire[0:0] mux_989_nl;
  wire[0:0] or_1357_nl;
  wire[0:0] or_1355_nl;
  wire[0:0] mux_988_nl;
  wire[0:0] or_1354_nl;
  wire[0:0] or_1352_nl;
  wire[0:0] mux_1018_nl;
  wire[0:0] nand_484_nl;
  wire[0:0] mux_1017_nl;
  wire[0:0] and_376_nl;
  wire[0:0] mux_1016_nl;
  wire[0:0] mux_1015_nl;
  wire[0:0] nor_637_nl;
  wire[0:0] nor_638_nl;
  wire[0:0] mux_1014_nl;
  wire[0:0] nor_639_nl;
  wire[0:0] nor_640_nl;
  wire[0:0] nor_641_nl;
  wire[0:0] mux_1013_nl;
  wire[0:0] mux_1012_nl;
  wire[0:0] or_1397_nl;
  wire[0:0] or_1395_nl;
  wire[0:0] mux_1011_nl;
  wire[0:0] or_1394_nl;
  wire[0:0] or_1392_nl;
  wire[0:0] or_2258_nl;
  wire[0:0] mux_1010_nl;
  wire[0:0] nand_129_nl;
  wire[0:0] mux_1009_nl;
  wire[0:0] mux_1008_nl;
  wire[0:0] nor_643_nl;
  wire[0:0] nor_644_nl;
  wire[0:0] nor_645_nl;
  wire[0:0] mux_1007_nl;
  wire[0:0] or_1386_nl;
  wire[0:0] or_1384_nl;
  wire[0:0] or_1383_nl;
  wire[0:0] mux_1006_nl;
  wire[0:0] mux_1005_nl;
  wire[0:0] or_1382_nl;
  wire[0:0] or_1380_nl;
  wire[0:0] or_1379_nl;
  wire[0:0] mux_1034_nl;
  wire[0:0] mux_1033_nl;
  wire[0:0] mux_1032_nl;
  wire[0:0] nor_630_nl;
  wire[0:0] nor_631_nl;
  wire[0:0] mux_1031_nl;
  wire[0:0] nor_632_nl;
  wire[0:0] mux_1027_nl;
  wire[0:0] nor_633_nl;
  wire[0:0] mux_1026_nl;
  wire[0:0] nor_634_nl;
  wire[0:0] nor_635_nl;
  wire[0:0] nor_636_nl;
  wire[0:0] mux_1025_nl;
  wire[0:0] mux_1024_nl;
  wire[0:0] mux_1023_nl;
  wire[0:0] or_1416_nl;
  wire[0:0] or_1414_nl;
  wire[0:0] mux_1022_nl;
  wire[0:0] or_1413_nl;
  wire[0:0] or_1411_nl;
  wire[0:0] mux_1021_nl;
  wire[0:0] mux_1020_nl;
  wire[0:0] or_1410_nl;
  wire[0:0] or_1408_nl;
  wire[0:0] mux_1019_nl;
  wire[0:0] or_1407_nl;
  wire[0:0] or_1405_nl;
  wire[0:0] mux_1049_nl;
  wire[0:0] nand_483_nl;
  wire[0:0] mux_1048_nl;
  wire[0:0] and_373_nl;
  wire[0:0] mux_1047_nl;
  wire[0:0] mux_1046_nl;
  wire[0:0] nor_618_nl;
  wire[0:0] nor_619_nl;
  wire[0:0] mux_1045_nl;
  wire[0:0] nor_620_nl;
  wire[0:0] nor_621_nl;
  wire[0:0] nor_622_nl;
  wire[0:0] mux_1044_nl;
  wire[0:0] mux_1043_nl;
  wire[0:0] or_1448_nl;
  wire[0:0] or_1446_nl;
  wire[0:0] mux_1042_nl;
  wire[0:0] or_1445_nl;
  wire[0:0] or_1443_nl;
  wire[0:0] or_2257_nl;
  wire[0:0] mux_1041_nl;
  wire[0:0] nand_135_nl;
  wire[0:0] mux_1040_nl;
  wire[0:0] mux_1039_nl;
  wire[0:0] nor_624_nl;
  wire[0:0] nor_625_nl;
  wire[0:0] and_374_nl;
  wire[0:0] mux_1038_nl;
  wire[0:0] nor_626_nl;
  wire[0:0] nor_627_nl;
  wire[0:0] or_1435_nl;
  wire[0:0] mux_1037_nl;
  wire[0:0] mux_1036_nl;
  wire[0:0] or_1434_nl;
  wire[0:0] or_1432_nl;
  wire[0:0] nand_133_nl;
  wire[0:0] mux_1065_nl;
  wire[0:0] mux_1064_nl;
  wire[0:0] mux_1063_nl;
  wire[0:0] nor_613_nl;
  wire[0:0] nor_614_nl;
  wire[0:0] mux_1062_nl;
  wire[0:0] and_370_nl;
  wire[0:0] mux_1058_nl;
  wire[0:0] and_371_nl;
  wire[0:0] mux_1057_nl;
  wire[0:0] and_526_nl;
  wire[0:0] nor_616_nl;
  wire[0:0] nor_617_nl;
  wire[0:0] mux_1056_nl;
  wire[0:0] mux_1055_nl;
  wire[0:0] mux_1054_nl;
  wire[0:0] or_1467_nl;
  wire[0:0] nand_307_nl;
  wire[0:0] mux_1053_nl;
  wire[0:0] nand_514_nl;
  wire[0:0] or_1462_nl;
  wire[0:0] mux_1052_nl;
  wire[0:0] mux_1051_nl;
  wire[0:0] or_1461_nl;
  wire[0:0] nand_310_nl;
  wire[0:0] mux_1050_nl;
  wire[0:0] nand_468_nl;
  wire[0:0] or_1456_nl;
  wire[0:0] mux_1080_nl;
  wire[0:0] nand_482_nl;
  wire[0:0] mux_1079_nl;
  wire[0:0] and_369_nl;
  wire[0:0] mux_1078_nl;
  wire[0:0] mux_1077_nl;
  wire[0:0] nor_604_nl;
  wire[0:0] nor_605_nl;
  wire[0:0] mux_1076_nl;
  wire[0:0] nor_606_nl;
  wire[0:0] nor_607_nl;
  wire[0:0] nor_608_nl;
  wire[0:0] mux_1075_nl;
  wire[0:0] mux_1074_nl;
  wire[0:0] or_1500_nl;
  wire[0:0] or_1498_nl;
  wire[0:0] mux_1073_nl;
  wire[0:0] or_1497_nl;
  wire[0:0] or_1495_nl;
  wire[0:0] or_2256_nl;
  wire[0:0] mux_1072_nl;
  wire[0:0] nand_140_nl;
  wire[0:0] mux_1071_nl;
  wire[0:0] mux_1070_nl;
  wire[0:0] nor_610_nl;
  wire[0:0] nor_611_nl;
  wire[0:0] nor_612_nl;
  wire[0:0] mux_1069_nl;
  wire[0:0] or_1489_nl;
  wire[0:0] or_1487_nl;
  wire[0:0] or_1486_nl;
  wire[0:0] mux_1068_nl;
  wire[0:0] mux_1067_nl;
  wire[0:0] or_1485_nl;
  wire[0:0] or_1483_nl;
  wire[0:0] or_1482_nl;
  wire[0:0] mux_1096_nl;
  wire[0:0] mux_1095_nl;
  wire[0:0] mux_1094_nl;
  wire[0:0] nor_597_nl;
  wire[0:0] nor_598_nl;
  wire[0:0] mux_1093_nl;
  wire[0:0] nor_599_nl;
  wire[0:0] mux_1089_nl;
  wire[0:0] nor_600_nl;
  wire[0:0] mux_1088_nl;
  wire[0:0] nor_601_nl;
  wire[0:0] nor_602_nl;
  wire[0:0] nor_603_nl;
  wire[0:0] mux_1087_nl;
  wire[0:0] mux_1086_nl;
  wire[0:0] mux_1085_nl;
  wire[0:0] or_1519_nl;
  wire[0:0] or_1517_nl;
  wire[0:0] mux_1084_nl;
  wire[0:0] or_1516_nl;
  wire[0:0] or_1514_nl;
  wire[0:0] mux_1083_nl;
  wire[0:0] mux_1082_nl;
  wire[0:0] or_1513_nl;
  wire[0:0] or_1511_nl;
  wire[0:0] mux_1081_nl;
  wire[0:0] or_1510_nl;
  wire[0:0] or_1508_nl;
  wire[0:0] mux_1111_nl;
  wire[0:0] nand_481_nl;
  wire[0:0] mux_1110_nl;
  wire[0:0] and_366_nl;
  wire[0:0] mux_1109_nl;
  wire[0:0] mux_1108_nl;
  wire[0:0] nor_585_nl;
  wire[0:0] nor_586_nl;
  wire[0:0] mux_1107_nl;
  wire[0:0] nor_587_nl;
  wire[0:0] nor_588_nl;
  wire[0:0] nor_589_nl;
  wire[0:0] mux_1106_nl;
  wire[0:0] mux_1105_nl;
  wire[0:0] or_1550_nl;
  wire[0:0] or_1548_nl;
  wire[0:0] mux_1104_nl;
  wire[0:0] or_1547_nl;
  wire[0:0] or_1545_nl;
  wire[0:0] or_2255_nl;
  wire[0:0] mux_1103_nl;
  wire[0:0] nand_146_nl;
  wire[0:0] mux_1102_nl;
  wire[0:0] mux_1101_nl;
  wire[0:0] nor_591_nl;
  wire[0:0] nor_592_nl;
  wire[0:0] and_367_nl;
  wire[0:0] mux_1100_nl;
  wire[0:0] nor_593_nl;
  wire[0:0] nor_594_nl;
  wire[0:0] or_1537_nl;
  wire[0:0] mux_1099_nl;
  wire[0:0] mux_1098_nl;
  wire[0:0] or_1536_nl;
  wire[0:0] or_1534_nl;
  wire[0:0] nand_144_nl;
  wire[0:0] mux_1127_nl;
  wire[0:0] mux_1126_nl;
  wire[0:0] mux_1125_nl;
  wire[0:0] nor_579_nl;
  wire[0:0] nor_580_nl;
  wire[0:0] mux_1124_nl;
  wire[0:0] and_364_nl;
  wire[0:0] mux_1120_nl;
  wire[0:0] nor_581_nl;
  wire[0:0] mux_1119_nl;
  wire[0:0] nor_582_nl;
  wire[0:0] nor_583_nl;
  wire[0:0] nor_584_nl;
  wire[0:0] mux_1118_nl;
  wire[0:0] mux_1117_nl;
  wire[0:0] mux_1116_nl;
  wire[0:0] or_1569_nl;
  wire[0:0] or_1567_nl;
  wire[0:0] mux_1115_nl;
  wire[0:0] or_1566_nl;
  wire[0:0] or_1564_nl;
  wire[0:0] mux_1114_nl;
  wire[0:0] mux_1113_nl;
  wire[0:0] or_1563_nl;
  wire[0:0] or_1561_nl;
  wire[0:0] mux_1112_nl;
  wire[0:0] or_1560_nl;
  wire[0:0] or_1558_nl;
  wire[0:0] mux_1142_nl;
  wire[0:0] nand_480_nl;
  wire[0:0] mux_1141_nl;
  wire[0:0] and_363_nl;
  wire[0:0] mux_1140_nl;
  wire[0:0] mux_1139_nl;
  wire[0:0] nor_570_nl;
  wire[0:0] nor_571_nl;
  wire[0:0] mux_1138_nl;
  wire[0:0] nor_572_nl;
  wire[0:0] nor_573_nl;
  wire[0:0] nor_574_nl;
  wire[0:0] mux_1137_nl;
  wire[0:0] mux_1136_nl;
  wire[0:0] or_1602_nl;
  wire[0:0] or_1600_nl;
  wire[0:0] mux_1135_nl;
  wire[0:0] or_1599_nl;
  wire[0:0] or_1597_nl;
  wire[0:0] or_2254_nl;
  wire[0:0] mux_1134_nl;
  wire[0:0] nand_151_nl;
  wire[0:0] mux_1133_nl;
  wire[0:0] mux_1132_nl;
  wire[0:0] nor_576_nl;
  wire[0:0] nor_577_nl;
  wire[0:0] nor_578_nl;
  wire[0:0] mux_1131_nl;
  wire[0:0] or_1591_nl;
  wire[0:0] or_1589_nl;
  wire[0:0] or_1588_nl;
  wire[0:0] mux_1130_nl;
  wire[0:0] mux_1129_nl;
  wire[0:0] or_1587_nl;
  wire[0:0] or_1585_nl;
  wire[0:0] or_1584_nl;
  wire[0:0] mux_1158_nl;
  wire[0:0] mux_1157_nl;
  wire[0:0] mux_1156_nl;
  wire[0:0] nor_563_nl;
  wire[0:0] nor_564_nl;
  wire[0:0] mux_1155_nl;
  wire[0:0] nor_565_nl;
  wire[0:0] mux_1151_nl;
  wire[0:0] nor_566_nl;
  wire[0:0] mux_1150_nl;
  wire[0:0] nor_567_nl;
  wire[0:0] nor_568_nl;
  wire[0:0] nor_569_nl;
  wire[0:0] mux_1149_nl;
  wire[0:0] mux_1148_nl;
  wire[0:0] mux_1147_nl;
  wire[0:0] or_1621_nl;
  wire[0:0] or_1619_nl;
  wire[0:0] mux_1146_nl;
  wire[0:0] or_1618_nl;
  wire[0:0] or_1616_nl;
  wire[0:0] mux_1145_nl;
  wire[0:0] mux_1144_nl;
  wire[0:0] or_1615_nl;
  wire[0:0] or_1613_nl;
  wire[0:0] mux_1143_nl;
  wire[0:0] or_1612_nl;
  wire[0:0] or_1610_nl;
  wire[0:0] mux_1173_nl;
  wire[0:0] nand_479_nl;
  wire[0:0] mux_1172_nl;
  wire[0:0] and_360_nl;
  wire[0:0] mux_1171_nl;
  wire[0:0] mux_1170_nl;
  wire[0:0] nor_551_nl;
  wire[0:0] nor_552_nl;
  wire[0:0] mux_1169_nl;
  wire[0:0] nor_553_nl;
  wire[0:0] nor_554_nl;
  wire[0:0] nor_555_nl;
  wire[0:0] mux_1168_nl;
  wire[0:0] mux_1167_nl;
  wire[0:0] or_1651_nl;
  wire[0:0] or_1649_nl;
  wire[0:0] mux_1166_nl;
  wire[0:0] or_1648_nl;
  wire[0:0] or_1647_nl;
  wire[0:0] or_2253_nl;
  wire[0:0] mux_1165_nl;
  wire[0:0] nand_157_nl;
  wire[0:0] mux_1164_nl;
  wire[0:0] mux_1163_nl;
  wire[0:0] nor_557_nl;
  wire[0:0] nor_558_nl;
  wire[0:0] and_361_nl;
  wire[0:0] mux_1162_nl;
  wire[0:0] nor_559_nl;
  wire[0:0] nor_560_nl;
  wire[0:0] or_1639_nl;
  wire[0:0] mux_1161_nl;
  wire[0:0] mux_1160_nl;
  wire[0:0] or_1638_nl;
  wire[0:0] or_1636_nl;
  wire[0:0] nand_155_nl;
  wire[0:0] mux_1189_nl;
  wire[0:0] mux_1188_nl;
  wire[0:0] mux_1187_nl;
  wire[0:0] nor_546_nl;
  wire[0:0] nor_547_nl;
  wire[0:0] mux_1186_nl;
  wire[0:0] and_357_nl;
  wire[0:0] mux_1182_nl;
  wire[0:0] and_358_nl;
  wire[0:0] mux_1181_nl;
  wire[0:0] and_525_nl;
  wire[0:0] nor_549_nl;
  wire[0:0] nor_550_nl;
  wire[0:0] mux_1180_nl;
  wire[0:0] mux_1179_nl;
  wire[0:0] mux_1178_nl;
  wire[0:0] or_1670_nl;
  wire[0:0] nand_273_nl;
  wire[0:0] mux_1177_nl;
  wire[0:0] nand_513_nl;
  wire[0:0] or_1665_nl;
  wire[0:0] mux_1176_nl;
  wire[0:0] mux_1175_nl;
  wire[0:0] or_1664_nl;
  wire[0:0] nand_276_nl;
  wire[0:0] mux_1174_nl;
  wire[0:0] nand_465_nl;
  wire[0:0] or_1659_nl;
  wire[0:0] mux_1204_nl;
  wire[0:0] nand_478_nl;
  wire[0:0] mux_1203_nl;
  wire[0:0] and_356_nl;
  wire[0:0] mux_1202_nl;
  wire[0:0] mux_1201_nl;
  wire[0:0] nor_537_nl;
  wire[0:0] nor_538_nl;
  wire[0:0] mux_1200_nl;
  wire[0:0] nor_539_nl;
  wire[0:0] nor_540_nl;
  wire[0:0] nor_541_nl;
  wire[0:0] mux_1199_nl;
  wire[0:0] mux_1198_nl;
  wire[0:0] or_1702_nl;
  wire[0:0] or_1700_nl;
  wire[0:0] mux_1197_nl;
  wire[0:0] or_1699_nl;
  wire[0:0] or_1697_nl;
  wire[0:0] or_2252_nl;
  wire[0:0] mux_1196_nl;
  wire[0:0] nand_162_nl;
  wire[0:0] mux_1195_nl;
  wire[0:0] mux_1194_nl;
  wire[0:0] nor_543_nl;
  wire[0:0] nor_544_nl;
  wire[0:0] nor_545_nl;
  wire[0:0] mux_1193_nl;
  wire[0:0] nand_519_nl;
  wire[0:0] or_1689_nl;
  wire[0:0] or_1688_nl;
  wire[0:0] mux_1192_nl;
  wire[0:0] mux_1191_nl;
  wire[0:0] or_1687_nl;
  wire[0:0] or_1685_nl;
  wire[0:0] or_1684_nl;
  wire[0:0] mux_1220_nl;
  wire[0:0] mux_1219_nl;
  wire[0:0] mux_1218_nl;
  wire[0:0] nor_530_nl;
  wire[0:0] nor_531_nl;
  wire[0:0] mux_1217_nl;
  wire[0:0] nor_532_nl;
  wire[0:0] mux_1213_nl;
  wire[0:0] nor_533_nl;
  wire[0:0] mux_1212_nl;
  wire[0:0] nor_534_nl;
  wire[0:0] nor_535_nl;
  wire[0:0] nor_536_nl;
  wire[0:0] mux_1211_nl;
  wire[0:0] mux_1210_nl;
  wire[0:0] mux_1209_nl;
  wire[0:0] or_1721_nl;
  wire[0:0] or_1719_nl;
  wire[0:0] mux_1208_nl;
  wire[0:0] or_1718_nl;
  wire[0:0] or_1716_nl;
  wire[0:0] mux_1207_nl;
  wire[0:0] mux_1206_nl;
  wire[0:0] or_1715_nl;
  wire[0:0] or_1713_nl;
  wire[0:0] mux_1205_nl;
  wire[0:0] or_1712_nl;
  wire[0:0] or_1710_nl;
  wire[0:0] mux_1235_nl;
  wire[0:0] nand_477_nl;
  wire[0:0] mux_1234_nl;
  wire[0:0] and_351_nl;
  wire[0:0] mux_1233_nl;
  wire[0:0] mux_1232_nl;
  wire[0:0] nor_520_nl;
  wire[0:0] nor_521_nl;
  wire[0:0] mux_1231_nl;
  wire[0:0] nor_522_nl;
  wire[0:0] nor_523_nl;
  wire[0:0] nor_524_nl;
  wire[0:0] mux_1230_nl;
  wire[0:0] mux_1229_nl;
  wire[0:0] or_1751_nl;
  wire[0:0] or_1749_nl;
  wire[0:0] mux_1228_nl;
  wire[0:0] or_1748_nl;
  wire[0:0] or_1746_nl;
  wire[0:0] or_2251_nl;
  wire[0:0] mux_1227_nl;
  wire[0:0] nand_168_nl;
  wire[0:0] mux_1226_nl;
  wire[0:0] mux_1225_nl;
  wire[0:0] nor_526_nl;
  wire[0:0] nor_527_nl;
  wire[0:0] and_352_nl;
  wire[0:0] mux_1224_nl;
  wire[0:0] and_524_nl;
  wire[0:0] nor_529_nl;
  wire[0:0] or_1738_nl;
  wire[0:0] mux_1223_nl;
  wire[0:0] mux_1222_nl;
  wire[0:0] nand_512_nl;
  wire[0:0] or_1735_nl;
  wire[0:0] nand_166_nl;
  wire[0:0] mux_1251_nl;
  wire[0:0] mux_1250_nl;
  wire[0:0] mux_1249_nl;
  wire[0:0] nor_515_nl;
  wire[0:0] nor_516_nl;
  wire[0:0] mux_1248_nl;
  wire[0:0] and_348_nl;
  wire[0:0] mux_1244_nl;
  wire[0:0] and_349_nl;
  wire[0:0] mux_1243_nl;
  wire[0:0] and_523_nl;
  wire[0:0] nor_518_nl;
  wire[0:0] nor_519_nl;
  wire[0:0] mux_1242_nl;
  wire[0:0] mux_1241_nl;
  wire[0:0] mux_1240_nl;
  wire[0:0] or_1768_nl;
  wire[0:0] nand_251_nl;
  wire[0:0] mux_1239_nl;
  wire[0:0] nand_511_nl;
  wire[0:0] or_1763_nl;
  wire[0:0] mux_1238_nl;
  wire[0:0] mux_1237_nl;
  wire[0:0] or_1762_nl;
  wire[0:0] nand_254_nl;
  wire[0:0] mux_1236_nl;
  wire[0:0] nand_462_nl;
  wire[0:0] or_1758_nl;
  wire[0:0] mux_1266_nl;
  wire[0:0] nand_476_nl;
  wire[0:0] mux_1265_nl;
  wire[0:0] and_347_nl;
  wire[0:0] mux_1264_nl;
  wire[0:0] mux_1263_nl;
  wire[0:0] and_529_nl;
  wire[0:0] nor_507_nl;
  wire[0:0] mux_1262_nl;
  wire[0:0] and_530_nl;
  wire[0:0] nor_509_nl;
  wire[0:0] nor_510_nl;
  wire[0:0] mux_1261_nl;
  wire[0:0] mux_1260_nl;
  wire[0:0] or_1796_nl;
  wire[0:0] or_1795_nl;
  wire[0:0] mux_1259_nl;
  wire[0:0] nand_510_nl;
  wire[0:0] or_1792_nl;
  wire[0:0] or_2250_nl;
  wire[0:0] mux_1258_nl;
  wire[0:0] nand_173_nl;
  wire[0:0] mux_1257_nl;
  wire[0:0] mux_1256_nl;
  wire[0:0] and_531_nl;
  wire[0:0] nor_513_nl;
  wire[0:0] nor_514_nl;
  wire[0:0] mux_1255_nl;
  wire[0:0] nand_243_nl;
  wire[0:0] nand_244_nl;
  wire[0:0] or_1785_nl;
  wire[0:0] mux_1254_nl;
  wire[0:0] mux_1253_nl;
  wire[0:0] or_1784_nl;
  wire[0:0] or_1783_nl;
  wire[0:0] or_1782_nl;
  wire[0:0] mux_1282_nl;
  wire[0:0] mux_1281_nl;
  wire[0:0] mux_1280_nl;
  wire[0:0] nor_500_nl;
  wire[0:0] nor_501_nl;
  wire[0:0] mux_1279_nl;
  wire[0:0] nor_502_nl;
  wire[0:0] mux_1275_nl;
  wire[0:0] and_345_nl;
  wire[0:0] mux_1274_nl;
  wire[0:0] and_522_nl;
  wire[0:0] nor_504_nl;
  wire[0:0] nor_505_nl;
  wire[0:0] mux_1273_nl;
  wire[0:0] mux_1272_nl;
  wire[0:0] mux_1271_nl;
  wire[0:0] or_1815_nl;
  wire[0:0] nand_231_nl;
  wire[0:0] mux_1270_nl;
  wire[0:0] nand_509_nl;
  wire[0:0] or_1810_nl;
  wire[0:0] mux_1269_nl;
  wire[0:0] mux_1268_nl;
  wire[0:0] or_1809_nl;
  wire[0:0] nand_234_nl;
  wire[0:0] mux_1267_nl;
  wire[0:0] nand_460_nl;
  wire[0:0] or_1804_nl;
  wire[0:0] mux_1297_nl;
  wire[0:0] nand_475_nl;
  wire[0:0] mux_1296_nl;
  wire[0:0] and_333_nl;
  wire[0:0] mux_1295_nl;
  wire[0:0] mux_1294_nl;
  wire[0:0] and_334_nl;
  wire[0:0] and_335_nl;
  wire[0:0] mux_1293_nl;
  wire[0:0] and_336_nl;
  wire[0:0] and_337_nl;
  wire[0:0] nor_498_nl;
  wire[0:0] mux_1292_nl;
  wire[0:0] mux_1291_nl;
  wire[0:0] nand_223_nl;
  wire[0:0] nand_224_nl;
  wire[0:0] mux_1290_nl;
  wire[0:0] nand_225_nl;
  wire[0:0] nand_226_nl;
  wire[0:0] or_2249_nl;
  wire[0:0] mux_1289_nl;
  wire[0:0] nand_179_nl;
  wire[0:0] mux_1288_nl;
  wire[0:0] mux_1287_nl;
  wire[0:0] and_338_nl;
  wire[0:0] and_339_nl;
  wire[0:0] and_340_nl;
  wire[0:0] mux_1286_nl;
  wire[0:0] and_341_nl;
  wire[0:0] and_342_nl;
  wire[0:0] or_1830_nl;
  wire[0:0] mux_1285_nl;
  wire[0:0] mux_1284_nl;
  wire[0:0] nand_227_nl;
  wire[0:0] nand_228_nl;
  wire[0:0] nand_177_nl;
  wire[0:0] mux_1313_nl;
  wire[0:0] mux_1312_nl;
  wire[0:0] mux_1311_nl;
  wire[0:0] nor_494_nl;
  wire[0:0] nor_495_nl;
  wire[0:0] mux_1310_nl;
  wire[0:0] and_329_nl;
  wire[0:0] mux_1306_nl;
  wire[0:0] and_330_nl;
  wire[0:0] mux_1305_nl;
  wire[0:0] and_521_nl;
  wire[0:0] and_331_nl;
  wire[0:0] nor_497_nl;
  wire[0:0] mux_1304_nl;
  wire[0:0] mux_1303_nl;
  wire[0:0] mux_1302_nl;
  wire[0:0] or_1848_nl;
  wire[0:0] nand_214_nl;
  wire[0:0] mux_1301_nl;
  wire[0:0] nand_508_nl;
  wire[0:0] nand_216_nl;
  wire[0:0] mux_1300_nl;
  wire[0:0] mux_1299_nl;
  wire[0:0] nand_217_nl;
  wire[0:0] nand_218_nl;
  wire[0:0] mux_1298_nl;
  wire[0:0] nand_458_nl;
  wire[0:0] nand_220_nl;
  wire[0:0] mux_1320_nl;
  wire[0:0] mux_1319_nl;
  wire[0:0] mux_1318_nl;
  wire[0:0] nor_486_nl;
  wire[0:0] nor_487_nl;
  wire[0:0] mux_1317_nl;
  wire[0:0] nor_488_nl;
  wire[0:0] mux_1316_nl;
  wire[0:0] mux_1315_nl;
  wire[0:0] nor_490_nl;
  wire[0:0] mux_1314_nl;
  wire[0:0] nor_492_nl;
  wire[0:0] nor_493_nl;
  wire[0:0] mux_1323_nl;
  wire[0:0] mux_1322_nl;
  wire[0:0] nor_483_nl;
  wire[0:0] nor_484_nl;
  wire[0:0] nor_485_nl;
  wire[0:0] mux_1321_nl;
  wire[0:0] or_1872_nl;
  wire[0:0] or_1870_nl;
  wire[0:0] mux_1328_nl;
  wire[0:0] mux_1327_nl;
  wire[0:0] nor_477_nl;
  wire[0:0] nor_478_nl;
  wire[0:0] mux_1326_nl;
  wire[0:0] mux_1325_nl;
  wire[0:0] mux_1324_nl;
  wire[0:0] mux_1331_nl;
  wire[0:0] mux_1330_nl;
  wire[0:0] nor_474_nl;
  wire[0:0] nor_475_nl;
  wire[0:0] nor_476_nl;
  wire[0:0] mux_1329_nl;
  wire[0:0] or_1886_nl;
  wire[0:0] or_1884_nl;
  wire[0:0] mux_1337_nl;
  wire[0:0] mux_1336_nl;
  wire[0:0] mux_1335_nl;
  wire[0:0] nor_467_nl;
  wire[0:0] nor_468_nl;
  wire[0:0] nor_469_nl;
  wire[0:0] mux_1334_nl;
  wire[0:0] mux_1333_nl;
  wire[0:0] nor_470_nl;
  wire[0:0] nor_471_nl;
  wire[0:0] mux_1332_nl;
  wire[0:0] nor_472_nl;
  wire[0:0] nor_473_nl;
  wire[0:0] mux_1340_nl;
  wire[0:0] mux_1339_nl;
  wire[0:0] nor_464_nl;
  wire[0:0] nor_465_nl;
  wire[0:0] nor_466_nl;
  wire[0:0] mux_1338_nl;
  wire[0:0] or_1902_nl;
  wire[0:0] or_1900_nl;
  wire[0:0] mux_1345_nl;
  wire[0:0] mux_1344_nl;
  wire[0:0] nor_458_nl;
  wire[0:0] nor_459_nl;
  wire[0:0] mux_1343_nl;
  wire[0:0] mux_1342_nl;
  wire[0:0] mux_1341_nl;
  wire[0:0] mux_1348_nl;
  wire[0:0] mux_1347_nl;
  wire[0:0] nor_455_nl;
  wire[0:0] nor_456_nl;
  wire[0:0] nor_457_nl;
  wire[0:0] mux_1346_nl;
  wire[0:0] or_1916_nl;
  wire[0:0] or_1914_nl;
  wire[0:0] mux_1355_nl;
  wire[0:0] mux_1354_nl;
  wire[0:0] mux_1353_nl;
  wire[0:0] nor_447_nl;
  wire[0:0] nor_448_nl;
  wire[0:0] mux_1352_nl;
  wire[0:0] nor_449_nl;
  wire[0:0] mux_1351_nl;
  wire[0:0] mux_1350_nl;
  wire[0:0] nor_451_nl;
  wire[0:0] mux_1349_nl;
  wire[0:0] nor_453_nl;
  wire[0:0] nor_454_nl;
  wire[0:0] mux_1358_nl;
  wire[0:0] mux_1357_nl;
  wire[0:0] nor_444_nl;
  wire[0:0] nor_445_nl;
  wire[0:0] nor_446_nl;
  wire[0:0] mux_1356_nl;
  wire[0:0] or_1933_nl;
  wire[0:0] or_1931_nl;
  wire[0:0] mux_1363_nl;
  wire[0:0] mux_1362_nl;
  wire[0:0] nor_438_nl;
  wire[0:0] nor_439_nl;
  wire[0:0] mux_1361_nl;
  wire[0:0] mux_1360_nl;
  wire[0:0] mux_1359_nl;
  wire[0:0] mux_1366_nl;
  wire[0:0] mux_1365_nl;
  wire[0:0] nor_435_nl;
  wire[0:0] nor_436_nl;
  wire[0:0] nor_437_nl;
  wire[0:0] mux_1364_nl;
  wire[0:0] or_1947_nl;
  wire[0:0] or_1945_nl;
  wire[0:0] mux_1372_nl;
  wire[0:0] mux_1371_nl;
  wire[0:0] mux_1370_nl;
  wire[0:0] nor_428_nl;
  wire[0:0] nor_429_nl;
  wire[0:0] nor_430_nl;
  wire[0:0] mux_1369_nl;
  wire[0:0] mux_1368_nl;
  wire[0:0] nor_431_nl;
  wire[0:0] nor_432_nl;
  wire[0:0] mux_1367_nl;
  wire[0:0] nor_433_nl;
  wire[0:0] nor_434_nl;
  wire[0:0] mux_1375_nl;
  wire[0:0] mux_1374_nl;
  wire[0:0] nor_425_nl;
  wire[0:0] nor_426_nl;
  wire[0:0] nor_427_nl;
  wire[0:0] mux_1373_nl;
  wire[0:0] or_1963_nl;
  wire[0:0] or_1961_nl;
  wire[0:0] mux_1380_nl;
  wire[0:0] mux_1379_nl;
  wire[0:0] nor_419_nl;
  wire[0:0] nor_420_nl;
  wire[0:0] mux_1378_nl;
  wire[0:0] mux_1377_nl;
  wire[0:0] mux_1376_nl;
  wire[0:0] mux_1383_nl;
  wire[0:0] mux_1382_nl;
  wire[0:0] nor_416_nl;
  wire[0:0] nor_417_nl;
  wire[0:0] nor_418_nl;
  wire[0:0] mux_1381_nl;
  wire[0:0] or_1977_nl;
  wire[0:0] or_1975_nl;
  wire[0:0] mux_1390_nl;
  wire[0:0] mux_1389_nl;
  wire[0:0] mux_1388_nl;
  wire[0:0] nor_408_nl;
  wire[0:0] nor_409_nl;
  wire[0:0] mux_1387_nl;
  wire[0:0] nor_410_nl;
  wire[0:0] mux_1386_nl;
  wire[0:0] mux_1385_nl;
  wire[0:0] nor_412_nl;
  wire[0:0] mux_1384_nl;
  wire[0:0] nor_414_nl;
  wire[0:0] nor_415_nl;
  wire[0:0] mux_1393_nl;
  wire[0:0] mux_1392_nl;
  wire[0:0] nor_405_nl;
  wire[0:0] nor_406_nl;
  wire[0:0] nor_407_nl;
  wire[0:0] mux_1391_nl;
  wire[0:0] or_1994_nl;
  wire[0:0] or_1992_nl;
  wire[0:0] mux_1398_nl;
  wire[0:0] mux_1397_nl;
  wire[0:0] nor_399_nl;
  wire[0:0] nor_400_nl;
  wire[0:0] mux_1396_nl;
  wire[0:0] mux_1395_nl;
  wire[0:0] mux_1394_nl;
  wire[0:0] mux_1401_nl;
  wire[0:0] mux_1400_nl;
  wire[0:0] nor_396_nl;
  wire[0:0] nor_397_nl;
  wire[0:0] nor_398_nl;
  wire[0:0] mux_1399_nl;
  wire[0:0] or_2008_nl;
  wire[0:0] or_2006_nl;
  wire[0:0] mux_1407_nl;
  wire[0:0] mux_1406_nl;
  wire[0:0] mux_1405_nl;
  wire[0:0] nor_389_nl;
  wire[0:0] nor_390_nl;
  wire[0:0] nor_391_nl;
  wire[0:0] mux_1404_nl;
  wire[0:0] mux_1403_nl;
  wire[0:0] nor_392_nl;
  wire[0:0] nor_393_nl;
  wire[0:0] mux_1402_nl;
  wire[0:0] nor_394_nl;
  wire[0:0] nor_395_nl;
  wire[0:0] mux_1410_nl;
  wire[0:0] mux_1409_nl;
  wire[0:0] nor_386_nl;
  wire[0:0] nor_387_nl;
  wire[0:0] nor_388_nl;
  wire[0:0] mux_1408_nl;
  wire[0:0] or_2024_nl;
  wire[0:0] or_2022_nl;
  wire[0:0] mux_1415_nl;
  wire[0:0] mux_1414_nl;
  wire[0:0] nor_380_nl;
  wire[0:0] nor_381_nl;
  wire[0:0] mux_1413_nl;
  wire[0:0] mux_1412_nl;
  wire[0:0] mux_1411_nl;
  wire[0:0] mux_1418_nl;
  wire[0:0] mux_1417_nl;
  wire[0:0] nor_377_nl;
  wire[0:0] nor_378_nl;
  wire[0:0] nor_379_nl;
  wire[0:0] mux_1416_nl;
  wire[0:0] or_2038_nl;
  wire[0:0] or_2036_nl;
  wire[0:0] mux_1425_nl;
  wire[0:0] mux_1424_nl;
  wire[0:0] mux_1423_nl;
  wire[0:0] nor_369_nl;
  wire[0:0] nor_370_nl;
  wire[0:0] mux_1422_nl;
  wire[0:0] nor_371_nl;
  wire[0:0] mux_1421_nl;
  wire[0:0] mux_1420_nl;
  wire[0:0] nor_373_nl;
  wire[0:0] mux_1419_nl;
  wire[0:0] nor_375_nl;
  wire[0:0] nor_376_nl;
  wire[0:0] mux_1428_nl;
  wire[0:0] mux_1427_nl;
  wire[0:0] nor_366_nl;
  wire[0:0] nor_367_nl;
  wire[0:0] nor_368_nl;
  wire[0:0] mux_1426_nl;
  wire[0:0] or_2054_nl;
  wire[0:0] or_2052_nl;
  wire[0:0] mux_1433_nl;
  wire[0:0] mux_1432_nl;
  wire[0:0] nor_360_nl;
  wire[0:0] nor_361_nl;
  wire[0:0] mux_1431_nl;
  wire[0:0] mux_1430_nl;
  wire[0:0] mux_1429_nl;
  wire[0:0] mux_1436_nl;
  wire[0:0] mux_1435_nl;
  wire[0:0] nor_357_nl;
  wire[0:0] nor_358_nl;
  wire[0:0] nor_359_nl;
  wire[0:0] mux_1434_nl;
  wire[0:0] or_2067_nl;
  wire[0:0] or_2066_nl;
  wire[0:0] mux_1442_nl;
  wire[0:0] mux_1441_nl;
  wire[0:0] mux_1440_nl;
  wire[0:0] nor_351_nl;
  wire[0:0] nor_352_nl;
  wire[0:0] nor_353_nl;
  wire[0:0] mux_1439_nl;
  wire[0:0] mux_1438_nl;
  wire[0:0] nor_354_nl;
  wire[0:0] nor_355_nl;
  wire[0:0] mux_1437_nl;
  wire[0:0] and_328_nl;
  wire[0:0] nor_356_nl;
  wire[0:0] mux_1445_nl;
  wire[0:0] mux_1444_nl;
  wire[0:0] and_327_nl;
  wire[0:0] nor_349_nl;
  wire[0:0] nor_350_nl;
  wire[0:0] mux_1443_nl;
  wire[0:0] nand_474_nl;
  wire[0:0] or_2080_nl;
  wire[0:0] mux_1450_nl;
  wire[0:0] mux_1449_nl;
  wire[0:0] and_323_nl;
  wire[0:0] and_324_nl;
  wire[0:0] mux_1448_nl;
  wire[0:0] mux_1447_nl;
  wire[0:0] mux_1446_nl;
  wire[0:0] mux_1453_nl;
  wire[0:0] mux_1452_nl;
  wire[0:0] and_321_nl;
  wire[0:0] and_322_nl;
  wire[0:0] nor_346_nl;
  wire[0:0] mux_1451_nl;
  wire[0:0] nand_192_nl;
  wire[0:0] nand_193_nl;
  wire[0:0] nand_520_nl;
  wire[0:0] mux_1600_nl;
  wire[6:0] COMP_LOOP_mux_382_nl;
  wire[0:0] and_755_nl;
  wire[11:0] acc_1_nl;
  wire[12:0] nl_acc_1_nl;
  wire[10:0] COMP_LOOP_mux_383_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_nand_1_nl;
  wire[9:0] COMP_LOOP_mux_384_nl;
  wire[3:0] STAGE_LOOP_mux_4_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_174_nl;
  wire[0:0] COMP_LOOP_tmp_mux_21_nl;
  wire[8:0] COMP_LOOP_tmp_mux1h_94_nl;
  wire[0:0] COMP_LOOP_tmp_or_76_nl;
  wire[0:0] COMP_LOOP_tmp_and_161_nl;
  wire[5:0] COMP_LOOP_tmp_mux1h_95_nl;
  wire[0:0] COMP_LOOP_tmp_or_77_nl;
  wire[0:0] COMP_LOOP_tmp_or_78_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_mux_18_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_or_1_nl;
  wire[63:0] COMP_LOOP_tmp_mux1h_96_nl;
  wire[0:0] and_756_nl;
  wire[63:0] COMP_LOOP_tmp_mux_22_nl;
  wire[0:0] COMP_LOOP_tmp_or_79_nl;
  wire[0:0] COMP_LOOP_mux1h_657_nl;
  wire[0:0] COMP_LOOP_mux1h_658_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_930_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_931_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_932_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_933_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_934_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_935_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_936_nl;
  wire[0:0] COMP_LOOP_mux1h_659_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_937_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_938_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_939_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_940_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_941_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_942_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_943_nl;
  wire[0:0] COMP_LOOP_mux1h_660_nl;
  wire[0:0] COMP_LOOP_mux1h_661_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_944_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_945_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_946_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_947_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_948_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_949_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_950_nl;
  wire[0:0] COMP_LOOP_mux1h_662_nl;
  wire[0:0] COMP_LOOP_mux1h_663_nl;
  wire[0:0] COMP_LOOP_mux1h_664_nl;
  wire[0:0] COMP_LOOP_mux1h_665_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_951_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_952_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_953_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_954_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_955_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_956_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_957_nl;
  wire[0:0] COMP_LOOP_mux1h_666_nl;
  wire[0:0] COMP_LOOP_mux1h_667_nl;
  wire[0:0] COMP_LOOP_mux1h_668_nl;
  wire[0:0] COMP_LOOP_mux1h_669_nl;
  wire[0:0] COMP_LOOP_mux1h_670_nl;
  wire[0:0] COMP_LOOP_mux1h_671_nl;
  wire[0:0] COMP_LOOP_mux1h_672_nl;
  wire[0:0] COMP_LOOP_mux1h_673_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_958_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_959_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_960_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_961_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_962_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_963_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_964_nl;
  wire[0:0] COMP_LOOP_mux1h_674_nl;
  wire[0:0] COMP_LOOP_mux1h_675_nl;
  wire[0:0] COMP_LOOP_mux1h_676_nl;
  wire[0:0] COMP_LOOP_mux1h_677_nl;
  wire[0:0] COMP_LOOP_mux1h_678_nl;
  wire[0:0] COMP_LOOP_mux1h_679_nl;
  wire[0:0] COMP_LOOP_mux1h_680_nl;
  wire[0:0] COMP_LOOP_mux1h_681_nl;
  wire[0:0] COMP_LOOP_mux1h_682_nl;
  wire[0:0] COMP_LOOP_mux1h_683_nl;
  wire[0:0] COMP_LOOP_mux1h_684_nl;
  wire[0:0] COMP_LOOP_mux1h_685_nl;
  wire[0:0] COMP_LOOP_mux1h_686_nl;
  wire[0:0] COMP_LOOP_mux1h_687_nl;
  wire[0:0] COMP_LOOP_mux1h_688_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[64:0] acc_4_nl;
  wire[65:0] nl_acc_4_nl;
  wire[63:0] COMP_LOOP_COMP_LOOP_mux_3_nl;
  wire[0:0] and_230_nl;
  wire[0:0] mux_1468_nl;
  wire[0:0] mux_1467_nl;
  wire[0:0] mux_1466_nl;
  wire[0:0] mux_1464_nl;
  wire[0:0] mux_1463_nl;
  wire[0:0] or_2103_nl;
  wire[0:0] COMP_LOOP_or_61_nl;
  wire [63:0] nl_COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat;
  assign COMP_LOOP_COMP_LOOP_mux_3_nl = MUX_v_64_2_2((~ COMP_LOOP_1_acc_8_itm), (~
      z_out_9), COMP_LOOP_or_33_itm);
  assign nl_acc_4_nl = ({COMP_LOOP_mux_385_cse , 1'b1}) + ({COMP_LOOP_COMP_LOOP_mux_3_nl
      , 1'b1});
  assign acc_4_nl = nl_acc_4_nl[64:0];
  assign mux_1466_nl = MUX_s_1_2_2((~ and_449_cse), mux_tmp_1430, fsm_output[4]);
  assign mux_1467_nl = MUX_s_1_2_2(mux_1466_nl, or_tmp_2025, fsm_output[2]);
  assign or_2103_nl = (~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[7]));
  assign mux_1463_nl = MUX_s_1_2_2(or_2103_nl, mux_tmp_1423, fsm_output[4]);
  assign mux_1464_nl = MUX_s_1_2_2(or_tmp_2025, mux_1463_nl, fsm_output[2]);
  assign mux_1468_nl = MUX_s_1_2_2(mux_1467_nl, mux_1464_nl, fsm_output[5]);
  assign and_230_nl = (~ mux_1468_nl) & and_dcpl_40;
  assign COMP_LOOP_or_61_nl = (and_dcpl_33 & and_dcpl_220) | (and_dcpl_33 & and_dcpl_223)
      | (and_dcpl_89 & and_dcpl_175) | (and_dcpl_89 & and_dcpl_36) | (and_dcpl_95
      & and_dcpl_30) | (and_dcpl_95 & and_dcpl_52) | (and_dcpl_95 & and_dcpl_56)
      | (and_dcpl_38 & and_dcpl_60);
  assign nl_COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat = MUX1HOT_v_64_3_2((readslicef_65_64_1(acc_4_nl)),
      COMP_LOOP_1_acc_8_itm, z_out_8, {COMP_LOOP_or_36_itm , and_230_nl , COMP_LOOP_or_61_nl});
  wire [63:0] nl_COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat;
  assign nl_COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat = p_sva;
  wire[0:0] mux_1478_nl;
  wire[0:0] mux_1477_nl;
  wire[0:0] mux_1476_nl;
  wire[0:0] or_2112_nl;
  wire[0:0] mux_1475_nl;
  wire[0:0] or_2111_nl;
  wire[0:0] mux_1474_nl;
  wire[0:0] mux_1473_nl;
  wire[0:0] or_2108_nl;
  wire[0:0] mux_1471_nl;
  wire[0:0] or_2106_nl;
  wire [0:0] nl_COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat;
  assign mux_1475_nl = MUX_s_1_2_2(or_145_cse, and_490_cse, fsm_output[0]);
  assign or_2112_nl = (fsm_output[3]) | (~ mux_1475_nl);
  assign mux_1476_nl = MUX_s_1_2_2(or_2112_nl, nand_tmp_184, fsm_output[6]);
  assign or_2111_nl = (fsm_output[6]) | mux_tmp_1437;
  assign mux_1477_nl = MUX_s_1_2_2(mux_1476_nl, or_2111_nl, fsm_output[5]);
  assign or_2108_nl = (fsm_output[3]) | (fsm_output[0]) | (~ and_490_cse);
  assign mux_1473_nl = MUX_s_1_2_2(mux_tmp_1437, or_2108_nl, fsm_output[6]);
  assign or_2106_nl = (fsm_output[3]) | (~((~ (fsm_output[0])) | (fsm_output[4])))
      | (fsm_output[7]);
  assign mux_1471_nl = MUX_s_1_2_2(nand_tmp_184, or_2106_nl, fsm_output[6]);
  assign mux_1474_nl = MUX_s_1_2_2(mux_1473_nl, mux_1471_nl, fsm_output[5]);
  assign mux_1478_nl = MUX_s_1_2_2(mux_1477_nl, mux_1474_nl, fsm_output[2]);
  assign nl_COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat = ~(mux_1478_nl |
      (fsm_output[1]));
  wire[0:0] and_541_nl;
  wire [3:0] nl_COMP_LOOP_5_tmp_lshift_rg_s;
  assign and_541_nl = (fsm_output==8'b00000010);
  assign nl_COMP_LOOP_5_tmp_lshift_rg_s = MUX_v_4_2_2(STAGE_LOOP_i_3_0_sva, z_out_4,
      and_541_nl);
  wire[0:0] COMP_LOOP_tmp_or_56_nl;
  wire [3:0] nl_COMP_LOOP_1_tmp_lshift_rg_s;
  assign COMP_LOOP_tmp_or_56_nl = (nor_1025_cse & (fsm_output[1:0]==2'b11) & and_dcpl_29
      & (~ (fsm_output[2])) & (~ (fsm_output[5]))) | (nor_1025_cse & (fsm_output[1:0]==2'b00)
      & and_dcpl_29 & (fsm_output[2]) & (~ (fsm_output[5])));
  assign nl_COMP_LOOP_1_tmp_lshift_rg_s = MUX_v_4_2_2(z_out_4, COMP_LOOP_1_tmp_acc_cse_sva,
      COMP_LOOP_tmp_or_56_nl);
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_28_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_28_tr0 = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_56_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_56_tr0 = ~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_84_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_84_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_112_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_112_tr0 = ~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_140_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_140_tr0 = ~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_168_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_168_tr0 = ~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_196_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_196_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_224_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_224_tr0 = ~ COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0 = z_out_3[10];
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0 = ~ (z_out_2[4]);
  ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd64)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_31_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_31_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_30_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_30_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_29_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_29_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_28_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_28_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_27_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_27_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_26_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_26_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_25_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_25_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_24_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_24_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_23_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_23_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_22_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_22_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_21_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_21_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_20_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_20_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_19_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_19_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_18_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_18_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_17_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_17_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_16_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_16_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_15_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_14_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_13_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_12_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_11_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_10_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_9_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_8_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_7_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_6_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_5_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_4_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_3_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_2_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_1_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(vec_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_31_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_31_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_30_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_30_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_29_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_29_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_28_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_28_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_27_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_27_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_26_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_26_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_25_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_25_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_24_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_24_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_23_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_23_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_22_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_22_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_21_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_21_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_20_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_20_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_19_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_19_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_18_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_18_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_17_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_17_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_16_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_16_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_15_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_14_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_13_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_12_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_11_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_10_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_9_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_8_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_7_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_6_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_5_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_4_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_3_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_2_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_1_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_0_lz)
    );
  modulo_dev  COMP_LOOP_1_modulo_dev_cmp (
      .base_rsc_dat(nl_COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat[63:0]),
      .m_rsc_dat(nl_COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat[63:0]),
      .return_rsc_z(COMP_LOOP_1_modulo_dev_cmp_return_rsc_z),
      .ccs_ccore_start_rsc_dat(nl_COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat[0:0]),
      .ccs_ccore_clk(clk),
      .ccs_ccore_srst(rst),
      .ccs_ccore_en(COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) COMP_LOOP_5_tmp_lshift_rg (
      .a(1'b1),
      .s(nl_COMP_LOOP_5_tmp_lshift_rg_s[3:0]),
      .z(z_out)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd10)) COMP_LOOP_1_tmp_lshift_rg (
      .a(1'b1),
      .s(nl_COMP_LOOP_1_tmp_lshift_rg_s[3:0]),
      .z(z_out_1)
    );
  inPlaceNTT_DIF_core_wait_dp inPlaceNTT_DIF_core_wait_dp_inst (
      .ensig_cgo_iro(mux_1462_rmff),
      .ensig_cgo(reg_ensig_cgo_cse),
      .COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en(COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en)
    );
  inPlaceNTT_DIF_core_core_fsm inPlaceNTT_DIF_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .COMP_LOOP_C_28_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_28_tr0[0:0]),
      .COMP_LOOP_C_56_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_56_tr0[0:0]),
      .COMP_LOOP_C_84_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_84_tr0[0:0]),
      .COMP_LOOP_C_112_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_112_tr0[0:0]),
      .COMP_LOOP_C_140_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_140_tr0[0:0]),
      .COMP_LOOP_C_168_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_168_tr0[0:0]),
      .COMP_LOOP_C_196_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_196_tr0[0:0]),
      .COMP_LOOP_C_224_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_224_tr0[0:0]),
      .VEC_LOOP_C_0_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0[0:0]),
      .STAGE_LOOP_C_1_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0[0:0])
    );
  assign and_449_cse = (fsm_output[3]) & (fsm_output[6]) & (fsm_output[7]);
  assign or_285_cse = (~ (fsm_output[4])) | (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b000)
      | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) | (fsm_output[7:6]!=2'b01);
  assign mux_347_nl = MUX_s_1_2_2(or_285_cse, mux_tmp_311, fsm_output[3]);
  assign nand_11_nl = ~((fsm_output[3]) & (~ mux_tmp_311));
  assign mux_348_cse = MUX_s_1_2_2(mux_347_nl, nand_11_nl, VEC_LOOP_j_10_0_sva_9_0[1]);
  assign nand_443_cse = ~((fsm_output[7:6]==2'b11));
  assign nand_444_cse = ~((COMP_LOOP_acc_10_cse_10_1_sva[0]) & (fsm_output[7:6]==2'b11));
  assign nand_22_nl = ~((fsm_output[3]) & (~ mux_tmp_373));
  assign mux_409_nl = MUX_s_1_2_2(or_285_cse, mux_tmp_373, fsm_output[3]);
  assign mux_410_cse = MUX_s_1_2_2(nand_22_nl, mux_409_nl, VEC_LOOP_j_10_0_sva_9_0[1]);
  assign or_493_cse = (~ (fsm_output[4])) | (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b001)
      | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) | (fsm_output[7:6]!=2'b01);
  assign mux_471_nl = MUX_s_1_2_2(or_493_cse, mux_tmp_435, fsm_output[3]);
  assign nand_33_nl = ~((fsm_output[3]) & (~ mux_tmp_435));
  assign mux_472_cse = MUX_s_1_2_2(mux_471_nl, nand_33_nl, VEC_LOOP_j_10_0_sva_9_0[1]);
  assign nand_44_nl = ~((fsm_output[3]) & (~ mux_tmp_497));
  assign mux_533_nl = MUX_s_1_2_2(or_493_cse, mux_tmp_497, fsm_output[3]);
  assign mux_534_cse = MUX_s_1_2_2(nand_44_nl, mux_533_nl, VEC_LOOP_j_10_0_sva_9_0[1]);
  assign or_701_cse = (~ (fsm_output[4])) | (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b010)
      | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) | (fsm_output[7:6]!=2'b01);
  assign mux_595_nl = MUX_s_1_2_2(or_701_cse, mux_tmp_559, fsm_output[3]);
  assign nand_55_nl = ~((fsm_output[3]) & (~ mux_tmp_559));
  assign mux_596_cse = MUX_s_1_2_2(mux_595_nl, nand_55_nl, VEC_LOOP_j_10_0_sva_9_0[1]);
  assign nand_66_nl = ~((fsm_output[3]) & (~ mux_tmp_621));
  assign mux_657_nl = MUX_s_1_2_2(or_701_cse, mux_tmp_621, fsm_output[3]);
  assign mux_658_cse = MUX_s_1_2_2(nand_66_nl, mux_657_nl, VEC_LOOP_j_10_0_sva_9_0[1]);
  assign nand_394_cse = ~((fsm_output[4]) & (COMP_LOOP_acc_13_psp_sva[2:0]==3'b011)
      & COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm & (fsm_output[7:6]==2'b01));
  assign mux_719_nl = MUX_s_1_2_2(nand_394_cse, mux_tmp_683, fsm_output[3]);
  assign nand_77_nl = ~((fsm_output[3]) & (~ mux_tmp_683));
  assign mux_720_cse = MUX_s_1_2_2(mux_719_nl, nand_77_nl, VEC_LOOP_j_10_0_sva_9_0[1]);
  assign nand_88_nl = ~((fsm_output[3]) & (~ mux_tmp_745));
  assign mux_781_nl = MUX_s_1_2_2(nand_394_cse, mux_tmp_745, fsm_output[3]);
  assign mux_782_cse = MUX_s_1_2_2(nand_88_nl, mux_781_nl, VEC_LOOP_j_10_0_sva_9_0[1]);
  assign nand_371_cse = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:1]==4'b0111));
  assign or_1066_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | nand_365_cse;
  assign or_1064_nl = (COMP_LOOP_acc_psp_sva[0]) | (VEC_LOOP_j_10_0_sva_9_0[2]) |
      (~ (COMP_LOOP_acc_psp_sva[1])) | (fsm_output[7]);
  assign mux_818_cse = MUX_s_1_2_2(or_1066_nl, or_1064_nl, fsm_output[4]);
  assign or_1113_cse = (~ (fsm_output[4])) | (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b100)
      | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) | (fsm_output[7:6]!=2'b01);
  assign mux_843_nl = MUX_s_1_2_2(or_1113_cse, mux_tmp_807, fsm_output[3]);
  assign nand_99_nl = ~((fsm_output[3]) & (~ mux_tmp_807));
  assign mux_844_cse = MUX_s_1_2_2(mux_843_nl, nand_99_nl, VEC_LOOP_j_10_0_sva_9_0[1]);
  assign nor_730_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | nand_365_cse);
  assign nor_731_nl = ~((COMP_LOOP_acc_psp_sva[0]) | (VEC_LOOP_j_10_0_sva_9_0[2])
      | (~ (COMP_LOOP_acc_psp_sva[1])) | (fsm_output[7]));
  assign mux_849_cse = MUX_s_1_2_2(nor_730_nl, nor_731_nl, fsm_output[4]);
  assign nand_356_cse = ~((COMP_LOOP_acc_10_cse_10_1_sva[4]) & (COMP_LOOP_acc_10_cse_10_1_sva[0])
      & (fsm_output[7:6]==2'b11));
  assign nand_110_nl = ~((fsm_output[3]) & (~ mux_tmp_869));
  assign mux_905_nl = MUX_s_1_2_2(or_1113_cse, mux_tmp_869, fsm_output[3]);
  assign mux_906_cse = MUX_s_1_2_2(nand_110_nl, mux_905_nl, VEC_LOOP_j_10_0_sva_9_0[1]);
  assign or_1274_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | nand_365_cse;
  assign or_1272_nl = (COMP_LOOP_acc_psp_sva[0]) | (~ (VEC_LOOP_j_10_0_sva_9_0[2]))
      | (~ (COMP_LOOP_acc_psp_sva[1])) | (fsm_output[7]);
  assign mux_942_cse = MUX_s_1_2_2(or_1274_nl, or_1272_nl, fsm_output[4]);
  assign nand_336_cse = ~((fsm_output[4]) & (COMP_LOOP_acc_13_psp_sva[2:0]==3'b101)
      & COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm & (fsm_output[7:6]==2'b01));
  assign mux_967_nl = MUX_s_1_2_2(nand_336_cse, mux_tmp_931, fsm_output[3]);
  assign nand_121_nl = ~((fsm_output[3]) & (~ mux_tmp_931));
  assign mux_968_cse = MUX_s_1_2_2(mux_967_nl, nand_121_nl, VEC_LOOP_j_10_0_sva_9_0[1]);
  assign nor_662_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | nand_365_cse);
  assign nor_663_nl = ~((COMP_LOOP_acc_psp_sva[0]) | (~ (VEC_LOOP_j_10_0_sva_9_0[2]))
      | (~ (COMP_LOOP_acc_psp_sva[1])) | (fsm_output[7]));
  assign mux_973_cse = MUX_s_1_2_2(nor_662_nl, nor_663_nl, fsm_output[4]);
  assign nand_132_nl = ~((fsm_output[3]) & (~ mux_tmp_993));
  assign mux_1029_nl = MUX_s_1_2_2(nand_336_cse, mux_tmp_993, fsm_output[3]);
  assign mux_1030_cse = MUX_s_1_2_2(nand_132_nl, mux_1029_nl, VEC_LOOP_j_10_0_sva_9_0[1]);
  assign or_1481_nl = (COMP_LOOP_acc_13_psp_sva[0]) | nand_303_cse;
  assign or_1480_nl = (~ (COMP_LOOP_acc_psp_sva[0])) | (VEC_LOOP_j_10_0_sva_9_0[2])
      | (~ (COMP_LOOP_acc_psp_sva[1])) | (fsm_output[7]);
  assign mux_1066_cse = MUX_s_1_2_2(or_1481_nl, or_1480_nl, fsm_output[4]);
  assign nand_300_cse = ~((fsm_output[4]) & (COMP_LOOP_acc_13_psp_sva[2:0]==3'b110)
      & COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm & (fsm_output[7:6]==2'b01));
  assign mux_1091_nl = MUX_s_1_2_2(nand_300_cse, mux_tmp_1055, fsm_output[3]);
  assign nand_143_nl = ~((fsm_output[3]) & (~ mux_tmp_1055));
  assign mux_1092_cse = MUX_s_1_2_2(mux_1091_nl, nand_143_nl, VEC_LOOP_j_10_0_sva_9_0[1]);
  assign nor_595_nl = ~((COMP_LOOP_acc_13_psp_sva[0]) | nand_303_cse);
  assign nor_596_nl = ~((~ (COMP_LOOP_acc_psp_sva[0])) | (VEC_LOOP_j_10_0_sva_9_0[2])
      | (~ (COMP_LOOP_acc_psp_sva[1])) | (fsm_output[7]));
  assign mux_1097_cse = MUX_s_1_2_2(nor_595_nl, nor_596_nl, fsm_output[4]);
  assign nand_293_cse = ~((COMP_LOOP_acc_10_cse_10_1_sva[3]) & (COMP_LOOP_acc_10_cse_10_1_sva[4])
      & (COMP_LOOP_acc_10_cse_10_1_sva[0]) & (fsm_output[7:6]==2'b11));
  assign nand_154_nl = ~((fsm_output[3]) & (~ mux_tmp_1117));
  assign mux_1153_nl = MUX_s_1_2_2(nand_300_cse, mux_tmp_1117, fsm_output[3]);
  assign mux_1154_cse = MUX_s_1_2_2(nand_154_nl, mux_1153_nl, VEC_LOOP_j_10_0_sva_9_0[1]);
  assign nand_264_cse = ~((fsm_output[4]) & (COMP_LOOP_acc_13_psp_sva[2:0]==3'b111)
      & COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm & (fsm_output[7:6]==2'b01));
  assign mux_1215_nl = MUX_s_1_2_2(nand_264_cse, mux_tmp_1179, fsm_output[3]);
  assign nand_165_nl = ~((fsm_output[3]) & (~ mux_tmp_1179));
  assign mux_1216_cse = MUX_s_1_2_2(mux_1215_nl, nand_165_nl, VEC_LOOP_j_10_0_sva_9_0[1]);
  assign nand_176_nl = ~((fsm_output[3]) & (~ mux_tmp_1241));
  assign mux_1277_nl = MUX_s_1_2_2(nand_264_cse, mux_tmp_1241, fsm_output[3]);
  assign mux_1278_cse = MUX_s_1_2_2(nand_176_nl, mux_1277_nl, VEC_LOOP_j_10_0_sva_9_0[1]);
  assign nand_204_cse = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[3]) & (fsm_output[3]));
  assign nand_205_cse = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[4]) & (fsm_output[3]));
  assign mux_1460_nl = MUX_s_1_2_2(mux_tmp_1424, mux_tmp_1423, fsm_output[4]);
  assign mux_1461_nl = MUX_s_1_2_2(or_tmp_2025, mux_1460_nl, fsm_output[2]);
  assign mux_1455_nl = MUX_s_1_2_2((fsm_output[6]), mux_189_cse, fsm_output[3]);
  assign mux_1456_nl = MUX_s_1_2_2(and_456_cse, mux_1455_nl, fsm_output[4]);
  assign mux_1457_nl = MUX_s_1_2_2(mux_1456_nl, and_464_cse, fsm_output[2]);
  assign mux_1462_rmff = MUX_s_1_2_2(mux_1461_nl, (~ mux_1457_nl), fsm_output[5]);
  assign or_220_cse = (fsm_output[4:2]!=3'b000);
  assign or_212_cse = (fsm_output[4:3]!=2'b00);
  assign and_316_cse = (fsm_output[1:0]==2'b11);
  assign nor_1023_cse = ~((fsm_output[2]) | (fsm_output[4]));
  assign and_496_cse = (fsm_output[1]) & (fsm_output[3]);
  assign or_32_cse = (fsm_output[1:0]!=2'b00);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse = ~((z_out_7[2:0]!=3'b000));
  assign and_491_cse = ((fsm_output[4]) | (fsm_output[6]) | (fsm_output[3])) & (fsm_output[7]);
  assign mux_189_cse = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[6]);
  assign and_33_cse = (fsm_output[6]) & or_212_cse & (fsm_output[7]);
  assign and_464_cse = (fsm_output[7:6]==2'b11);
  assign COMP_LOOP_tmp_or_cse = and_dcpl_46 | and_dcpl_49 | and_dcpl_171 | and_dcpl_172
      | and_dcpl_173 | and_dcpl_176;
  assign COMP_LOOP_or_59_cse = and_dcpl_172 | and_dcpl_176;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse = (z_out_7[4:0]==5'b01001);
  assign COMP_LOOP_tmp_nor_27_cse = ~((z_out_7[3:2]!=2'b00));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse = (z_out_7[4:0]==5'b01110);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse = (z_out_7[4:0]==5'b00011);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_36_cse = (z_out_7[1:0]==2'b11) & COMP_LOOP_tmp_nor_27_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse = (z_out_7[4:0]==5'b01010);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_cse = (z_out_7[4:0]==5'b01111);
  assign COMP_LOOP_tmp_nor_29_cse = ~((z_out_7[3]) | (z_out_7[1]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse = (z_out_7[4:0]==5'b00101);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_38_cse = (z_out_7[2]) & (z_out_7[0]) & COMP_LOOP_tmp_nor_29_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse = (z_out_7[4:0]==5'b01011);
  assign COMP_LOOP_tmp_nor_78_cse = ~((z_out_7[3:1]!=3'b000));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse = (z_out_7[4]) & (z_out_7[0]) &
      COMP_LOOP_tmp_nor_78_cse;
  assign COMP_LOOP_tmp_nor_30_cse = ~((z_out_7[3]) | (z_out_7[0]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse = (z_out_7[4:0]==5'b00110);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_39_cse = (z_out_7[2:1]==2'b11) & COMP_LOOP_tmp_nor_30_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse = (z_out_7[4:0]==5'b01100);
  assign COMP_LOOP_tmp_nor_79_cse = ~((z_out_7[3]) | (z_out_7[2]) | (z_out_7[0]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_cse = (z_out_7[4]) & (z_out_7[1]) &
      COMP_LOOP_tmp_nor_79_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_40_cse = (z_out_7[3:0]==4'b0111);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse = (z_out_7[4:0]==5'b00111);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse = (z_out_7[4:0]==5'b01101);
  assign COMP_LOOP_tmp_nor_32_cse = ~((z_out_7[2:1]!=2'b00));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_cse = (z_out_7[4]) & (z_out_7[1]) &
      (z_out_7[0]) & COMP_LOOP_tmp_nor_27_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_42_cse = (z_out_7[3]) & (z_out_7[0]) & COMP_LOOP_tmp_nor_32_cse;
  assign COMP_LOOP_tmp_nor_81_cse = ~((z_out_7[3]) | (z_out_7[1]) | (z_out_7[0]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_cse = (z_out_7[4]) & (z_out_7[2]) &
      COMP_LOOP_tmp_nor_81_cse;
  assign COMP_LOOP_tmp_nor_33_cse = ~((z_out_7[2]) | (z_out_7[0]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_43_cse = (z_out_7[3]) & (z_out_7[1]) & COMP_LOOP_tmp_nor_33_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_44_cse = (z_out_7[3:0]==4'b1011);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_cse = (z_out_7[4]) & (z_out_7[2]) &
      (z_out_7[0]) & COMP_LOOP_tmp_nor_29_cse;
  assign COMP_LOOP_tmp_nor_34_cse = ~((z_out_7[1:0]!=2'b00));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_cse = (z_out_7[4]) & (z_out_7[2]) &
      (z_out_7[1]) & COMP_LOOP_tmp_nor_30_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_45_cse = (z_out_7[3:2]==2'b11) & COMP_LOOP_tmp_nor_34_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_cse = (z_out_7[4:0]==5'b10111);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_46_cse = (z_out_7[3:0]==4'b1101);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_47_cse = (z_out_7[3:0]==4'b1110);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse = (z_out_7[4:3]==2'b11) & COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_48_cse = (z_out_7[3:0]==4'b1111);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_cse = (z_out_7[4]) & (z_out_7[3]) &
      (z_out_7[0]) & COMP_LOOP_tmp_nor_32_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse = ~((z_out_7[3:0]!=4'b0000));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_cse = (z_out_7[4]) & (z_out_7[3]) &
      (z_out_7[1]) & COMP_LOOP_tmp_nor_33_cse;
  assign COMP_LOOP_tmp_or_12_cse = and_dcpl_46 | and_dcpl_49 | and_dcpl_172 | and_dcpl_173
      | and_dcpl_176;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_cse = (z_out_7[4:0]==5'b11011);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_cse = (z_out_7[4:2]==3'b111) & COMP_LOOP_tmp_nor_34_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_cse = (z_out_7[4:0]==5'b11101);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_cse = (z_out_7[4:0]==5'b11110);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_cse = (z_out_7[4:0]==5'b11111);
  assign COMP_LOOP_tmp_or_17_cse = and_dcpl_46 | and_dcpl_49 | and_dcpl_172 | and_dcpl_174;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_cse = ~((z_out_7[4:0]!=5'b00000));
  assign COMP_LOOP_or_42_cse = and_dcpl_49 | and_dcpl_172;
  assign COMP_LOOP_tmp_nor_1_cse = ~((z_out_7[4]) | (z_out_7[3]) | (z_out_7[2]) |
      (z_out_7[0]));
  assign COMP_LOOP_or_41_cse = and_dcpl_172 | and_dcpl_173;
  assign COMP_LOOP_tmp_nor_101_cse = ~((z_out_7[4]) | (z_out_7[3]) | (z_out_7[1])
      | (z_out_7[0]));
  assign COMP_LOOP_tmp_nor_35_cse = ~((z_out_7[4:1]!=4'b0000));
  assign COMP_LOOP_tmp_nor_105_cse = ~((z_out_7[4]) | (z_out_7[2]) | (z_out_7[1])
      | (z_out_7[0]));
  assign COMP_LOOP_or_39_cse = and_dcpl_49 | and_dcpl_172 | and_dcpl_173;
  assign COMP_LOOP_or_36_itm = and_dcpl_171 | and_dcpl_222 | and_dcpl_226 | and_dcpl_229
      | and_dcpl_232 | and_dcpl_234 | and_dcpl_236 | and_dcpl_238;
  assign COMP_LOOP_tmp_or_35_cse = and_dcpl_171 | and_dcpl_174;
  assign COMP_LOOP_tmp_or_40_cse = and_dcpl_173 | and_dcpl_176;
  assign and_298_m1c = and_dcpl_45 & and_dcpl_175;
  assign and_1_cse = (COMP_LOOP_2_tmp_mul_idiv_sva[0]) & COMP_LOOP_tmp_nor_1_itm;
  assign nor_1025_cse = ~((fsm_output[7:6]!=2'b00));
  assign and_456_cse = ((fsm_output[3]) | (fsm_output[6])) & (fsm_output[7]);
  assign mux_1588_nl = MUX_s_1_2_2(mux_189_cse, and_464_cse, or_32_cse);
  assign mux_1589_nl = MUX_s_1_2_2(mux_189_cse, mux_1588_nl, fsm_output[3]);
  assign mux_1590_nl = MUX_s_1_2_2(mux_1589_nl, and_464_cse, fsm_output[4]);
  assign mux_1586_nl = MUX_s_1_2_2(mux_189_cse, and_464_cse, fsm_output[3]);
  assign mux_1587_nl = MUX_s_1_2_2(mux_1586_nl, and_456_cse, fsm_output[4]);
  assign mux_1591_nl = MUX_s_1_2_2(mux_1590_nl, mux_1587_nl, fsm_output[2]);
  assign mux_1592_tmp = MUX_s_1_2_2(mux_1591_nl, (fsm_output[7]), fsm_output[5]);
  assign and_490_cse = (fsm_output[4]) & (fsm_output[7]);
  assign or_167_cse = (fsm_output[7:6]!=2'b01);
  assign nl_COMP_LOOP_1_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_3_sva_6_0
      , 3'b000}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_1_acc_10_nl = nl_COMP_LOOP_1_acc_10_nl[10:0];
  assign COMP_LOOP_1_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_1_acc_10_nl);
  assign nl_COMP_LOOP_acc_psp_sva_mx0w0 = (VEC_LOOP_j_10_0_sva_9_0[9:3]) + COMP_LOOP_k_10_3_sva_6_0;
  assign COMP_LOOP_acc_psp_sva_mx0w0 = nl_COMP_LOOP_acc_psp_sva_mx0w0[6:0];
  assign nl_COMP_LOOP_acc_1_cse_6_sva_1 = VEC_LOOP_j_10_0_sva_9_0 + ({COMP_LOOP_k_10_3_sva_6_0
      , 3'b101});
  assign COMP_LOOP_acc_1_cse_6_sva_1 = nl_COMP_LOOP_acc_1_cse_6_sva_1[9:0];
  assign nl_COMP_LOOP_acc_1_cse_4_sva_1 = VEC_LOOP_j_10_0_sva_9_0 + ({COMP_LOOP_k_10_3_sva_6_0
      , 3'b011});
  assign COMP_LOOP_acc_1_cse_4_sva_1 = nl_COMP_LOOP_acc_1_cse_4_sva_1[9:0];
  assign nl_COMP_LOOP_acc_1_cse_2_sva_1 = VEC_LOOP_j_10_0_sva_9_0 + ({COMP_LOOP_k_10_3_sva_6_0
      , 3'b001});
  assign COMP_LOOP_acc_1_cse_2_sva_1 = nl_COMP_LOOP_acc_1_cse_2_sva_1[9:0];
  assign nl_COMP_LOOP_2_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_3_sva_6_0
      , 3'b001}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_2_acc_10_nl = nl_COMP_LOOP_2_acc_10_nl[10:0];
  assign COMP_LOOP_2_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_2_acc_10_nl);
  assign nl_COMP_LOOP_3_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_3_sva_6_0
      , 3'b010}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_3_acc_10_nl = nl_COMP_LOOP_3_acc_10_nl[10:0];
  assign COMP_LOOP_3_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_3_acc_10_nl);
  assign nl_COMP_LOOP_4_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_3_sva_6_0
      , 3'b011}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_4_acc_10_nl = nl_COMP_LOOP_4_acc_10_nl[10:0];
  assign COMP_LOOP_4_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_4_acc_10_nl);
  assign nl_COMP_LOOP_5_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_3_sva_6_0
      , 3'b100}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_5_acc_10_nl = nl_COMP_LOOP_5_acc_10_nl[10:0];
  assign COMP_LOOP_5_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_5_acc_10_nl);
  assign nl_COMP_LOOP_6_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_3_sva_6_0
      , 3'b101}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_6_acc_10_nl = nl_COMP_LOOP_6_acc_10_nl[10:0];
  assign COMP_LOOP_6_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_6_acc_10_nl);
  assign nl_COMP_LOOP_7_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_3_sva_6_0
      , 3'b110}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_7_acc_10_nl = nl_COMP_LOOP_7_acc_10_nl[10:0];
  assign COMP_LOOP_7_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_7_acc_10_nl);
  assign nl_COMP_LOOP_8_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_3_sva_6_0
      , 3'b111}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_8_acc_10_nl = nl_COMP_LOOP_8_acc_10_nl[10:0];
  assign COMP_LOOP_8_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_8_acc_10_nl);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_rgt = (COMP_LOOP_2_tmp_lshift_ncse_sva[1])
      & COMP_LOOP_tmp_nor_49_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_rgt = (COMP_LOOP_2_tmp_lshift_ncse_sva[2])
      & COMP_LOOP_tmp_nor_1_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_rgt = (COMP_LOOP_2_tmp_lshift_ncse_sva[3])
      & COMP_LOOP_tmp_nor_14_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_rgt = (COMP_LOOP_2_tmp_lshift_ncse_sva[4])
      & COMP_LOOP_tmp_nor_3_itm;
  assign and_4_cse = (COMP_LOOP_2_tmp_mul_idiv_sva[1]) & COMP_LOOP_tmp_nor_14_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_119_rgt = (COMP_LOOP_3_tmp_lshift_ncse_sva[1])
      & COMP_LOOP_tmp_nor_26_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_121_rgt = (COMP_LOOP_3_tmp_lshift_ncse_sva[2])
      & COMP_LOOP_tmp_nor_28_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_125_rgt = (COMP_LOOP_3_tmp_lshift_ncse_sva[3])
      & COMP_LOOP_tmp_nor_31_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_165 = (COMP_LOOP_2_tmp_mul_idiv_sva[4])
      & COMP_LOOP_tmp_nor_49_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_167 = (COMP_LOOP_2_tmp_mul_idiv_sva[3])
      & COMP_LOOP_tmp_nor_42_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_169 = (COMP_LOOP_2_tmp_mul_idiv_sva[2])
      & COMP_LOOP_tmp_nor_3_itm;
  assign nor_tmp_53 = ((fsm_output[6]) | (fsm_output[4])) & (fsm_output[7]);
  assign or_145_cse = (fsm_output[4]) | (fsm_output[7]);
  assign and_485_cse = (fsm_output[6]) & (fsm_output[4]);
  assign and_479_cse = (fsm_output[4:3]==2'b11);
  assign or_tmp_142 = (fsm_output[7:6]!=2'b00);
  assign and_dcpl_28 = ~((fsm_output[2]) | (fsm_output[5]));
  assign and_dcpl_29 = ~((fsm_output[4:3]!=2'b00));
  assign and_dcpl_30 = and_dcpl_29 & and_dcpl_28;
  assign and_dcpl_31 = ~((fsm_output[1:0]!=2'b00));
  assign and_dcpl_33 = nor_1025_cse & and_dcpl_31;
  assign and_dcpl_35 = (fsm_output[2]) & (fsm_output[5]);
  assign and_dcpl_36 = and_dcpl_29 & and_dcpl_35;
  assign and_dcpl_38 = and_464_cse & and_dcpl_31;
  assign nor_tmp_95 = ((fsm_output[4]) | (fsm_output[3]) | (fsm_output[0]) | (fsm_output[1]))
      & (fsm_output[7:6]==2'b11);
  assign and_dcpl_40 = (fsm_output[1:0]==2'b01);
  assign and_dcpl_44 = (fsm_output[1:0]==2'b10);
  assign and_dcpl_45 = nor_1025_cse & and_dcpl_44;
  assign and_dcpl_46 = and_dcpl_45 & and_dcpl_30;
  assign and_dcpl_48 = nor_1025_cse & and_316_cse;
  assign and_dcpl_49 = and_dcpl_48 & and_dcpl_30;
  assign and_dcpl_50 = (fsm_output[2]) & (~ (fsm_output[5]));
  assign and_dcpl_52 = and_479_cse & and_dcpl_50;
  assign and_dcpl_54 = and_dcpl_48 & and_dcpl_52;
  assign and_dcpl_55 = (~ (fsm_output[2])) & (fsm_output[5]);
  assign and_dcpl_56 = and_479_cse & and_dcpl_55;
  assign and_dcpl_58 = and_dcpl_48 & and_dcpl_56;
  assign and_dcpl_59 = (fsm_output[4:3]==2'b10);
  assign and_dcpl_60 = and_dcpl_59 & and_dcpl_50;
  assign and_dcpl_61 = (fsm_output[7:6]==2'b01);
  assign and_dcpl_62 = and_dcpl_61 & and_dcpl_44;
  assign and_dcpl_64 = and_dcpl_61 & and_316_cse;
  assign and_dcpl_65 = and_dcpl_64 & and_dcpl_60;
  assign and_dcpl_66 = and_dcpl_59 & and_dcpl_55;
  assign and_dcpl_68 = and_dcpl_64 & and_dcpl_66;
  assign and_dcpl_69 = (fsm_output[4:3]==2'b01);
  assign and_dcpl_70 = and_dcpl_69 & and_dcpl_50;
  assign and_dcpl_71 = (fsm_output[7:6]==2'b10);
  assign and_dcpl_72 = and_dcpl_71 & and_dcpl_44;
  assign and_dcpl_74 = and_dcpl_71 & and_316_cse;
  assign and_dcpl_75 = and_dcpl_74 & and_dcpl_70;
  assign and_dcpl_76 = and_dcpl_69 & and_dcpl_55;
  assign and_dcpl_78 = and_dcpl_74 & and_dcpl_76;
  assign and_dcpl_79 = and_dcpl_29 & and_dcpl_50;
  assign and_dcpl_82 = and_464_cse & and_316_cse;
  assign and_dcpl_83 = and_dcpl_82 & and_dcpl_79;
  assign and_dcpl_85 = nor_1025_cse & and_dcpl_40;
  assign and_dcpl_89 = and_dcpl_61 & and_dcpl_31;
  assign and_dcpl_91 = and_dcpl_61 & and_dcpl_40;
  assign and_dcpl_95 = and_dcpl_71 & and_dcpl_31;
  assign and_dcpl_97 = and_dcpl_71 & and_dcpl_40;
  assign and_dcpl_102 = and_464_cse & and_dcpl_40;
  assign and_dcpl_104 = and_dcpl_29 & and_dcpl_55;
  assign or_238_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b000) | (~ (fsm_output[7]));
  assign or_236_nl = (COMP_LOOP_acc_psp_sva[0]) | (VEC_LOOP_j_10_0_sva_9_0[2]) |
      (COMP_LOOP_acc_psp_sva[1]) | (fsm_output[7]);
  assign mux_322_cse = MUX_s_1_2_2(or_238_nl, or_236_nl, fsm_output[4]);
  assign or_284_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b0000) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_282_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0000) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_tmp_311 = MUX_s_1_2_2(or_284_nl, or_282_nl, fsm_output[4]);
  assign nand_445_cse = ~((COMP_LOOP_acc_10_cse_10_1_sva[0]) & (fsm_output[7]));
  assign nand_447_cse = ~((COMP_LOOP_acc_1_cse_6_sva[0]) & (fsm_output[7]));
  assign nor_1001_nl = ~((COMP_LOOP_acc_13_psp_sva[2:0]!=3'b000) | (~ (fsm_output[7])));
  assign nor_1002_nl = ~((COMP_LOOP_acc_psp_sva[0]) | (VEC_LOOP_j_10_0_sva_9_0[2])
      | (COMP_LOOP_acc_psp_sva[1]) | (fsm_output[7]));
  assign mux_353_cse = MUX_s_1_2_2(nor_1001_nl, nor_1002_nl, fsm_output[4]);
  assign nand_446_cse = ~((COMP_LOOP_acc_1_cse_sva[0]) & (fsm_output[7]));
  assign nand_448_cse = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[0]) & (fsm_output[7]));
  assign nor_98_cse = ~((VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01));
  assign nand_441_cse = ~((COMP_LOOP_acc_14_psp_sva[0]) & (fsm_output[7]));
  assign nand_442_cse = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[1]) & (fsm_output[7]));
  assign or_388_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b0001) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_386_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0001) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_tmp_373 = MUX_s_1_2_2(or_388_nl, or_386_nl, fsm_output[4]);
  assign nand_435_cse = ~((COMP_LOOP_acc_1_cse_sva[1:0]==2'b11) & (fsm_output[7]));
  assign nand_437_cse = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[1:0]==2'b11) & (fsm_output[7]));
  assign or_446_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b001) | (~ (fsm_output[7]));
  assign or_444_nl = (COMP_LOOP_acc_psp_sva[0]) | (~ (VEC_LOOP_j_10_0_sva_9_0[2]))
      | (COMP_LOOP_acc_psp_sva[1]) | (fsm_output[7]);
  assign mux_446_cse = MUX_s_1_2_2(or_446_nl, or_444_nl, fsm_output[4]);
  assign or_492_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b0010) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_490_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0010) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_tmp_435 = MUX_s_1_2_2(or_492_nl, or_490_nl, fsm_output[4]);
  assign nor_933_nl = ~((COMP_LOOP_acc_13_psp_sva[2:0]!=3'b001) | (~ (fsm_output[7])));
  assign nor_934_nl = ~((COMP_LOOP_acc_psp_sva[0]) | (~ (VEC_LOOP_j_10_0_sva_9_0[2]))
      | (COMP_LOOP_acc_psp_sva[1]) | (fsm_output[7]));
  assign mux_477_cse = MUX_s_1_2_2(nor_933_nl, nor_934_nl, fsm_output[4]);
  assign nand_423_cse = ~((COMP_LOOP_acc_14_psp_sva[1:0]==2'b11) & (fsm_output[7]));
  assign or_596_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b0011) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_594_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0011) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_tmp_497 = MUX_s_1_2_2(or_596_nl, or_594_nl, fsm_output[4]);
  assign nand_417_cse = ~((COMP_LOOP_acc_1_cse_sva[2:0]==3'b111) & (fsm_output[7]));
  assign nand_419_cse = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[2:0]==3'b111) & (fsm_output[7]));
  assign or_654_nl = (COMP_LOOP_acc_13_psp_sva[2:0]!=3'b010) | (~ (fsm_output[7]));
  assign or_652_nl = (~ (COMP_LOOP_acc_psp_sva[0])) | (VEC_LOOP_j_10_0_sva_9_0[2])
      | (COMP_LOOP_acc_psp_sva[1]) | (fsm_output[7]);
  assign mux_570_cse = MUX_s_1_2_2(or_654_nl, or_652_nl, fsm_output[4]);
  assign or_700_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b0100) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_698_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0100) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_tmp_559 = MUX_s_1_2_2(or_700_nl, or_698_nl, fsm_output[4]);
  assign nand_411_cse = ~((COMP_LOOP_acc_1_cse_6_sva[3]) & (COMP_LOOP_acc_1_cse_6_sva[0])
      & (fsm_output[7]));
  assign nor_865_nl = ~((COMP_LOOP_acc_13_psp_sva[2:0]!=3'b010) | (~ (fsm_output[7])));
  assign nor_866_nl = ~((~ (COMP_LOOP_acc_psp_sva[0])) | (VEC_LOOP_j_10_0_sva_9_0[2])
      | (COMP_LOOP_acc_psp_sva[1]) | (fsm_output[7]));
  assign mux_601_cse = MUX_s_1_2_2(nor_865_nl, nor_866_nl, fsm_output[4]);
  assign or_804_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b0101) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_802_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0101) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_tmp_621 = MUX_s_1_2_2(or_804_nl, or_802_nl, fsm_output[4]);
  assign nand_518_nl = ~((COMP_LOOP_acc_13_psp_sva[2:0]==3'b011) & (fsm_output[7]));
  assign or_860_nl = (~ (COMP_LOOP_acc_psp_sva[0])) | (~ (VEC_LOOP_j_10_0_sva_9_0[2]))
      | (COMP_LOOP_acc_psp_sva[1]) | (fsm_output[7]);
  assign mux_694_cse = MUX_s_1_2_2(nand_518_nl, or_860_nl, fsm_output[4]);
  assign or_908_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b0110) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_906_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0110) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_tmp_683 = MUX_s_1_2_2(or_908_nl, or_906_nl, fsm_output[4]);
  assign and_532_nl = (COMP_LOOP_acc_13_psp_sva[2:0]==3'b011) & (fsm_output[7]);
  assign nor_798_nl = ~((~ (COMP_LOOP_acc_psp_sva[0])) | (~ (VEC_LOOP_j_10_0_sva_9_0[2]))
      | (COMP_LOOP_acc_psp_sva[1]) | (fsm_output[7]));
  assign mux_725_cse = MUX_s_1_2_2(and_532_nl, nor_798_nl, fsm_output[4]);
  assign nand_385_cse = ~((COMP_LOOP_acc_14_psp_sva[2:0]==3'b111) & (fsm_output[7]));
  assign nand_472_nl = ~((COMP_LOOP_acc_14_psp_sva[3:0]==4'b0111) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[7:6]==2'b10));
  assign or_1009_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0111) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_tmp_745 = MUX_s_1_2_2(nand_472_nl, or_1009_nl, fsm_output[4]);
  assign nand_364_cse = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[4]) & (fsm_output[7]));
  assign nand_365_cse = ~((COMP_LOOP_acc_13_psp_sva[2]) & (fsm_output[7]));
  assign or_1112_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b1000) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_1110_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1000) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_tmp_807 = MUX_s_1_2_2(or_1112_nl, or_1110_nl, fsm_output[4]);
  assign nand_357_cse = ~((COMP_LOOP_acc_10_cse_10_1_sva[4]) & (COMP_LOOP_acc_10_cse_10_1_sva[0])
      & (fsm_output[7]));
  assign nand_353_cse = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4]) & (COMP_LOOP_acc_10_cse_10_1_5_sva[1])
      & (fsm_output[7]));
  assign or_1216_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b1001) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_1214_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1001) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_tmp_869 = MUX_s_1_2_2(or_1216_nl, or_1214_nl, fsm_output[4]);
  assign or_1320_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b1010) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_1318_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1010) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_tmp_931 = MUX_s_1_2_2(or_1320_nl, or_1318_nl, fsm_output[4]);
  assign nand_469_nl = ~((COMP_LOOP_acc_14_psp_sva[3:0]==4'b1011) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[7:6]==2'b10));
  assign or_1422_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1011) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_tmp_993 = MUX_s_1_2_2(nand_469_nl, or_1422_nl, fsm_output[4]);
  assign nand_302_cse = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[4:3]==2'b11) & (fsm_output[7]));
  assign nand_303_cse = ~((COMP_LOOP_acc_13_psp_sva[2:1]==2'b11) & (fsm_output[7]));
  assign or_1527_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b1100) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_1525_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1100) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_tmp_1055 = MUX_s_1_2_2(or_1527_nl, or_1525_nl, fsm_output[4]);
  assign nand_294_cse = ~((COMP_LOOP_acc_10_cse_10_1_sva[3]) & (COMP_LOOP_acc_10_cse_10_1_sva[4])
      & (COMP_LOOP_acc_10_cse_10_1_sva[0]) & (fsm_output[7]));
  assign nand_297_cse = ~((COMP_LOOP_acc_1_cse_6_sva[4]) & (COMP_LOOP_acc_1_cse_6_sva[3])
      & (COMP_LOOP_acc_1_cse_6_sva[0]) & (fsm_output[7]));
  assign nand_289_cse = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3]) & (COMP_LOOP_acc_10_cse_10_1_5_sva[4])
      & (COMP_LOOP_acc_10_cse_10_1_5_sva[1]) & (fsm_output[7]));
  assign nand_466_nl = ~((COMP_LOOP_acc_14_psp_sva[3:0]==4'b1101) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[7:6]==2'b10));
  assign or_1627_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1101) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_tmp_1117 = MUX_s_1_2_2(nand_466_nl, or_1627_nl, fsm_output[4]);
  assign nand_266_cse = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[4:2]==3'b111) & (fsm_output[7]));
  assign nand_268_nl = ~((COMP_LOOP_acc_13_psp_sva[2:0]==3'b111) & (fsm_output[7]));
  assign nand_269_nl = ~((COMP_LOOP_acc_psp_sva[0]) & (VEC_LOOP_j_10_0_sva_9_0[2])
      & (COMP_LOOP_acc_psp_sva[1]) & (~ (fsm_output[7])));
  assign mux_1190_cse = MUX_s_1_2_2(nand_268_nl, nand_269_nl, fsm_output[4]);
  assign nand_463_nl = ~((COMP_LOOP_acc_14_psp_sva[3:0]==4'b1110) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[7:6]==2'b10));
  assign or_1727_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1110) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_tmp_1179 = MUX_s_1_2_2(nand_463_nl, or_1727_nl, fsm_output[4]);
  assign and_353_nl = (COMP_LOOP_acc_13_psp_sva[2:0]==3'b111) & (fsm_output[7]);
  assign and_354_nl = (COMP_LOOP_acc_psp_sva[0]) & (VEC_LOOP_j_10_0_sva_9_0[2]) &
      (COMP_LOOP_acc_psp_sva[1]) & (~ (fsm_output[7]));
  assign mux_1221_cse = MUX_s_1_2_2(and_353_nl, and_354_nl, fsm_output[4]);
  assign nand_459_nl = ~((COMP_LOOP_acc_14_psp_sva[3:0]==4'b1111) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[7:6]==2'b10));
  assign nand_236_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]==4'b1111) & COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[7:6]==2'b00));
  assign mux_tmp_1241 = MUX_s_1_2_2(nand_459_nl, nand_236_nl, fsm_output[4]);
  assign and_dcpl_171 = and_dcpl_33 & and_dcpl_79;
  assign and_dcpl_172 = and_dcpl_85 & and_dcpl_79;
  assign and_dcpl_173 = and_dcpl_45 & and_dcpl_79;
  assign and_dcpl_174 = and_dcpl_48 & and_dcpl_79;
  assign and_dcpl_175 = and_dcpl_69 & and_dcpl_28;
  assign and_dcpl_176 = and_dcpl_33 & and_dcpl_175;
  assign and_dcpl_177 = and_dcpl_85 & and_dcpl_175;
  assign and_dcpl_178 = ~((fsm_output[5:4]!=2'b00));
  assign and_dcpl_179 = nor_1025_cse & and_dcpl_178;
  assign not_tmp_617 = ~((z_out_7[1:0]==2'b11) & (fsm_output[1]));
  assign not_tmp_618 = ~((z_out_7[1]) & (fsm_output[1:0]==2'b11));
  assign not_tmp_625 = ~((z_out_7[2:0]==3'b111) & (fsm_output[1:0]==2'b11));
  assign not_tmp_632 = ~((z_out_7[3]) & (z_out_7[0]) & (z_out_7[1]) & (fsm_output[1]));
  assign mux_tmp_1423 = MUX_s_1_2_2(or_167_cse, or_tmp_142, fsm_output[3]);
  assign or_tmp_2024 = (fsm_output[7:6]!=2'b10);
  assign mux_tmp_1424 = MUX_s_1_2_2((~ and_464_cse), or_tmp_2024, fsm_output[3]);
  assign or_tmp_2025 = (fsm_output[4]) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[7]);
  assign mux_tmp_1430 = MUX_s_1_2_2(or_tmp_2024, or_167_cse, fsm_output[3]);
  assign and_dcpl_220 = and_dcpl_59 & and_dcpl_28;
  assign and_dcpl_222 = and_dcpl_33 & and_dcpl_104;
  assign and_dcpl_223 = and_dcpl_69 & and_dcpl_35;
  assign and_dcpl_226 = and_dcpl_33 & and_479_cse & and_dcpl_35;
  assign and_dcpl_229 = and_dcpl_89 & and_479_cse & and_dcpl_28;
  assign and_dcpl_232 = and_dcpl_89 & and_dcpl_59 & and_dcpl_35;
  assign and_dcpl_234 = and_dcpl_95 & and_dcpl_220;
  assign and_dcpl_236 = and_dcpl_95 & and_dcpl_223;
  assign and_dcpl_238 = and_dcpl_38 & and_dcpl_175;
  assign mux_240_nl = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[4]);
  assign mux_1470_nl = MUX_s_1_2_2(and_490_cse, mux_240_nl, fsm_output[0]);
  assign nand_tmp_184 = ~((fsm_output[3]) & (~ mux_1470_nl));
  assign or_2109_nl = (fsm_output[0]) | (~ and_490_cse);
  assign mux_tmp_1437 = MUX_s_1_2_2(or_145_cse, or_2109_nl, fsm_output[3]);
  assign and_dcpl_244 = (fsm_output[0]) & (~ (fsm_output[3]));
  assign or_dcpl_84 = or_tmp_142 | (fsm_output[1:0]!=2'b10) | or_212_cse | (fsm_output[2])
      | (fsm_output[5]);
  assign or_tmp_2048 = and_316_cse | (fsm_output[7:6]!=2'b00);
  assign mux_tmp_1452 = MUX_s_1_2_2((~ or_tmp_2048), and_464_cse, or_212_cse);
  assign mux_1486_nl = MUX_s_1_2_2(and_dcpl_82, and_464_cse, or_212_cse);
  assign mux_1488_nl = MUX_s_1_2_2(mux_tmp_1452, mux_1486_nl, fsm_output[2]);
  assign mux_1489_itm = MUX_s_1_2_2(mux_1488_nl, and_464_cse, fsm_output[5]);
  assign and_448_nl = ((fsm_output[0]) | (fsm_output[1]) | (fsm_output[6])) & (fsm_output[7]);
  assign mux_1490_nl = MUX_s_1_2_2(and_464_cse, and_448_nl, fsm_output[3]);
  assign mux_tmp_1456 = MUX_s_1_2_2(mux_1490_nl, (fsm_output[7]), fsm_output[4]);
  assign mux_1606_nl = MUX_s_1_2_2(mux_189_cse, and_464_cse, and_316_cse);
  assign mux_tmp_1459 = MUX_s_1_2_2(mux_1606_nl, and_464_cse, or_220_cse);
  assign and_tmp_11 = (fsm_output[4]) & ((fsm_output[3]) | (fsm_output[0]) | (fsm_output[1]))
      & (fsm_output[6]);
  assign or_tmp_2054 = and_316_cse | (fsm_output[6]);
  assign not_tmp_692 = ~((fsm_output[4:2]!=3'b000) | or_tmp_2054);
  assign or_tmp_2057 = (fsm_output[4:2]!=3'b000) | and_316_cse;
  assign and_dcpl_252 = or_tmp_2057 & nor_1025_cse & (~ (fsm_output[5]));
  assign nor_340_nl = ~((fsm_output[3]) | or_tmp_2054);
  assign and_511_nl = (fsm_output[3]) & (fsm_output[6]);
  assign mux_tmp_1468 = MUX_s_1_2_2(nor_340_nl, and_511_nl, fsm_output[4]);
  assign and_tmp_13 = (fsm_output[4]) & ((fsm_output[3]) | (fsm_output[1])) & (fsm_output[6]);
  assign nand_188_nl = ~((fsm_output[4:2]==3'b111));
  assign mux_1510_nl = MUX_s_1_2_2(or_tmp_2057, nand_188_nl, fsm_output[5]);
  assign and_dcpl_256 = mux_1510_nl & nor_1025_cse;
  assign nor_tmp_324 = (fsm_output[4]) & (fsm_output[3]) & (fsm_output[6]);
  assign mux_1514_nl = MUX_s_1_2_2(mux_tmp_1468, nor_tmp_324, fsm_output[2]);
  assign mux_1515_nl = MUX_s_1_2_2(mux_1514_nl, (fsm_output[6]), fsm_output[5]);
  assign and_dcpl_259 = ~(mux_1515_nl | (fsm_output[7]));
  assign mux_1599_nl = MUX_s_1_2_2(mux_189_cse, and_464_cse, and_316_cse);
  assign mux_1516_nl = MUX_s_1_2_2(mux_1599_nl, and_464_cse, fsm_output[3]);
  assign mux_tmp_1482 = MUX_s_1_2_2(mux_1516_nl, (fsm_output[7]), fsm_output[4]);
  assign and_446_nl = (and_496_cse | (fsm_output[6])) & (fsm_output[7]);
  assign mux_tmp_1487 = MUX_s_1_2_2(and_446_nl, (fsm_output[7]), fsm_output[4]);
  assign mux_1525_nl = MUX_s_1_2_2(nor_tmp_324, and_485_cse, fsm_output[2]);
  assign mux_1526_nl = MUX_s_1_2_2(not_tmp_692, mux_1525_nl, fsm_output[5]);
  assign and_dcpl_260 = ~(mux_1526_nl | (fsm_output[7]));
  assign mux_1530_nl = MUX_s_1_2_2(mux_tmp_1482, nor_tmp_53, fsm_output[2]);
  assign mux_1531_itm = MUX_s_1_2_2(mux_1530_nl, (fsm_output[7]), fsm_output[5]);
  assign and_306_nl = ((fsm_output[4]) | (fsm_output[3]) | (fsm_output[1])) & (fsm_output[7:6]==2'b11);
  assign mux_1535_nl = MUX_s_1_2_2(mux_tmp_1452, and_306_nl, fsm_output[2]);
  assign mux_1536_itm = MUX_s_1_2_2(mux_1535_nl, and_464_cse, fsm_output[5]);
  assign mux_1537_nl = MUX_s_1_2_2(nor_tmp_53, and_491_cse, fsm_output[2]);
  assign mux_1538_itm = MUX_s_1_2_2(mux_tmp_1459, mux_1537_nl, fsm_output[5]);
  assign not_tmp_717 = ~((fsm_output[4:2]!=3'b000) | or_tmp_2048);
  assign mux_1542_nl = MUX_s_1_2_2(mux_tmp_1452, and_33_cse, fsm_output[2]);
  assign mux_1543_itm = MUX_s_1_2_2(mux_1542_nl, and_464_cse, fsm_output[5]);
  assign and_dcpl_262 = nor_1023_cse & (~ (fsm_output[5]));
  assign and_dcpl_264 = (~((~ (fsm_output[1])) | (fsm_output[6]) | (fsm_output[7])))
      & and_dcpl_244;
  assign nor_1128_nl = ~((~ (fsm_output[3])) | (fsm_output[1]));
  assign nor_1129_nl = ~((fsm_output[3]) | (~ (fsm_output[1])));
  assign mux_1551_nl = MUX_s_1_2_2(nor_1128_nl, nor_1129_nl, fsm_output[2]);
  assign and_dcpl_278 = mux_1551_nl & (~ (fsm_output[7])) & (~ (fsm_output[6])) &
      (fsm_output[0]) & and_dcpl_178;
  assign or_tmp_2075 = (fsm_output[3]) | (fsm_output[6]) | (fsm_output[7]);
  assign or_dcpl_109 = or_tmp_142 | (~ and_316_cse) | or_212_cse | (~ (fsm_output[2]))
      | (fsm_output[5]);
  assign STAGE_LOOP_i_3_0_sva_mx0c1 = and_dcpl_38 & and_dcpl_36;
  assign VEC_LOOP_j_10_0_sva_9_0_mx0c0 = and_dcpl_85 & and_dcpl_30;
  assign COMP_LOOP_tmp_mux1h_itm_mx0c0 = and_dcpl_264 & and_dcpl_262 & (COMP_LOOP_1_tmp_mul_idiv_sva_1_0==2'b00);
  assign COMP_LOOP_tmp_mux1h_itm_mx0c1 = and_dcpl_264 & and_dcpl_262 & (COMP_LOOP_1_tmp_mul_idiv_sva_1_0==2'b01);
  assign COMP_LOOP_tmp_mux1h_itm_mx0c2 = and_dcpl_264 & and_dcpl_262 & (COMP_LOOP_1_tmp_mul_idiv_sva_1_0==2'b10);
  assign COMP_LOOP_tmp_mux1h_itm_mx0c3 = and_dcpl_264 & and_dcpl_262 & (COMP_LOOP_1_tmp_mul_idiv_sva_1_0==2'b11);
  assign mux_1553_nl = MUX_s_1_2_2(mux_tmp_1430, or_tmp_2075, fsm_output[4]);
  assign nand_185_nl = ~((fsm_output[4]) & (~ mux_tmp_1424));
  assign mux_1554_nl = MUX_s_1_2_2(mux_1553_nl, nand_185_nl, fsm_output[2]);
  assign nand_473_nl = ~((fsm_output[4]) & (fsm_output[3]) & (~ (fsm_output[6]))
      & (fsm_output[7]));
  assign or_2171_nl = (fsm_output[4]) | mux_tmp_1423;
  assign mux_1552_nl = MUX_s_1_2_2(nand_473_nl, or_2171_nl, fsm_output[2]);
  assign mux_1555_nl = MUX_s_1_2_2(mux_1554_nl, mux_1552_nl, fsm_output[5]);
  assign COMP_LOOP_1_acc_8_itm_mx0c4 = (~ mux_1555_nl) & and_dcpl_40;
  assign or_229_nl = or_32_cse | or_212_cse;
  assign mux_1574_nl = MUX_s_1_2_2(or_212_cse, or_229_nl, fsm_output[2]);
  assign mux_1573_nl = MUX_s_1_2_2((fsm_output[4]), or_212_cse, fsm_output[2]);
  assign mux_1575_nl = MUX_s_1_2_2(mux_1574_nl, (~ mux_1573_nl), fsm_output[5]);
  assign and_294_tmp = mux_1575_nl & nor_1025_cse;
  assign mux_1577_nl = MUX_s_1_2_2((~ (fsm_output[6])), (fsm_output[6]), or_212_cse);
  assign nor_1059_nl = ~((fsm_output[1]) | (fsm_output[6]));
  assign mux_1576_nl = MUX_s_1_2_2(nor_1059_nl, (fsm_output[6]), or_212_cse);
  assign mux_1578_nl = MUX_s_1_2_2(mux_1577_nl, mux_1576_nl, fsm_output[2]);
  assign mux_1579_nl = MUX_s_1_2_2(mux_1578_nl, (fsm_output[6]), fsm_output[5]);
  assign nor_1119_tmp = ~(mux_1579_nl | (fsm_output[7]));
  assign nor_1062_nl = ~((fsm_output[4]) | (fsm_output[3]) | (fsm_output[6]));
  assign nor_1063_nl = ~((fsm_output[4:3]!=2'b00) | or_tmp_2054);
  assign mux_1580_nl = MUX_s_1_2_2(nor_1062_nl, nor_1063_nl, fsm_output[2]);
  assign and_520_nl = or_220_cse & (fsm_output[6]);
  assign mux_1581_nl = MUX_s_1_2_2(mux_1580_nl, and_520_nl, fsm_output[5]);
  assign nor_tmp = ~(mux_1581_nl | (fsm_output[7]));
  assign nor_1117_tmp = ~((~((fsm_output[6:3]!=4'b0000))) | (fsm_output[7]));
  assign and_54_nl = ((fsm_output[6]) ^ (fsm_output[3])) & ((fsm_output[7]) ^ (fsm_output[4]))
      & and_dcpl_40 & ((fsm_output[2]) ^ (fsm_output[5]));
  assign vec_rsc_0_0_i_d_d_pff = MUX_v_64_2_2(COMP_LOOP_1_modulo_dev_cmp_return_rsc_z,
      COMP_LOOP_1_acc_8_itm, and_54_nl);
  assign and_64_nl = and_dcpl_45 & and_dcpl_52;
  assign and_68_nl = and_dcpl_45 & and_dcpl_56;
  assign and_74_nl = and_dcpl_62 & and_dcpl_60;
  assign and_78_nl = and_dcpl_62 & and_dcpl_66;
  assign and_84_nl = and_dcpl_72 & and_dcpl_70;
  assign and_88_nl = and_dcpl_72 & and_dcpl_76;
  assign and_92_nl = and_464_cse & and_dcpl_44 & and_dcpl_79;
  assign vec_rsc_0_0_i_radr_d_pff = MUX1HOT_v_5_16_2((COMP_LOOP_1_acc_10_itm_10_1_1[9:5]),
      (COMP_LOOP_acc_psp_sva[6:2]), (COMP_LOOP_acc_1_cse_2_sva[9:5]), (COMP_LOOP_acc_10_cse_10_1_2_sva[9:5]),
      (COMP_LOOP_acc_11_psp_sva[8:4]), (COMP_LOOP_acc_10_cse_10_1_3_sva[9:5]), (COMP_LOOP_acc_1_cse_4_sva[9:5]),
      (COMP_LOOP_acc_10_cse_10_1_4_sva[9:5]), (COMP_LOOP_acc_13_psp_sva[7:3]), (COMP_LOOP_acc_10_cse_10_1_5_sva[9:5]),
      (COMP_LOOP_acc_1_cse_6_sva[9:5]), (COMP_LOOP_acc_10_cse_10_1_6_sva[9:5]), (COMP_LOOP_acc_14_psp_sva[8:4]),
      (COMP_LOOP_acc_10_cse_10_1_7_sva[9:5]), (COMP_LOOP_acc_1_cse_sva[9:5]), (COMP_LOOP_acc_10_cse_10_1_sva[9:5]),
      {and_dcpl_46 , and_dcpl_49 , and_64_nl , and_dcpl_54 , and_68_nl , and_dcpl_58
      , and_74_nl , and_dcpl_65 , and_78_nl , and_dcpl_68 , and_84_nl , and_dcpl_75
      , and_88_nl , and_dcpl_78 , and_92_nl , and_dcpl_83});
  assign and_95_nl = and_dcpl_33 & and_dcpl_52;
  assign and_97_nl = and_dcpl_85 & and_dcpl_52;
  assign and_98_nl = and_dcpl_33 & and_dcpl_56;
  assign and_99_nl = and_dcpl_85 & and_dcpl_56;
  assign and_101_nl = and_dcpl_89 & and_dcpl_60;
  assign and_103_nl = and_dcpl_91 & and_dcpl_60;
  assign and_104_nl = and_dcpl_89 & and_dcpl_66;
  assign and_105_nl = and_dcpl_91 & and_dcpl_66;
  assign and_107_nl = and_dcpl_95 & and_dcpl_70;
  assign and_109_nl = and_dcpl_97 & and_dcpl_70;
  assign and_110_nl = and_dcpl_95 & and_dcpl_76;
  assign and_111_nl = and_dcpl_97 & and_dcpl_76;
  assign and_112_nl = and_dcpl_38 & and_dcpl_79;
  assign and_114_nl = and_dcpl_102 & and_dcpl_79;
  assign and_116_nl = and_dcpl_38 & and_dcpl_104;
  assign and_117_nl = and_dcpl_102 & and_dcpl_104;
  assign vec_rsc_0_0_i_wadr_d_pff = MUX1HOT_v_5_16_2((COMP_LOOP_acc_10_cse_10_1_1_sva[9:5]),
      (COMP_LOOP_acc_psp_sva[6:2]), (COMP_LOOP_acc_10_cse_10_1_2_sva[9:5]), (COMP_LOOP_acc_1_cse_2_sva[9:5]),
      (COMP_LOOP_acc_10_cse_10_1_3_sva[9:5]), (COMP_LOOP_acc_11_psp_sva[8:4]), (COMP_LOOP_acc_10_cse_10_1_4_sva[9:5]),
      (COMP_LOOP_acc_1_cse_4_sva[9:5]), (COMP_LOOP_acc_10_cse_10_1_5_sva[9:5]), (COMP_LOOP_acc_13_psp_sva[7:3]),
      (COMP_LOOP_acc_10_cse_10_1_6_sva[9:5]), (COMP_LOOP_acc_1_cse_6_sva[9:5]), (COMP_LOOP_acc_10_cse_10_1_7_sva[9:5]),
      (COMP_LOOP_acc_14_psp_sva[8:4]), (COMP_LOOP_acc_10_cse_10_1_sva[9:5]), (COMP_LOOP_acc_1_cse_sva[9:5]),
      {and_95_nl , and_97_nl , and_98_nl , and_99_nl , and_101_nl , and_103_nl ,
      and_104_nl , and_105_nl , and_107_nl , and_109_nl , and_110_nl , and_111_nl
      , and_112_nl , and_114_nl , and_116_nl , and_117_nl});
  assign nor_1010_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b00000) | (~ (fsm_output[7])));
  assign nor_1011_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b00000) | (fsm_output[7]));
  assign mux_333_nl = MUX_s_1_2_2(nor_1010_nl, nor_1011_nl, fsm_output[4]);
  assign nor_1012_nl = ~((COMP_LOOP_acc_1_cse_sva[4:0]!=5'b00000) | (~ (fsm_output[7])));
  assign nor_1013_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b00000) | (fsm_output[7]));
  assign mux_332_nl = MUX_s_1_2_2(nor_1012_nl, nor_1013_nl, fsm_output[4]);
  assign mux_334_nl = MUX_s_1_2_2(mux_333_nl, mux_332_nl, fsm_output[0]);
  assign and_443_nl = (fsm_output[6]) & mux_334_nl;
  assign or_257_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00000) | (~ (fsm_output[7]));
  assign or_255_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b00000) | (fsm_output[7]);
  assign mux_330_nl = MUX_s_1_2_2(or_257_nl, or_255_nl, fsm_output[4]);
  assign or_254_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00000) | (~ (fsm_output[7]));
  assign or_252_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b00000) | (fsm_output[7]);
  assign mux_329_nl = MUX_s_1_2_2(or_254_nl, or_252_nl, fsm_output[4]);
  assign mux_331_nl = MUX_s_1_2_2(mux_330_nl, mux_329_nl, fsm_output[0]);
  assign nor_1014_nl = ~((fsm_output[6]) | mux_331_nl);
  assign mux_335_nl = MUX_s_1_2_2(and_443_nl, nor_1014_nl, fsm_output[3]);
  assign nand_506_nl = ~((fsm_output[5]) & mux_335_nl);
  assign nor_1016_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b00000) | (~ (fsm_output[7])));
  assign nor_1017_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b00000) | (fsm_output[7]));
  assign mux_326_nl = MUX_s_1_2_2(nor_1016_nl, nor_1017_nl, fsm_output[4]);
  assign or_246_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b0000) | (~ (fsm_output[7]));
  assign or_244_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0000) | (fsm_output[7]);
  assign mux_325_nl = MUX_s_1_2_2(or_246_nl, or_244_nl, fsm_output[4]);
  assign nor_1018_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_325_nl);
  assign mux_327_nl = MUX_s_1_2_2(mux_326_nl, nor_1018_nl, fsm_output[0]);
  assign nand_8_nl = ~((fsm_output[6]) & mux_327_nl);
  assign or_242_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b00000) | (~ (fsm_output[7]));
  assign or_240_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b00000) | (fsm_output[7]);
  assign mux_323_nl = MUX_s_1_2_2(or_242_nl, or_240_nl, fsm_output[4]);
  assign or_239_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | mux_322_cse;
  assign mux_324_nl = MUX_s_1_2_2(mux_323_nl, or_239_nl, fsm_output[0]);
  assign or_243_nl = (fsm_output[6]) | mux_324_nl;
  assign mux_328_nl = MUX_s_1_2_2(nand_8_nl, or_243_nl, fsm_output[3]);
  assign or_2280_nl = (fsm_output[5]) | mux_328_nl;
  assign mux_336_nl = MUX_s_1_2_2(nand_506_nl, or_2280_nl, fsm_output[2]);
  assign vec_rsc_0_0_i_we_d_pff = ~(mux_336_nl | (fsm_output[1]));
  assign nor_1003_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b00000) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_1004_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_350_nl = MUX_s_1_2_2(nor_1003_nl, nor_1004_nl, fsm_output[0]);
  assign nor_1005_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_348_cse);
  assign nor_1006_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b00000) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_1007_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b00000) | (fsm_output[7:6]!=2'b10));
  assign nor_1008_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b00000) | (fsm_output[7:6]!=2'b00));
  assign mux_344_nl = MUX_s_1_2_2(nor_1007_nl, nor_1008_nl, fsm_output[4]);
  assign mux_345_nl = MUX_s_1_2_2(nor_1006_nl, mux_344_nl, fsm_output[3]);
  assign mux_349_nl = MUX_s_1_2_2(nor_1005_nl, mux_345_nl, fsm_output[0]);
  assign mux_351_nl = MUX_s_1_2_2(mux_350_nl, mux_349_nl, fsm_output[5]);
  assign or_276_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b00000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_274_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b00000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_341_nl = MUX_s_1_2_2(or_276_nl, or_274_nl, fsm_output[4]);
  assign or_273_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00000) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_271_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b00000) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_340_nl = MUX_s_1_2_2(or_273_nl, or_271_nl, fsm_output[4]);
  assign mux_342_nl = MUX_s_1_2_2(mux_341_nl, mux_340_nl, fsm_output[3]);
  assign or_270_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b00000) | nand_443_cse;
  assign or_268_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b00000) | (fsm_output[7:6]!=2'b01);
  assign mux_338_nl = MUX_s_1_2_2(or_270_nl, or_268_nl, fsm_output[4]);
  assign or_267_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00000) | (fsm_output[7:6]!=2'b10);
  assign or_265_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b00000) | (fsm_output[7:6]!=2'b00);
  assign mux_337_nl = MUX_s_1_2_2(or_267_nl, or_265_nl, fsm_output[4]);
  assign mux_339_nl = MUX_s_1_2_2(mux_338_nl, mux_337_nl, fsm_output[3]);
  assign mux_343_nl = MUX_s_1_2_2(mux_342_nl, mux_339_nl, fsm_output[0]);
  assign nor_1009_nl = ~((fsm_output[5]) | mux_343_nl);
  assign mux_352_nl = MUX_s_1_2_2(mux_351_nl, nor_1009_nl, fsm_output[2]);
  assign vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d = mux_352_nl & (fsm_output[1]);
  assign nor_991_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:1]!=4'b0000) | nand_445_cse);
  assign nor_992_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b00001) | (fsm_output[7]));
  assign mux_364_nl = MUX_s_1_2_2(nor_991_nl, nor_992_nl, fsm_output[4]);
  assign nor_993_nl = ~((COMP_LOOP_acc_1_cse_sva[4:1]!=4'b0000) | nand_446_cse);
  assign nor_994_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b00001) | (fsm_output[7]));
  assign mux_363_nl = MUX_s_1_2_2(nor_993_nl, nor_994_nl, fsm_output[4]);
  assign mux_365_nl = MUX_s_1_2_2(mux_364_nl, mux_363_nl, fsm_output[0]);
  assign and_440_nl = (fsm_output[6]) & mux_365_nl;
  assign or_308_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00001) | (~ (fsm_output[7]));
  assign or_306_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b00001) | (fsm_output[7]);
  assign mux_361_nl = MUX_s_1_2_2(or_308_nl, or_306_nl, fsm_output[4]);
  assign or_305_nl = (COMP_LOOP_acc_1_cse_6_sva[4:1]!=4'b0000) | nand_447_cse;
  assign or_303_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b00001) | (fsm_output[7]);
  assign mux_360_nl = MUX_s_1_2_2(or_305_nl, or_303_nl, fsm_output[4]);
  assign mux_362_nl = MUX_s_1_2_2(mux_361_nl, mux_360_nl, fsm_output[0]);
  assign nor_995_nl = ~((fsm_output[6]) | mux_362_nl);
  assign mux_366_nl = MUX_s_1_2_2(and_440_nl, nor_995_nl, fsm_output[3]);
  assign nand_505_nl = ~((fsm_output[5]) & mux_366_nl);
  assign nor_997_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:1]!=4'b0000) | nand_448_cse);
  assign nor_998_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b00001) | (fsm_output[7]));
  assign mux_357_nl = MUX_s_1_2_2(nor_997_nl, nor_998_nl, fsm_output[4]);
  assign nor_999_nl = ~((COMP_LOOP_acc_14_psp_sva[3:0]!=4'b0000) | (~ (fsm_output[7])));
  assign nor_1000_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0000) | (fsm_output[7]));
  assign mux_356_nl = MUX_s_1_2_2(nor_999_nl, nor_1000_nl, fsm_output[4]);
  assign and_441_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_356_nl;
  assign mux_358_nl = MUX_s_1_2_2(mux_357_nl, and_441_nl, fsm_output[0]);
  assign nand_14_nl = ~((fsm_output[6]) & mux_358_nl);
  assign or_294_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b00001) | (~ (fsm_output[7]));
  assign or_292_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b00001) | (fsm_output[7]);
  assign mux_354_nl = MUX_s_1_2_2(or_294_nl, or_292_nl, fsm_output[4]);
  assign nand_12_nl = ~(nor_98_cse & mux_353_cse);
  assign mux_355_nl = MUX_s_1_2_2(mux_354_nl, nand_12_nl, fsm_output[0]);
  assign or_295_nl = (fsm_output[6]) | mux_355_nl;
  assign mux_359_nl = MUX_s_1_2_2(nand_14_nl, or_295_nl, fsm_output[3]);
  assign or_2279_nl = (fsm_output[5]) | mux_359_nl;
  assign mux_367_nl = MUX_s_1_2_2(nand_505_nl, or_2279_nl, fsm_output[2]);
  assign vec_rsc_0_1_i_we_d_pff = ~(mux_367_nl | (fsm_output[1]));
  assign nor_985_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b00001) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_986_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_381_nl = MUX_s_1_2_2(nor_985_nl, nor_986_nl, fsm_output[0]);
  assign and_438_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (~ mux_348_cse);
  assign nor_987_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b00001) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_988_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b00001) | (fsm_output[7:6]!=2'b10));
  assign nor_989_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b00001) | (fsm_output[7:6]!=2'b00));
  assign mux_375_nl = MUX_s_1_2_2(nor_988_nl, nor_989_nl, fsm_output[4]);
  assign mux_376_nl = MUX_s_1_2_2(nor_987_nl, mux_375_nl, fsm_output[3]);
  assign mux_380_nl = MUX_s_1_2_2(and_438_nl, mux_376_nl, fsm_output[0]);
  assign mux_382_nl = MUX_s_1_2_2(mux_381_nl, mux_380_nl, fsm_output[5]);
  assign or_327_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b00001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_325_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b00001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_372_nl = MUX_s_1_2_2(or_327_nl, or_325_nl, fsm_output[4]);
  assign or_324_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00001) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_322_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b00001) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_371_nl = MUX_s_1_2_2(or_324_nl, or_322_nl, fsm_output[4]);
  assign mux_373_nl = MUX_s_1_2_2(mux_372_nl, mux_371_nl, fsm_output[3]);
  assign or_321_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:1]!=4'b0000) | nand_444_cse;
  assign or_319_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b00001) | (fsm_output[7:6]!=2'b01);
  assign mux_369_nl = MUX_s_1_2_2(or_321_nl, or_319_nl, fsm_output[4]);
  assign or_318_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00001) | (fsm_output[7:6]!=2'b10);
  assign or_316_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b00001) | (fsm_output[7:6]!=2'b00);
  assign mux_368_nl = MUX_s_1_2_2(or_318_nl, or_316_nl, fsm_output[4]);
  assign mux_370_nl = MUX_s_1_2_2(mux_369_nl, mux_368_nl, fsm_output[3]);
  assign mux_374_nl = MUX_s_1_2_2(mux_373_nl, mux_370_nl, fsm_output[0]);
  assign nor_990_nl = ~((fsm_output[5]) | mux_374_nl);
  assign mux_383_nl = MUX_s_1_2_2(mux_382_nl, nor_990_nl, fsm_output[2]);
  assign vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d = mux_383_nl & (fsm_output[1]);
  assign nor_976_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b00010) | (~ (fsm_output[7])));
  assign nor_977_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b00010) | (fsm_output[7]));
  assign mux_395_nl = MUX_s_1_2_2(nor_976_nl, nor_977_nl, fsm_output[4]);
  assign nor_978_nl = ~((COMP_LOOP_acc_1_cse_sva[4:0]!=5'b00010) | (~ (fsm_output[7])));
  assign nor_979_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b00010) | (fsm_output[7]));
  assign mux_394_nl = MUX_s_1_2_2(nor_978_nl, nor_979_nl, fsm_output[4]);
  assign mux_396_nl = MUX_s_1_2_2(mux_395_nl, mux_394_nl, fsm_output[0]);
  assign and_437_nl = (fsm_output[6]) & mux_396_nl;
  assign or_361_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00010) | (~ (fsm_output[7]));
  assign or_359_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b00010) | (fsm_output[7]);
  assign mux_392_nl = MUX_s_1_2_2(or_361_nl, or_359_nl, fsm_output[4]);
  assign or_358_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00010) | (~ (fsm_output[7]));
  assign or_356_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b00010) | (fsm_output[7]);
  assign mux_391_nl = MUX_s_1_2_2(or_358_nl, or_356_nl, fsm_output[4]);
  assign mux_393_nl = MUX_s_1_2_2(mux_392_nl, mux_391_nl, fsm_output[0]);
  assign nor_980_nl = ~((fsm_output[6]) | mux_393_nl);
  assign mux_397_nl = MUX_s_1_2_2(and_437_nl, nor_980_nl, fsm_output[3]);
  assign nand_504_nl = ~((fsm_output[5]) & mux_397_nl);
  assign nor_982_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b00010) | (~ (fsm_output[7])));
  assign nor_983_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b00010) | (fsm_output[7]));
  assign mux_388_nl = MUX_s_1_2_2(nor_982_nl, nor_983_nl, fsm_output[4]);
  assign or_350_nl = (COMP_LOOP_acc_14_psp_sva[3:1]!=3'b000) | nand_441_cse;
  assign or_348_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0001) | (fsm_output[7]);
  assign mux_387_nl = MUX_s_1_2_2(or_350_nl, or_348_nl, fsm_output[4]);
  assign nor_984_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_387_nl);
  assign mux_389_nl = MUX_s_1_2_2(mux_388_nl, nor_984_nl, fsm_output[0]);
  assign nand_19_nl = ~((fsm_output[6]) & mux_389_nl);
  assign or_346_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[3]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[4])
      | nand_442_cse;
  assign or_344_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b00010) | (fsm_output[7]);
  assign mux_385_nl = MUX_s_1_2_2(or_346_nl, or_344_nl, fsm_output[4]);
  assign or_343_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | mux_322_cse;
  assign mux_386_nl = MUX_s_1_2_2(mux_385_nl, or_343_nl, fsm_output[0]);
  assign or_347_nl = (fsm_output[6]) | mux_386_nl;
  assign mux_390_nl = MUX_s_1_2_2(nand_19_nl, or_347_nl, fsm_output[3]);
  assign or_2278_nl = (fsm_output[5]) | mux_390_nl;
  assign mux_398_nl = MUX_s_1_2_2(nand_504_nl, or_2278_nl, fsm_output[2]);
  assign vec_rsc_0_2_i_we_d_pff = ~(mux_398_nl | (fsm_output[1]));
  assign nor_969_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b00010) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_970_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_412_nl = MUX_s_1_2_2(nor_969_nl, nor_970_nl, fsm_output[0]);
  assign nor_971_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_410_cse);
  assign nor_972_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b00010) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_973_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b00010) | (fsm_output[7:6]!=2'b10));
  assign nor_974_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b00010) | (fsm_output[7:6]!=2'b00));
  assign mux_406_nl = MUX_s_1_2_2(nor_973_nl, nor_974_nl, fsm_output[4]);
  assign mux_407_nl = MUX_s_1_2_2(nor_972_nl, mux_406_nl, fsm_output[3]);
  assign mux_411_nl = MUX_s_1_2_2(nor_971_nl, mux_407_nl, fsm_output[0]);
  assign mux_413_nl = MUX_s_1_2_2(mux_412_nl, mux_411_nl, fsm_output[5]);
  assign or_380_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b00010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_378_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b00010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_403_nl = MUX_s_1_2_2(or_380_nl, or_378_nl, fsm_output[4]);
  assign or_377_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00010) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_375_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b00010) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_402_nl = MUX_s_1_2_2(or_377_nl, or_375_nl, fsm_output[4]);
  assign mux_404_nl = MUX_s_1_2_2(mux_403_nl, mux_402_nl, fsm_output[3]);
  assign or_374_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b00010) | nand_443_cse;
  assign or_372_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b00010) | (fsm_output[7:6]!=2'b01);
  assign mux_400_nl = MUX_s_1_2_2(or_374_nl, or_372_nl, fsm_output[4]);
  assign or_371_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00010) | (fsm_output[7:6]!=2'b10);
  assign or_369_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b00010) | (fsm_output[7:6]!=2'b00);
  assign mux_399_nl = MUX_s_1_2_2(or_371_nl, or_369_nl, fsm_output[4]);
  assign mux_401_nl = MUX_s_1_2_2(mux_400_nl, mux_399_nl, fsm_output[3]);
  assign mux_405_nl = MUX_s_1_2_2(mux_404_nl, mux_401_nl, fsm_output[0]);
  assign nor_975_nl = ~((fsm_output[5]) | mux_405_nl);
  assign mux_414_nl = MUX_s_1_2_2(mux_413_nl, nor_975_nl, fsm_output[2]);
  assign vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d = mux_414_nl & (fsm_output[1]);
  assign nor_957_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:1]!=4'b0001) | nand_445_cse);
  assign nor_958_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b00011) | (fsm_output[7]));
  assign mux_426_nl = MUX_s_1_2_2(nor_957_nl, nor_958_nl, fsm_output[4]);
  assign nor_959_nl = ~((COMP_LOOP_acc_1_cse_sva[4:2]!=3'b000) | nand_435_cse);
  assign nor_960_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b00011) | (fsm_output[7]));
  assign mux_425_nl = MUX_s_1_2_2(nor_959_nl, nor_960_nl, fsm_output[4]);
  assign mux_427_nl = MUX_s_1_2_2(mux_426_nl, mux_425_nl, fsm_output[0]);
  assign and_434_nl = (fsm_output[6]) & mux_427_nl;
  assign or_412_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00011) | (~ (fsm_output[7]));
  assign or_410_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b00011) | (fsm_output[7]);
  assign mux_423_nl = MUX_s_1_2_2(or_412_nl, or_410_nl, fsm_output[4]);
  assign or_409_nl = (COMP_LOOP_acc_1_cse_6_sva[4:1]!=4'b0001) | nand_447_cse;
  assign or_407_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b00011) | (fsm_output[7]);
  assign mux_422_nl = MUX_s_1_2_2(or_409_nl, or_407_nl, fsm_output[4]);
  assign mux_424_nl = MUX_s_1_2_2(mux_423_nl, mux_422_nl, fsm_output[0]);
  assign nor_961_nl = ~((fsm_output[6]) | mux_424_nl);
  assign mux_428_nl = MUX_s_1_2_2(and_434_nl, nor_961_nl, fsm_output[3]);
  assign nand_503_nl = ~((fsm_output[5]) & mux_428_nl);
  assign nor_963_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:2]!=3'b000) | nand_437_cse);
  assign nor_964_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b00011) | (fsm_output[7]));
  assign mux_419_nl = MUX_s_1_2_2(nor_963_nl, nor_964_nl, fsm_output[4]);
  assign nor_965_nl = ~((COMP_LOOP_acc_14_psp_sva[3:1]!=3'b000) | nand_441_cse);
  assign nor_966_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0001) | (fsm_output[7]));
  assign mux_418_nl = MUX_s_1_2_2(nor_965_nl, nor_966_nl, fsm_output[4]);
  assign and_435_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_418_nl;
  assign mux_420_nl = MUX_s_1_2_2(mux_419_nl, and_435_nl, fsm_output[0]);
  assign nand_25_nl = ~((fsm_output[6]) & mux_420_nl);
  assign or_398_nl = (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[0])) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[3]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[4])
      | nand_442_cse;
  assign or_396_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b00011) | (fsm_output[7]);
  assign mux_416_nl = MUX_s_1_2_2(or_398_nl, or_396_nl, fsm_output[4]);
  assign nand_23_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & mux_353_cse);
  assign mux_417_nl = MUX_s_1_2_2(mux_416_nl, nand_23_nl, fsm_output[0]);
  assign or_399_nl = (fsm_output[6]) | mux_417_nl;
  assign mux_421_nl = MUX_s_1_2_2(nand_25_nl, or_399_nl, fsm_output[3]);
  assign or_2277_nl = (fsm_output[5]) | mux_421_nl;
  assign mux_429_nl = MUX_s_1_2_2(nand_503_nl, or_2277_nl, fsm_output[2]);
  assign vec_rsc_0_3_i_we_d_pff = ~(mux_429_nl | (fsm_output[1]));
  assign nor_951_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b00011) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_952_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_443_nl = MUX_s_1_2_2(nor_951_nl, nor_952_nl, fsm_output[0]);
  assign and_432_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (~ mux_410_cse);
  assign nor_953_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b00011) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_954_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b00011) | (fsm_output[7:6]!=2'b10));
  assign nor_955_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b00011) | (fsm_output[7:6]!=2'b00));
  assign mux_437_nl = MUX_s_1_2_2(nor_954_nl, nor_955_nl, fsm_output[4]);
  assign mux_438_nl = MUX_s_1_2_2(nor_953_nl, mux_437_nl, fsm_output[3]);
  assign mux_442_nl = MUX_s_1_2_2(and_432_nl, mux_438_nl, fsm_output[0]);
  assign mux_444_nl = MUX_s_1_2_2(mux_443_nl, mux_442_nl, fsm_output[5]);
  assign or_431_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b00011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_429_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b00011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_434_nl = MUX_s_1_2_2(or_431_nl, or_429_nl, fsm_output[4]);
  assign or_428_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00011) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_426_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b00011) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_433_nl = MUX_s_1_2_2(or_428_nl, or_426_nl, fsm_output[4]);
  assign mux_435_nl = MUX_s_1_2_2(mux_434_nl, mux_433_nl, fsm_output[3]);
  assign or_425_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:1]!=4'b0001) | nand_444_cse;
  assign or_423_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b00011) | (fsm_output[7:6]!=2'b01);
  assign mux_431_nl = MUX_s_1_2_2(or_425_nl, or_423_nl, fsm_output[4]);
  assign or_422_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00011) | (fsm_output[7:6]!=2'b10);
  assign or_420_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b00011) | (fsm_output[7:6]!=2'b00);
  assign mux_430_nl = MUX_s_1_2_2(or_422_nl, or_420_nl, fsm_output[4]);
  assign mux_432_nl = MUX_s_1_2_2(mux_431_nl, mux_430_nl, fsm_output[3]);
  assign mux_436_nl = MUX_s_1_2_2(mux_435_nl, mux_432_nl, fsm_output[0]);
  assign nor_956_nl = ~((fsm_output[5]) | mux_436_nl);
  assign mux_445_nl = MUX_s_1_2_2(mux_444_nl, nor_956_nl, fsm_output[2]);
  assign vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d = mux_445_nl & (fsm_output[1]);
  assign nor_942_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b00100) | (~ (fsm_output[7])));
  assign nor_943_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b00100) | (fsm_output[7]));
  assign mux_457_nl = MUX_s_1_2_2(nor_942_nl, nor_943_nl, fsm_output[4]);
  assign nor_944_nl = ~((COMP_LOOP_acc_1_cse_sva[4:0]!=5'b00100) | (~ (fsm_output[7])));
  assign nor_945_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b00100) | (fsm_output[7]));
  assign mux_456_nl = MUX_s_1_2_2(nor_944_nl, nor_945_nl, fsm_output[4]);
  assign mux_458_nl = MUX_s_1_2_2(mux_457_nl, mux_456_nl, fsm_output[0]);
  assign and_431_nl = (fsm_output[6]) & mux_458_nl;
  assign or_465_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00100) | (~ (fsm_output[7]));
  assign or_463_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b00100) | (fsm_output[7]);
  assign mux_454_nl = MUX_s_1_2_2(or_465_nl, or_463_nl, fsm_output[4]);
  assign or_462_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00100) | (~ (fsm_output[7]));
  assign or_460_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b00100) | (fsm_output[7]);
  assign mux_453_nl = MUX_s_1_2_2(or_462_nl, or_460_nl, fsm_output[4]);
  assign mux_455_nl = MUX_s_1_2_2(mux_454_nl, mux_453_nl, fsm_output[0]);
  assign nor_946_nl = ~((fsm_output[6]) | mux_455_nl);
  assign mux_459_nl = MUX_s_1_2_2(and_431_nl, nor_946_nl, fsm_output[3]);
  assign nand_502_nl = ~((fsm_output[5]) & mux_459_nl);
  assign nor_948_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b00100) | (~ (fsm_output[7])));
  assign nor_949_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b00100) | (fsm_output[7]));
  assign mux_450_nl = MUX_s_1_2_2(nor_948_nl, nor_949_nl, fsm_output[4]);
  assign or_454_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b0010) | (~ (fsm_output[7]));
  assign or_452_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0010) | (fsm_output[7]);
  assign mux_449_nl = MUX_s_1_2_2(or_454_nl, or_452_nl, fsm_output[4]);
  assign nor_950_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_449_nl);
  assign mux_451_nl = MUX_s_1_2_2(mux_450_nl, nor_950_nl, fsm_output[0]);
  assign nand_30_nl = ~((fsm_output[6]) & mux_451_nl);
  assign or_450_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b00100) | (~ (fsm_output[7]));
  assign or_448_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b00100) | (fsm_output[7]);
  assign mux_447_nl = MUX_s_1_2_2(or_450_nl, or_448_nl, fsm_output[4]);
  assign or_447_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | mux_446_cse;
  assign mux_448_nl = MUX_s_1_2_2(mux_447_nl, or_447_nl, fsm_output[0]);
  assign or_451_nl = (fsm_output[6]) | mux_448_nl;
  assign mux_452_nl = MUX_s_1_2_2(nand_30_nl, or_451_nl, fsm_output[3]);
  assign or_2276_nl = (fsm_output[5]) | mux_452_nl;
  assign mux_460_nl = MUX_s_1_2_2(nand_502_nl, or_2276_nl, fsm_output[2]);
  assign vec_rsc_0_4_i_we_d_pff = ~(mux_460_nl | (fsm_output[1]));
  assign nor_935_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b00100) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_936_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_474_nl = MUX_s_1_2_2(nor_935_nl, nor_936_nl, fsm_output[0]);
  assign nor_937_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_472_cse);
  assign nor_938_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b00100) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_939_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b00100) | (fsm_output[7:6]!=2'b10));
  assign nor_940_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b00100) | (fsm_output[7:6]!=2'b00));
  assign mux_468_nl = MUX_s_1_2_2(nor_939_nl, nor_940_nl, fsm_output[4]);
  assign mux_469_nl = MUX_s_1_2_2(nor_938_nl, mux_468_nl, fsm_output[3]);
  assign mux_473_nl = MUX_s_1_2_2(nor_937_nl, mux_469_nl, fsm_output[0]);
  assign mux_475_nl = MUX_s_1_2_2(mux_474_nl, mux_473_nl, fsm_output[5]);
  assign or_484_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b00100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_482_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b00100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_465_nl = MUX_s_1_2_2(or_484_nl, or_482_nl, fsm_output[4]);
  assign or_481_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00100) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_479_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b00100) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_464_nl = MUX_s_1_2_2(or_481_nl, or_479_nl, fsm_output[4]);
  assign mux_466_nl = MUX_s_1_2_2(mux_465_nl, mux_464_nl, fsm_output[3]);
  assign or_478_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b00100) | nand_443_cse;
  assign or_476_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b00100) | (fsm_output[7:6]!=2'b01);
  assign mux_462_nl = MUX_s_1_2_2(or_478_nl, or_476_nl, fsm_output[4]);
  assign or_475_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00100) | (fsm_output[7:6]!=2'b10);
  assign or_473_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b00100) | (fsm_output[7:6]!=2'b00);
  assign mux_461_nl = MUX_s_1_2_2(or_475_nl, or_473_nl, fsm_output[4]);
  assign mux_463_nl = MUX_s_1_2_2(mux_462_nl, mux_461_nl, fsm_output[3]);
  assign mux_467_nl = MUX_s_1_2_2(mux_466_nl, mux_463_nl, fsm_output[0]);
  assign nor_941_nl = ~((fsm_output[5]) | mux_467_nl);
  assign mux_476_nl = MUX_s_1_2_2(mux_475_nl, nor_941_nl, fsm_output[2]);
  assign vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d = mux_476_nl & (fsm_output[1]);
  assign nor_923_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:1]!=4'b0010) | nand_445_cse);
  assign nor_924_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b00101) | (fsm_output[7]));
  assign mux_488_nl = MUX_s_1_2_2(nor_923_nl, nor_924_nl, fsm_output[4]);
  assign nor_925_nl = ~((COMP_LOOP_acc_1_cse_sva[4:1]!=4'b0010) | nand_446_cse);
  assign nor_926_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b00101) | (fsm_output[7]));
  assign mux_487_nl = MUX_s_1_2_2(nor_925_nl, nor_926_nl, fsm_output[4]);
  assign mux_489_nl = MUX_s_1_2_2(mux_488_nl, mux_487_nl, fsm_output[0]);
  assign and_428_nl = (fsm_output[6]) & mux_489_nl;
  assign or_516_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00101) | (~ (fsm_output[7]));
  assign or_514_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b00101) | (fsm_output[7]);
  assign mux_485_nl = MUX_s_1_2_2(or_516_nl, or_514_nl, fsm_output[4]);
  assign or_513_nl = (COMP_LOOP_acc_1_cse_6_sva[4:1]!=4'b0010) | nand_447_cse;
  assign or_511_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b00101) | (fsm_output[7]);
  assign mux_484_nl = MUX_s_1_2_2(or_513_nl, or_511_nl, fsm_output[4]);
  assign mux_486_nl = MUX_s_1_2_2(mux_485_nl, mux_484_nl, fsm_output[0]);
  assign nor_927_nl = ~((fsm_output[6]) | mux_486_nl);
  assign mux_490_nl = MUX_s_1_2_2(and_428_nl, nor_927_nl, fsm_output[3]);
  assign nand_501_nl = ~((fsm_output[5]) & mux_490_nl);
  assign nor_929_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:1]!=4'b0010) | nand_448_cse);
  assign nor_930_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b00101) | (fsm_output[7]));
  assign mux_481_nl = MUX_s_1_2_2(nor_929_nl, nor_930_nl, fsm_output[4]);
  assign nor_931_nl = ~((COMP_LOOP_acc_14_psp_sva[3:0]!=4'b0010) | (~ (fsm_output[7])));
  assign nor_932_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0010) | (fsm_output[7]));
  assign mux_480_nl = MUX_s_1_2_2(nor_931_nl, nor_932_nl, fsm_output[4]);
  assign and_429_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_480_nl;
  assign mux_482_nl = MUX_s_1_2_2(mux_481_nl, and_429_nl, fsm_output[0]);
  assign nand_36_nl = ~((fsm_output[6]) & mux_482_nl);
  assign or_502_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b00101) | (~ (fsm_output[7]));
  assign or_500_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b00101) | (fsm_output[7]);
  assign mux_478_nl = MUX_s_1_2_2(or_502_nl, or_500_nl, fsm_output[4]);
  assign nand_34_nl = ~(nor_98_cse & mux_477_cse);
  assign mux_479_nl = MUX_s_1_2_2(mux_478_nl, nand_34_nl, fsm_output[0]);
  assign or_503_nl = (fsm_output[6]) | mux_479_nl;
  assign mux_483_nl = MUX_s_1_2_2(nand_36_nl, or_503_nl, fsm_output[3]);
  assign or_2275_nl = (fsm_output[5]) | mux_483_nl;
  assign mux_491_nl = MUX_s_1_2_2(nand_501_nl, or_2275_nl, fsm_output[2]);
  assign vec_rsc_0_5_i_we_d_pff = ~(mux_491_nl | (fsm_output[1]));
  assign nor_917_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b00101) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_918_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_505_nl = MUX_s_1_2_2(nor_917_nl, nor_918_nl, fsm_output[0]);
  assign and_426_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (~ mux_472_cse);
  assign nor_919_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b00101) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_920_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b00101) | (fsm_output[7:6]!=2'b10));
  assign nor_921_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b00101) | (fsm_output[7:6]!=2'b00));
  assign mux_499_nl = MUX_s_1_2_2(nor_920_nl, nor_921_nl, fsm_output[4]);
  assign mux_500_nl = MUX_s_1_2_2(nor_919_nl, mux_499_nl, fsm_output[3]);
  assign mux_504_nl = MUX_s_1_2_2(and_426_nl, mux_500_nl, fsm_output[0]);
  assign mux_506_nl = MUX_s_1_2_2(mux_505_nl, mux_504_nl, fsm_output[5]);
  assign or_535_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b00101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_533_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b00101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_496_nl = MUX_s_1_2_2(or_535_nl, or_533_nl, fsm_output[4]);
  assign or_532_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00101) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_530_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b00101) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_495_nl = MUX_s_1_2_2(or_532_nl, or_530_nl, fsm_output[4]);
  assign mux_497_nl = MUX_s_1_2_2(mux_496_nl, mux_495_nl, fsm_output[3]);
  assign or_529_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:1]!=4'b0010) | nand_444_cse;
  assign or_527_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b00101) | (fsm_output[7:6]!=2'b01);
  assign mux_493_nl = MUX_s_1_2_2(or_529_nl, or_527_nl, fsm_output[4]);
  assign or_526_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00101) | (fsm_output[7:6]!=2'b10);
  assign or_524_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b00101) | (fsm_output[7:6]!=2'b00);
  assign mux_492_nl = MUX_s_1_2_2(or_526_nl, or_524_nl, fsm_output[4]);
  assign mux_494_nl = MUX_s_1_2_2(mux_493_nl, mux_492_nl, fsm_output[3]);
  assign mux_498_nl = MUX_s_1_2_2(mux_497_nl, mux_494_nl, fsm_output[0]);
  assign nor_922_nl = ~((fsm_output[5]) | mux_498_nl);
  assign mux_507_nl = MUX_s_1_2_2(mux_506_nl, nor_922_nl, fsm_output[2]);
  assign vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d = mux_507_nl & (fsm_output[1]);
  assign nor_908_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b00110) | (~ (fsm_output[7])));
  assign nor_909_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b00110) | (fsm_output[7]));
  assign mux_519_nl = MUX_s_1_2_2(nor_908_nl, nor_909_nl, fsm_output[4]);
  assign nor_910_nl = ~((COMP_LOOP_acc_1_cse_sva[4:0]!=5'b00110) | (~ (fsm_output[7])));
  assign nor_911_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b00110) | (fsm_output[7]));
  assign mux_518_nl = MUX_s_1_2_2(nor_910_nl, nor_911_nl, fsm_output[4]);
  assign mux_520_nl = MUX_s_1_2_2(mux_519_nl, mux_518_nl, fsm_output[0]);
  assign and_425_nl = (fsm_output[6]) & mux_520_nl;
  assign or_569_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00110) | (~ (fsm_output[7]));
  assign or_567_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b00110) | (fsm_output[7]);
  assign mux_516_nl = MUX_s_1_2_2(or_569_nl, or_567_nl, fsm_output[4]);
  assign or_566_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00110) | (~ (fsm_output[7]));
  assign or_564_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b00110) | (fsm_output[7]);
  assign mux_515_nl = MUX_s_1_2_2(or_566_nl, or_564_nl, fsm_output[4]);
  assign mux_517_nl = MUX_s_1_2_2(mux_516_nl, mux_515_nl, fsm_output[0]);
  assign nor_912_nl = ~((fsm_output[6]) | mux_517_nl);
  assign mux_521_nl = MUX_s_1_2_2(and_425_nl, nor_912_nl, fsm_output[3]);
  assign nand_500_nl = ~((fsm_output[5]) & mux_521_nl);
  assign nor_914_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b00110) | (~ (fsm_output[7])));
  assign nor_915_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b00110) | (fsm_output[7]));
  assign mux_512_nl = MUX_s_1_2_2(nor_914_nl, nor_915_nl, fsm_output[4]);
  assign or_558_nl = (COMP_LOOP_acc_14_psp_sva[3:2]!=2'b00) | nand_423_cse;
  assign or_556_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0011) | (fsm_output[7]);
  assign mux_511_nl = MUX_s_1_2_2(or_558_nl, or_556_nl, fsm_output[4]);
  assign nor_916_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_511_nl);
  assign mux_513_nl = MUX_s_1_2_2(mux_512_nl, nor_916_nl, fsm_output[0]);
  assign nand_41_nl = ~((fsm_output[6]) & mux_513_nl);
  assign or_554_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[2]))
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[3]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[4])
      | nand_442_cse;
  assign or_552_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b00110) | (fsm_output[7]);
  assign mux_509_nl = MUX_s_1_2_2(or_554_nl, or_552_nl, fsm_output[4]);
  assign or_551_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | mux_446_cse;
  assign mux_510_nl = MUX_s_1_2_2(mux_509_nl, or_551_nl, fsm_output[0]);
  assign or_555_nl = (fsm_output[6]) | mux_510_nl;
  assign mux_514_nl = MUX_s_1_2_2(nand_41_nl, or_555_nl, fsm_output[3]);
  assign or_2274_nl = (fsm_output[5]) | mux_514_nl;
  assign mux_522_nl = MUX_s_1_2_2(nand_500_nl, or_2274_nl, fsm_output[2]);
  assign vec_rsc_0_6_i_we_d_pff = ~(mux_522_nl | (fsm_output[1]));
  assign nor_901_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b00110) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_902_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_536_nl = MUX_s_1_2_2(nor_901_nl, nor_902_nl, fsm_output[0]);
  assign nor_903_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_534_cse);
  assign nor_904_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b00110) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_905_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b00110) | (fsm_output[7:6]!=2'b10));
  assign nor_906_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b00110) | (fsm_output[7:6]!=2'b00));
  assign mux_530_nl = MUX_s_1_2_2(nor_905_nl, nor_906_nl, fsm_output[4]);
  assign mux_531_nl = MUX_s_1_2_2(nor_904_nl, mux_530_nl, fsm_output[3]);
  assign mux_535_nl = MUX_s_1_2_2(nor_903_nl, mux_531_nl, fsm_output[0]);
  assign mux_537_nl = MUX_s_1_2_2(mux_536_nl, mux_535_nl, fsm_output[5]);
  assign or_588_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b00110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_586_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b00110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_527_nl = MUX_s_1_2_2(or_588_nl, or_586_nl, fsm_output[4]);
  assign or_585_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00110) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_583_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b00110) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_526_nl = MUX_s_1_2_2(or_585_nl, or_583_nl, fsm_output[4]);
  assign mux_528_nl = MUX_s_1_2_2(mux_527_nl, mux_526_nl, fsm_output[3]);
  assign or_582_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b00110) | nand_443_cse;
  assign or_580_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b00110) | (fsm_output[7:6]!=2'b01);
  assign mux_524_nl = MUX_s_1_2_2(or_582_nl, or_580_nl, fsm_output[4]);
  assign or_579_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00110) | (fsm_output[7:6]!=2'b10);
  assign or_577_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b00110) | (fsm_output[7:6]!=2'b00);
  assign mux_523_nl = MUX_s_1_2_2(or_579_nl, or_577_nl, fsm_output[4]);
  assign mux_525_nl = MUX_s_1_2_2(mux_524_nl, mux_523_nl, fsm_output[3]);
  assign mux_529_nl = MUX_s_1_2_2(mux_528_nl, mux_525_nl, fsm_output[0]);
  assign nor_907_nl = ~((fsm_output[5]) | mux_529_nl);
  assign mux_538_nl = MUX_s_1_2_2(mux_537_nl, nor_907_nl, fsm_output[2]);
  assign vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d = mux_538_nl & (fsm_output[1]);
  assign nor_889_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:1]!=4'b0011) | nand_445_cse);
  assign nor_890_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b00111) | (fsm_output[7]));
  assign mux_550_nl = MUX_s_1_2_2(nor_889_nl, nor_890_nl, fsm_output[4]);
  assign nor_891_nl = ~((COMP_LOOP_acc_1_cse_sva[4:3]!=2'b00) | nand_417_cse);
  assign nor_892_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b00111) | (fsm_output[7]));
  assign mux_549_nl = MUX_s_1_2_2(nor_891_nl, nor_892_nl, fsm_output[4]);
  assign mux_551_nl = MUX_s_1_2_2(mux_550_nl, mux_549_nl, fsm_output[0]);
  assign and_422_nl = (fsm_output[6]) & mux_551_nl;
  assign or_620_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00111) | (~ (fsm_output[7]));
  assign or_618_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b00111) | (fsm_output[7]);
  assign mux_547_nl = MUX_s_1_2_2(or_620_nl, or_618_nl, fsm_output[4]);
  assign or_617_nl = (COMP_LOOP_acc_1_cse_6_sva[4:1]!=4'b0011) | nand_447_cse;
  assign or_615_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b00111) | (fsm_output[7]);
  assign mux_546_nl = MUX_s_1_2_2(or_617_nl, or_615_nl, fsm_output[4]);
  assign mux_548_nl = MUX_s_1_2_2(mux_547_nl, mux_546_nl, fsm_output[0]);
  assign nor_893_nl = ~((fsm_output[6]) | mux_548_nl);
  assign mux_552_nl = MUX_s_1_2_2(and_422_nl, nor_893_nl, fsm_output[3]);
  assign nand_499_nl = ~((fsm_output[5]) & mux_552_nl);
  assign nor_895_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:3]!=2'b00) | nand_419_cse);
  assign nor_896_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b00111) | (fsm_output[7]));
  assign mux_543_nl = MUX_s_1_2_2(nor_895_nl, nor_896_nl, fsm_output[4]);
  assign nor_897_nl = ~((COMP_LOOP_acc_14_psp_sva[3:2]!=2'b00) | nand_423_cse);
  assign nor_898_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0011) | (fsm_output[7]));
  assign mux_542_nl = MUX_s_1_2_2(nor_897_nl, nor_898_nl, fsm_output[4]);
  assign and_423_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_542_nl;
  assign mux_544_nl = MUX_s_1_2_2(mux_543_nl, and_423_nl, fsm_output[0]);
  assign nand_47_nl = ~((fsm_output[6]) & mux_544_nl);
  assign or_606_nl = (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[0])) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[2]))
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[3]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[4])
      | nand_442_cse;
  assign or_604_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b00111) | (fsm_output[7]);
  assign mux_540_nl = MUX_s_1_2_2(or_606_nl, or_604_nl, fsm_output[4]);
  assign nand_45_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & mux_477_cse);
  assign mux_541_nl = MUX_s_1_2_2(mux_540_nl, nand_45_nl, fsm_output[0]);
  assign or_607_nl = (fsm_output[6]) | mux_541_nl;
  assign mux_545_nl = MUX_s_1_2_2(nand_47_nl, or_607_nl, fsm_output[3]);
  assign or_2273_nl = (fsm_output[5]) | mux_545_nl;
  assign mux_553_nl = MUX_s_1_2_2(nand_499_nl, or_2273_nl, fsm_output[2]);
  assign vec_rsc_0_7_i_we_d_pff = ~(mux_553_nl | (fsm_output[1]));
  assign nor_883_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b00111) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_884_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_567_nl = MUX_s_1_2_2(nor_883_nl, nor_884_nl, fsm_output[0]);
  assign and_420_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (~ mux_534_cse);
  assign nor_885_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b00111) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_886_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b00111) | (fsm_output[7:6]!=2'b10));
  assign nor_887_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b00111) | (fsm_output[7:6]!=2'b00));
  assign mux_561_nl = MUX_s_1_2_2(nor_886_nl, nor_887_nl, fsm_output[4]);
  assign mux_562_nl = MUX_s_1_2_2(nor_885_nl, mux_561_nl, fsm_output[3]);
  assign mux_566_nl = MUX_s_1_2_2(and_420_nl, mux_562_nl, fsm_output[0]);
  assign mux_568_nl = MUX_s_1_2_2(mux_567_nl, mux_566_nl, fsm_output[5]);
  assign or_639_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b00111) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_637_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b00111) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_558_nl = MUX_s_1_2_2(or_639_nl, or_637_nl, fsm_output[4]);
  assign or_636_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00111) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_634_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b00111) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_557_nl = MUX_s_1_2_2(or_636_nl, or_634_nl, fsm_output[4]);
  assign mux_559_nl = MUX_s_1_2_2(mux_558_nl, mux_557_nl, fsm_output[3]);
  assign or_633_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:1]!=4'b0011) | nand_444_cse;
  assign or_631_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b00111) | (fsm_output[7:6]!=2'b01);
  assign mux_555_nl = MUX_s_1_2_2(or_633_nl, or_631_nl, fsm_output[4]);
  assign or_630_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00111) | (fsm_output[7:6]!=2'b10);
  assign or_628_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b00111) | (fsm_output[7:6]!=2'b00);
  assign mux_554_nl = MUX_s_1_2_2(or_630_nl, or_628_nl, fsm_output[4]);
  assign mux_556_nl = MUX_s_1_2_2(mux_555_nl, mux_554_nl, fsm_output[3]);
  assign mux_560_nl = MUX_s_1_2_2(mux_559_nl, mux_556_nl, fsm_output[0]);
  assign nor_888_nl = ~((fsm_output[5]) | mux_560_nl);
  assign mux_569_nl = MUX_s_1_2_2(mux_568_nl, nor_888_nl, fsm_output[2]);
  assign vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d = mux_569_nl & (fsm_output[1]);
  assign nor_874_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b01000) | (~ (fsm_output[7])));
  assign nor_875_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b01000) | (fsm_output[7]));
  assign mux_581_nl = MUX_s_1_2_2(nor_874_nl, nor_875_nl, fsm_output[4]);
  assign nor_876_nl = ~((COMP_LOOP_acc_1_cse_sva[4:0]!=5'b01000) | (~ (fsm_output[7])));
  assign nor_877_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b01000) | (fsm_output[7]));
  assign mux_580_nl = MUX_s_1_2_2(nor_876_nl, nor_877_nl, fsm_output[4]);
  assign mux_582_nl = MUX_s_1_2_2(mux_581_nl, mux_580_nl, fsm_output[0]);
  assign and_419_nl = (fsm_output[6]) & mux_582_nl;
  assign or_673_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01000) | (~ (fsm_output[7]));
  assign or_671_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b01000) | (fsm_output[7]);
  assign mux_578_nl = MUX_s_1_2_2(or_673_nl, or_671_nl, fsm_output[4]);
  assign or_670_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01000) | (~ (fsm_output[7]));
  assign or_668_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b01000) | (fsm_output[7]);
  assign mux_577_nl = MUX_s_1_2_2(or_670_nl, or_668_nl, fsm_output[4]);
  assign mux_579_nl = MUX_s_1_2_2(mux_578_nl, mux_577_nl, fsm_output[0]);
  assign nor_878_nl = ~((fsm_output[6]) | mux_579_nl);
  assign mux_583_nl = MUX_s_1_2_2(and_419_nl, nor_878_nl, fsm_output[3]);
  assign nand_498_nl = ~((fsm_output[5]) & mux_583_nl);
  assign nor_880_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b01000) | (~ (fsm_output[7])));
  assign nor_881_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b01000) | (fsm_output[7]));
  assign mux_574_nl = MUX_s_1_2_2(nor_880_nl, nor_881_nl, fsm_output[4]);
  assign or_662_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b0100) | (~ (fsm_output[7]));
  assign or_660_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0100) | (fsm_output[7]);
  assign mux_573_nl = MUX_s_1_2_2(or_662_nl, or_660_nl, fsm_output[4]);
  assign nor_882_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_573_nl);
  assign mux_575_nl = MUX_s_1_2_2(mux_574_nl, nor_882_nl, fsm_output[0]);
  assign nand_52_nl = ~((fsm_output[6]) & mux_575_nl);
  assign or_658_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b01000) | (~ (fsm_output[7]));
  assign or_656_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b01000) | (fsm_output[7]);
  assign mux_571_nl = MUX_s_1_2_2(or_658_nl, or_656_nl, fsm_output[4]);
  assign or_655_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | mux_570_cse;
  assign mux_572_nl = MUX_s_1_2_2(mux_571_nl, or_655_nl, fsm_output[0]);
  assign or_659_nl = (fsm_output[6]) | mux_572_nl;
  assign mux_576_nl = MUX_s_1_2_2(nand_52_nl, or_659_nl, fsm_output[3]);
  assign or_2272_nl = (fsm_output[5]) | mux_576_nl;
  assign mux_584_nl = MUX_s_1_2_2(nand_498_nl, or_2272_nl, fsm_output[2]);
  assign vec_rsc_0_8_i_we_d_pff = ~(mux_584_nl | (fsm_output[1]));
  assign nor_867_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b01000) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_868_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_598_nl = MUX_s_1_2_2(nor_867_nl, nor_868_nl, fsm_output[0]);
  assign nor_869_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_596_cse);
  assign nor_870_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b01000) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_871_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b01000) | (fsm_output[7:6]!=2'b10));
  assign nor_872_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b01000) | (fsm_output[7:6]!=2'b00));
  assign mux_592_nl = MUX_s_1_2_2(nor_871_nl, nor_872_nl, fsm_output[4]);
  assign mux_593_nl = MUX_s_1_2_2(nor_870_nl, mux_592_nl, fsm_output[3]);
  assign mux_597_nl = MUX_s_1_2_2(nor_869_nl, mux_593_nl, fsm_output[0]);
  assign mux_599_nl = MUX_s_1_2_2(mux_598_nl, mux_597_nl, fsm_output[5]);
  assign or_692_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b01000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_690_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b01000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_589_nl = MUX_s_1_2_2(or_692_nl, or_690_nl, fsm_output[4]);
  assign or_689_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01000) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_687_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b01000) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_588_nl = MUX_s_1_2_2(or_689_nl, or_687_nl, fsm_output[4]);
  assign mux_590_nl = MUX_s_1_2_2(mux_589_nl, mux_588_nl, fsm_output[3]);
  assign or_686_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b01000) | nand_443_cse;
  assign or_684_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b01000) | (fsm_output[7:6]!=2'b01);
  assign mux_586_nl = MUX_s_1_2_2(or_686_nl, or_684_nl, fsm_output[4]);
  assign or_683_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01000) | (fsm_output[7:6]!=2'b10);
  assign or_681_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b01000) | (fsm_output[7:6]!=2'b00);
  assign mux_585_nl = MUX_s_1_2_2(or_683_nl, or_681_nl, fsm_output[4]);
  assign mux_587_nl = MUX_s_1_2_2(mux_586_nl, mux_585_nl, fsm_output[3]);
  assign mux_591_nl = MUX_s_1_2_2(mux_590_nl, mux_587_nl, fsm_output[0]);
  assign nor_873_nl = ~((fsm_output[5]) | mux_591_nl);
  assign mux_600_nl = MUX_s_1_2_2(mux_599_nl, nor_873_nl, fsm_output[2]);
  assign vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d = mux_600_nl & (fsm_output[1]);
  assign nor_855_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:1]!=4'b0100) | nand_445_cse);
  assign nor_856_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b01001) | (fsm_output[7]));
  assign mux_612_nl = MUX_s_1_2_2(nor_855_nl, nor_856_nl, fsm_output[4]);
  assign nor_857_nl = ~((COMP_LOOP_acc_1_cse_sva[4:1]!=4'b0100) | nand_446_cse);
  assign nor_858_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b01001) | (fsm_output[7]));
  assign mux_611_nl = MUX_s_1_2_2(nor_857_nl, nor_858_nl, fsm_output[4]);
  assign mux_613_nl = MUX_s_1_2_2(mux_612_nl, mux_611_nl, fsm_output[0]);
  assign and_416_nl = (fsm_output[6]) & mux_613_nl;
  assign or_724_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01001) | (~ (fsm_output[7]));
  assign or_722_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b01001) | (fsm_output[7]);
  assign mux_609_nl = MUX_s_1_2_2(or_724_nl, or_722_nl, fsm_output[4]);
  assign or_721_nl = (COMP_LOOP_acc_1_cse_6_sva[2]) | (COMP_LOOP_acc_1_cse_6_sva[1])
      | (COMP_LOOP_acc_1_cse_6_sva[4]) | nand_411_cse;
  assign or_719_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b01001) | (fsm_output[7]);
  assign mux_608_nl = MUX_s_1_2_2(or_721_nl, or_719_nl, fsm_output[4]);
  assign mux_610_nl = MUX_s_1_2_2(mux_609_nl, mux_608_nl, fsm_output[0]);
  assign nor_859_nl = ~((fsm_output[6]) | mux_610_nl);
  assign mux_614_nl = MUX_s_1_2_2(and_416_nl, nor_859_nl, fsm_output[3]);
  assign nand_497_nl = ~((fsm_output[5]) & mux_614_nl);
  assign nor_861_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:1]!=4'b0100) | nand_448_cse);
  assign nor_862_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b01001) | (fsm_output[7]));
  assign mux_605_nl = MUX_s_1_2_2(nor_861_nl, nor_862_nl, fsm_output[4]);
  assign nor_863_nl = ~((COMP_LOOP_acc_14_psp_sva[3:0]!=4'b0100) | (~ (fsm_output[7])));
  assign nor_864_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0100) | (fsm_output[7]));
  assign mux_604_nl = MUX_s_1_2_2(nor_863_nl, nor_864_nl, fsm_output[4]);
  assign and_417_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_604_nl;
  assign mux_606_nl = MUX_s_1_2_2(mux_605_nl, and_417_nl, fsm_output[0]);
  assign nand_58_nl = ~((fsm_output[6]) & mux_606_nl);
  assign or_710_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b01001) | (~ (fsm_output[7]));
  assign or_708_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b01001) | (fsm_output[7]);
  assign mux_602_nl = MUX_s_1_2_2(or_710_nl, or_708_nl, fsm_output[4]);
  assign nand_56_nl = ~(nor_98_cse & mux_601_cse);
  assign mux_603_nl = MUX_s_1_2_2(mux_602_nl, nand_56_nl, fsm_output[0]);
  assign or_711_nl = (fsm_output[6]) | mux_603_nl;
  assign mux_607_nl = MUX_s_1_2_2(nand_58_nl, or_711_nl, fsm_output[3]);
  assign or_2271_nl = (fsm_output[5]) | mux_607_nl;
  assign mux_615_nl = MUX_s_1_2_2(nand_497_nl, or_2271_nl, fsm_output[2]);
  assign vec_rsc_0_9_i_we_d_pff = ~(mux_615_nl | (fsm_output[1]));
  assign nor_849_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b01001) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_850_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_629_nl = MUX_s_1_2_2(nor_849_nl, nor_850_nl, fsm_output[0]);
  assign and_414_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (~ mux_596_cse);
  assign nor_851_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b01001) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_852_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b01001) | (fsm_output[7:6]!=2'b10));
  assign nor_853_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b01001) | (fsm_output[7:6]!=2'b00));
  assign mux_623_nl = MUX_s_1_2_2(nor_852_nl, nor_853_nl, fsm_output[4]);
  assign mux_624_nl = MUX_s_1_2_2(nor_851_nl, mux_623_nl, fsm_output[3]);
  assign mux_628_nl = MUX_s_1_2_2(and_414_nl, mux_624_nl, fsm_output[0]);
  assign mux_630_nl = MUX_s_1_2_2(mux_629_nl, mux_628_nl, fsm_output[5]);
  assign or_743_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b01001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_741_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b01001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_620_nl = MUX_s_1_2_2(or_743_nl, or_741_nl, fsm_output[4]);
  assign or_740_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01001) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_738_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b01001) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_619_nl = MUX_s_1_2_2(or_740_nl, or_738_nl, fsm_output[4]);
  assign mux_621_nl = MUX_s_1_2_2(mux_620_nl, mux_619_nl, fsm_output[3]);
  assign or_737_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:1]!=4'b0100) | nand_444_cse;
  assign or_735_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b01001) | (fsm_output[7:6]!=2'b01);
  assign mux_617_nl = MUX_s_1_2_2(or_737_nl, or_735_nl, fsm_output[4]);
  assign or_734_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01001) | (fsm_output[7:6]!=2'b10);
  assign or_732_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b01001) | (fsm_output[7:6]!=2'b00);
  assign mux_616_nl = MUX_s_1_2_2(or_734_nl, or_732_nl, fsm_output[4]);
  assign mux_618_nl = MUX_s_1_2_2(mux_617_nl, mux_616_nl, fsm_output[3]);
  assign mux_622_nl = MUX_s_1_2_2(mux_621_nl, mux_618_nl, fsm_output[0]);
  assign nor_854_nl = ~((fsm_output[5]) | mux_622_nl);
  assign mux_631_nl = MUX_s_1_2_2(mux_630_nl, nor_854_nl, fsm_output[2]);
  assign vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d = mux_631_nl & (fsm_output[1]);
  assign nor_840_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b01010) | (~ (fsm_output[7])));
  assign nor_841_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b01010) | (fsm_output[7]));
  assign mux_643_nl = MUX_s_1_2_2(nor_840_nl, nor_841_nl, fsm_output[4]);
  assign nor_842_nl = ~((COMP_LOOP_acc_1_cse_sva[4:0]!=5'b01010) | (~ (fsm_output[7])));
  assign nor_843_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b01010) | (fsm_output[7]));
  assign mux_642_nl = MUX_s_1_2_2(nor_842_nl, nor_843_nl, fsm_output[4]);
  assign mux_644_nl = MUX_s_1_2_2(mux_643_nl, mux_642_nl, fsm_output[0]);
  assign and_413_nl = (fsm_output[6]) & mux_644_nl;
  assign or_777_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01010) | (~ (fsm_output[7]));
  assign or_775_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b01010) | (fsm_output[7]);
  assign mux_640_nl = MUX_s_1_2_2(or_777_nl, or_775_nl, fsm_output[4]);
  assign or_774_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01010) | (~ (fsm_output[7]));
  assign or_772_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b01010) | (fsm_output[7]);
  assign mux_639_nl = MUX_s_1_2_2(or_774_nl, or_772_nl, fsm_output[4]);
  assign mux_641_nl = MUX_s_1_2_2(mux_640_nl, mux_639_nl, fsm_output[0]);
  assign nor_844_nl = ~((fsm_output[6]) | mux_641_nl);
  assign mux_645_nl = MUX_s_1_2_2(and_413_nl, nor_844_nl, fsm_output[3]);
  assign nand_496_nl = ~((fsm_output[5]) & mux_645_nl);
  assign nor_846_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b01010) | (~ (fsm_output[7])));
  assign nor_847_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b01010) | (fsm_output[7]));
  assign mux_636_nl = MUX_s_1_2_2(nor_846_nl, nor_847_nl, fsm_output[4]);
  assign or_766_nl = (COMP_LOOP_acc_14_psp_sva[3:1]!=3'b010) | nand_441_cse;
  assign or_764_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0101) | (fsm_output[7]);
  assign mux_635_nl = MUX_s_1_2_2(or_766_nl, or_764_nl, fsm_output[4]);
  assign nor_848_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_635_nl);
  assign mux_637_nl = MUX_s_1_2_2(mux_636_nl, nor_848_nl, fsm_output[0]);
  assign nand_63_nl = ~((fsm_output[6]) & mux_637_nl);
  assign or_762_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[3])) | (COMP_LOOP_acc_10_cse_10_1_5_sva[4])
      | nand_442_cse;
  assign or_760_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b01010) | (fsm_output[7]);
  assign mux_633_nl = MUX_s_1_2_2(or_762_nl, or_760_nl, fsm_output[4]);
  assign or_759_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | mux_570_cse;
  assign mux_634_nl = MUX_s_1_2_2(mux_633_nl, or_759_nl, fsm_output[0]);
  assign or_763_nl = (fsm_output[6]) | mux_634_nl;
  assign mux_638_nl = MUX_s_1_2_2(nand_63_nl, or_763_nl, fsm_output[3]);
  assign or_2270_nl = (fsm_output[5]) | mux_638_nl;
  assign mux_646_nl = MUX_s_1_2_2(nand_496_nl, or_2270_nl, fsm_output[2]);
  assign vec_rsc_0_10_i_we_d_pff = ~(mux_646_nl | (fsm_output[1]));
  assign nor_833_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b01010) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_834_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_660_nl = MUX_s_1_2_2(nor_833_nl, nor_834_nl, fsm_output[0]);
  assign nor_835_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_658_cse);
  assign nor_836_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b01010) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_837_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b01010) | (fsm_output[7:6]!=2'b10));
  assign nor_838_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b01010) | (fsm_output[7:6]!=2'b00));
  assign mux_654_nl = MUX_s_1_2_2(nor_837_nl, nor_838_nl, fsm_output[4]);
  assign mux_655_nl = MUX_s_1_2_2(nor_836_nl, mux_654_nl, fsm_output[3]);
  assign mux_659_nl = MUX_s_1_2_2(nor_835_nl, mux_655_nl, fsm_output[0]);
  assign mux_661_nl = MUX_s_1_2_2(mux_660_nl, mux_659_nl, fsm_output[5]);
  assign or_796_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b01010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_794_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b01010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_651_nl = MUX_s_1_2_2(or_796_nl, or_794_nl, fsm_output[4]);
  assign or_793_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01010) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_791_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b01010) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_650_nl = MUX_s_1_2_2(or_793_nl, or_791_nl, fsm_output[4]);
  assign mux_652_nl = MUX_s_1_2_2(mux_651_nl, mux_650_nl, fsm_output[3]);
  assign or_790_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b01010) | nand_443_cse;
  assign or_788_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b01010) | (fsm_output[7:6]!=2'b01);
  assign mux_648_nl = MUX_s_1_2_2(or_790_nl, or_788_nl, fsm_output[4]);
  assign or_787_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01010) | (fsm_output[7:6]!=2'b10);
  assign or_785_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b01010) | (fsm_output[7:6]!=2'b00);
  assign mux_647_nl = MUX_s_1_2_2(or_787_nl, or_785_nl, fsm_output[4]);
  assign mux_649_nl = MUX_s_1_2_2(mux_648_nl, mux_647_nl, fsm_output[3]);
  assign mux_653_nl = MUX_s_1_2_2(mux_652_nl, mux_649_nl, fsm_output[0]);
  assign nor_839_nl = ~((fsm_output[5]) | mux_653_nl);
  assign mux_662_nl = MUX_s_1_2_2(mux_661_nl, nor_839_nl, fsm_output[2]);
  assign vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d = mux_662_nl & (fsm_output[1]);
  assign nor_821_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:1]!=4'b0101) | nand_445_cse);
  assign nor_822_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b01011) | (fsm_output[7]));
  assign mux_674_nl = MUX_s_1_2_2(nor_821_nl, nor_822_nl, fsm_output[4]);
  assign nor_823_nl = ~((COMP_LOOP_acc_1_cse_sva[4:2]!=3'b010) | nand_435_cse);
  assign nor_824_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b01011) | (fsm_output[7]));
  assign mux_673_nl = MUX_s_1_2_2(nor_823_nl, nor_824_nl, fsm_output[4]);
  assign mux_675_nl = MUX_s_1_2_2(mux_674_nl, mux_673_nl, fsm_output[0]);
  assign and_410_nl = (fsm_output[6]) & mux_675_nl;
  assign or_828_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01011) | (~ (fsm_output[7]));
  assign or_826_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b01011) | (fsm_output[7]);
  assign mux_671_nl = MUX_s_1_2_2(or_828_nl, or_826_nl, fsm_output[4]);
  assign or_825_nl = (COMP_LOOP_acc_1_cse_6_sva[2]) | (~ (COMP_LOOP_acc_1_cse_6_sva[1]))
      | (COMP_LOOP_acc_1_cse_6_sva[4]) | nand_411_cse;
  assign or_823_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b01011) | (fsm_output[7]);
  assign mux_670_nl = MUX_s_1_2_2(or_825_nl, or_823_nl, fsm_output[4]);
  assign mux_672_nl = MUX_s_1_2_2(mux_671_nl, mux_670_nl, fsm_output[0]);
  assign nor_825_nl = ~((fsm_output[6]) | mux_672_nl);
  assign mux_676_nl = MUX_s_1_2_2(and_410_nl, nor_825_nl, fsm_output[3]);
  assign nand_495_nl = ~((fsm_output[5]) & mux_676_nl);
  assign nor_827_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:2]!=3'b010) | nand_437_cse);
  assign nor_828_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b01011) | (fsm_output[7]));
  assign mux_667_nl = MUX_s_1_2_2(nor_827_nl, nor_828_nl, fsm_output[4]);
  assign nor_829_nl = ~((COMP_LOOP_acc_14_psp_sva[3:1]!=3'b010) | nand_441_cse);
  assign nor_830_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0101) | (fsm_output[7]));
  assign mux_666_nl = MUX_s_1_2_2(nor_829_nl, nor_830_nl, fsm_output[4]);
  assign and_411_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_666_nl;
  assign mux_668_nl = MUX_s_1_2_2(mux_667_nl, and_411_nl, fsm_output[0]);
  assign nand_69_nl = ~((fsm_output[6]) & mux_668_nl);
  assign or_814_nl = (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[0])) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[3])) | (COMP_LOOP_acc_10_cse_10_1_5_sva[4])
      | nand_442_cse;
  assign or_812_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b01011) | (fsm_output[7]);
  assign mux_664_nl = MUX_s_1_2_2(or_814_nl, or_812_nl, fsm_output[4]);
  assign nand_67_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & mux_601_cse);
  assign mux_665_nl = MUX_s_1_2_2(mux_664_nl, nand_67_nl, fsm_output[0]);
  assign or_815_nl = (fsm_output[6]) | mux_665_nl;
  assign mux_669_nl = MUX_s_1_2_2(nand_69_nl, or_815_nl, fsm_output[3]);
  assign or_2269_nl = (fsm_output[5]) | mux_669_nl;
  assign mux_677_nl = MUX_s_1_2_2(nand_495_nl, or_2269_nl, fsm_output[2]);
  assign vec_rsc_0_11_i_we_d_pff = ~(mux_677_nl | (fsm_output[1]));
  assign nor_815_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b01011) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_816_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_691_nl = MUX_s_1_2_2(nor_815_nl, nor_816_nl, fsm_output[0]);
  assign and_408_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (~ mux_658_cse);
  assign nor_817_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b01011) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_818_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b01011) | (fsm_output[7:6]!=2'b10));
  assign nor_819_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b01011) | (fsm_output[7:6]!=2'b00));
  assign mux_685_nl = MUX_s_1_2_2(nor_818_nl, nor_819_nl, fsm_output[4]);
  assign mux_686_nl = MUX_s_1_2_2(nor_817_nl, mux_685_nl, fsm_output[3]);
  assign mux_690_nl = MUX_s_1_2_2(and_408_nl, mux_686_nl, fsm_output[0]);
  assign mux_692_nl = MUX_s_1_2_2(mux_691_nl, mux_690_nl, fsm_output[5]);
  assign or_847_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b01011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_845_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b01011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_682_nl = MUX_s_1_2_2(or_847_nl, or_845_nl, fsm_output[4]);
  assign or_844_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01011) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_842_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b01011) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_681_nl = MUX_s_1_2_2(or_844_nl, or_842_nl, fsm_output[4]);
  assign mux_683_nl = MUX_s_1_2_2(mux_682_nl, mux_681_nl, fsm_output[3]);
  assign or_841_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:1]!=4'b0101) | nand_444_cse;
  assign or_839_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b01011) | (fsm_output[7:6]!=2'b01);
  assign mux_679_nl = MUX_s_1_2_2(or_841_nl, or_839_nl, fsm_output[4]);
  assign or_838_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01011) | (fsm_output[7:6]!=2'b10);
  assign or_836_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b01011) | (fsm_output[7:6]!=2'b00);
  assign mux_678_nl = MUX_s_1_2_2(or_838_nl, or_836_nl, fsm_output[4]);
  assign mux_680_nl = MUX_s_1_2_2(mux_679_nl, mux_678_nl, fsm_output[3]);
  assign mux_684_nl = MUX_s_1_2_2(mux_683_nl, mux_680_nl, fsm_output[0]);
  assign nor_820_nl = ~((fsm_output[5]) | mux_684_nl);
  assign mux_693_nl = MUX_s_1_2_2(mux_692_nl, nor_820_nl, fsm_output[2]);
  assign vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d = mux_693_nl & (fsm_output[1]);
  assign nor_806_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b01100) | (~ (fsm_output[7])));
  assign nor_807_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b01100) | (fsm_output[7]));
  assign mux_705_nl = MUX_s_1_2_2(nor_806_nl, nor_807_nl, fsm_output[4]);
  assign nor_808_nl = ~((COMP_LOOP_acc_1_cse_sva[4:0]!=5'b01100) | (~ (fsm_output[7])));
  assign nor_809_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b01100) | (fsm_output[7]));
  assign mux_704_nl = MUX_s_1_2_2(nor_808_nl, nor_809_nl, fsm_output[4]);
  assign mux_706_nl = MUX_s_1_2_2(mux_705_nl, mux_704_nl, fsm_output[0]);
  assign and_407_nl = (fsm_output[6]) & mux_706_nl;
  assign or_881_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01100) | (~ (fsm_output[7]));
  assign or_879_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b01100) | (fsm_output[7]);
  assign mux_702_nl = MUX_s_1_2_2(or_881_nl, or_879_nl, fsm_output[4]);
  assign or_878_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01100) | (~ (fsm_output[7]));
  assign or_876_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b01100) | (fsm_output[7]);
  assign mux_701_nl = MUX_s_1_2_2(or_878_nl, or_876_nl, fsm_output[4]);
  assign mux_703_nl = MUX_s_1_2_2(mux_702_nl, mux_701_nl, fsm_output[0]);
  assign nor_810_nl = ~((fsm_output[6]) | mux_703_nl);
  assign mux_707_nl = MUX_s_1_2_2(and_407_nl, nor_810_nl, fsm_output[3]);
  assign nand_494_nl = ~((fsm_output[5]) & mux_707_nl);
  assign nor_812_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b01100) | (~ (fsm_output[7])));
  assign nor_813_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b01100) | (fsm_output[7]));
  assign mux_698_nl = MUX_s_1_2_2(nor_812_nl, nor_813_nl, fsm_output[4]);
  assign or_870_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b0110) | (~ (fsm_output[7]));
  assign or_868_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0110) | (fsm_output[7]);
  assign mux_697_nl = MUX_s_1_2_2(or_870_nl, or_868_nl, fsm_output[4]);
  assign nor_814_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_697_nl);
  assign mux_699_nl = MUX_s_1_2_2(mux_698_nl, nor_814_nl, fsm_output[0]);
  assign nand_74_nl = ~((fsm_output[6]) & mux_699_nl);
  assign or_866_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b01100) | (~ (fsm_output[7]));
  assign or_864_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b01100) | (fsm_output[7]);
  assign mux_695_nl = MUX_s_1_2_2(or_866_nl, or_864_nl, fsm_output[4]);
  assign or_863_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | mux_694_cse;
  assign mux_696_nl = MUX_s_1_2_2(mux_695_nl, or_863_nl, fsm_output[0]);
  assign or_867_nl = (fsm_output[6]) | mux_696_nl;
  assign mux_700_nl = MUX_s_1_2_2(nand_74_nl, or_867_nl, fsm_output[3]);
  assign or_2268_nl = (fsm_output[5]) | mux_700_nl;
  assign mux_708_nl = MUX_s_1_2_2(nand_494_nl, or_2268_nl, fsm_output[2]);
  assign vec_rsc_0_12_i_we_d_pff = ~(mux_708_nl | (fsm_output[1]));
  assign nor_799_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b01100) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_800_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_722_nl = MUX_s_1_2_2(nor_799_nl, nor_800_nl, fsm_output[0]);
  assign nor_801_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_720_cse);
  assign nor_802_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b01100) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_803_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b01100) | (fsm_output[7:6]!=2'b10));
  assign nor_804_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b01100) | (fsm_output[7:6]!=2'b00));
  assign mux_716_nl = MUX_s_1_2_2(nor_803_nl, nor_804_nl, fsm_output[4]);
  assign mux_717_nl = MUX_s_1_2_2(nor_802_nl, mux_716_nl, fsm_output[3]);
  assign mux_721_nl = MUX_s_1_2_2(nor_801_nl, mux_717_nl, fsm_output[0]);
  assign mux_723_nl = MUX_s_1_2_2(mux_722_nl, mux_721_nl, fsm_output[5]);
  assign or_900_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b01100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_898_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b01100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_713_nl = MUX_s_1_2_2(or_900_nl, or_898_nl, fsm_output[4]);
  assign or_897_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01100) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_895_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b01100) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_712_nl = MUX_s_1_2_2(or_897_nl, or_895_nl, fsm_output[4]);
  assign mux_714_nl = MUX_s_1_2_2(mux_713_nl, mux_712_nl, fsm_output[3]);
  assign or_894_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b01100) | nand_443_cse;
  assign or_892_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b01100) | (fsm_output[7:6]!=2'b01);
  assign mux_710_nl = MUX_s_1_2_2(or_894_nl, or_892_nl, fsm_output[4]);
  assign or_891_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01100) | (fsm_output[7:6]!=2'b10);
  assign or_889_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b01100) | (fsm_output[7:6]!=2'b00);
  assign mux_709_nl = MUX_s_1_2_2(or_891_nl, or_889_nl, fsm_output[4]);
  assign mux_711_nl = MUX_s_1_2_2(mux_710_nl, mux_709_nl, fsm_output[3]);
  assign mux_715_nl = MUX_s_1_2_2(mux_714_nl, mux_711_nl, fsm_output[0]);
  assign nor_805_nl = ~((fsm_output[5]) | mux_715_nl);
  assign mux_724_nl = MUX_s_1_2_2(mux_723_nl, nor_805_nl, fsm_output[2]);
  assign vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d = mux_724_nl & (fsm_output[1]);
  assign nor_787_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:1]!=4'b0110) | nand_445_cse);
  assign nor_788_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b01101) | (fsm_output[7]));
  assign mux_736_nl = MUX_s_1_2_2(nor_787_nl, nor_788_nl, fsm_output[4]);
  assign nor_789_nl = ~((COMP_LOOP_acc_1_cse_sva[4:1]!=4'b0110) | nand_446_cse);
  assign nor_790_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b01101) | (fsm_output[7]));
  assign mux_735_nl = MUX_s_1_2_2(nor_789_nl, nor_790_nl, fsm_output[4]);
  assign mux_737_nl = MUX_s_1_2_2(mux_736_nl, mux_735_nl, fsm_output[0]);
  assign and_404_nl = (fsm_output[6]) & mux_737_nl;
  assign or_932_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01101) | (~ (fsm_output[7]));
  assign or_930_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b01101) | (fsm_output[7]);
  assign mux_733_nl = MUX_s_1_2_2(or_932_nl, or_930_nl, fsm_output[4]);
  assign or_929_nl = (~ (COMP_LOOP_acc_1_cse_6_sva[2])) | (COMP_LOOP_acc_1_cse_6_sva[1])
      | (COMP_LOOP_acc_1_cse_6_sva[4]) | nand_411_cse;
  assign or_927_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b01101) | (fsm_output[7]);
  assign mux_732_nl = MUX_s_1_2_2(or_929_nl, or_927_nl, fsm_output[4]);
  assign mux_734_nl = MUX_s_1_2_2(mux_733_nl, mux_732_nl, fsm_output[0]);
  assign nor_791_nl = ~((fsm_output[6]) | mux_734_nl);
  assign mux_738_nl = MUX_s_1_2_2(and_404_nl, nor_791_nl, fsm_output[3]);
  assign nand_493_nl = ~((fsm_output[5]) & mux_738_nl);
  assign nor_793_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:1]!=4'b0110) | nand_448_cse);
  assign nor_794_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b01101) | (fsm_output[7]));
  assign mux_729_nl = MUX_s_1_2_2(nor_793_nl, nor_794_nl, fsm_output[4]);
  assign nor_795_nl = ~((COMP_LOOP_acc_14_psp_sva[3:0]!=4'b0110) | (~ (fsm_output[7])));
  assign nor_796_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0110) | (fsm_output[7]));
  assign mux_728_nl = MUX_s_1_2_2(nor_795_nl, nor_796_nl, fsm_output[4]);
  assign and_405_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_728_nl;
  assign mux_730_nl = MUX_s_1_2_2(mux_729_nl, and_405_nl, fsm_output[0]);
  assign nand_80_nl = ~((fsm_output[6]) & mux_730_nl);
  assign or_918_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b01101) | (~ (fsm_output[7]));
  assign or_916_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b01101) | (fsm_output[7]);
  assign mux_726_nl = MUX_s_1_2_2(or_918_nl, or_916_nl, fsm_output[4]);
  assign nand_78_nl = ~(nor_98_cse & mux_725_cse);
  assign mux_727_nl = MUX_s_1_2_2(mux_726_nl, nand_78_nl, fsm_output[0]);
  assign or_919_nl = (fsm_output[6]) | mux_727_nl;
  assign mux_731_nl = MUX_s_1_2_2(nand_80_nl, or_919_nl, fsm_output[3]);
  assign or_2267_nl = (fsm_output[5]) | mux_731_nl;
  assign mux_739_nl = MUX_s_1_2_2(nand_493_nl, or_2267_nl, fsm_output[2]);
  assign vec_rsc_0_13_i_we_d_pff = ~(mux_739_nl | (fsm_output[1]));
  assign nor_781_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b01101) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_782_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_753_nl = MUX_s_1_2_2(nor_781_nl, nor_782_nl, fsm_output[0]);
  assign and_402_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (~ mux_720_cse);
  assign nor_783_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b01101) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_784_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b01101) | (fsm_output[7:6]!=2'b10));
  assign nor_785_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b01101) | (fsm_output[7:6]!=2'b00));
  assign mux_747_nl = MUX_s_1_2_2(nor_784_nl, nor_785_nl, fsm_output[4]);
  assign mux_748_nl = MUX_s_1_2_2(nor_783_nl, mux_747_nl, fsm_output[3]);
  assign mux_752_nl = MUX_s_1_2_2(and_402_nl, mux_748_nl, fsm_output[0]);
  assign mux_754_nl = MUX_s_1_2_2(mux_753_nl, mux_752_nl, fsm_output[5]);
  assign or_951_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b01101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_949_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b01101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_744_nl = MUX_s_1_2_2(or_951_nl, or_949_nl, fsm_output[4]);
  assign or_948_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01101) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_946_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b01101) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_743_nl = MUX_s_1_2_2(or_948_nl, or_946_nl, fsm_output[4]);
  assign mux_745_nl = MUX_s_1_2_2(mux_744_nl, mux_743_nl, fsm_output[3]);
  assign or_945_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:1]!=4'b0110) | nand_444_cse;
  assign or_943_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b01101) | (fsm_output[7:6]!=2'b01);
  assign mux_741_nl = MUX_s_1_2_2(or_945_nl, or_943_nl, fsm_output[4]);
  assign or_942_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01101) | (fsm_output[7:6]!=2'b10);
  assign or_940_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b01101) | (fsm_output[7:6]!=2'b00);
  assign mux_740_nl = MUX_s_1_2_2(or_942_nl, or_940_nl, fsm_output[4]);
  assign mux_742_nl = MUX_s_1_2_2(mux_741_nl, mux_740_nl, fsm_output[3]);
  assign mux_746_nl = MUX_s_1_2_2(mux_745_nl, mux_742_nl, fsm_output[0]);
  assign nor_786_nl = ~((fsm_output[5]) | mux_746_nl);
  assign mux_755_nl = MUX_s_1_2_2(mux_754_nl, nor_786_nl, fsm_output[2]);
  assign vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d = mux_755_nl & (fsm_output[1]);
  assign nor_772_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b01110) | (~ (fsm_output[7])));
  assign nor_773_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b01110) | (fsm_output[7]));
  assign mux_767_nl = MUX_s_1_2_2(nor_772_nl, nor_773_nl, fsm_output[4]);
  assign nor_774_nl = ~((COMP_LOOP_acc_1_cse_sva[4:0]!=5'b01110) | (~ (fsm_output[7])));
  assign nor_775_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b01110) | (fsm_output[7]));
  assign mux_766_nl = MUX_s_1_2_2(nor_774_nl, nor_775_nl, fsm_output[4]);
  assign mux_768_nl = MUX_s_1_2_2(mux_767_nl, mux_766_nl, fsm_output[0]);
  assign and_401_nl = (fsm_output[6]) & mux_768_nl;
  assign or_984_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01110) | (~ (fsm_output[7]));
  assign or_982_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b01110) | (fsm_output[7]);
  assign mux_764_nl = MUX_s_1_2_2(or_984_nl, or_982_nl, fsm_output[4]);
  assign or_981_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01110) | (~ (fsm_output[7]));
  assign or_979_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b01110) | (fsm_output[7]);
  assign mux_763_nl = MUX_s_1_2_2(or_981_nl, or_979_nl, fsm_output[4]);
  assign mux_765_nl = MUX_s_1_2_2(mux_764_nl, mux_763_nl, fsm_output[0]);
  assign nor_776_nl = ~((fsm_output[6]) | mux_765_nl);
  assign mux_769_nl = MUX_s_1_2_2(and_401_nl, nor_776_nl, fsm_output[3]);
  assign nand_492_nl = ~((fsm_output[5]) & mux_769_nl);
  assign nor_778_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b01110) | (~ (fsm_output[7])));
  assign nor_779_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b01110) | (fsm_output[7]));
  assign mux_760_nl = MUX_s_1_2_2(nor_778_nl, nor_779_nl, fsm_output[4]);
  assign or_973_nl = (COMP_LOOP_acc_14_psp_sva[3]) | nand_385_cse;
  assign or_972_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0111) | (fsm_output[7]);
  assign mux_759_nl = MUX_s_1_2_2(or_973_nl, or_972_nl, fsm_output[4]);
  assign nor_780_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_759_nl);
  assign mux_761_nl = MUX_s_1_2_2(mux_760_nl, nor_780_nl, fsm_output[0]);
  assign nand_85_nl = ~((fsm_output[6]) & mux_761_nl);
  assign or_970_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[2]))
      | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[3])) | (COMP_LOOP_acc_10_cse_10_1_5_sva[4])
      | nand_442_cse;
  assign or_968_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b01110) | (fsm_output[7]);
  assign mux_757_nl = MUX_s_1_2_2(or_970_nl, or_968_nl, fsm_output[4]);
  assign or_967_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | mux_694_cse;
  assign mux_758_nl = MUX_s_1_2_2(mux_757_nl, or_967_nl, fsm_output[0]);
  assign or_971_nl = (fsm_output[6]) | mux_758_nl;
  assign mux_762_nl = MUX_s_1_2_2(nand_85_nl, or_971_nl, fsm_output[3]);
  assign or_2266_nl = (fsm_output[5]) | mux_762_nl;
  assign mux_770_nl = MUX_s_1_2_2(nand_492_nl, or_2266_nl, fsm_output[2]);
  assign vec_rsc_0_14_i_we_d_pff = ~(mux_770_nl | (fsm_output[1]));
  assign nor_765_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b01110) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_766_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_784_nl = MUX_s_1_2_2(nor_765_nl, nor_766_nl, fsm_output[0]);
  assign nor_767_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_782_cse);
  assign nor_768_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b01110) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_769_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b01110) | (fsm_output[7:6]!=2'b10));
  assign nor_770_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b01110) | (fsm_output[7:6]!=2'b00));
  assign mux_778_nl = MUX_s_1_2_2(nor_769_nl, nor_770_nl, fsm_output[4]);
  assign mux_779_nl = MUX_s_1_2_2(nor_768_nl, mux_778_nl, fsm_output[3]);
  assign mux_783_nl = MUX_s_1_2_2(nor_767_nl, mux_779_nl, fsm_output[0]);
  assign mux_785_nl = MUX_s_1_2_2(mux_784_nl, mux_783_nl, fsm_output[5]);
  assign or_1003_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b01110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_1001_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b01110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_775_nl = MUX_s_1_2_2(or_1003_nl, or_1001_nl, fsm_output[4]);
  assign or_1000_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01110) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_998_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b01110) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_774_nl = MUX_s_1_2_2(or_1000_nl, or_998_nl, fsm_output[4]);
  assign mux_776_nl = MUX_s_1_2_2(mux_775_nl, mux_774_nl, fsm_output[3]);
  assign or_997_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b01110) | nand_443_cse;
  assign or_995_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b01110) | (fsm_output[7:6]!=2'b01);
  assign mux_772_nl = MUX_s_1_2_2(or_997_nl, or_995_nl, fsm_output[4]);
  assign or_994_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01110) | (fsm_output[7:6]!=2'b10);
  assign or_992_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b01110) | (fsm_output[7:6]!=2'b00);
  assign mux_771_nl = MUX_s_1_2_2(or_994_nl, or_992_nl, fsm_output[4]);
  assign mux_773_nl = MUX_s_1_2_2(mux_772_nl, mux_771_nl, fsm_output[3]);
  assign mux_777_nl = MUX_s_1_2_2(mux_776_nl, mux_773_nl, fsm_output[0]);
  assign nor_771_nl = ~((fsm_output[5]) | mux_777_nl);
  assign mux_786_nl = MUX_s_1_2_2(mux_785_nl, nor_771_nl, fsm_output[2]);
  assign vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d = mux_786_nl & (fsm_output[1]);
  assign nor_753_nl = ~(nand_371_cse | nand_445_cse);
  assign nor_754_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b01111) | (fsm_output[7]));
  assign mux_798_nl = MUX_s_1_2_2(nor_753_nl, nor_754_nl, fsm_output[4]);
  assign nor_755_nl = ~((COMP_LOOP_acc_1_cse_sva[4]) | (~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1111)
      & (fsm_output[7]))));
  assign nor_756_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b01111) | (fsm_output[7]));
  assign mux_797_nl = MUX_s_1_2_2(nor_755_nl, nor_756_nl, fsm_output[4]);
  assign mux_799_nl = MUX_s_1_2_2(mux_798_nl, mux_797_nl, fsm_output[0]);
  assign and_398_nl = (fsm_output[6]) & mux_799_nl;
  assign nand_516_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]==5'b01111) & (fsm_output[7]));
  assign or_1031_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b01111) | (fsm_output[7]);
  assign mux_795_nl = MUX_s_1_2_2(nand_516_nl, or_1031_nl, fsm_output[4]);
  assign or_1030_nl = (~ (COMP_LOOP_acc_1_cse_6_sva[2])) | (~ (COMP_LOOP_acc_1_cse_6_sva[1]))
      | (COMP_LOOP_acc_1_cse_6_sva[4]) | nand_411_cse;
  assign or_1028_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b01111) | (fsm_output[7]);
  assign mux_794_nl = MUX_s_1_2_2(or_1030_nl, or_1028_nl, fsm_output[4]);
  assign mux_796_nl = MUX_s_1_2_2(mux_795_nl, mux_794_nl, fsm_output[0]);
  assign nor_757_nl = ~((fsm_output[6]) | mux_796_nl);
  assign mux_800_nl = MUX_s_1_2_2(and_398_nl, nor_757_nl, fsm_output[3]);
  assign nand_491_nl = ~((fsm_output[5]) & mux_800_nl);
  assign nor_759_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4]) | (~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]==4'b1111)
      & (fsm_output[7]))));
  assign nor_760_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b01111) | (fsm_output[7]));
  assign mux_791_nl = MUX_s_1_2_2(nor_759_nl, nor_760_nl, fsm_output[4]);
  assign nor_761_nl = ~((COMP_LOOP_acc_14_psp_sva[3]) | nand_385_cse);
  assign nor_762_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]!=4'b0111) | (fsm_output[7]));
  assign mux_790_nl = MUX_s_1_2_2(nor_761_nl, nor_762_nl, fsm_output[4]);
  assign and_399_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_790_nl;
  assign mux_792_nl = MUX_s_1_2_2(mux_791_nl, and_399_nl, fsm_output[0]);
  assign nand_91_nl = ~((fsm_output[6]) & mux_792_nl);
  assign or_1021_nl = (~((COMP_LOOP_acc_10_cse_10_1_5_sva[0]) & (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      & (COMP_LOOP_acc_10_cse_10_1_5_sva[3]) & (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[4]))))
      | nand_442_cse;
  assign or_1019_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b01111) | (fsm_output[7]);
  assign mux_788_nl = MUX_s_1_2_2(or_1021_nl, or_1019_nl, fsm_output[4]);
  assign nand_89_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & mux_725_cse);
  assign mux_789_nl = MUX_s_1_2_2(mux_788_nl, nand_89_nl, fsm_output[0]);
  assign or_1022_nl = (fsm_output[6]) | mux_789_nl;
  assign mux_793_nl = MUX_s_1_2_2(nand_91_nl, or_1022_nl, fsm_output[3]);
  assign or_2265_nl = (fsm_output[5]) | mux_793_nl;
  assign mux_801_nl = MUX_s_1_2_2(nand_491_nl, or_2265_nl, fsm_output[2]);
  assign vec_rsc_0_15_i_we_d_pff = ~(mux_801_nl | (fsm_output[1]));
  assign nor_748_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b01111) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_749_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_815_nl = MUX_s_1_2_2(nor_748_nl, nor_749_nl, fsm_output[0]);
  assign and_395_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (~ mux_782_cse);
  assign and_396_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]==5'b01111) & (fsm_output[4])
      & (fsm_output[6]) & (~ (fsm_output[7]));
  assign and_527_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]==5'b01111) & (fsm_output[7:6]==2'b10);
  assign nor_751_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b01111) | (fsm_output[7:6]!=2'b00));
  assign mux_809_nl = MUX_s_1_2_2(and_527_nl, nor_751_nl, fsm_output[4]);
  assign mux_810_nl = MUX_s_1_2_2(and_396_nl, mux_809_nl, fsm_output[3]);
  assign mux_814_nl = MUX_s_1_2_2(and_395_nl, mux_810_nl, fsm_output[0]);
  assign mux_816_nl = MUX_s_1_2_2(mux_815_nl, mux_814_nl, fsm_output[5]);
  assign or_1051_nl = (~((COMP_LOOP_acc_1_cse_sva[4:0]==5'b01111) & COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm))
      | nand_443_cse;
  assign nand_369_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]==5'b01111) & COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm
      & (fsm_output[7:6]==2'b01));
  assign mux_806_nl = MUX_s_1_2_2(or_1051_nl, nand_369_nl, fsm_output[4]);
  assign nand_515_nl = ~((COMP_LOOP_acc_1_cse_6_sva[4:0]==5'b01111) & COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[7:6]==2'b10));
  assign or_1046_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b01111) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_805_nl = MUX_s_1_2_2(nand_515_nl, or_1046_nl, fsm_output[4]);
  assign mux_807_nl = MUX_s_1_2_2(mux_806_nl, mux_805_nl, fsm_output[3]);
  assign or_1045_nl = nand_371_cse | nand_444_cse;
  assign nand_373_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]==5'b01111) & (fsm_output[7:6]==2'b01));
  assign mux_803_nl = MUX_s_1_2_2(or_1045_nl, nand_373_nl, fsm_output[4]);
  assign nand_471_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]==5'b01111) & (fsm_output[7:6]==2'b10));
  assign or_1040_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b01111) | (fsm_output[7:6]!=2'b00);
  assign mux_802_nl = MUX_s_1_2_2(nand_471_nl, or_1040_nl, fsm_output[4]);
  assign mux_804_nl = MUX_s_1_2_2(mux_803_nl, mux_802_nl, fsm_output[3]);
  assign mux_808_nl = MUX_s_1_2_2(mux_807_nl, mux_804_nl, fsm_output[0]);
  assign nor_752_nl = ~((fsm_output[5]) | mux_808_nl);
  assign mux_817_nl = MUX_s_1_2_2(mux_816_nl, nor_752_nl, fsm_output[2]);
  assign vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d = mux_817_nl & (fsm_output[1]);
  assign nor_739_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b10000) | (~ (fsm_output[7])));
  assign nor_740_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b10000) | (fsm_output[7]));
  assign mux_829_nl = MUX_s_1_2_2(nor_739_nl, nor_740_nl, fsm_output[4]);
  assign nor_741_nl = ~((COMP_LOOP_acc_1_cse_sva[4:0]!=5'b10000) | (~ (fsm_output[7])));
  assign nor_742_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b10000) | (fsm_output[7]));
  assign mux_828_nl = MUX_s_1_2_2(nor_741_nl, nor_742_nl, fsm_output[4]);
  assign mux_830_nl = MUX_s_1_2_2(mux_829_nl, mux_828_nl, fsm_output[0]);
  assign and_394_nl = (fsm_output[6]) & mux_830_nl;
  assign or_1085_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0000) | nand_364_cse;
  assign or_1083_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b10000) | (fsm_output[7]);
  assign mux_826_nl = MUX_s_1_2_2(or_1085_nl, or_1083_nl, fsm_output[4]);
  assign or_1082_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b10000) | (~ (fsm_output[7]));
  assign or_1080_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b10000) | (fsm_output[7]);
  assign mux_825_nl = MUX_s_1_2_2(or_1082_nl, or_1080_nl, fsm_output[4]);
  assign mux_827_nl = MUX_s_1_2_2(mux_826_nl, mux_825_nl, fsm_output[0]);
  assign nor_743_nl = ~((fsm_output[6]) | mux_827_nl);
  assign mux_831_nl = MUX_s_1_2_2(and_394_nl, nor_743_nl, fsm_output[3]);
  assign nand_490_nl = ~((fsm_output[5]) & mux_831_nl);
  assign nor_745_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b10000) | (~ (fsm_output[7])));
  assign nor_746_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b10000) | (fsm_output[7]));
  assign mux_822_nl = MUX_s_1_2_2(nor_745_nl, nor_746_nl, fsm_output[4]);
  assign or_1074_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b1000) | (~ (fsm_output[7]));
  assign or_1072_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1000) | (fsm_output[7]);
  assign mux_821_nl = MUX_s_1_2_2(or_1074_nl, or_1072_nl, fsm_output[4]);
  assign nor_747_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_821_nl);
  assign mux_823_nl = MUX_s_1_2_2(mux_822_nl, nor_747_nl, fsm_output[0]);
  assign nand_96_nl = ~((fsm_output[6]) & mux_823_nl);
  assign or_1070_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b10000) | (~ (fsm_output[7]));
  assign or_1068_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b10000) | (fsm_output[7]);
  assign mux_819_nl = MUX_s_1_2_2(or_1070_nl, or_1068_nl, fsm_output[4]);
  assign or_1067_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | mux_818_cse;
  assign mux_820_nl = MUX_s_1_2_2(mux_819_nl, or_1067_nl, fsm_output[0]);
  assign or_1071_nl = (fsm_output[6]) | mux_820_nl;
  assign mux_824_nl = MUX_s_1_2_2(nand_96_nl, or_1071_nl, fsm_output[3]);
  assign or_2264_nl = (fsm_output[5]) | mux_824_nl;
  assign mux_832_nl = MUX_s_1_2_2(nand_490_nl, or_2264_nl, fsm_output[2]);
  assign vec_rsc_0_16_i_we_d_pff = ~(mux_832_nl | (fsm_output[1]));
  assign nor_732_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b10000) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_733_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_846_nl = MUX_s_1_2_2(nor_732_nl, nor_733_nl, fsm_output[0]);
  assign nor_734_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_844_cse);
  assign nor_735_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b10000) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_736_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b10000) | (fsm_output[7:6]!=2'b10));
  assign nor_737_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b10000) | (fsm_output[7:6]!=2'b00));
  assign mux_840_nl = MUX_s_1_2_2(nor_736_nl, nor_737_nl, fsm_output[4]);
  assign mux_841_nl = MUX_s_1_2_2(nor_735_nl, mux_840_nl, fsm_output[3]);
  assign mux_845_nl = MUX_s_1_2_2(nor_734_nl, mux_841_nl, fsm_output[0]);
  assign mux_847_nl = MUX_s_1_2_2(mux_846_nl, mux_845_nl, fsm_output[5]);
  assign or_1104_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b10000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_1102_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b10000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_837_nl = MUX_s_1_2_2(or_1104_nl, or_1102_nl, fsm_output[4]);
  assign or_1101_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b10000) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_1099_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b10000) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_836_nl = MUX_s_1_2_2(or_1101_nl, or_1099_nl, fsm_output[4]);
  assign mux_838_nl = MUX_s_1_2_2(mux_837_nl, mux_836_nl, fsm_output[3]);
  assign or_1098_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b10000) | nand_443_cse;
  assign or_1096_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b10000) | (fsm_output[7:6]!=2'b01);
  assign mux_834_nl = MUX_s_1_2_2(or_1098_nl, or_1096_nl, fsm_output[4]);
  assign or_1095_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b10000) | (fsm_output[7:6]!=2'b10);
  assign or_1093_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b10000) | (fsm_output[7:6]!=2'b00);
  assign mux_833_nl = MUX_s_1_2_2(or_1095_nl, or_1093_nl, fsm_output[4]);
  assign mux_835_nl = MUX_s_1_2_2(mux_834_nl, mux_833_nl, fsm_output[3]);
  assign mux_839_nl = MUX_s_1_2_2(mux_838_nl, mux_835_nl, fsm_output[0]);
  assign nor_738_nl = ~((fsm_output[5]) | mux_839_nl);
  assign mux_848_nl = MUX_s_1_2_2(mux_847_nl, nor_738_nl, fsm_output[2]);
  assign vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d = mux_848_nl & (fsm_output[1]);
  assign nor_720_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:1]!=3'b000) | nand_357_cse);
  assign nor_721_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b10001) | (fsm_output[7]));
  assign mux_860_nl = MUX_s_1_2_2(nor_720_nl, nor_721_nl, fsm_output[4]);
  assign nor_722_nl = ~((COMP_LOOP_acc_1_cse_sva[4:1]!=4'b1000) | nand_446_cse);
  assign nor_723_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b10001) | (fsm_output[7]));
  assign mux_859_nl = MUX_s_1_2_2(nor_722_nl, nor_723_nl, fsm_output[4]);
  assign mux_861_nl = MUX_s_1_2_2(mux_860_nl, mux_859_nl, fsm_output[0]);
  assign and_391_nl = (fsm_output[6]) & mux_861_nl;
  assign or_1136_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0001) | nand_364_cse;
  assign or_1134_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b10001) | (fsm_output[7]);
  assign mux_857_nl = MUX_s_1_2_2(or_1136_nl, or_1134_nl, fsm_output[4]);
  assign or_1133_nl = (COMP_LOOP_acc_1_cse_6_sva[4:1]!=4'b1000) | nand_447_cse;
  assign or_1131_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b10001) | (fsm_output[7]);
  assign mux_856_nl = MUX_s_1_2_2(or_1133_nl, or_1131_nl, fsm_output[4]);
  assign mux_858_nl = MUX_s_1_2_2(mux_857_nl, mux_856_nl, fsm_output[0]);
  assign nor_724_nl = ~((fsm_output[6]) | mux_858_nl);
  assign mux_862_nl = MUX_s_1_2_2(and_391_nl, nor_724_nl, fsm_output[3]);
  assign nand_489_nl = ~((fsm_output[5]) & mux_862_nl);
  assign nor_726_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:1]!=4'b1000) | nand_448_cse);
  assign nor_727_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b10001) | (fsm_output[7]));
  assign mux_853_nl = MUX_s_1_2_2(nor_726_nl, nor_727_nl, fsm_output[4]);
  assign nor_728_nl = ~((COMP_LOOP_acc_14_psp_sva[3:0]!=4'b1000) | (~ (fsm_output[7])));
  assign nor_729_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1000) | (fsm_output[7]));
  assign mux_852_nl = MUX_s_1_2_2(nor_728_nl, nor_729_nl, fsm_output[4]);
  assign and_392_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_852_nl;
  assign mux_854_nl = MUX_s_1_2_2(mux_853_nl, and_392_nl, fsm_output[0]);
  assign nand_102_nl = ~((fsm_output[6]) & mux_854_nl);
  assign or_1122_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b10001) | (~ (fsm_output[7]));
  assign or_1120_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b10001) | (fsm_output[7]);
  assign mux_850_nl = MUX_s_1_2_2(or_1122_nl, or_1120_nl, fsm_output[4]);
  assign nand_100_nl = ~(nor_98_cse & mux_849_cse);
  assign mux_851_nl = MUX_s_1_2_2(mux_850_nl, nand_100_nl, fsm_output[0]);
  assign or_1123_nl = (fsm_output[6]) | mux_851_nl;
  assign mux_855_nl = MUX_s_1_2_2(nand_102_nl, or_1123_nl, fsm_output[3]);
  assign or_2263_nl = (fsm_output[5]) | mux_855_nl;
  assign mux_863_nl = MUX_s_1_2_2(nand_489_nl, or_2263_nl, fsm_output[2]);
  assign vec_rsc_0_17_i_we_d_pff = ~(mux_863_nl | (fsm_output[1]));
  assign nor_714_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b10001) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_715_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_877_nl = MUX_s_1_2_2(nor_714_nl, nor_715_nl, fsm_output[0]);
  assign and_389_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (~ mux_844_cse);
  assign nor_716_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b10001) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_717_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b10001) | (fsm_output[7:6]!=2'b10));
  assign nor_718_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b10001) | (fsm_output[7:6]!=2'b00));
  assign mux_871_nl = MUX_s_1_2_2(nor_717_nl, nor_718_nl, fsm_output[4]);
  assign mux_872_nl = MUX_s_1_2_2(nor_716_nl, mux_871_nl, fsm_output[3]);
  assign mux_876_nl = MUX_s_1_2_2(and_389_nl, mux_872_nl, fsm_output[0]);
  assign mux_878_nl = MUX_s_1_2_2(mux_877_nl, mux_876_nl, fsm_output[5]);
  assign or_1155_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b10001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_1153_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b10001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_868_nl = MUX_s_1_2_2(or_1155_nl, or_1153_nl, fsm_output[4]);
  assign or_1152_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b10001) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_1150_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b10001) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_867_nl = MUX_s_1_2_2(or_1152_nl, or_1150_nl, fsm_output[4]);
  assign mux_869_nl = MUX_s_1_2_2(mux_868_nl, mux_867_nl, fsm_output[3]);
  assign or_1149_nl = (COMP_LOOP_acc_10_cse_10_1_sva[3:1]!=3'b000) | nand_356_cse;
  assign or_1147_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b10001) | (fsm_output[7:6]!=2'b01);
  assign mux_865_nl = MUX_s_1_2_2(or_1149_nl, or_1147_nl, fsm_output[4]);
  assign or_1146_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b10001) | (fsm_output[7:6]!=2'b10);
  assign or_1144_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b10001) | (fsm_output[7:6]!=2'b00);
  assign mux_864_nl = MUX_s_1_2_2(or_1146_nl, or_1144_nl, fsm_output[4]);
  assign mux_866_nl = MUX_s_1_2_2(mux_865_nl, mux_864_nl, fsm_output[3]);
  assign mux_870_nl = MUX_s_1_2_2(mux_869_nl, mux_866_nl, fsm_output[0]);
  assign nor_719_nl = ~((fsm_output[5]) | mux_870_nl);
  assign mux_879_nl = MUX_s_1_2_2(mux_878_nl, nor_719_nl, fsm_output[2]);
  assign vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d = mux_879_nl & (fsm_output[1]);
  assign nor_705_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b10010) | (~ (fsm_output[7])));
  assign nor_706_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b10010) | (fsm_output[7]));
  assign mux_891_nl = MUX_s_1_2_2(nor_705_nl, nor_706_nl, fsm_output[4]);
  assign nor_707_nl = ~((COMP_LOOP_acc_1_cse_sva[4:0]!=5'b10010) | (~ (fsm_output[7])));
  assign nor_708_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b10010) | (fsm_output[7]));
  assign mux_890_nl = MUX_s_1_2_2(nor_707_nl, nor_708_nl, fsm_output[4]);
  assign mux_892_nl = MUX_s_1_2_2(mux_891_nl, mux_890_nl, fsm_output[0]);
  assign and_388_nl = (fsm_output[6]) & mux_892_nl;
  assign or_1189_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0010) | nand_364_cse;
  assign or_1187_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b10010) | (fsm_output[7]);
  assign mux_888_nl = MUX_s_1_2_2(or_1189_nl, or_1187_nl, fsm_output[4]);
  assign or_1186_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b10010) | (~ (fsm_output[7]));
  assign or_1184_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b10010) | (fsm_output[7]);
  assign mux_887_nl = MUX_s_1_2_2(or_1186_nl, or_1184_nl, fsm_output[4]);
  assign mux_889_nl = MUX_s_1_2_2(mux_888_nl, mux_887_nl, fsm_output[0]);
  assign nor_709_nl = ~((fsm_output[6]) | mux_889_nl);
  assign mux_893_nl = MUX_s_1_2_2(and_388_nl, nor_709_nl, fsm_output[3]);
  assign nand_488_nl = ~((fsm_output[5]) & mux_893_nl);
  assign nor_711_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b10010) | (~ (fsm_output[7])));
  assign nor_712_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b10010) | (fsm_output[7]));
  assign mux_884_nl = MUX_s_1_2_2(nor_711_nl, nor_712_nl, fsm_output[4]);
  assign or_1178_nl = (COMP_LOOP_acc_14_psp_sva[3:1]!=3'b100) | nand_441_cse;
  assign or_1176_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1001) | (fsm_output[7]);
  assign mux_883_nl = MUX_s_1_2_2(or_1178_nl, or_1176_nl, fsm_output[4]);
  assign nor_713_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_883_nl);
  assign mux_885_nl = MUX_s_1_2_2(mux_884_nl, nor_713_nl, fsm_output[0]);
  assign nand_107_nl = ~((fsm_output[6]) & mux_885_nl);
  assign or_1174_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[3]) | nand_353_cse;
  assign or_1172_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b10010) | (fsm_output[7]);
  assign mux_881_nl = MUX_s_1_2_2(or_1174_nl, or_1172_nl, fsm_output[4]);
  assign or_1171_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | mux_818_cse;
  assign mux_882_nl = MUX_s_1_2_2(mux_881_nl, or_1171_nl, fsm_output[0]);
  assign or_1175_nl = (fsm_output[6]) | mux_882_nl;
  assign mux_886_nl = MUX_s_1_2_2(nand_107_nl, or_1175_nl, fsm_output[3]);
  assign or_2262_nl = (fsm_output[5]) | mux_886_nl;
  assign mux_894_nl = MUX_s_1_2_2(nand_488_nl, or_2262_nl, fsm_output[2]);
  assign vec_rsc_0_18_i_we_d_pff = ~(mux_894_nl | (fsm_output[1]));
  assign nor_698_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b10010) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_699_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_908_nl = MUX_s_1_2_2(nor_698_nl, nor_699_nl, fsm_output[0]);
  assign nor_700_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_906_cse);
  assign nor_701_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b10010) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_702_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b10010) | (fsm_output[7:6]!=2'b10));
  assign nor_703_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b10010) | (fsm_output[7:6]!=2'b00));
  assign mux_902_nl = MUX_s_1_2_2(nor_702_nl, nor_703_nl, fsm_output[4]);
  assign mux_903_nl = MUX_s_1_2_2(nor_701_nl, mux_902_nl, fsm_output[3]);
  assign mux_907_nl = MUX_s_1_2_2(nor_700_nl, mux_903_nl, fsm_output[0]);
  assign mux_909_nl = MUX_s_1_2_2(mux_908_nl, mux_907_nl, fsm_output[5]);
  assign or_1208_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b10010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_1206_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b10010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_899_nl = MUX_s_1_2_2(or_1208_nl, or_1206_nl, fsm_output[4]);
  assign or_1205_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b10010) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_1203_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b10010) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_898_nl = MUX_s_1_2_2(or_1205_nl, or_1203_nl, fsm_output[4]);
  assign mux_900_nl = MUX_s_1_2_2(mux_899_nl, mux_898_nl, fsm_output[3]);
  assign or_1202_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b10010) | nand_443_cse;
  assign or_1200_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b10010) | (fsm_output[7:6]!=2'b01);
  assign mux_896_nl = MUX_s_1_2_2(or_1202_nl, or_1200_nl, fsm_output[4]);
  assign or_1199_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b10010) | (fsm_output[7:6]!=2'b10);
  assign or_1197_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b10010) | (fsm_output[7:6]!=2'b00);
  assign mux_895_nl = MUX_s_1_2_2(or_1199_nl, or_1197_nl, fsm_output[4]);
  assign mux_897_nl = MUX_s_1_2_2(mux_896_nl, mux_895_nl, fsm_output[3]);
  assign mux_901_nl = MUX_s_1_2_2(mux_900_nl, mux_897_nl, fsm_output[0]);
  assign nor_704_nl = ~((fsm_output[5]) | mux_901_nl);
  assign mux_910_nl = MUX_s_1_2_2(mux_909_nl, nor_704_nl, fsm_output[2]);
  assign vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d = mux_910_nl & (fsm_output[1]);
  assign nor_686_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:1]!=3'b001) | nand_357_cse);
  assign nor_687_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b10011) | (fsm_output[7]));
  assign mux_922_nl = MUX_s_1_2_2(nor_686_nl, nor_687_nl, fsm_output[4]);
  assign nor_688_nl = ~((COMP_LOOP_acc_1_cse_sva[4:2]!=3'b100) | nand_435_cse);
  assign nor_689_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b10011) | (fsm_output[7]));
  assign mux_921_nl = MUX_s_1_2_2(nor_688_nl, nor_689_nl, fsm_output[4]);
  assign mux_923_nl = MUX_s_1_2_2(mux_922_nl, mux_921_nl, fsm_output[0]);
  assign and_385_nl = (fsm_output[6]) & mux_923_nl;
  assign or_1240_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0011) | nand_364_cse;
  assign or_1238_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b10011) | (fsm_output[7]);
  assign mux_919_nl = MUX_s_1_2_2(or_1240_nl, or_1238_nl, fsm_output[4]);
  assign or_1237_nl = (COMP_LOOP_acc_1_cse_6_sva[4:1]!=4'b1001) | nand_447_cse;
  assign or_1235_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b10011) | (fsm_output[7]);
  assign mux_918_nl = MUX_s_1_2_2(or_1237_nl, or_1235_nl, fsm_output[4]);
  assign mux_920_nl = MUX_s_1_2_2(mux_919_nl, mux_918_nl, fsm_output[0]);
  assign nor_690_nl = ~((fsm_output[6]) | mux_920_nl);
  assign mux_924_nl = MUX_s_1_2_2(and_385_nl, nor_690_nl, fsm_output[3]);
  assign nand_487_nl = ~((fsm_output[5]) & mux_924_nl);
  assign nor_692_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:2]!=3'b100) | nand_437_cse);
  assign nor_693_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b10011) | (fsm_output[7]));
  assign mux_915_nl = MUX_s_1_2_2(nor_692_nl, nor_693_nl, fsm_output[4]);
  assign nor_694_nl = ~((COMP_LOOP_acc_14_psp_sva[3:1]!=3'b100) | nand_441_cse);
  assign nor_695_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1001) | (fsm_output[7]));
  assign mux_914_nl = MUX_s_1_2_2(nor_694_nl, nor_695_nl, fsm_output[4]);
  assign and_386_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_914_nl;
  assign mux_916_nl = MUX_s_1_2_2(mux_915_nl, and_386_nl, fsm_output[0]);
  assign nand_113_nl = ~((fsm_output[6]) & mux_916_nl);
  assign or_1226_nl = (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[0])) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[3]) | nand_353_cse;
  assign or_1224_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b10011) | (fsm_output[7]);
  assign mux_912_nl = MUX_s_1_2_2(or_1226_nl, or_1224_nl, fsm_output[4]);
  assign nand_111_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & mux_849_cse);
  assign mux_913_nl = MUX_s_1_2_2(mux_912_nl, nand_111_nl, fsm_output[0]);
  assign or_1227_nl = (fsm_output[6]) | mux_913_nl;
  assign mux_917_nl = MUX_s_1_2_2(nand_113_nl, or_1227_nl, fsm_output[3]);
  assign or_2261_nl = (fsm_output[5]) | mux_917_nl;
  assign mux_925_nl = MUX_s_1_2_2(nand_487_nl, or_2261_nl, fsm_output[2]);
  assign vec_rsc_0_19_i_we_d_pff = ~(mux_925_nl | (fsm_output[1]));
  assign nor_680_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b10011) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_681_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_939_nl = MUX_s_1_2_2(nor_680_nl, nor_681_nl, fsm_output[0]);
  assign and_383_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (~ mux_906_cse);
  assign nor_682_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b10011) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_683_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b10011) | (fsm_output[7:6]!=2'b10));
  assign nor_684_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b10011) | (fsm_output[7:6]!=2'b00));
  assign mux_933_nl = MUX_s_1_2_2(nor_683_nl, nor_684_nl, fsm_output[4]);
  assign mux_934_nl = MUX_s_1_2_2(nor_682_nl, mux_933_nl, fsm_output[3]);
  assign mux_938_nl = MUX_s_1_2_2(and_383_nl, mux_934_nl, fsm_output[0]);
  assign mux_940_nl = MUX_s_1_2_2(mux_939_nl, mux_938_nl, fsm_output[5]);
  assign or_1259_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b10011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_1257_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b10011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_930_nl = MUX_s_1_2_2(or_1259_nl, or_1257_nl, fsm_output[4]);
  assign or_1256_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b10011) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_1254_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b10011) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_929_nl = MUX_s_1_2_2(or_1256_nl, or_1254_nl, fsm_output[4]);
  assign mux_931_nl = MUX_s_1_2_2(mux_930_nl, mux_929_nl, fsm_output[3]);
  assign or_1253_nl = (COMP_LOOP_acc_10_cse_10_1_sva[3:1]!=3'b001) | nand_356_cse;
  assign or_1251_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b10011) | (fsm_output[7:6]!=2'b01);
  assign mux_927_nl = MUX_s_1_2_2(or_1253_nl, or_1251_nl, fsm_output[4]);
  assign or_1250_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b10011) | (fsm_output[7:6]!=2'b10);
  assign or_1248_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b10011) | (fsm_output[7:6]!=2'b00);
  assign mux_926_nl = MUX_s_1_2_2(or_1250_nl, or_1248_nl, fsm_output[4]);
  assign mux_928_nl = MUX_s_1_2_2(mux_927_nl, mux_926_nl, fsm_output[3]);
  assign mux_932_nl = MUX_s_1_2_2(mux_931_nl, mux_928_nl, fsm_output[0]);
  assign nor_685_nl = ~((fsm_output[5]) | mux_932_nl);
  assign mux_941_nl = MUX_s_1_2_2(mux_940_nl, nor_685_nl, fsm_output[2]);
  assign vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d = mux_941_nl & (fsm_output[1]);
  assign nor_671_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b10100) | (~ (fsm_output[7])));
  assign nor_672_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b10100) | (fsm_output[7]));
  assign mux_953_nl = MUX_s_1_2_2(nor_671_nl, nor_672_nl, fsm_output[4]);
  assign nor_673_nl = ~((COMP_LOOP_acc_1_cse_sva[4:0]!=5'b10100) | (~ (fsm_output[7])));
  assign nor_674_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b10100) | (fsm_output[7]));
  assign mux_952_nl = MUX_s_1_2_2(nor_673_nl, nor_674_nl, fsm_output[4]);
  assign mux_954_nl = MUX_s_1_2_2(mux_953_nl, mux_952_nl, fsm_output[0]);
  assign and_382_nl = (fsm_output[6]) & mux_954_nl;
  assign or_1293_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0100) | nand_364_cse;
  assign or_1291_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b10100) | (fsm_output[7]);
  assign mux_950_nl = MUX_s_1_2_2(or_1293_nl, or_1291_nl, fsm_output[4]);
  assign or_1290_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b10100) | (~ (fsm_output[7]));
  assign or_1288_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b10100) | (fsm_output[7]);
  assign mux_949_nl = MUX_s_1_2_2(or_1290_nl, or_1288_nl, fsm_output[4]);
  assign mux_951_nl = MUX_s_1_2_2(mux_950_nl, mux_949_nl, fsm_output[0]);
  assign nor_675_nl = ~((fsm_output[6]) | mux_951_nl);
  assign mux_955_nl = MUX_s_1_2_2(and_382_nl, nor_675_nl, fsm_output[3]);
  assign nand_486_nl = ~((fsm_output[5]) & mux_955_nl);
  assign nor_677_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b10100) | (~ (fsm_output[7])));
  assign nor_678_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b10100) | (fsm_output[7]));
  assign mux_946_nl = MUX_s_1_2_2(nor_677_nl, nor_678_nl, fsm_output[4]);
  assign or_1282_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b1010) | (~ (fsm_output[7]));
  assign or_1280_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1010) | (fsm_output[7]);
  assign mux_945_nl = MUX_s_1_2_2(or_1282_nl, or_1280_nl, fsm_output[4]);
  assign nor_679_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_945_nl);
  assign mux_947_nl = MUX_s_1_2_2(mux_946_nl, nor_679_nl, fsm_output[0]);
  assign nand_118_nl = ~((fsm_output[6]) & mux_947_nl);
  assign or_1278_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b10100) | (~ (fsm_output[7]));
  assign or_1276_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b10100) | (fsm_output[7]);
  assign mux_943_nl = MUX_s_1_2_2(or_1278_nl, or_1276_nl, fsm_output[4]);
  assign or_1275_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | mux_942_cse;
  assign mux_944_nl = MUX_s_1_2_2(mux_943_nl, or_1275_nl, fsm_output[0]);
  assign or_1279_nl = (fsm_output[6]) | mux_944_nl;
  assign mux_948_nl = MUX_s_1_2_2(nand_118_nl, or_1279_nl, fsm_output[3]);
  assign or_2260_nl = (fsm_output[5]) | mux_948_nl;
  assign mux_956_nl = MUX_s_1_2_2(nand_486_nl, or_2260_nl, fsm_output[2]);
  assign vec_rsc_0_20_i_we_d_pff = ~(mux_956_nl | (fsm_output[1]));
  assign nor_664_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b10100) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_665_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_970_nl = MUX_s_1_2_2(nor_664_nl, nor_665_nl, fsm_output[0]);
  assign nor_666_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_968_cse);
  assign nor_667_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b10100) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_668_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b10100) | (fsm_output[7:6]!=2'b10));
  assign nor_669_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b10100) | (fsm_output[7:6]!=2'b00));
  assign mux_964_nl = MUX_s_1_2_2(nor_668_nl, nor_669_nl, fsm_output[4]);
  assign mux_965_nl = MUX_s_1_2_2(nor_667_nl, mux_964_nl, fsm_output[3]);
  assign mux_969_nl = MUX_s_1_2_2(nor_666_nl, mux_965_nl, fsm_output[0]);
  assign mux_971_nl = MUX_s_1_2_2(mux_970_nl, mux_969_nl, fsm_output[5]);
  assign or_1312_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b10100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_1310_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b10100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_961_nl = MUX_s_1_2_2(or_1312_nl, or_1310_nl, fsm_output[4]);
  assign or_1309_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b10100) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_1307_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b10100) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_960_nl = MUX_s_1_2_2(or_1309_nl, or_1307_nl, fsm_output[4]);
  assign mux_962_nl = MUX_s_1_2_2(mux_961_nl, mux_960_nl, fsm_output[3]);
  assign or_1306_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b10100) | nand_443_cse;
  assign or_1304_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b10100) | (fsm_output[7:6]!=2'b01);
  assign mux_958_nl = MUX_s_1_2_2(or_1306_nl, or_1304_nl, fsm_output[4]);
  assign or_1303_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b10100) | (fsm_output[7:6]!=2'b10);
  assign or_1301_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b10100) | (fsm_output[7:6]!=2'b00);
  assign mux_957_nl = MUX_s_1_2_2(or_1303_nl, or_1301_nl, fsm_output[4]);
  assign mux_959_nl = MUX_s_1_2_2(mux_958_nl, mux_957_nl, fsm_output[3]);
  assign mux_963_nl = MUX_s_1_2_2(mux_962_nl, mux_959_nl, fsm_output[0]);
  assign nor_670_nl = ~((fsm_output[5]) | mux_963_nl);
  assign mux_972_nl = MUX_s_1_2_2(mux_971_nl, nor_670_nl, fsm_output[2]);
  assign vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d = mux_972_nl & (fsm_output[1]);
  assign nor_652_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:1]!=3'b010) | nand_357_cse);
  assign nor_653_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b10101) | (fsm_output[7]));
  assign mux_984_nl = MUX_s_1_2_2(nor_652_nl, nor_653_nl, fsm_output[4]);
  assign nor_654_nl = ~((COMP_LOOP_acc_1_cse_sva[4:1]!=4'b1010) | nand_446_cse);
  assign nor_655_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b10101) | (fsm_output[7]));
  assign mux_983_nl = MUX_s_1_2_2(nor_654_nl, nor_655_nl, fsm_output[4]);
  assign mux_985_nl = MUX_s_1_2_2(mux_984_nl, mux_983_nl, fsm_output[0]);
  assign and_379_nl = (fsm_output[6]) & mux_985_nl;
  assign or_1344_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0101) | nand_364_cse;
  assign or_1342_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b10101) | (fsm_output[7]);
  assign mux_981_nl = MUX_s_1_2_2(or_1344_nl, or_1342_nl, fsm_output[4]);
  assign or_1341_nl = (COMP_LOOP_acc_1_cse_6_sva[4:1]!=4'b1010) | nand_447_cse;
  assign or_1339_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b10101) | (fsm_output[7]);
  assign mux_980_nl = MUX_s_1_2_2(or_1341_nl, or_1339_nl, fsm_output[4]);
  assign mux_982_nl = MUX_s_1_2_2(mux_981_nl, mux_980_nl, fsm_output[0]);
  assign nor_656_nl = ~((fsm_output[6]) | mux_982_nl);
  assign mux_986_nl = MUX_s_1_2_2(and_379_nl, nor_656_nl, fsm_output[3]);
  assign nand_485_nl = ~((fsm_output[5]) & mux_986_nl);
  assign nor_658_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:1]!=4'b1010) | nand_448_cse);
  assign nor_659_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b10101) | (fsm_output[7]));
  assign mux_977_nl = MUX_s_1_2_2(nor_658_nl, nor_659_nl, fsm_output[4]);
  assign nor_660_nl = ~((COMP_LOOP_acc_14_psp_sva[3:0]!=4'b1010) | (~ (fsm_output[7])));
  assign nor_661_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1010) | (fsm_output[7]));
  assign mux_976_nl = MUX_s_1_2_2(nor_660_nl, nor_661_nl, fsm_output[4]);
  assign and_380_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_976_nl;
  assign mux_978_nl = MUX_s_1_2_2(mux_977_nl, and_380_nl, fsm_output[0]);
  assign nand_124_nl = ~((fsm_output[6]) & mux_978_nl);
  assign or_1330_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b10101) | (~ (fsm_output[7]));
  assign or_1328_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b10101) | (fsm_output[7]);
  assign mux_974_nl = MUX_s_1_2_2(or_1330_nl, or_1328_nl, fsm_output[4]);
  assign nand_122_nl = ~(nor_98_cse & mux_973_cse);
  assign mux_975_nl = MUX_s_1_2_2(mux_974_nl, nand_122_nl, fsm_output[0]);
  assign or_1331_nl = (fsm_output[6]) | mux_975_nl;
  assign mux_979_nl = MUX_s_1_2_2(nand_124_nl, or_1331_nl, fsm_output[3]);
  assign or_2259_nl = (fsm_output[5]) | mux_979_nl;
  assign mux_987_nl = MUX_s_1_2_2(nand_485_nl, or_2259_nl, fsm_output[2]);
  assign vec_rsc_0_21_i_we_d_pff = ~(mux_987_nl | (fsm_output[1]));
  assign nor_646_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b10101) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_647_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_1001_nl = MUX_s_1_2_2(nor_646_nl, nor_647_nl, fsm_output[0]);
  assign and_377_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (~ mux_968_cse);
  assign nor_648_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b10101) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_649_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b10101) | (fsm_output[7:6]!=2'b10));
  assign nor_650_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b10101) | (fsm_output[7:6]!=2'b00));
  assign mux_995_nl = MUX_s_1_2_2(nor_649_nl, nor_650_nl, fsm_output[4]);
  assign mux_996_nl = MUX_s_1_2_2(nor_648_nl, mux_995_nl, fsm_output[3]);
  assign mux_1000_nl = MUX_s_1_2_2(and_377_nl, mux_996_nl, fsm_output[0]);
  assign mux_1002_nl = MUX_s_1_2_2(mux_1001_nl, mux_1000_nl, fsm_output[5]);
  assign or_1363_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b10101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_1361_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b10101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_992_nl = MUX_s_1_2_2(or_1363_nl, or_1361_nl, fsm_output[4]);
  assign or_1360_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b10101) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_1358_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b10101) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_991_nl = MUX_s_1_2_2(or_1360_nl, or_1358_nl, fsm_output[4]);
  assign mux_993_nl = MUX_s_1_2_2(mux_992_nl, mux_991_nl, fsm_output[3]);
  assign or_1357_nl = (COMP_LOOP_acc_10_cse_10_1_sva[3:1]!=3'b010) | nand_356_cse;
  assign or_1355_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b10101) | (fsm_output[7:6]!=2'b01);
  assign mux_989_nl = MUX_s_1_2_2(or_1357_nl, or_1355_nl, fsm_output[4]);
  assign or_1354_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b10101) | (fsm_output[7:6]!=2'b10);
  assign or_1352_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b10101) | (fsm_output[7:6]!=2'b00);
  assign mux_988_nl = MUX_s_1_2_2(or_1354_nl, or_1352_nl, fsm_output[4]);
  assign mux_990_nl = MUX_s_1_2_2(mux_989_nl, mux_988_nl, fsm_output[3]);
  assign mux_994_nl = MUX_s_1_2_2(mux_993_nl, mux_990_nl, fsm_output[0]);
  assign nor_651_nl = ~((fsm_output[5]) | mux_994_nl);
  assign mux_1003_nl = MUX_s_1_2_2(mux_1002_nl, nor_651_nl, fsm_output[2]);
  assign vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1003_nl & (fsm_output[1]);
  assign nor_637_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b10110) | (~ (fsm_output[7])));
  assign nor_638_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b10110) | (fsm_output[7]));
  assign mux_1015_nl = MUX_s_1_2_2(nor_637_nl, nor_638_nl, fsm_output[4]);
  assign nor_639_nl = ~((COMP_LOOP_acc_1_cse_sva[4:0]!=5'b10110) | (~ (fsm_output[7])));
  assign nor_640_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b10110) | (fsm_output[7]));
  assign mux_1014_nl = MUX_s_1_2_2(nor_639_nl, nor_640_nl, fsm_output[4]);
  assign mux_1016_nl = MUX_s_1_2_2(mux_1015_nl, mux_1014_nl, fsm_output[0]);
  assign and_376_nl = (fsm_output[6]) & mux_1016_nl;
  assign or_1397_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]!=4'b0110) | nand_364_cse;
  assign or_1395_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b10110) | (fsm_output[7]);
  assign mux_1012_nl = MUX_s_1_2_2(or_1397_nl, or_1395_nl, fsm_output[4]);
  assign or_1394_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b10110) | (~ (fsm_output[7]));
  assign or_1392_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b10110) | (fsm_output[7]);
  assign mux_1011_nl = MUX_s_1_2_2(or_1394_nl, or_1392_nl, fsm_output[4]);
  assign mux_1013_nl = MUX_s_1_2_2(mux_1012_nl, mux_1011_nl, fsm_output[0]);
  assign nor_641_nl = ~((fsm_output[6]) | mux_1013_nl);
  assign mux_1017_nl = MUX_s_1_2_2(and_376_nl, nor_641_nl, fsm_output[3]);
  assign nand_484_nl = ~((fsm_output[5]) & mux_1017_nl);
  assign nor_643_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b10110) | (~ (fsm_output[7])));
  assign nor_644_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b10110) | (fsm_output[7]));
  assign mux_1008_nl = MUX_s_1_2_2(nor_643_nl, nor_644_nl, fsm_output[4]);
  assign or_1386_nl = (COMP_LOOP_acc_14_psp_sva[3:2]!=2'b10) | nand_423_cse;
  assign or_1384_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1011) | (fsm_output[7]);
  assign mux_1007_nl = MUX_s_1_2_2(or_1386_nl, or_1384_nl, fsm_output[4]);
  assign nor_645_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1007_nl);
  assign mux_1009_nl = MUX_s_1_2_2(mux_1008_nl, nor_645_nl, fsm_output[0]);
  assign nand_129_nl = ~((fsm_output[6]) & mux_1009_nl);
  assign or_1382_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[2]))
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[3]) | nand_353_cse;
  assign or_1380_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b10110) | (fsm_output[7]);
  assign mux_1005_nl = MUX_s_1_2_2(or_1382_nl, or_1380_nl, fsm_output[4]);
  assign or_1379_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | mux_942_cse;
  assign mux_1006_nl = MUX_s_1_2_2(mux_1005_nl, or_1379_nl, fsm_output[0]);
  assign or_1383_nl = (fsm_output[6]) | mux_1006_nl;
  assign mux_1010_nl = MUX_s_1_2_2(nand_129_nl, or_1383_nl, fsm_output[3]);
  assign or_2258_nl = (fsm_output[5]) | mux_1010_nl;
  assign mux_1018_nl = MUX_s_1_2_2(nand_484_nl, or_2258_nl, fsm_output[2]);
  assign vec_rsc_0_22_i_we_d_pff = ~(mux_1018_nl | (fsm_output[1]));
  assign nor_630_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b10110) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_631_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_1032_nl = MUX_s_1_2_2(nor_630_nl, nor_631_nl, fsm_output[0]);
  assign nor_632_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1030_cse);
  assign nor_633_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b10110) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_634_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b10110) | (fsm_output[7:6]!=2'b10));
  assign nor_635_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b10110) | (fsm_output[7:6]!=2'b00));
  assign mux_1026_nl = MUX_s_1_2_2(nor_634_nl, nor_635_nl, fsm_output[4]);
  assign mux_1027_nl = MUX_s_1_2_2(nor_633_nl, mux_1026_nl, fsm_output[3]);
  assign mux_1031_nl = MUX_s_1_2_2(nor_632_nl, mux_1027_nl, fsm_output[0]);
  assign mux_1033_nl = MUX_s_1_2_2(mux_1032_nl, mux_1031_nl, fsm_output[5]);
  assign or_1416_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b10110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_1414_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b10110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_1023_nl = MUX_s_1_2_2(or_1416_nl, or_1414_nl, fsm_output[4]);
  assign or_1413_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b10110) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_1411_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b10110) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_1022_nl = MUX_s_1_2_2(or_1413_nl, or_1411_nl, fsm_output[4]);
  assign mux_1024_nl = MUX_s_1_2_2(mux_1023_nl, mux_1022_nl, fsm_output[3]);
  assign or_1410_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b10110) | nand_443_cse;
  assign or_1408_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b10110) | (fsm_output[7:6]!=2'b01);
  assign mux_1020_nl = MUX_s_1_2_2(or_1410_nl, or_1408_nl, fsm_output[4]);
  assign or_1407_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b10110) | (fsm_output[7:6]!=2'b10);
  assign or_1405_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b10110) | (fsm_output[7:6]!=2'b00);
  assign mux_1019_nl = MUX_s_1_2_2(or_1407_nl, or_1405_nl, fsm_output[4]);
  assign mux_1021_nl = MUX_s_1_2_2(mux_1020_nl, mux_1019_nl, fsm_output[3]);
  assign mux_1025_nl = MUX_s_1_2_2(mux_1024_nl, mux_1021_nl, fsm_output[0]);
  assign nor_636_nl = ~((fsm_output[5]) | mux_1025_nl);
  assign mux_1034_nl = MUX_s_1_2_2(mux_1033_nl, nor_636_nl, fsm_output[2]);
  assign vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1034_nl & (fsm_output[1]);
  assign nor_618_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[3:1]!=3'b011) | nand_357_cse);
  assign nor_619_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b10111) | (fsm_output[7]));
  assign mux_1046_nl = MUX_s_1_2_2(nor_618_nl, nor_619_nl, fsm_output[4]);
  assign nor_620_nl = ~((COMP_LOOP_acc_1_cse_sva[4:3]!=2'b10) | nand_417_cse);
  assign nor_621_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b10111) | (fsm_output[7]));
  assign mux_1045_nl = MUX_s_1_2_2(nor_620_nl, nor_621_nl, fsm_output[4]);
  assign mux_1047_nl = MUX_s_1_2_2(mux_1046_nl, mux_1045_nl, fsm_output[0]);
  assign and_373_nl = (fsm_output[6]) & mux_1047_nl;
  assign or_1448_nl = (~((COMP_LOOP_acc_10_cse_10_1_6_sva[3:0]==4'b0111))) | nand_364_cse;
  assign or_1446_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b10111) | (fsm_output[7]);
  assign mux_1043_nl = MUX_s_1_2_2(or_1448_nl, or_1446_nl, fsm_output[4]);
  assign or_1445_nl = (~((COMP_LOOP_acc_1_cse_6_sva[4:1]==4'b1011))) | nand_447_cse;
  assign or_1443_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b10111) | (fsm_output[7]);
  assign mux_1042_nl = MUX_s_1_2_2(or_1445_nl, or_1443_nl, fsm_output[4]);
  assign mux_1044_nl = MUX_s_1_2_2(mux_1043_nl, mux_1042_nl, fsm_output[0]);
  assign nor_622_nl = ~((fsm_output[6]) | mux_1044_nl);
  assign mux_1048_nl = MUX_s_1_2_2(and_373_nl, nor_622_nl, fsm_output[3]);
  assign nand_483_nl = ~((fsm_output[5]) & mux_1048_nl);
  assign nor_624_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:3]!=2'b10) | nand_419_cse);
  assign nor_625_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b10111) | (fsm_output[7]));
  assign mux_1039_nl = MUX_s_1_2_2(nor_624_nl, nor_625_nl, fsm_output[4]);
  assign nor_626_nl = ~((COMP_LOOP_acc_14_psp_sva[3:2]!=2'b10) | nand_423_cse);
  assign nor_627_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1011) | (fsm_output[7]));
  assign mux_1038_nl = MUX_s_1_2_2(nor_626_nl, nor_627_nl, fsm_output[4]);
  assign and_374_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1038_nl;
  assign mux_1040_nl = MUX_s_1_2_2(mux_1039_nl, and_374_nl, fsm_output[0]);
  assign nand_135_nl = ~((fsm_output[6]) & mux_1040_nl);
  assign or_1434_nl = (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[0])) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[2]))
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[3]) | nand_353_cse;
  assign or_1432_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b10111) | (fsm_output[7]);
  assign mux_1036_nl = MUX_s_1_2_2(or_1434_nl, or_1432_nl, fsm_output[4]);
  assign nand_133_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & mux_973_cse);
  assign mux_1037_nl = MUX_s_1_2_2(mux_1036_nl, nand_133_nl, fsm_output[0]);
  assign or_1435_nl = (fsm_output[6]) | mux_1037_nl;
  assign mux_1041_nl = MUX_s_1_2_2(nand_135_nl, or_1435_nl, fsm_output[3]);
  assign or_2257_nl = (fsm_output[5]) | mux_1041_nl;
  assign mux_1049_nl = MUX_s_1_2_2(nand_483_nl, or_2257_nl, fsm_output[2]);
  assign vec_rsc_0_23_i_we_d_pff = ~(mux_1049_nl | (fsm_output[1]));
  assign nor_613_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b10111) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_614_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_1063_nl = MUX_s_1_2_2(nor_613_nl, nor_614_nl, fsm_output[0]);
  assign and_370_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (~ mux_1030_cse);
  assign and_371_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]==5'b10111) & (fsm_output[4])
      & (fsm_output[6]) & (~ (fsm_output[7]));
  assign and_526_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]==5'b10111) & (fsm_output[7:6]==2'b10);
  assign nor_616_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b10111) | (fsm_output[7:6]!=2'b00));
  assign mux_1057_nl = MUX_s_1_2_2(and_526_nl, nor_616_nl, fsm_output[4]);
  assign mux_1058_nl = MUX_s_1_2_2(and_371_nl, mux_1057_nl, fsm_output[3]);
  assign mux_1062_nl = MUX_s_1_2_2(and_370_nl, mux_1058_nl, fsm_output[0]);
  assign mux_1064_nl = MUX_s_1_2_2(mux_1063_nl, mux_1062_nl, fsm_output[5]);
  assign or_1467_nl = (~((COMP_LOOP_acc_1_cse_sva[4:0]==5'b10111) & COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm))
      | nand_443_cse;
  assign nand_307_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]==5'b10111) & COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm
      & (fsm_output[7:6]==2'b01));
  assign mux_1054_nl = MUX_s_1_2_2(or_1467_nl, nand_307_nl, fsm_output[4]);
  assign nand_514_nl = ~((COMP_LOOP_acc_1_cse_6_sva[4:0]==5'b10111) & COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[7:6]==2'b10));
  assign or_1462_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b10111) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_1053_nl = MUX_s_1_2_2(nand_514_nl, or_1462_nl, fsm_output[4]);
  assign mux_1055_nl = MUX_s_1_2_2(mux_1054_nl, mux_1053_nl, fsm_output[3]);
  assign or_1461_nl = (COMP_LOOP_acc_10_cse_10_1_sva[3:1]!=3'b011) | nand_356_cse;
  assign nand_310_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]==5'b10111) & (fsm_output[7:6]==2'b01));
  assign mux_1051_nl = MUX_s_1_2_2(or_1461_nl, nand_310_nl, fsm_output[4]);
  assign nand_468_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]==5'b10111) & (fsm_output[7:6]==2'b10));
  assign or_1456_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b10111) | (fsm_output[7:6]!=2'b00);
  assign mux_1050_nl = MUX_s_1_2_2(nand_468_nl, or_1456_nl, fsm_output[4]);
  assign mux_1052_nl = MUX_s_1_2_2(mux_1051_nl, mux_1050_nl, fsm_output[3]);
  assign mux_1056_nl = MUX_s_1_2_2(mux_1055_nl, mux_1052_nl, fsm_output[0]);
  assign nor_617_nl = ~((fsm_output[5]) | mux_1056_nl);
  assign mux_1065_nl = MUX_s_1_2_2(mux_1064_nl, nor_617_nl, fsm_output[2]);
  assign vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1065_nl & (fsm_output[1]);
  assign nor_604_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b11000) | (~ (fsm_output[7])));
  assign nor_605_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b11000) | (fsm_output[7]));
  assign mux_1077_nl = MUX_s_1_2_2(nor_604_nl, nor_605_nl, fsm_output[4]);
  assign nor_606_nl = ~((COMP_LOOP_acc_1_cse_sva[4:0]!=5'b11000) | (~ (fsm_output[7])));
  assign nor_607_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b11000) | (fsm_output[7]));
  assign mux_1076_nl = MUX_s_1_2_2(nor_606_nl, nor_607_nl, fsm_output[4]);
  assign mux_1078_nl = MUX_s_1_2_2(mux_1077_nl, mux_1076_nl, fsm_output[0]);
  assign and_369_nl = (fsm_output[6]) & mux_1078_nl;
  assign or_1500_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[2:0]!=3'b000) | nand_302_cse;
  assign or_1498_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b11000) | (fsm_output[7]);
  assign mux_1074_nl = MUX_s_1_2_2(or_1500_nl, or_1498_nl, fsm_output[4]);
  assign or_1497_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b11000) | (~ (fsm_output[7]));
  assign or_1495_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b11000) | (fsm_output[7]);
  assign mux_1073_nl = MUX_s_1_2_2(or_1497_nl, or_1495_nl, fsm_output[4]);
  assign mux_1075_nl = MUX_s_1_2_2(mux_1074_nl, mux_1073_nl, fsm_output[0]);
  assign nor_608_nl = ~((fsm_output[6]) | mux_1075_nl);
  assign mux_1079_nl = MUX_s_1_2_2(and_369_nl, nor_608_nl, fsm_output[3]);
  assign nand_482_nl = ~((fsm_output[5]) & mux_1079_nl);
  assign nor_610_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b11000) | (~ (fsm_output[7])));
  assign nor_611_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b11000) | (fsm_output[7]));
  assign mux_1070_nl = MUX_s_1_2_2(nor_610_nl, nor_611_nl, fsm_output[4]);
  assign or_1489_nl = (COMP_LOOP_acc_14_psp_sva[3:0]!=4'b1100) | (~ (fsm_output[7]));
  assign or_1487_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1100) | (fsm_output[7]);
  assign mux_1069_nl = MUX_s_1_2_2(or_1489_nl, or_1487_nl, fsm_output[4]);
  assign nor_612_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1069_nl);
  assign mux_1071_nl = MUX_s_1_2_2(mux_1070_nl, nor_612_nl, fsm_output[0]);
  assign nand_140_nl = ~((fsm_output[6]) & mux_1071_nl);
  assign or_1485_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b11000) | (~ (fsm_output[7]));
  assign or_1483_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b11000) | (fsm_output[7]);
  assign mux_1067_nl = MUX_s_1_2_2(or_1485_nl, or_1483_nl, fsm_output[4]);
  assign or_1482_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | mux_1066_cse;
  assign mux_1068_nl = MUX_s_1_2_2(mux_1067_nl, or_1482_nl, fsm_output[0]);
  assign or_1486_nl = (fsm_output[6]) | mux_1068_nl;
  assign mux_1072_nl = MUX_s_1_2_2(nand_140_nl, or_1486_nl, fsm_output[3]);
  assign or_2256_nl = (fsm_output[5]) | mux_1072_nl;
  assign mux_1080_nl = MUX_s_1_2_2(nand_482_nl, or_2256_nl, fsm_output[2]);
  assign vec_rsc_0_24_i_we_d_pff = ~(mux_1080_nl | (fsm_output[1]));
  assign nor_597_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b11000) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_598_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_1094_nl = MUX_s_1_2_2(nor_597_nl, nor_598_nl, fsm_output[0]);
  assign nor_599_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1092_cse);
  assign nor_600_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b11000) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_601_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b11000) | (fsm_output[7:6]!=2'b10));
  assign nor_602_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b11000) | (fsm_output[7:6]!=2'b00));
  assign mux_1088_nl = MUX_s_1_2_2(nor_601_nl, nor_602_nl, fsm_output[4]);
  assign mux_1089_nl = MUX_s_1_2_2(nor_600_nl, mux_1088_nl, fsm_output[3]);
  assign mux_1093_nl = MUX_s_1_2_2(nor_599_nl, mux_1089_nl, fsm_output[0]);
  assign mux_1095_nl = MUX_s_1_2_2(mux_1094_nl, mux_1093_nl, fsm_output[5]);
  assign or_1519_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b11000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_1517_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b11000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_1085_nl = MUX_s_1_2_2(or_1519_nl, or_1517_nl, fsm_output[4]);
  assign or_1516_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b11000) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_1514_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b11000) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_1084_nl = MUX_s_1_2_2(or_1516_nl, or_1514_nl, fsm_output[4]);
  assign mux_1086_nl = MUX_s_1_2_2(mux_1085_nl, mux_1084_nl, fsm_output[3]);
  assign or_1513_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b11000) | nand_443_cse;
  assign or_1511_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b11000) | (fsm_output[7:6]!=2'b01);
  assign mux_1082_nl = MUX_s_1_2_2(or_1513_nl, or_1511_nl, fsm_output[4]);
  assign or_1510_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b11000) | (fsm_output[7:6]!=2'b10);
  assign or_1508_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b11000) | (fsm_output[7:6]!=2'b00);
  assign mux_1081_nl = MUX_s_1_2_2(or_1510_nl, or_1508_nl, fsm_output[4]);
  assign mux_1083_nl = MUX_s_1_2_2(mux_1082_nl, mux_1081_nl, fsm_output[3]);
  assign mux_1087_nl = MUX_s_1_2_2(mux_1086_nl, mux_1083_nl, fsm_output[0]);
  assign nor_603_nl = ~((fsm_output[5]) | mux_1087_nl);
  assign mux_1096_nl = MUX_s_1_2_2(mux_1095_nl, nor_603_nl, fsm_output[2]);
  assign vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1096_nl & (fsm_output[1]);
  assign nor_585_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[2:1]!=2'b00) | nand_294_cse);
  assign nor_586_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b11001) | (fsm_output[7]));
  assign mux_1108_nl = MUX_s_1_2_2(nor_585_nl, nor_586_nl, fsm_output[4]);
  assign nor_587_nl = ~((COMP_LOOP_acc_1_cse_sva[4:1]!=4'b1100) | nand_446_cse);
  assign nor_588_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b11001) | (fsm_output[7]));
  assign mux_1107_nl = MUX_s_1_2_2(nor_587_nl, nor_588_nl, fsm_output[4]);
  assign mux_1109_nl = MUX_s_1_2_2(mux_1108_nl, mux_1107_nl, fsm_output[0]);
  assign and_366_nl = (fsm_output[6]) & mux_1109_nl;
  assign or_1550_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[2:0]!=3'b001) | nand_302_cse;
  assign or_1548_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b11001) | (fsm_output[7]);
  assign mux_1105_nl = MUX_s_1_2_2(or_1550_nl, or_1548_nl, fsm_output[4]);
  assign or_1547_nl = (COMP_LOOP_acc_1_cse_6_sva[2:1]!=2'b00) | nand_297_cse;
  assign or_1545_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b11001) | (fsm_output[7]);
  assign mux_1104_nl = MUX_s_1_2_2(or_1547_nl, or_1545_nl, fsm_output[4]);
  assign mux_1106_nl = MUX_s_1_2_2(mux_1105_nl, mux_1104_nl, fsm_output[0]);
  assign nor_589_nl = ~((fsm_output[6]) | mux_1106_nl);
  assign mux_1110_nl = MUX_s_1_2_2(and_366_nl, nor_589_nl, fsm_output[3]);
  assign nand_481_nl = ~((fsm_output[5]) & mux_1110_nl);
  assign nor_591_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:1]!=4'b1100) | nand_448_cse);
  assign nor_592_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b11001) | (fsm_output[7]));
  assign mux_1101_nl = MUX_s_1_2_2(nor_591_nl, nor_592_nl, fsm_output[4]);
  assign nor_593_nl = ~((COMP_LOOP_acc_14_psp_sva[3:0]!=4'b1100) | (~ (fsm_output[7])));
  assign nor_594_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1100) | (fsm_output[7]));
  assign mux_1100_nl = MUX_s_1_2_2(nor_593_nl, nor_594_nl, fsm_output[4]);
  assign and_367_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1100_nl;
  assign mux_1102_nl = MUX_s_1_2_2(mux_1101_nl, and_367_nl, fsm_output[0]);
  assign nand_146_nl = ~((fsm_output[6]) & mux_1102_nl);
  assign or_1536_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b11001) | (~ (fsm_output[7]));
  assign or_1534_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b11001) | (fsm_output[7]);
  assign mux_1098_nl = MUX_s_1_2_2(or_1536_nl, or_1534_nl, fsm_output[4]);
  assign nand_144_nl = ~(nor_98_cse & mux_1097_cse);
  assign mux_1099_nl = MUX_s_1_2_2(mux_1098_nl, nand_144_nl, fsm_output[0]);
  assign or_1537_nl = (fsm_output[6]) | mux_1099_nl;
  assign mux_1103_nl = MUX_s_1_2_2(nand_146_nl, or_1537_nl, fsm_output[3]);
  assign or_2255_nl = (fsm_output[5]) | mux_1103_nl;
  assign mux_1111_nl = MUX_s_1_2_2(nand_481_nl, or_2255_nl, fsm_output[2]);
  assign vec_rsc_0_25_i_we_d_pff = ~(mux_1111_nl | (fsm_output[1]));
  assign nor_579_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b11001) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_580_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_1125_nl = MUX_s_1_2_2(nor_579_nl, nor_580_nl, fsm_output[0]);
  assign and_364_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (~ mux_1092_cse);
  assign nor_581_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b11001) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_582_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b11001) | (fsm_output[7:6]!=2'b10));
  assign nor_583_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b11001) | (fsm_output[7:6]!=2'b00));
  assign mux_1119_nl = MUX_s_1_2_2(nor_582_nl, nor_583_nl, fsm_output[4]);
  assign mux_1120_nl = MUX_s_1_2_2(nor_581_nl, mux_1119_nl, fsm_output[3]);
  assign mux_1124_nl = MUX_s_1_2_2(and_364_nl, mux_1120_nl, fsm_output[0]);
  assign mux_1126_nl = MUX_s_1_2_2(mux_1125_nl, mux_1124_nl, fsm_output[5]);
  assign or_1569_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b11001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_1567_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b11001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_1116_nl = MUX_s_1_2_2(or_1569_nl, or_1567_nl, fsm_output[4]);
  assign or_1566_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b11001) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_1564_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b11001) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_1115_nl = MUX_s_1_2_2(or_1566_nl, or_1564_nl, fsm_output[4]);
  assign mux_1117_nl = MUX_s_1_2_2(mux_1116_nl, mux_1115_nl, fsm_output[3]);
  assign or_1563_nl = (COMP_LOOP_acc_10_cse_10_1_sva[2:1]!=2'b00) | nand_293_cse;
  assign or_1561_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b11001) | (fsm_output[7:6]!=2'b01);
  assign mux_1113_nl = MUX_s_1_2_2(or_1563_nl, or_1561_nl, fsm_output[4]);
  assign or_1560_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b11001) | (fsm_output[7:6]!=2'b10);
  assign or_1558_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b11001) | (fsm_output[7:6]!=2'b00);
  assign mux_1112_nl = MUX_s_1_2_2(or_1560_nl, or_1558_nl, fsm_output[4]);
  assign mux_1114_nl = MUX_s_1_2_2(mux_1113_nl, mux_1112_nl, fsm_output[3]);
  assign mux_1118_nl = MUX_s_1_2_2(mux_1117_nl, mux_1114_nl, fsm_output[0]);
  assign nor_584_nl = ~((fsm_output[5]) | mux_1118_nl);
  assign mux_1127_nl = MUX_s_1_2_2(mux_1126_nl, nor_584_nl, fsm_output[2]);
  assign vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1127_nl & (fsm_output[1]);
  assign nor_570_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b11010) | (~ (fsm_output[7])));
  assign nor_571_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b11010) | (fsm_output[7]));
  assign mux_1139_nl = MUX_s_1_2_2(nor_570_nl, nor_571_nl, fsm_output[4]);
  assign nor_572_nl = ~((COMP_LOOP_acc_1_cse_sva[4:0]!=5'b11010) | (~ (fsm_output[7])));
  assign nor_573_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b11010) | (fsm_output[7]));
  assign mux_1138_nl = MUX_s_1_2_2(nor_572_nl, nor_573_nl, fsm_output[4]);
  assign mux_1140_nl = MUX_s_1_2_2(mux_1139_nl, mux_1138_nl, fsm_output[0]);
  assign and_363_nl = (fsm_output[6]) & mux_1140_nl;
  assign or_1602_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[2:0]!=3'b010) | nand_302_cse;
  assign or_1600_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b11010) | (fsm_output[7]);
  assign mux_1136_nl = MUX_s_1_2_2(or_1602_nl, or_1600_nl, fsm_output[4]);
  assign or_1599_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b11010) | (~ (fsm_output[7]));
  assign or_1597_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b11010) | (fsm_output[7]);
  assign mux_1135_nl = MUX_s_1_2_2(or_1599_nl, or_1597_nl, fsm_output[4]);
  assign mux_1137_nl = MUX_s_1_2_2(mux_1136_nl, mux_1135_nl, fsm_output[0]);
  assign nor_574_nl = ~((fsm_output[6]) | mux_1137_nl);
  assign mux_1141_nl = MUX_s_1_2_2(and_363_nl, nor_574_nl, fsm_output[3]);
  assign nand_480_nl = ~((fsm_output[5]) & mux_1141_nl);
  assign nor_576_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b11010) | (~ (fsm_output[7])));
  assign nor_577_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b11010) | (fsm_output[7]));
  assign mux_1132_nl = MUX_s_1_2_2(nor_576_nl, nor_577_nl, fsm_output[4]);
  assign or_1591_nl = (COMP_LOOP_acc_14_psp_sva[3:1]!=3'b110) | nand_441_cse;
  assign or_1589_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1101) | (fsm_output[7]);
  assign mux_1131_nl = MUX_s_1_2_2(or_1591_nl, or_1589_nl, fsm_output[4]);
  assign nor_578_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1131_nl);
  assign mux_1133_nl = MUX_s_1_2_2(mux_1132_nl, nor_578_nl, fsm_output[0]);
  assign nand_151_nl = ~((fsm_output[6]) & mux_1133_nl);
  assign or_1587_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | nand_289_cse;
  assign or_1585_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b11010) | (fsm_output[7]);
  assign mux_1129_nl = MUX_s_1_2_2(or_1587_nl, or_1585_nl, fsm_output[4]);
  assign or_1584_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | mux_1066_cse;
  assign mux_1130_nl = MUX_s_1_2_2(mux_1129_nl, or_1584_nl, fsm_output[0]);
  assign or_1588_nl = (fsm_output[6]) | mux_1130_nl;
  assign mux_1134_nl = MUX_s_1_2_2(nand_151_nl, or_1588_nl, fsm_output[3]);
  assign or_2254_nl = (fsm_output[5]) | mux_1134_nl;
  assign mux_1142_nl = MUX_s_1_2_2(nand_480_nl, or_2254_nl, fsm_output[2]);
  assign vec_rsc_0_26_i_we_d_pff = ~(mux_1142_nl | (fsm_output[1]));
  assign nor_563_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b11010) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_564_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_1156_nl = MUX_s_1_2_2(nor_563_nl, nor_564_nl, fsm_output[0]);
  assign nor_565_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1154_cse);
  assign nor_566_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b11010) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_567_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b11010) | (fsm_output[7:6]!=2'b10));
  assign nor_568_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b11010) | (fsm_output[7:6]!=2'b00));
  assign mux_1150_nl = MUX_s_1_2_2(nor_567_nl, nor_568_nl, fsm_output[4]);
  assign mux_1151_nl = MUX_s_1_2_2(nor_566_nl, mux_1150_nl, fsm_output[3]);
  assign mux_1155_nl = MUX_s_1_2_2(nor_565_nl, mux_1151_nl, fsm_output[0]);
  assign mux_1157_nl = MUX_s_1_2_2(mux_1156_nl, mux_1155_nl, fsm_output[5]);
  assign or_1621_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b11010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_1619_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b11010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_1147_nl = MUX_s_1_2_2(or_1621_nl, or_1619_nl, fsm_output[4]);
  assign or_1618_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b11010) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_1616_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b11010) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_1146_nl = MUX_s_1_2_2(or_1618_nl, or_1616_nl, fsm_output[4]);
  assign mux_1148_nl = MUX_s_1_2_2(mux_1147_nl, mux_1146_nl, fsm_output[3]);
  assign or_1615_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b11010) | nand_443_cse;
  assign or_1613_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b11010) | (fsm_output[7:6]!=2'b01);
  assign mux_1144_nl = MUX_s_1_2_2(or_1615_nl, or_1613_nl, fsm_output[4]);
  assign or_1612_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b11010) | (fsm_output[7:6]!=2'b10);
  assign or_1610_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b11010) | (fsm_output[7:6]!=2'b00);
  assign mux_1143_nl = MUX_s_1_2_2(or_1612_nl, or_1610_nl, fsm_output[4]);
  assign mux_1145_nl = MUX_s_1_2_2(mux_1144_nl, mux_1143_nl, fsm_output[3]);
  assign mux_1149_nl = MUX_s_1_2_2(mux_1148_nl, mux_1145_nl, fsm_output[0]);
  assign nor_569_nl = ~((fsm_output[5]) | mux_1149_nl);
  assign mux_1158_nl = MUX_s_1_2_2(mux_1157_nl, nor_569_nl, fsm_output[2]);
  assign vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1158_nl & (fsm_output[1]);
  assign nor_551_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[2:1]!=2'b01) | nand_294_cse);
  assign nor_552_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b11011) | (fsm_output[7]));
  assign mux_1170_nl = MUX_s_1_2_2(nor_551_nl, nor_552_nl, fsm_output[4]);
  assign nor_553_nl = ~((COMP_LOOP_acc_1_cse_sva[4:2]!=3'b110) | nand_435_cse);
  assign nor_554_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b11011) | (fsm_output[7]));
  assign mux_1169_nl = MUX_s_1_2_2(nor_553_nl, nor_554_nl, fsm_output[4]);
  assign mux_1171_nl = MUX_s_1_2_2(mux_1170_nl, mux_1169_nl, fsm_output[0]);
  assign and_360_nl = (fsm_output[6]) & mux_1171_nl;
  assign or_1651_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[2:0]!=3'b011) | nand_302_cse;
  assign or_1649_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b11011) | (fsm_output[7]);
  assign mux_1167_nl = MUX_s_1_2_2(or_1651_nl, or_1649_nl, fsm_output[4]);
  assign or_1648_nl = (COMP_LOOP_acc_1_cse_6_sva[2]) | (~((COMP_LOOP_acc_1_cse_6_sva[1])
      & (COMP_LOOP_acc_1_cse_6_sva[4]) & (COMP_LOOP_acc_1_cse_6_sva[3]) & (COMP_LOOP_acc_1_cse_6_sva[0])
      & (fsm_output[7])));
  assign or_1647_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b11011) | (fsm_output[7]);
  assign mux_1166_nl = MUX_s_1_2_2(or_1648_nl, or_1647_nl, fsm_output[4]);
  assign mux_1168_nl = MUX_s_1_2_2(mux_1167_nl, mux_1166_nl, fsm_output[0]);
  assign nor_555_nl = ~((fsm_output[6]) | mux_1168_nl);
  assign mux_1172_nl = MUX_s_1_2_2(and_360_nl, nor_555_nl, fsm_output[3]);
  assign nand_479_nl = ~((fsm_output[5]) & mux_1172_nl);
  assign nor_557_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:2]!=3'b110) | nand_437_cse);
  assign nor_558_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b11011) | (fsm_output[7]));
  assign mux_1163_nl = MUX_s_1_2_2(nor_557_nl, nor_558_nl, fsm_output[4]);
  assign nor_559_nl = ~((COMP_LOOP_acc_14_psp_sva[3:1]!=3'b110) | nand_441_cse);
  assign nor_560_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1101) | (fsm_output[7]));
  assign mux_1162_nl = MUX_s_1_2_2(nor_559_nl, nor_560_nl, fsm_output[4]);
  assign and_361_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1162_nl;
  assign mux_1164_nl = MUX_s_1_2_2(mux_1163_nl, and_361_nl, fsm_output[0]);
  assign nand_157_nl = ~((fsm_output[6]) & mux_1164_nl);
  assign or_1638_nl = (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[0])) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | nand_289_cse;
  assign or_1636_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b11011) | (fsm_output[7]);
  assign mux_1160_nl = MUX_s_1_2_2(or_1638_nl, or_1636_nl, fsm_output[4]);
  assign nand_155_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & mux_1097_cse);
  assign mux_1161_nl = MUX_s_1_2_2(mux_1160_nl, nand_155_nl, fsm_output[0]);
  assign or_1639_nl = (fsm_output[6]) | mux_1161_nl;
  assign mux_1165_nl = MUX_s_1_2_2(nand_157_nl, or_1639_nl, fsm_output[3]);
  assign or_2253_nl = (fsm_output[5]) | mux_1165_nl;
  assign mux_1173_nl = MUX_s_1_2_2(nand_479_nl, or_2253_nl, fsm_output[2]);
  assign vec_rsc_0_27_i_we_d_pff = ~(mux_1173_nl | (fsm_output[1]));
  assign nor_546_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b11011) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_547_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_1187_nl = MUX_s_1_2_2(nor_546_nl, nor_547_nl, fsm_output[0]);
  assign and_357_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (~ mux_1154_cse);
  assign and_358_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]==5'b11011) & (fsm_output[4])
      & (fsm_output[6]) & (~ (fsm_output[7]));
  assign and_525_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]==5'b11011) & (fsm_output[7:6]==2'b10);
  assign nor_549_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b11011) | (fsm_output[7:6]!=2'b00));
  assign mux_1181_nl = MUX_s_1_2_2(and_525_nl, nor_549_nl, fsm_output[4]);
  assign mux_1182_nl = MUX_s_1_2_2(and_358_nl, mux_1181_nl, fsm_output[3]);
  assign mux_1186_nl = MUX_s_1_2_2(and_357_nl, mux_1182_nl, fsm_output[0]);
  assign mux_1188_nl = MUX_s_1_2_2(mux_1187_nl, mux_1186_nl, fsm_output[5]);
  assign or_1670_nl = (~((COMP_LOOP_acc_1_cse_sva[4:0]==5'b11011) & COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm))
      | nand_443_cse;
  assign nand_273_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]==5'b11011) & COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm
      & (fsm_output[7:6]==2'b01));
  assign mux_1178_nl = MUX_s_1_2_2(or_1670_nl, nand_273_nl, fsm_output[4]);
  assign nand_513_nl = ~((COMP_LOOP_acc_1_cse_6_sva[4:0]==5'b11011) & COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[7:6]==2'b10));
  assign or_1665_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b11011) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_1177_nl = MUX_s_1_2_2(nand_513_nl, or_1665_nl, fsm_output[4]);
  assign mux_1179_nl = MUX_s_1_2_2(mux_1178_nl, mux_1177_nl, fsm_output[3]);
  assign or_1664_nl = (COMP_LOOP_acc_10_cse_10_1_sva[2:1]!=2'b01) | nand_293_cse;
  assign nand_276_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]==5'b11011) & (fsm_output[7:6]==2'b01));
  assign mux_1175_nl = MUX_s_1_2_2(or_1664_nl, nand_276_nl, fsm_output[4]);
  assign nand_465_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]==5'b11011) & (fsm_output[7:6]==2'b10));
  assign or_1659_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b11011) | (fsm_output[7:6]!=2'b00);
  assign mux_1174_nl = MUX_s_1_2_2(nand_465_nl, or_1659_nl, fsm_output[4]);
  assign mux_1176_nl = MUX_s_1_2_2(mux_1175_nl, mux_1174_nl, fsm_output[3]);
  assign mux_1180_nl = MUX_s_1_2_2(mux_1179_nl, mux_1176_nl, fsm_output[0]);
  assign nor_550_nl = ~((fsm_output[5]) | mux_1180_nl);
  assign mux_1189_nl = MUX_s_1_2_2(mux_1188_nl, nor_550_nl, fsm_output[2]);
  assign vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1189_nl & (fsm_output[1]);
  assign nor_537_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b11100) | (~ (fsm_output[7])));
  assign nor_538_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b11100) | (fsm_output[7]));
  assign mux_1201_nl = MUX_s_1_2_2(nor_537_nl, nor_538_nl, fsm_output[4]);
  assign nor_539_nl = ~((COMP_LOOP_acc_1_cse_sva[4:0]!=5'b11100) | (~ (fsm_output[7])));
  assign nor_540_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b11100) | (fsm_output[7]));
  assign mux_1200_nl = MUX_s_1_2_2(nor_539_nl, nor_540_nl, fsm_output[4]);
  assign mux_1202_nl = MUX_s_1_2_2(mux_1201_nl, mux_1200_nl, fsm_output[0]);
  assign and_356_nl = (fsm_output[6]) & mux_1202_nl;
  assign or_1702_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[1:0]!=2'b00) | nand_266_cse;
  assign or_1700_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b11100) | (fsm_output[7]);
  assign mux_1198_nl = MUX_s_1_2_2(or_1702_nl, or_1700_nl, fsm_output[4]);
  assign or_1699_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b11100) | (~ (fsm_output[7]));
  assign or_1697_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b11100) | (fsm_output[7]);
  assign mux_1197_nl = MUX_s_1_2_2(or_1699_nl, or_1697_nl, fsm_output[4]);
  assign mux_1199_nl = MUX_s_1_2_2(mux_1198_nl, mux_1197_nl, fsm_output[0]);
  assign nor_541_nl = ~((fsm_output[6]) | mux_1199_nl);
  assign mux_1203_nl = MUX_s_1_2_2(and_356_nl, nor_541_nl, fsm_output[3]);
  assign nand_478_nl = ~((fsm_output[5]) & mux_1203_nl);
  assign nor_543_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b11100) | (~ (fsm_output[7])));
  assign nor_544_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b11100) | (fsm_output[7]));
  assign mux_1194_nl = MUX_s_1_2_2(nor_543_nl, nor_544_nl, fsm_output[4]);
  assign nand_519_nl = ~((COMP_LOOP_acc_14_psp_sva[3:0]==4'b1110) & (fsm_output[7]));
  assign or_1689_nl = (COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1110) | (fsm_output[7]);
  assign mux_1193_nl = MUX_s_1_2_2(nand_519_nl, or_1689_nl, fsm_output[4]);
  assign nor_545_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1193_nl);
  assign mux_1195_nl = MUX_s_1_2_2(mux_1194_nl, nor_545_nl, fsm_output[0]);
  assign nand_162_nl = ~((fsm_output[6]) & mux_1195_nl);
  assign or_1687_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b11100) | (~ (fsm_output[7]));
  assign or_1685_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b11100) | (fsm_output[7]);
  assign mux_1191_nl = MUX_s_1_2_2(or_1687_nl, or_1685_nl, fsm_output[4]);
  assign or_1684_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | mux_1190_cse;
  assign mux_1192_nl = MUX_s_1_2_2(mux_1191_nl, or_1684_nl, fsm_output[0]);
  assign or_1688_nl = (fsm_output[6]) | mux_1192_nl;
  assign mux_1196_nl = MUX_s_1_2_2(nand_162_nl, or_1688_nl, fsm_output[3]);
  assign or_2252_nl = (fsm_output[5]) | mux_1196_nl;
  assign mux_1204_nl = MUX_s_1_2_2(nand_478_nl, or_2252_nl, fsm_output[2]);
  assign vec_rsc_0_28_i_we_d_pff = ~(mux_1204_nl | (fsm_output[1]));
  assign nor_530_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b11100) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_531_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_1218_nl = MUX_s_1_2_2(nor_530_nl, nor_531_nl, fsm_output[0]);
  assign nor_532_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1216_cse);
  assign nor_533_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]!=5'b11100) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[7]));
  assign nor_534_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]!=5'b11100) | (fsm_output[7:6]!=2'b10));
  assign nor_535_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b11100) | (fsm_output[7:6]!=2'b00));
  assign mux_1212_nl = MUX_s_1_2_2(nor_534_nl, nor_535_nl, fsm_output[4]);
  assign mux_1213_nl = MUX_s_1_2_2(nor_533_nl, mux_1212_nl, fsm_output[3]);
  assign mux_1217_nl = MUX_s_1_2_2(nor_532_nl, mux_1213_nl, fsm_output[0]);
  assign mux_1219_nl = MUX_s_1_2_2(mux_1218_nl, mux_1217_nl, fsm_output[5]);
  assign or_1721_nl = (COMP_LOOP_acc_1_cse_sva[4:0]!=5'b11100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)
      | nand_443_cse;
  assign or_1719_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b11100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm)
      | (fsm_output[7:6]!=2'b01);
  assign mux_1209_nl = MUX_s_1_2_2(or_1721_nl, or_1719_nl, fsm_output[4]);
  assign or_1718_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b11100) | (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b10);
  assign or_1716_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b11100) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_1208_nl = MUX_s_1_2_2(or_1718_nl, or_1716_nl, fsm_output[4]);
  assign mux_1210_nl = MUX_s_1_2_2(mux_1209_nl, mux_1208_nl, fsm_output[3]);
  assign or_1715_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]!=5'b11100) | nand_443_cse;
  assign or_1713_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b11100) | (fsm_output[7:6]!=2'b01);
  assign mux_1206_nl = MUX_s_1_2_2(or_1715_nl, or_1713_nl, fsm_output[4]);
  assign or_1712_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b11100) | (fsm_output[7:6]!=2'b10);
  assign or_1710_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b11100) | (fsm_output[7:6]!=2'b00);
  assign mux_1205_nl = MUX_s_1_2_2(or_1712_nl, or_1710_nl, fsm_output[4]);
  assign mux_1207_nl = MUX_s_1_2_2(mux_1206_nl, mux_1205_nl, fsm_output[3]);
  assign mux_1211_nl = MUX_s_1_2_2(mux_1210_nl, mux_1207_nl, fsm_output[0]);
  assign nor_536_nl = ~((fsm_output[5]) | mux_1211_nl);
  assign mux_1220_nl = MUX_s_1_2_2(mux_1219_nl, nor_536_nl, fsm_output[2]);
  assign vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1220_nl & (fsm_output[1]);
  assign nor_520_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[1]) | (~((COMP_LOOP_acc_10_cse_10_1_sva[2])
      & (COMP_LOOP_acc_10_cse_10_1_sva[3]) & (COMP_LOOP_acc_10_cse_10_1_sva[4]) &
      (COMP_LOOP_acc_10_cse_10_1_sva[0]) & (fsm_output[7]))));
  assign nor_521_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b11101) | (fsm_output[7]));
  assign mux_1232_nl = MUX_s_1_2_2(nor_520_nl, nor_521_nl, fsm_output[4]);
  assign nor_522_nl = ~((~((COMP_LOOP_acc_1_cse_sva[4:1]==4'b1110))) | nand_446_cse);
  assign nor_523_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b11101) | (fsm_output[7]));
  assign mux_1231_nl = MUX_s_1_2_2(nor_522_nl, nor_523_nl, fsm_output[4]);
  assign mux_1233_nl = MUX_s_1_2_2(mux_1232_nl, mux_1231_nl, fsm_output[0]);
  assign and_351_nl = (fsm_output[6]) & mux_1233_nl;
  assign or_1751_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[1:0]!=2'b01) | nand_266_cse;
  assign or_1749_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b11101) | (fsm_output[7]);
  assign mux_1229_nl = MUX_s_1_2_2(or_1751_nl, or_1749_nl, fsm_output[4]);
  assign or_1748_nl = (COMP_LOOP_acc_1_cse_6_sva[2:1]!=2'b10) | nand_297_cse;
  assign or_1746_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b11101) | (fsm_output[7]);
  assign mux_1228_nl = MUX_s_1_2_2(or_1748_nl, or_1746_nl, fsm_output[4]);
  assign mux_1230_nl = MUX_s_1_2_2(mux_1229_nl, mux_1228_nl, fsm_output[0]);
  assign nor_524_nl = ~((fsm_output[6]) | mux_1230_nl);
  assign mux_1234_nl = MUX_s_1_2_2(and_351_nl, nor_524_nl, fsm_output[3]);
  assign nand_477_nl = ~((fsm_output[5]) & mux_1234_nl);
  assign nor_526_nl = ~((~((COMP_LOOP_acc_10_cse_10_1_7_sva[4:1]==4'b1110))) | nand_448_cse);
  assign nor_527_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b11101) | (fsm_output[7]));
  assign mux_1225_nl = MUX_s_1_2_2(nor_526_nl, nor_527_nl, fsm_output[4]);
  assign and_524_nl = (COMP_LOOP_acc_14_psp_sva[3:0]==4'b1110) & (fsm_output[7]);
  assign nor_529_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]!=4'b1110) | (fsm_output[7]));
  assign mux_1224_nl = MUX_s_1_2_2(and_524_nl, nor_529_nl, fsm_output[4]);
  assign and_352_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1224_nl;
  assign mux_1226_nl = MUX_s_1_2_2(mux_1225_nl, and_352_nl, fsm_output[0]);
  assign nand_168_nl = ~((fsm_output[6]) & mux_1226_nl);
  assign nand_512_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]==5'b11101) & (fsm_output[7]));
  assign or_1735_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b11101) | (fsm_output[7]);
  assign mux_1222_nl = MUX_s_1_2_2(nand_512_nl, or_1735_nl, fsm_output[4]);
  assign nand_166_nl = ~(nor_98_cse & mux_1221_cse);
  assign mux_1223_nl = MUX_s_1_2_2(mux_1222_nl, nand_166_nl, fsm_output[0]);
  assign or_1738_nl = (fsm_output[6]) | mux_1223_nl;
  assign mux_1227_nl = MUX_s_1_2_2(nand_168_nl, or_1738_nl, fsm_output[3]);
  assign or_2251_nl = (fsm_output[5]) | mux_1227_nl;
  assign mux_1235_nl = MUX_s_1_2_2(nand_477_nl, or_2251_nl, fsm_output[2]);
  assign vec_rsc_0_29_i_we_d_pff = ~(mux_1235_nl | (fsm_output[1]));
  assign nor_515_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b11101) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_516_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_1249_nl = MUX_s_1_2_2(nor_515_nl, nor_516_nl, fsm_output[0]);
  assign and_348_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (~ mux_1216_cse);
  assign and_349_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]==5'b11101) & (fsm_output[4])
      & (fsm_output[6]) & (~ (fsm_output[7]));
  assign and_523_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]==5'b11101) & (fsm_output[7:6]==2'b10);
  assign nor_518_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b11101) | (fsm_output[7:6]!=2'b00));
  assign mux_1243_nl = MUX_s_1_2_2(and_523_nl, nor_518_nl, fsm_output[4]);
  assign mux_1244_nl = MUX_s_1_2_2(and_349_nl, mux_1243_nl, fsm_output[3]);
  assign mux_1248_nl = MUX_s_1_2_2(and_348_nl, mux_1244_nl, fsm_output[0]);
  assign mux_1250_nl = MUX_s_1_2_2(mux_1249_nl, mux_1248_nl, fsm_output[5]);
  assign or_1768_nl = (~((COMP_LOOP_acc_1_cse_sva[4:0]==5'b11101) & COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm))
      | nand_443_cse;
  assign nand_251_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]==5'b11101) & COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm
      & (fsm_output[7:6]==2'b01));
  assign mux_1240_nl = MUX_s_1_2_2(or_1768_nl, nand_251_nl, fsm_output[4]);
  assign nand_511_nl = ~((COMP_LOOP_acc_1_cse_6_sva[4:0]==5'b11101) & COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[7:6]==2'b10));
  assign or_1763_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b11101) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_1239_nl = MUX_s_1_2_2(nand_511_nl, or_1763_nl, fsm_output[4]);
  assign mux_1241_nl = MUX_s_1_2_2(mux_1240_nl, mux_1239_nl, fsm_output[3]);
  assign or_1762_nl = (COMP_LOOP_acc_10_cse_10_1_sva[1]) | (~((COMP_LOOP_acc_10_cse_10_1_sva[2])
      & (COMP_LOOP_acc_10_cse_10_1_sva[3]) & (COMP_LOOP_acc_10_cse_10_1_sva[4]) &
      (COMP_LOOP_acc_10_cse_10_1_sva[0]) & (fsm_output[7:6]==2'b11)));
  assign nand_254_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]==5'b11101) & (fsm_output[7:6]==2'b01));
  assign mux_1237_nl = MUX_s_1_2_2(or_1762_nl, nand_254_nl, fsm_output[4]);
  assign nand_462_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]==5'b11101) & (fsm_output[7:6]==2'b10));
  assign or_1758_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b11101) | (fsm_output[7:6]!=2'b00);
  assign mux_1236_nl = MUX_s_1_2_2(nand_462_nl, or_1758_nl, fsm_output[4]);
  assign mux_1238_nl = MUX_s_1_2_2(mux_1237_nl, mux_1236_nl, fsm_output[3]);
  assign mux_1242_nl = MUX_s_1_2_2(mux_1241_nl, mux_1238_nl, fsm_output[0]);
  assign nor_519_nl = ~((fsm_output[5]) | mux_1242_nl);
  assign mux_1251_nl = MUX_s_1_2_2(mux_1250_nl, nor_519_nl, fsm_output[2]);
  assign vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1251_nl & (fsm_output[1]);
  assign and_529_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]==5'b11110) & (fsm_output[7]);
  assign nor_507_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]!=5'b11110) | (fsm_output[7]));
  assign mux_1263_nl = MUX_s_1_2_2(and_529_nl, nor_507_nl, fsm_output[4]);
  assign and_530_nl = (COMP_LOOP_acc_1_cse_sva[4:0]==5'b11110) & (fsm_output[7]);
  assign nor_509_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]!=5'b11110) | (fsm_output[7]));
  assign mux_1262_nl = MUX_s_1_2_2(and_530_nl, nor_509_nl, fsm_output[4]);
  assign mux_1264_nl = MUX_s_1_2_2(mux_1263_nl, mux_1262_nl, fsm_output[0]);
  assign and_347_nl = (fsm_output[6]) & mux_1264_nl;
  assign or_1796_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[0]) | (~((COMP_LOOP_acc_10_cse_10_1_6_sva[4:1]==4'b1111)
      & (fsm_output[7])));
  assign or_1795_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b11110) | (fsm_output[7]);
  assign mux_1260_nl = MUX_s_1_2_2(or_1796_nl, or_1795_nl, fsm_output[4]);
  assign nand_510_nl = ~((COMP_LOOP_acc_1_cse_6_sva[4:0]==5'b11110) & (fsm_output[7]));
  assign or_1792_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b11110) | (fsm_output[7]);
  assign mux_1259_nl = MUX_s_1_2_2(nand_510_nl, or_1792_nl, fsm_output[4]);
  assign mux_1261_nl = MUX_s_1_2_2(mux_1260_nl, mux_1259_nl, fsm_output[0]);
  assign nor_510_nl = ~((fsm_output[6]) | mux_1261_nl);
  assign mux_1265_nl = MUX_s_1_2_2(and_347_nl, nor_510_nl, fsm_output[3]);
  assign nand_476_nl = ~((fsm_output[5]) & mux_1265_nl);
  assign and_531_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]==5'b11110) & (fsm_output[7]);
  assign nor_513_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b11110) | (fsm_output[7]));
  assign mux_1256_nl = MUX_s_1_2_2(and_531_nl, nor_513_nl, fsm_output[4]);
  assign nand_243_nl = ~((COMP_LOOP_acc_14_psp_sva[3:0]==4'b1111) & (fsm_output[7]));
  assign nand_244_nl = ~((COMP_LOOP_acc_11_psp_sva[3:0]==4'b1111) & (~ (fsm_output[7])));
  assign mux_1255_nl = MUX_s_1_2_2(nand_243_nl, nand_244_nl, fsm_output[4]);
  assign nor_514_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1255_nl);
  assign mux_1257_nl = MUX_s_1_2_2(mux_1256_nl, nor_514_nl, fsm_output[0]);
  assign nand_173_nl = ~((fsm_output[6]) & mux_1257_nl);
  assign or_1784_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:1]==4'b1111)
      & (fsm_output[7])));
  assign or_1783_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]!=5'b11110) | (fsm_output[7]);
  assign mux_1253_nl = MUX_s_1_2_2(or_1784_nl, or_1783_nl, fsm_output[4]);
  assign or_1782_nl = (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | mux_1190_cse;
  assign mux_1254_nl = MUX_s_1_2_2(mux_1253_nl, or_1782_nl, fsm_output[0]);
  assign or_1785_nl = (fsm_output[6]) | mux_1254_nl;
  assign mux_1258_nl = MUX_s_1_2_2(nand_173_nl, or_1785_nl, fsm_output[3]);
  assign or_2250_nl = (fsm_output[5]) | mux_1258_nl;
  assign mux_1266_nl = MUX_s_1_2_2(nand_476_nl, or_2250_nl, fsm_output[2]);
  assign vec_rsc_0_30_i_we_d_pff = ~(mux_1266_nl | (fsm_output[1]));
  assign nor_500_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b11110) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_501_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_1280_nl = MUX_s_1_2_2(nor_500_nl, nor_501_nl, fsm_output[0]);
  assign nor_502_nl = ~((VEC_LOOP_j_10_0_sva_9_0[0]) | mux_1278_cse);
  assign and_345_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]==5'b11110) & (fsm_output[4])
      & (fsm_output[6]) & (~ (fsm_output[7]));
  assign and_522_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]==5'b11110) & (fsm_output[7:6]==2'b10);
  assign nor_504_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]!=5'b11110) | (fsm_output[7:6]!=2'b00));
  assign mux_1274_nl = MUX_s_1_2_2(and_522_nl, nor_504_nl, fsm_output[4]);
  assign mux_1275_nl = MUX_s_1_2_2(and_345_nl, mux_1274_nl, fsm_output[3]);
  assign mux_1279_nl = MUX_s_1_2_2(nor_502_nl, mux_1275_nl, fsm_output[0]);
  assign mux_1281_nl = MUX_s_1_2_2(mux_1280_nl, mux_1279_nl, fsm_output[5]);
  assign or_1815_nl = (~((COMP_LOOP_acc_1_cse_sva[4:0]==5'b11110) & COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm))
      | nand_443_cse;
  assign nand_231_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]==5'b11110) & COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm
      & (fsm_output[7:6]==2'b01));
  assign mux_1271_nl = MUX_s_1_2_2(or_1815_nl, nand_231_nl, fsm_output[4]);
  assign nand_509_nl = ~((COMP_LOOP_acc_1_cse_6_sva[4:0]==5'b11110) & COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[7:6]==2'b10));
  assign or_1810_nl = (COMP_LOOP_acc_1_cse_2_sva[4:0]!=5'b11110) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm)
      | (fsm_output[7:6]!=2'b00);
  assign mux_1270_nl = MUX_s_1_2_2(nand_509_nl, or_1810_nl, fsm_output[4]);
  assign mux_1272_nl = MUX_s_1_2_2(mux_1271_nl, mux_1270_nl, fsm_output[3]);
  assign or_1809_nl = (~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]==5'b11110))) | nand_443_cse;
  assign nand_234_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]==5'b11110) & (fsm_output[7:6]==2'b01));
  assign mux_1268_nl = MUX_s_1_2_2(or_1809_nl, nand_234_nl, fsm_output[4]);
  assign nand_460_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]==5'b11110) & (fsm_output[7:6]==2'b10));
  assign or_1804_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]!=5'b11110) | (fsm_output[7:6]!=2'b00);
  assign mux_1267_nl = MUX_s_1_2_2(nand_460_nl, or_1804_nl, fsm_output[4]);
  assign mux_1269_nl = MUX_s_1_2_2(mux_1268_nl, mux_1267_nl, fsm_output[3]);
  assign mux_1273_nl = MUX_s_1_2_2(mux_1272_nl, mux_1269_nl, fsm_output[0]);
  assign nor_505_nl = ~((fsm_output[5]) | mux_1273_nl);
  assign mux_1282_nl = MUX_s_1_2_2(mux_1281_nl, nor_505_nl, fsm_output[2]);
  assign vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1282_nl & (fsm_output[1]);
  assign and_334_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:0]==5'b11111) & (fsm_output[7]);
  assign and_335_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]==5'b11111) & (~ (fsm_output[7]));
  assign mux_1294_nl = MUX_s_1_2_2(and_334_nl, and_335_nl, fsm_output[4]);
  assign and_336_nl = (COMP_LOOP_acc_1_cse_sva[4:0]==5'b11111) & (fsm_output[7]);
  assign and_337_nl = (COMP_LOOP_acc_1_cse_4_sva[4:0]==5'b11111) & (~ (fsm_output[7]));
  assign mux_1293_nl = MUX_s_1_2_2(and_336_nl, and_337_nl, fsm_output[4]);
  assign mux_1295_nl = MUX_s_1_2_2(mux_1294_nl, mux_1293_nl, fsm_output[0]);
  assign and_333_nl = (fsm_output[6]) & mux_1295_nl;
  assign nand_223_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]==5'b11111) & (fsm_output[7]));
  assign nand_224_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]==5'b11111) & (~ (fsm_output[7])));
  assign mux_1291_nl = MUX_s_1_2_2(nand_223_nl, nand_224_nl, fsm_output[4]);
  assign nand_225_nl = ~((COMP_LOOP_acc_1_cse_6_sva[4:0]==5'b11111) & (fsm_output[7]));
  assign nand_226_nl = ~((COMP_LOOP_acc_1_cse_2_sva[4:0]==5'b11111) & (~ (fsm_output[7])));
  assign mux_1290_nl = MUX_s_1_2_2(nand_225_nl, nand_226_nl, fsm_output[4]);
  assign mux_1292_nl = MUX_s_1_2_2(mux_1291_nl, mux_1290_nl, fsm_output[0]);
  assign nor_498_nl = ~((fsm_output[6]) | mux_1292_nl);
  assign mux_1296_nl = MUX_s_1_2_2(and_333_nl, nor_498_nl, fsm_output[3]);
  assign nand_475_nl = ~((fsm_output[5]) & mux_1296_nl);
  assign and_338_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]==5'b11111) & (fsm_output[7]);
  assign and_339_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]==5'b11111) & (~ (fsm_output[7]));
  assign mux_1287_nl = MUX_s_1_2_2(and_338_nl, and_339_nl, fsm_output[4]);
  assign and_341_nl = (COMP_LOOP_acc_14_psp_sva[3:0]==4'b1111) & (fsm_output[7]);
  assign and_342_nl = (COMP_LOOP_acc_11_psp_sva[3:0]==4'b1111) & (~ (fsm_output[7]));
  assign mux_1286_nl = MUX_s_1_2_2(and_341_nl, and_342_nl, fsm_output[4]);
  assign and_340_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & mux_1286_nl;
  assign mux_1288_nl = MUX_s_1_2_2(mux_1287_nl, and_340_nl, fsm_output[0]);
  assign nand_179_nl = ~((fsm_output[6]) & mux_1288_nl);
  assign nand_227_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]==5'b11111) & (fsm_output[7]));
  assign nand_228_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[4:0]==5'b11111) & (~ (fsm_output[7])));
  assign mux_1284_nl = MUX_s_1_2_2(nand_227_nl, nand_228_nl, fsm_output[4]);
  assign nand_177_nl = ~((VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & mux_1221_cse);
  assign mux_1285_nl = MUX_s_1_2_2(mux_1284_nl, nand_177_nl, fsm_output[0]);
  assign or_1830_nl = (fsm_output[6]) | mux_1285_nl;
  assign mux_1289_nl = MUX_s_1_2_2(nand_179_nl, or_1830_nl, fsm_output[3]);
  assign or_2249_nl = (fsm_output[5]) | mux_1289_nl;
  assign mux_1297_nl = MUX_s_1_2_2(nand_475_nl, or_2249_nl, fsm_output[2]);
  assign vec_rsc_0_31_i_we_d_pff = ~(mux_1297_nl | (fsm_output[1]));
  assign nor_494_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b11111) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_495_nl = ~((COMP_LOOP_acc_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_1311_nl = MUX_s_1_2_2(nor_494_nl, nor_495_nl, fsm_output[0]);
  assign and_329_nl = (VEC_LOOP_j_10_0_sva_9_0[0]) & (~ mux_1278_cse);
  assign and_330_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:0]==5'b11111) & (fsm_output[4])
      & (fsm_output[6]) & (~ (fsm_output[7]));
  assign and_521_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[4:0]==5'b11111) & (fsm_output[7:6]==2'b10);
  assign and_331_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[4:0]==5'b11111) & (fsm_output[7:6]==2'b00);
  assign mux_1305_nl = MUX_s_1_2_2(and_521_nl, and_331_nl, fsm_output[4]);
  assign mux_1306_nl = MUX_s_1_2_2(and_330_nl, mux_1305_nl, fsm_output[3]);
  assign mux_1310_nl = MUX_s_1_2_2(and_329_nl, mux_1306_nl, fsm_output[0]);
  assign mux_1312_nl = MUX_s_1_2_2(mux_1311_nl, mux_1310_nl, fsm_output[5]);
  assign or_1848_nl = (~((COMP_LOOP_acc_1_cse_sva[4:0]==5'b11111) & COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm))
      | nand_443_cse;
  assign nand_214_nl = ~((COMP_LOOP_acc_1_cse_4_sva[4:0]==5'b11111) & COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm
      & (fsm_output[7:6]==2'b01));
  assign mux_1302_nl = MUX_s_1_2_2(or_1848_nl, nand_214_nl, fsm_output[4]);
  assign nand_508_nl = ~((COMP_LOOP_acc_1_cse_6_sva[4:0]==5'b11111) & COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[7:6]==2'b10));
  assign nand_216_nl = ~((COMP_LOOP_acc_1_cse_2_sva[4:0]==5'b11111) & COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm
      & (fsm_output[7:6]==2'b00));
  assign mux_1301_nl = MUX_s_1_2_2(nand_508_nl, nand_216_nl, fsm_output[4]);
  assign mux_1303_nl = MUX_s_1_2_2(mux_1302_nl, mux_1301_nl, fsm_output[3]);
  assign nand_217_nl = ~((COMP_LOOP_acc_10_cse_10_1_sva[4:0]==5'b11111) & (fsm_output[7:6]==2'b11));
  assign nand_218_nl = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[4:0]==5'b11111) & (fsm_output[7:6]==2'b01));
  assign mux_1299_nl = MUX_s_1_2_2(nand_217_nl, nand_218_nl, fsm_output[4]);
  assign nand_458_nl = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]==5'b11111) & (fsm_output[7:6]==2'b10));
  assign nand_220_nl = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[4:0]==5'b11111) & (fsm_output[7:6]==2'b00));
  assign mux_1298_nl = MUX_s_1_2_2(nand_458_nl, nand_220_nl, fsm_output[4]);
  assign mux_1300_nl = MUX_s_1_2_2(mux_1299_nl, mux_1298_nl, fsm_output[3]);
  assign mux_1304_nl = MUX_s_1_2_2(mux_1303_nl, mux_1300_nl, fsm_output[0]);
  assign nor_497_nl = ~((fsm_output[5]) | mux_1304_nl);
  assign mux_1313_nl = MUX_s_1_2_2(mux_1312_nl, nor_497_nl, fsm_output[2]);
  assign vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1313_nl & (fsm_output[1]);
  assign twiddle_rsc_0_0_i_radr_d_pff = MUX1HOT_v_5_7_2((z_out_8[6:2]), (z_out_7[9:5]),
      (z_out_7[8:4]), (COMP_LOOP_5_tmp_mul_idiv_sva[7:3]), (COMP_LOOP_2_tmp_mul_idiv_sva[9:5]),
      (COMP_LOOP_3_tmp_lshift_ncse_sva[8:4]), (COMP_LOOP_2_tmp_lshift_ncse_sva[9:5]),
      {and_dcpl_46 , COMP_LOOP_or_42_cse , and_dcpl_171 , and_dcpl_173 , and_dcpl_174
      , and_dcpl_176 , and_dcpl_177});
  assign nor_489_cse = ~((z_out_7[4:0]!=5'b00000) | (fsm_output[3]));
  assign nor_486_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[3:0]!=4'b0000) | (~ (fsm_output[3])));
  assign nor_487_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[4:0]!=5'b00000) | (~ (fsm_output[3])));
  assign mux_1318_nl = MUX_s_1_2_2(nor_486_nl, nor_487_nl, fsm_output[0]);
  assign nor_488_nl = ~((z_out_8[1:0]!=2'b00) | (fsm_output[3]));
  assign mux_1317_nl = MUX_s_1_2_2(nor_488_nl, nor_489_cse, fsm_output[0]);
  assign mux_1319_nl = MUX_s_1_2_2(mux_1318_nl, mux_1317_nl, fsm_output[1]);
  assign nor_490_nl = ~((z_out_7[3:0]!=4'b0000) | (fsm_output[3]));
  assign mux_1315_nl = MUX_s_1_2_2(nor_490_nl, nor_489_cse, fsm_output[0]);
  assign nor_492_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[2:0]!=3'b000) | (fsm_output[3]));
  assign nor_493_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[4:0]!=5'b00000) | (fsm_output[3]));
  assign mux_1314_nl = MUX_s_1_2_2(nor_492_nl, nor_493_nl, fsm_output[0]);
  assign mux_1316_nl = MUX_s_1_2_2(mux_1315_nl, mux_1314_nl, fsm_output[1]);
  assign mux_1320_nl = MUX_s_1_2_2(mux_1319_nl, mux_1316_nl, fsm_output[2]);
  assign twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1320_nl & and_dcpl_179;
  assign twiddle_rsc_0_1_i_radr_d_pff = z_out_7[9:5];
  assign nor_483_nl = ~((z_out_7[4:0]!=5'b00001) | (~ and_316_cse));
  assign nor_484_nl = ~((z_out_7[4:0]!=5'b00001) | (fsm_output[1:0]!=2'b00));
  assign mux_1322_nl = MUX_s_1_2_2(nor_483_nl, nor_484_nl, fsm_output[3]);
  assign or_1872_nl = (z_out_7[4:0]!=5'b00001) | (~ (fsm_output[1]));
  assign or_1870_nl = (z_out_7[4:0]!=5'b00001) | (fsm_output[1]);
  assign mux_1321_nl = MUX_s_1_2_2(or_1872_nl, or_1870_nl, fsm_output[0]);
  assign nor_485_nl = ~((fsm_output[3]) | mux_1321_nl);
  assign mux_1323_nl = MUX_s_1_2_2(mux_1322_nl, nor_485_nl, fsm_output[2]);
  assign twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1323_nl & and_dcpl_179;
  assign twiddle_rsc_0_2_i_radr_d_pff = MUX_v_5_2_2((z_out_7[9:5]), (z_out_7[8:4]),
      COMP_LOOP_tmp_or_35_cse);
  assign nor_480_cse = ~((z_out_7[4:0]!=5'b00010) | (fsm_output[3]));
  assign nor_479_cse = ~((z_out_7[3:0]!=4'b0001) | (fsm_output[3]));
  assign nor_477_nl = ~((fsm_output[0]) | (z_out_7[4:0]!=5'b00010) | (~ (fsm_output[3])));
  assign nor_478_nl = ~((~ (fsm_output[0])) | (z_out_7[4:0]!=5'b00010) | (fsm_output[3]));
  assign mux_1327_nl = MUX_s_1_2_2(nor_477_nl, nor_478_nl, fsm_output[1]);
  assign mux_1325_nl = MUX_s_1_2_2(nor_479_cse, nor_480_cse, fsm_output[0]);
  assign mux_1324_nl = MUX_s_1_2_2(nor_480_cse, nor_479_cse, fsm_output[0]);
  assign mux_1326_nl = MUX_s_1_2_2(mux_1325_nl, mux_1324_nl, fsm_output[1]);
  assign mux_1328_nl = MUX_s_1_2_2(mux_1327_nl, mux_1326_nl, fsm_output[2]);
  assign twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1328_nl & and_dcpl_179;
  assign nor_474_nl = ~((z_out_7[3]) | (z_out_7[4]) | (~ (z_out_7[0])) | (z_out_7[2])
      | not_tmp_618);
  assign nor_475_nl = ~((z_out_7[4:0]!=5'b00011) | (fsm_output[1:0]!=2'b00));
  assign mux_1330_nl = MUX_s_1_2_2(nor_474_nl, nor_475_nl, fsm_output[3]);
  assign or_1886_nl = (z_out_7[4:2]!=3'b000) | not_tmp_617;
  assign or_1884_nl = (z_out_7[4:0]!=5'b00011) | (fsm_output[1]);
  assign mux_1329_nl = MUX_s_1_2_2(or_1886_nl, or_1884_nl, fsm_output[0]);
  assign nor_476_nl = ~((fsm_output[3]) | mux_1329_nl);
  assign mux_1331_nl = MUX_s_1_2_2(mux_1330_nl, nor_476_nl, fsm_output[2]);
  assign twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1331_nl & and_dcpl_179;
  assign twiddle_rsc_0_4_i_radr_d_pff = MUX1HOT_v_5_6_2((z_out_7[9:5]), (z_out_7[8:4]),
      (COMP_LOOP_5_tmp_mul_idiv_sva[7:3]), (COMP_LOOP_2_tmp_mul_idiv_sva[9:5]), (COMP_LOOP_3_tmp_lshift_ncse_sva[8:4]),
      (COMP_LOOP_2_tmp_lshift_ncse_sva[9:5]), {COMP_LOOP_or_42_cse , and_dcpl_171
      , and_dcpl_173 , and_dcpl_174 , and_dcpl_176 , and_dcpl_177});
  assign nor_467_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[3:0]!=4'b0010) | (~ (fsm_output[3])));
  assign nor_468_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[4:0]!=5'b00100) | (~ (fsm_output[3])));
  assign mux_1335_nl = MUX_s_1_2_2(nor_467_nl, nor_468_nl, fsm_output[0]);
  assign nor_469_nl = ~((~ (fsm_output[0])) | (z_out_7[4:0]!=5'b00100) | (fsm_output[3]));
  assign mux_1336_nl = MUX_s_1_2_2(mux_1335_nl, nor_469_nl, fsm_output[1]);
  assign nor_470_nl = ~((z_out_7[3:0]!=4'b0010) | (fsm_output[3]));
  assign nor_471_nl = ~((z_out_7[4:0]!=5'b00100) | (fsm_output[3]));
  assign mux_1333_nl = MUX_s_1_2_2(nor_470_nl, nor_471_nl, fsm_output[0]);
  assign nor_472_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[2:0]!=3'b001) | (fsm_output[3]));
  assign nor_473_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[4:0]!=5'b00100) | (fsm_output[3]));
  assign mux_1332_nl = MUX_s_1_2_2(nor_472_nl, nor_473_nl, fsm_output[0]);
  assign mux_1334_nl = MUX_s_1_2_2(mux_1333_nl, mux_1332_nl, fsm_output[1]);
  assign mux_1337_nl = MUX_s_1_2_2(mux_1336_nl, mux_1334_nl, fsm_output[2]);
  assign twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1337_nl & and_dcpl_179;
  assign nor_464_nl = ~((z_out_7[4:0]!=5'b00101) | (~ and_316_cse));
  assign nor_465_nl = ~((z_out_7[4:0]!=5'b00101) | (fsm_output[1:0]!=2'b00));
  assign mux_1339_nl = MUX_s_1_2_2(nor_464_nl, nor_465_nl, fsm_output[3]);
  assign or_1902_nl = (z_out_7[4:0]!=5'b00101) | (~ (fsm_output[1]));
  assign or_1900_nl = (z_out_7[4:0]!=5'b00101) | (fsm_output[1]);
  assign mux_1338_nl = MUX_s_1_2_2(or_1902_nl, or_1900_nl, fsm_output[0]);
  assign nor_466_nl = ~((fsm_output[3]) | mux_1338_nl);
  assign mux_1340_nl = MUX_s_1_2_2(mux_1339_nl, nor_466_nl, fsm_output[2]);
  assign twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1340_nl & and_dcpl_179;
  assign nor_461_cse = ~((z_out_7[4:0]!=5'b00110) | (fsm_output[3]));
  assign nor_460_cse = ~((z_out_7[3:0]!=4'b0011) | (fsm_output[3]));
  assign nor_458_nl = ~((fsm_output[0]) | (z_out_7[4:0]!=5'b00110) | (~ (fsm_output[3])));
  assign nor_459_nl = ~((~ (fsm_output[0])) | (z_out_7[4:0]!=5'b00110) | (fsm_output[3]));
  assign mux_1344_nl = MUX_s_1_2_2(nor_458_nl, nor_459_nl, fsm_output[1]);
  assign mux_1342_nl = MUX_s_1_2_2(nor_460_cse, nor_461_cse, fsm_output[0]);
  assign mux_1341_nl = MUX_s_1_2_2(nor_461_cse, nor_460_cse, fsm_output[0]);
  assign mux_1343_nl = MUX_s_1_2_2(mux_1342_nl, mux_1341_nl, fsm_output[1]);
  assign mux_1345_nl = MUX_s_1_2_2(mux_1344_nl, mux_1343_nl, fsm_output[2]);
  assign twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1345_nl & and_dcpl_179;
  assign nor_455_nl = ~((z_out_7[4:3]!=2'b00) | not_tmp_625);
  assign nor_456_nl = ~((z_out_7[4:0]!=5'b00111) | (fsm_output[1:0]!=2'b00));
  assign mux_1347_nl = MUX_s_1_2_2(nor_455_nl, nor_456_nl, fsm_output[3]);
  assign or_1916_nl = (z_out_7[4:2]!=3'b001) | not_tmp_617;
  assign or_1914_nl = (z_out_7[4:0]!=5'b00111) | (fsm_output[1]);
  assign mux_1346_nl = MUX_s_1_2_2(or_1916_nl, or_1914_nl, fsm_output[0]);
  assign nor_457_nl = ~((fsm_output[3]) | mux_1346_nl);
  assign mux_1348_nl = MUX_s_1_2_2(mux_1347_nl, nor_457_nl, fsm_output[2]);
  assign twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1348_nl & and_dcpl_179;
  assign nor_450_cse = ~((z_out_7[4:0]!=5'b01000) | (fsm_output[3]));
  assign nor_447_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[3:0]!=4'b0100) | (~ (fsm_output[3])));
  assign nor_448_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[4:0]!=5'b01000) | (~ (fsm_output[3])));
  assign mux_1353_nl = MUX_s_1_2_2(nor_447_nl, nor_448_nl, fsm_output[0]);
  assign nor_449_nl = ~((z_out_8[1:0]!=2'b01) | (fsm_output[3]));
  assign mux_1352_nl = MUX_s_1_2_2(nor_449_nl, nor_450_cse, fsm_output[0]);
  assign mux_1354_nl = MUX_s_1_2_2(mux_1353_nl, mux_1352_nl, fsm_output[1]);
  assign nor_451_nl = ~((z_out_7[3:0]!=4'b0100) | (fsm_output[3]));
  assign mux_1350_nl = MUX_s_1_2_2(nor_451_nl, nor_450_cse, fsm_output[0]);
  assign nor_453_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[2:0]!=3'b010) | (fsm_output[3]));
  assign nor_454_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[4:0]!=5'b01000) | (fsm_output[3]));
  assign mux_1349_nl = MUX_s_1_2_2(nor_453_nl, nor_454_nl, fsm_output[0]);
  assign mux_1351_nl = MUX_s_1_2_2(mux_1350_nl, mux_1349_nl, fsm_output[1]);
  assign mux_1355_nl = MUX_s_1_2_2(mux_1354_nl, mux_1351_nl, fsm_output[2]);
  assign twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1355_nl & and_dcpl_179;
  assign nor_444_nl = ~((z_out_7[4:0]!=5'b01001) | (~ and_316_cse));
  assign nor_445_nl = ~((z_out_7[4:0]!=5'b01001) | (fsm_output[1:0]!=2'b00));
  assign mux_1357_nl = MUX_s_1_2_2(nor_444_nl, nor_445_nl, fsm_output[3]);
  assign or_1933_nl = (z_out_7[4:0]!=5'b01001) | (~ (fsm_output[1]));
  assign or_1931_nl = (z_out_7[4:0]!=5'b01001) | (fsm_output[1]);
  assign mux_1356_nl = MUX_s_1_2_2(or_1933_nl, or_1931_nl, fsm_output[0]);
  assign nor_446_nl = ~((fsm_output[3]) | mux_1356_nl);
  assign mux_1358_nl = MUX_s_1_2_2(mux_1357_nl, nor_446_nl, fsm_output[2]);
  assign twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1358_nl & and_dcpl_179;
  assign nor_441_cse = ~((z_out_7[4:0]!=5'b01010) | (fsm_output[3]));
  assign nor_440_cse = ~((z_out_7[3:0]!=4'b0101) | (fsm_output[3]));
  assign nor_438_nl = ~((fsm_output[0]) | (z_out_7[4:0]!=5'b01010) | (~ (fsm_output[3])));
  assign nor_439_nl = ~((~ (fsm_output[0])) | (z_out_7[4:0]!=5'b01010) | (fsm_output[3]));
  assign mux_1362_nl = MUX_s_1_2_2(nor_438_nl, nor_439_nl, fsm_output[1]);
  assign mux_1360_nl = MUX_s_1_2_2(nor_440_cse, nor_441_cse, fsm_output[0]);
  assign mux_1359_nl = MUX_s_1_2_2(nor_441_cse, nor_440_cse, fsm_output[0]);
  assign mux_1361_nl = MUX_s_1_2_2(mux_1360_nl, mux_1359_nl, fsm_output[1]);
  assign mux_1363_nl = MUX_s_1_2_2(mux_1362_nl, mux_1361_nl, fsm_output[2]);
  assign twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1363_nl & and_dcpl_179;
  assign nor_435_nl = ~((~ (z_out_7[3])) | (z_out_7[4]) | (~ (z_out_7[0])) | (z_out_7[2])
      | not_tmp_618);
  assign nor_436_nl = ~((z_out_7[4:0]!=5'b01011) | (fsm_output[1:0]!=2'b00));
  assign mux_1365_nl = MUX_s_1_2_2(nor_435_nl, nor_436_nl, fsm_output[3]);
  assign or_1947_nl = (z_out_7[2]) | (z_out_7[4]) | not_tmp_632;
  assign or_1945_nl = (z_out_7[4:0]!=5'b01011) | (fsm_output[1]);
  assign mux_1364_nl = MUX_s_1_2_2(or_1947_nl, or_1945_nl, fsm_output[0]);
  assign nor_437_nl = ~((fsm_output[3]) | mux_1364_nl);
  assign mux_1366_nl = MUX_s_1_2_2(mux_1365_nl, nor_437_nl, fsm_output[2]);
  assign twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1366_nl & and_dcpl_179;
  assign nor_428_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[3:0]!=4'b0110) | (~ (fsm_output[3])));
  assign nor_429_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[4:0]!=5'b01100) | (~ (fsm_output[3])));
  assign mux_1370_nl = MUX_s_1_2_2(nor_428_nl, nor_429_nl, fsm_output[0]);
  assign nor_430_nl = ~((~ (fsm_output[0])) | (z_out_7[4:0]!=5'b01100) | (fsm_output[3]));
  assign mux_1371_nl = MUX_s_1_2_2(mux_1370_nl, nor_430_nl, fsm_output[1]);
  assign nor_431_nl = ~((z_out_7[3:0]!=4'b0110) | (fsm_output[3]));
  assign nor_432_nl = ~((z_out_7[4:0]!=5'b01100) | (fsm_output[3]));
  assign mux_1368_nl = MUX_s_1_2_2(nor_431_nl, nor_432_nl, fsm_output[0]);
  assign nor_433_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[2:0]!=3'b011) | (fsm_output[3]));
  assign nor_434_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[4:0]!=5'b01100) | (fsm_output[3]));
  assign mux_1367_nl = MUX_s_1_2_2(nor_433_nl, nor_434_nl, fsm_output[0]);
  assign mux_1369_nl = MUX_s_1_2_2(mux_1368_nl, mux_1367_nl, fsm_output[1]);
  assign mux_1372_nl = MUX_s_1_2_2(mux_1371_nl, mux_1369_nl, fsm_output[2]);
  assign twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1372_nl & and_dcpl_179;
  assign nor_425_nl = ~((z_out_7[4:0]!=5'b01101) | (~ and_316_cse));
  assign nor_426_nl = ~((z_out_7[4:0]!=5'b01101) | (fsm_output[1:0]!=2'b00));
  assign mux_1374_nl = MUX_s_1_2_2(nor_425_nl, nor_426_nl, fsm_output[3]);
  assign or_1963_nl = (z_out_7[4:0]!=5'b01101) | (~ (fsm_output[1]));
  assign or_1961_nl = (z_out_7[4:0]!=5'b01101) | (fsm_output[1]);
  assign mux_1373_nl = MUX_s_1_2_2(or_1963_nl, or_1961_nl, fsm_output[0]);
  assign nor_427_nl = ~((fsm_output[3]) | mux_1373_nl);
  assign mux_1375_nl = MUX_s_1_2_2(mux_1374_nl, nor_427_nl, fsm_output[2]);
  assign twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1375_nl & and_dcpl_179;
  assign nor_422_cse = ~((z_out_7[4:0]!=5'b01110) | (fsm_output[3]));
  assign nor_421_cse = ~((z_out_7[3:0]!=4'b0111) | (fsm_output[3]));
  assign nor_419_nl = ~((fsm_output[0]) | (z_out_7[4:0]!=5'b01110) | (~ (fsm_output[3])));
  assign nor_420_nl = ~((~ (fsm_output[0])) | (z_out_7[4:0]!=5'b01110) | (fsm_output[3]));
  assign mux_1379_nl = MUX_s_1_2_2(nor_419_nl, nor_420_nl, fsm_output[1]);
  assign mux_1377_nl = MUX_s_1_2_2(nor_421_cse, nor_422_cse, fsm_output[0]);
  assign mux_1376_nl = MUX_s_1_2_2(nor_422_cse, nor_421_cse, fsm_output[0]);
  assign mux_1378_nl = MUX_s_1_2_2(mux_1377_nl, mux_1376_nl, fsm_output[1]);
  assign mux_1380_nl = MUX_s_1_2_2(mux_1379_nl, mux_1378_nl, fsm_output[2]);
  assign twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1380_nl & and_dcpl_179;
  assign nor_416_nl = ~((z_out_7[4:3]!=2'b01) | not_tmp_625);
  assign nor_417_nl = ~((z_out_7[4:0]!=5'b01111) | (fsm_output[1:0]!=2'b00));
  assign mux_1382_nl = MUX_s_1_2_2(nor_416_nl, nor_417_nl, fsm_output[3]);
  assign or_1977_nl = (~ (z_out_7[2])) | (z_out_7[4]) | not_tmp_632;
  assign or_1975_nl = (z_out_7[4:0]!=5'b01111) | (fsm_output[1]);
  assign mux_1381_nl = MUX_s_1_2_2(or_1977_nl, or_1975_nl, fsm_output[0]);
  assign nor_418_nl = ~((fsm_output[3]) | mux_1381_nl);
  assign mux_1383_nl = MUX_s_1_2_2(mux_1382_nl, nor_418_nl, fsm_output[2]);
  assign twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1383_nl & and_dcpl_179;
  assign nor_411_cse = ~((z_out_7[4:0]!=5'b10000) | (fsm_output[3]));
  assign nor_408_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[2:0]!=3'b000) | nand_204_cse);
  assign nor_409_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[3:0]!=4'b0000) | nand_205_cse);
  assign mux_1388_nl = MUX_s_1_2_2(nor_408_nl, nor_409_nl, fsm_output[0]);
  assign nor_410_nl = ~((z_out_8[1:0]!=2'b10) | (fsm_output[3]));
  assign mux_1387_nl = MUX_s_1_2_2(nor_410_nl, nor_411_cse, fsm_output[0]);
  assign mux_1389_nl = MUX_s_1_2_2(mux_1388_nl, mux_1387_nl, fsm_output[1]);
  assign nor_412_nl = ~((z_out_7[3:0]!=4'b1000) | (fsm_output[3]));
  assign mux_1385_nl = MUX_s_1_2_2(nor_412_nl, nor_411_cse, fsm_output[0]);
  assign nor_414_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[2:0]!=3'b100) | (fsm_output[3]));
  assign nor_415_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[4:0]!=5'b10000) | (fsm_output[3]));
  assign mux_1384_nl = MUX_s_1_2_2(nor_414_nl, nor_415_nl, fsm_output[0]);
  assign mux_1386_nl = MUX_s_1_2_2(mux_1385_nl, mux_1384_nl, fsm_output[1]);
  assign mux_1390_nl = MUX_s_1_2_2(mux_1389_nl, mux_1386_nl, fsm_output[2]);
  assign twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1390_nl & and_dcpl_179;
  assign nor_405_nl = ~((z_out_7[4:0]!=5'b10001) | (~ and_316_cse));
  assign nor_406_nl = ~((z_out_7[4:0]!=5'b10001) | (fsm_output[1:0]!=2'b00));
  assign mux_1392_nl = MUX_s_1_2_2(nor_405_nl, nor_406_nl, fsm_output[3]);
  assign or_1994_nl = (z_out_7[4:0]!=5'b10001) | (~ (fsm_output[1]));
  assign or_1992_nl = (z_out_7[4:0]!=5'b10001) | (fsm_output[1]);
  assign mux_1391_nl = MUX_s_1_2_2(or_1994_nl, or_1992_nl, fsm_output[0]);
  assign nor_407_nl = ~((fsm_output[3]) | mux_1391_nl);
  assign mux_1393_nl = MUX_s_1_2_2(mux_1392_nl, nor_407_nl, fsm_output[2]);
  assign twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1393_nl & and_dcpl_179;
  assign nor_402_cse = ~((z_out_7[4:0]!=5'b10010) | (fsm_output[3]));
  assign nor_401_cse = ~((z_out_7[3:0]!=4'b1001) | (fsm_output[3]));
  assign nor_399_nl = ~((fsm_output[0]) | (z_out_7[4:0]!=5'b10010) | (~ (fsm_output[3])));
  assign nor_400_nl = ~((~ (fsm_output[0])) | (z_out_7[4:0]!=5'b10010) | (fsm_output[3]));
  assign mux_1397_nl = MUX_s_1_2_2(nor_399_nl, nor_400_nl, fsm_output[1]);
  assign mux_1395_nl = MUX_s_1_2_2(nor_401_cse, nor_402_cse, fsm_output[0]);
  assign mux_1394_nl = MUX_s_1_2_2(nor_402_cse, nor_401_cse, fsm_output[0]);
  assign mux_1396_nl = MUX_s_1_2_2(mux_1395_nl, mux_1394_nl, fsm_output[1]);
  assign mux_1398_nl = MUX_s_1_2_2(mux_1397_nl, mux_1396_nl, fsm_output[2]);
  assign twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1398_nl & and_dcpl_179;
  assign nor_396_nl = ~((z_out_7[3]) | (~ (z_out_7[4])) | (~ (z_out_7[0])) | (z_out_7[2])
      | not_tmp_618);
  assign nor_397_nl = ~((z_out_7[4:0]!=5'b10011) | (fsm_output[1:0]!=2'b00));
  assign mux_1400_nl = MUX_s_1_2_2(nor_396_nl, nor_397_nl, fsm_output[3]);
  assign or_2008_nl = (z_out_7[4:2]!=3'b100) | not_tmp_617;
  assign or_2006_nl = (z_out_7[4:0]!=5'b10011) | (fsm_output[1]);
  assign mux_1399_nl = MUX_s_1_2_2(or_2008_nl, or_2006_nl, fsm_output[0]);
  assign nor_398_nl = ~((fsm_output[3]) | mux_1399_nl);
  assign mux_1401_nl = MUX_s_1_2_2(mux_1400_nl, nor_398_nl, fsm_output[2]);
  assign twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1401_nl & and_dcpl_179;
  assign nor_389_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[2:0]!=3'b010) | nand_204_cse);
  assign nor_390_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[3:0]!=4'b0100) | nand_205_cse);
  assign mux_1405_nl = MUX_s_1_2_2(nor_389_nl, nor_390_nl, fsm_output[0]);
  assign nor_391_nl = ~((~ (fsm_output[0])) | (z_out_7[4:0]!=5'b10100) | (fsm_output[3]));
  assign mux_1406_nl = MUX_s_1_2_2(mux_1405_nl, nor_391_nl, fsm_output[1]);
  assign nor_392_nl = ~((z_out_7[3:0]!=4'b1010) | (fsm_output[3]));
  assign nor_393_nl = ~((z_out_7[4:0]!=5'b10100) | (fsm_output[3]));
  assign mux_1403_nl = MUX_s_1_2_2(nor_392_nl, nor_393_nl, fsm_output[0]);
  assign nor_394_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[2:0]!=3'b101) | (fsm_output[3]));
  assign nor_395_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[4:0]!=5'b10100) | (fsm_output[3]));
  assign mux_1402_nl = MUX_s_1_2_2(nor_394_nl, nor_395_nl, fsm_output[0]);
  assign mux_1404_nl = MUX_s_1_2_2(mux_1403_nl, mux_1402_nl, fsm_output[1]);
  assign mux_1407_nl = MUX_s_1_2_2(mux_1406_nl, mux_1404_nl, fsm_output[2]);
  assign twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1407_nl & and_dcpl_179;
  assign nor_386_nl = ~((z_out_7[4:0]!=5'b10101) | (~ and_316_cse));
  assign nor_387_nl = ~((z_out_7[4:0]!=5'b10101) | (fsm_output[1:0]!=2'b00));
  assign mux_1409_nl = MUX_s_1_2_2(nor_386_nl, nor_387_nl, fsm_output[3]);
  assign or_2024_nl = (z_out_7[4:0]!=5'b10101) | (~ (fsm_output[1]));
  assign or_2022_nl = (z_out_7[4:0]!=5'b10101) | (fsm_output[1]);
  assign mux_1408_nl = MUX_s_1_2_2(or_2024_nl, or_2022_nl, fsm_output[0]);
  assign nor_388_nl = ~((fsm_output[3]) | mux_1408_nl);
  assign mux_1410_nl = MUX_s_1_2_2(mux_1409_nl, nor_388_nl, fsm_output[2]);
  assign twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1410_nl & and_dcpl_179;
  assign nor_383_cse = ~((z_out_7[4:0]!=5'b10110) | (fsm_output[3]));
  assign nor_382_cse = ~((z_out_7[3:0]!=4'b1011) | (fsm_output[3]));
  assign nor_380_nl = ~((fsm_output[0]) | (z_out_7[4:0]!=5'b10110) | (~ (fsm_output[3])));
  assign nor_381_nl = ~((~ (fsm_output[0])) | (z_out_7[4:0]!=5'b10110) | (fsm_output[3]));
  assign mux_1414_nl = MUX_s_1_2_2(nor_380_nl, nor_381_nl, fsm_output[1]);
  assign mux_1412_nl = MUX_s_1_2_2(nor_382_cse, nor_383_cse, fsm_output[0]);
  assign mux_1411_nl = MUX_s_1_2_2(nor_383_cse, nor_382_cse, fsm_output[0]);
  assign mux_1413_nl = MUX_s_1_2_2(mux_1412_nl, mux_1411_nl, fsm_output[1]);
  assign mux_1415_nl = MUX_s_1_2_2(mux_1414_nl, mux_1413_nl, fsm_output[2]);
  assign twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1415_nl & and_dcpl_179;
  assign nor_377_nl = ~((z_out_7[3]) | (~((z_out_7[4]) & (z_out_7[0]) & (z_out_7[2])
      & (z_out_7[1]) & (fsm_output[1:0]==2'b11))));
  assign nor_378_nl = ~((z_out_7[4:0]!=5'b10111) | (fsm_output[1:0]!=2'b00));
  assign mux_1417_nl = MUX_s_1_2_2(nor_377_nl, nor_378_nl, fsm_output[3]);
  assign or_2038_nl = (z_out_7[4:2]!=3'b101) | not_tmp_617;
  assign or_2036_nl = (z_out_7[4:0]!=5'b10111) | (fsm_output[1]);
  assign mux_1416_nl = MUX_s_1_2_2(or_2038_nl, or_2036_nl, fsm_output[0]);
  assign nor_379_nl = ~((fsm_output[3]) | mux_1416_nl);
  assign mux_1418_nl = MUX_s_1_2_2(mux_1417_nl, nor_379_nl, fsm_output[2]);
  assign twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1418_nl & and_dcpl_179;
  assign nor_372_cse = ~((z_out_7[4:0]!=5'b11000) | (fsm_output[3]));
  assign nor_369_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[1:0]!=2'b00) | (~((COMP_LOOP_3_tmp_lshift_ncse_sva[3:2]==2'b11)
      & (fsm_output[3]))));
  assign nor_370_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[2:0]!=3'b000) | (~((COMP_LOOP_2_tmp_lshift_ncse_sva[4:3]==2'b11)
      & (fsm_output[3]))));
  assign mux_1423_nl = MUX_s_1_2_2(nor_369_nl, nor_370_nl, fsm_output[0]);
  assign nor_371_nl = ~((z_out_8[1:0]!=2'b11) | (fsm_output[3]));
  assign mux_1422_nl = MUX_s_1_2_2(nor_371_nl, nor_372_cse, fsm_output[0]);
  assign mux_1424_nl = MUX_s_1_2_2(mux_1423_nl, mux_1422_nl, fsm_output[1]);
  assign nor_373_nl = ~((z_out_7[3:0]!=4'b1100) | (fsm_output[3]));
  assign mux_1420_nl = MUX_s_1_2_2(nor_373_nl, nor_372_cse, fsm_output[0]);
  assign nor_375_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[2:0]!=3'b110) | (fsm_output[3]));
  assign nor_376_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[4:0]!=5'b11000) | (fsm_output[3]));
  assign mux_1419_nl = MUX_s_1_2_2(nor_375_nl, nor_376_nl, fsm_output[0]);
  assign mux_1421_nl = MUX_s_1_2_2(mux_1420_nl, mux_1419_nl, fsm_output[1]);
  assign mux_1425_nl = MUX_s_1_2_2(mux_1424_nl, mux_1421_nl, fsm_output[2]);
  assign twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1425_nl & and_dcpl_179;
  assign nor_366_nl = ~((z_out_7[4:0]!=5'b11001) | (~ and_316_cse));
  assign nor_367_nl = ~((z_out_7[4:0]!=5'b11001) | (fsm_output[1:0]!=2'b00));
  assign mux_1427_nl = MUX_s_1_2_2(nor_366_nl, nor_367_nl, fsm_output[3]);
  assign or_2054_nl = (z_out_7[4:0]!=5'b11001) | (~ (fsm_output[1]));
  assign or_2052_nl = (z_out_7[4:0]!=5'b11001) | (fsm_output[1]);
  assign mux_1426_nl = MUX_s_1_2_2(or_2054_nl, or_2052_nl, fsm_output[0]);
  assign nor_368_nl = ~((fsm_output[3]) | mux_1426_nl);
  assign mux_1428_nl = MUX_s_1_2_2(mux_1427_nl, nor_368_nl, fsm_output[2]);
  assign twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1428_nl & and_dcpl_179;
  assign nor_363_cse = ~((z_out_7[4:0]!=5'b11010) | (fsm_output[3]));
  assign nor_362_cse = ~((z_out_7[3:0]!=4'b1101) | (fsm_output[3]));
  assign nor_360_nl = ~((fsm_output[0]) | (z_out_7[4:0]!=5'b11010) | (~ (fsm_output[3])));
  assign nor_361_nl = ~((~ (fsm_output[0])) | (z_out_7[4:0]!=5'b11010) | (fsm_output[3]));
  assign mux_1432_nl = MUX_s_1_2_2(nor_360_nl, nor_361_nl, fsm_output[1]);
  assign mux_1430_nl = MUX_s_1_2_2(nor_362_cse, nor_363_cse, fsm_output[0]);
  assign mux_1429_nl = MUX_s_1_2_2(nor_363_cse, nor_362_cse, fsm_output[0]);
  assign mux_1431_nl = MUX_s_1_2_2(mux_1430_nl, mux_1429_nl, fsm_output[1]);
  assign mux_1433_nl = MUX_s_1_2_2(mux_1432_nl, mux_1431_nl, fsm_output[2]);
  assign twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1433_nl & and_dcpl_179;
  assign nor_357_nl = ~((~((z_out_7[3]) & (z_out_7[4]) & (z_out_7[0]) & (~ (z_out_7[2]))))
      | not_tmp_618);
  assign nor_358_nl = ~((z_out_7[4:0]!=5'b11011) | (fsm_output[1:0]!=2'b00));
  assign mux_1435_nl = MUX_s_1_2_2(nor_357_nl, nor_358_nl, fsm_output[3]);
  assign or_2067_nl = (z_out_7[2]) | (~((z_out_7[4]) & (z_out_7[3]) & (z_out_7[0])
      & (z_out_7[1]) & (fsm_output[1])));
  assign or_2066_nl = (z_out_7[4:0]!=5'b11011) | (fsm_output[1]);
  assign mux_1434_nl = MUX_s_1_2_2(or_2067_nl, or_2066_nl, fsm_output[0]);
  assign nor_359_nl = ~((fsm_output[3]) | mux_1434_nl);
  assign mux_1436_nl = MUX_s_1_2_2(mux_1435_nl, nor_359_nl, fsm_output[2]);
  assign twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1436_nl & and_dcpl_179;
  assign nor_351_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[0]) | (~((COMP_LOOP_3_tmp_lshift_ncse_sva[3:1]==3'b111)
      & (fsm_output[3]))));
  assign nor_352_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[1:0]!=2'b00) | (~((COMP_LOOP_2_tmp_lshift_ncse_sva[4:2]==3'b111)
      & (fsm_output[3]))));
  assign mux_1440_nl = MUX_s_1_2_2(nor_351_nl, nor_352_nl, fsm_output[0]);
  assign nor_353_nl = ~((~ (fsm_output[0])) | (z_out_7[4:0]!=5'b11100) | (fsm_output[3]));
  assign mux_1441_nl = MUX_s_1_2_2(mux_1440_nl, nor_353_nl, fsm_output[1]);
  assign nor_354_nl = ~((z_out_7[3:0]!=4'b1110) | (fsm_output[3]));
  assign nor_355_nl = ~((z_out_7[4:0]!=5'b11100) | (fsm_output[3]));
  assign mux_1438_nl = MUX_s_1_2_2(nor_354_nl, nor_355_nl, fsm_output[0]);
  assign and_328_nl = (COMP_LOOP_5_tmp_mul_idiv_sva[2:0]==3'b111) & (~ (fsm_output[3]));
  assign nor_356_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[4:0]!=5'b11100) | (fsm_output[3]));
  assign mux_1437_nl = MUX_s_1_2_2(and_328_nl, nor_356_nl, fsm_output[0]);
  assign mux_1439_nl = MUX_s_1_2_2(mux_1438_nl, mux_1437_nl, fsm_output[1]);
  assign mux_1442_nl = MUX_s_1_2_2(mux_1441_nl, mux_1439_nl, fsm_output[2]);
  assign twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1442_nl & and_dcpl_179;
  assign and_327_nl = (z_out_7[4:0]==5'b11101) & and_316_cse;
  assign nor_349_nl = ~((z_out_7[4:0]!=5'b11101) | (fsm_output[1:0]!=2'b00));
  assign mux_1444_nl = MUX_s_1_2_2(and_327_nl, nor_349_nl, fsm_output[3]);
  assign nand_474_nl = ~((z_out_7[4:0]==5'b11101) & (fsm_output[1]));
  assign or_2080_nl = (z_out_7[4:0]!=5'b11101) | (fsm_output[1]);
  assign mux_1443_nl = MUX_s_1_2_2(nand_474_nl, or_2080_nl, fsm_output[0]);
  assign nor_350_nl = ~((fsm_output[3]) | mux_1443_nl);
  assign mux_1445_nl = MUX_s_1_2_2(mux_1444_nl, nor_350_nl, fsm_output[2]);
  assign twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1445_nl & and_dcpl_179;
  assign nor_347_cse = ~((z_out_7[4:0]!=5'b11110) | (fsm_output[3]));
  assign and_325_cse = (z_out_7[3:0]==4'b1111) & (~ (fsm_output[3]));
  assign and_323_nl = (~ (fsm_output[0])) & (z_out_7[4:0]==5'b11110) & (fsm_output[3]);
  assign and_324_nl = (fsm_output[0]) & (z_out_7[4:0]==5'b11110) & (~ (fsm_output[3]));
  assign mux_1449_nl = MUX_s_1_2_2(and_323_nl, and_324_nl, fsm_output[1]);
  assign mux_1447_nl = MUX_s_1_2_2(and_325_cse, nor_347_cse, fsm_output[0]);
  assign mux_1446_nl = MUX_s_1_2_2(nor_347_cse, and_325_cse, fsm_output[0]);
  assign mux_1448_nl = MUX_s_1_2_2(mux_1447_nl, mux_1446_nl, fsm_output[1]);
  assign mux_1450_nl = MUX_s_1_2_2(mux_1449_nl, mux_1448_nl, fsm_output[2]);
  assign twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1450_nl & and_dcpl_179;
  assign and_321_nl = (z_out_7[4:0]==5'b11111) & (fsm_output[1:0]==2'b11);
  assign and_322_nl = (z_out_7[4:0]==5'b11111) & (fsm_output[1:0]==2'b00);
  assign mux_1452_nl = MUX_s_1_2_2(and_321_nl, and_322_nl, fsm_output[3]);
  assign nand_192_nl = ~((z_out_7[4:0]==5'b11111) & (fsm_output[1]));
  assign nand_193_nl = ~((z_out_7[4:0]==5'b11111) & (~ (fsm_output[1])));
  assign mux_1451_nl = MUX_s_1_2_2(nand_192_nl, nand_193_nl, fsm_output[0]);
  assign nor_346_nl = ~((fsm_output[3]) | mux_1451_nl);
  assign mux_1453_nl = MUX_s_1_2_2(mux_1452_nl, nor_346_nl, fsm_output[2]);
  assign twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d = mux_1453_nl & and_dcpl_179;
  assign and_dcpl_334 = (fsm_output[6]) & (fsm_output[7]) & (fsm_output[1]) & (fsm_output[0])
      & and_dcpl_29 & (~ (fsm_output[2])) & (fsm_output[5]);
  assign and_dcpl_347 = nor_1025_cse & (fsm_output[1:0]==2'b10) & and_dcpl_29 & and_dcpl_28;
  assign and_dcpl_353 = (fsm_output[7:6]==2'b00) & and_dcpl_31;
  assign and_605_cse = and_dcpl_353 & and_dcpl_29 & (~ (fsm_output[2])) & (fsm_output[5]);
  assign and_609_cse = and_dcpl_353 & and_479_cse & and_dcpl_35;
  assign and_dcpl_365 = (fsm_output[7:6]==2'b01) & and_dcpl_31;
  assign and_614_cse = and_dcpl_365 & and_479_cse & and_dcpl_28;
  assign and_617_cse = and_dcpl_365 & and_dcpl_59 & and_dcpl_35;
  assign and_dcpl_372 = (fsm_output[7:6]==2'b10) & and_dcpl_31;
  assign and_621_cse = and_dcpl_372 & and_dcpl_59 & and_dcpl_28;
  assign and_624_cse = and_dcpl_372 & and_dcpl_69 & and_dcpl_35;
  assign and_628_cse = (fsm_output[7:6]==2'b11) & and_dcpl_31 & and_dcpl_69 & and_dcpl_28;
  assign and_dcpl_419 = nor_1025_cse & (fsm_output[1:0]==2'b10);
  assign and_dcpl_420 = and_dcpl_419 & and_dcpl_30;
  assign and_dcpl_422 = nor_1025_cse & (fsm_output[1:0]==2'b11);
  assign and_dcpl_423 = and_dcpl_422 & and_dcpl_30;
  assign and_dcpl_425 = and_dcpl_29 & (fsm_output[2]) & (~ (fsm_output[5]));
  assign and_dcpl_428 = nor_1025_cse & (fsm_output[1:0]==2'b01) & and_dcpl_425;
  assign and_dcpl_429 = and_dcpl_419 & and_dcpl_425;
  assign and_dcpl_433 = nor_1025_cse & (fsm_output[1:0]==2'b00);
  assign and_dcpl_434 = and_dcpl_433 & (fsm_output[4:3]==2'b01) & and_dcpl_28;
  assign and_dcpl_435 = and_dcpl_433 & and_dcpl_425;
  assign and_dcpl_436 = and_dcpl_422 & and_dcpl_425;
  assign and_dcpl_448 = and_dcpl_33 & and_dcpl_59 & and_dcpl_28;
  assign and_dcpl_452 = and_dcpl_33 & and_dcpl_69 & and_dcpl_35;
  assign and_dcpl_456 = and_dcpl_365 & and_dcpl_69 & and_dcpl_28;
  assign and_dcpl_458 = and_dcpl_365 & and_dcpl_29 & and_dcpl_35;
  assign and_dcpl_461 = and_dcpl_372 & and_dcpl_30;
  assign and_dcpl_465 = and_dcpl_372 & and_479_cse & and_dcpl_50;
  assign and_dcpl_468 = and_dcpl_372 & and_479_cse & (~ (fsm_output[2])) & (fsm_output[5]);
  assign and_dcpl_472 = (fsm_output[7:6]==2'b11) & and_dcpl_31 & and_dcpl_59 & and_dcpl_50;
  assign and_dcpl_479 = and_dcpl_353 & and_dcpl_29 & (fsm_output[2]) & (~ (fsm_output[5]));
  assign or_tmp_2098 = (~ (fsm_output[7])) | (fsm_output[5]) | (~ or_212_cse);
  assign mux_1600_nl = MUX_s_1_2_2(or_212_cse, (~ or_212_cse), fsm_output[5]);
  assign nand_520_nl = ~((fsm_output[7]) & mux_1600_nl);
  assign mux_tmp_1564 = MUX_s_1_2_2(nand_520_nl, or_tmp_2098, fsm_output[2]);
  assign COMP_LOOP_or_33_itm = and_605_cse | and_609_cse | and_614_cse | and_617_cse
      | and_621_cse | and_624_cse | and_628_cse;
  assign COMP_LOOP_tmp_or_71_itm = and_dcpl_435 | and_dcpl_436;
  assign COMP_LOOP_tmp_or_54_ssc = and_dcpl_428 | and_dcpl_429 | and_dcpl_434;
  always @(posedge clk) begin
    if ( (and_dcpl_33 & and_dcpl_30) | STAGE_LOOP_i_3_0_sva_mx0c1 ) begin
      STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(4'b1010, z_out_4, STAGE_LOOP_i_3_0_sva_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(nor_1019_nl, mux_320_nl, fsm_output[5]) ) begin
      p_sva <= p_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_vec_rsc_triosy_0_31_obj_ld_cse <= 1'b0;
      reg_ensig_cgo_cse <= 1'b0;
      COMP_LOOP_1_tmp_mul_idiv_sva_1_0 <= 2'b00;
      COMP_LOOP_3_tmp_mul_idiv_sva_3_0 <= 4'b0000;
    end
    else begin
      reg_vec_rsc_triosy_0_31_obj_ld_cse <= and_464_cse & (fsm_output[5:0]==6'b100100)
          & (~ (z_out_2[4]));
      reg_ensig_cgo_cse <= mux_1462_rmff;
      COMP_LOOP_1_tmp_mul_idiv_sva_1_0 <= z_out_8[1:0];
      COMP_LOOP_3_tmp_mul_idiv_sva_3_0 <= z_out_7[3:0];
    end
  end
  always @(posedge clk) begin
    tmp_21_sva_2 <= twiddle_rsc_0_2_i_q_d;
    tmp_21_sva_6 <= twiddle_rsc_0_6_i_q_d;
    tmp_21_sva_11 <= MUX_v_64_2_2(twiddle_rsc_0_11_i_q_d, twiddle_rsc_0_30_i_q_d,
        and_dcpl_176);
    tmp_21_sva_13 <= MUX_v_64_2_2(twiddle_rsc_0_13_i_q_d, twiddle_rsc_0_6_i_q_d,
        and_dcpl_176);
    tmp_21_sva_14 <= MUX_v_64_2_2(twiddle_rsc_0_14_i_q_d, twiddle_rsc_0_10_i_q_d,
        and_dcpl_176);
    tmp_21_sva_15 <= MUX_v_64_2_2(twiddle_rsc_0_15_i_q_d, twiddle_rsc_0_14_i_q_d,
        and_dcpl_176);
    tmp_21_sva_17 <= MUX_v_64_2_2(twiddle_rsc_0_17_i_q_d, twiddle_rsc_0_18_i_q_d,
        and_dcpl_176);
    tmp_21_sva_18 <= twiddle_rsc_0_18_i_q_d;
    tmp_21_sva_22 <= twiddle_rsc_0_22_i_q_d;
    tmp_21_sva_26 <= twiddle_rsc_0_26_i_q_d;
    tmp_21_sva_30 <= twiddle_rsc_0_30_i_q_d;
  end
  always @(posedge clk) begin
    if ( rst ) begin
      VEC_LOOP_j_10_0_sva_9_0 <= 10'b0000000000;
    end
    else if ( VEC_LOOP_j_10_0_sva_9_0_mx0c0 | (and_dcpl_82 & and_dcpl_104) ) begin
      VEC_LOOP_j_10_0_sva_9_0 <= MUX_v_10_2_2(10'b0000000000, (z_out_3[9:0]), VEC_LOOP_j_not_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(nor_1160_nl, and_nl, fsm_output[5]) ) begin
      STAGE_LOOP_lshift_psp_sva <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_1604_nl, mux_1603_nl, fsm_output[1]) ) begin
      COMP_LOOP_k_10_3_sva_6_0 <= MUX_v_7_2_2(7'b0000000, reg_COMP_LOOP_k_10_3_ftd,
          nand_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_1_sva <= 10'b0000000000;
    end
    else if ( ~ or_dcpl_84 ) begin
      COMP_LOOP_acc_10_cse_10_1_1_sva <= COMP_LOOP_1_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_psp_sva <= 7'b0000000;
    end
    else if ( ~ or_dcpl_84 ) begin
      COMP_LOOP_acc_psp_sva <= COMP_LOOP_acc_psp_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_5_tmp_mul_idiv_sva <= 8'b00000000;
    end
    else if ( ~ or_dcpl_84 ) begin
      COMP_LOOP_5_tmp_mul_idiv_sva <= z_out_7[7:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ or_dcpl_84 ) begin
      COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm <= z_out_3[10];
    end
  end
  always @(posedge clk) begin
    if ( ~ or_dcpl_84 ) begin
      COMP_LOOP_1_tmp_acc_cse_sva <= z_out_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_625_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_126_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_377_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_128_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_129_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_130_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_6_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_132_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_133_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_134_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_10_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_136_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_12_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_13_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_14_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_140_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_141_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_142_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_18_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_144_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_20_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_21_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_22_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_23_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_24_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_25_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_26_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_27_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_28_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_29_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_30_itm <= 1'b0;
    end
    else if ( mux_1489_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_itm <= ~((COMP_LOOP_acc_psp_sva_mx0w0[1:0]!=2'b00)
          | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_625_itm <= (COMP_LOOP_acc_1_cse_6_sva_1[4:0]==5'b00110);
      COMP_LOOP_COMP_LOOP_and_126_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[4:0]==5'b00011);
      COMP_LOOP_COMP_LOOP_and_377_itm <= (COMP_LOOP_acc_1_cse_4_sva_1[4:0]==5'b00110);
      COMP_LOOP_COMP_LOOP_and_128_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[4:0]==5'b00101);
      COMP_LOOP_COMP_LOOP_and_129_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[4:0]==5'b00110);
      COMP_LOOP_COMP_LOOP_and_130_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[4:0]==5'b00111);
      COMP_LOOP_COMP_LOOP_and_6_itm <= (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111) & (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b00);
      COMP_LOOP_COMP_LOOP_and_132_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[4:0]==5'b01001);
      COMP_LOOP_COMP_LOOP_and_133_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[4:0]==5'b01010);
      COMP_LOOP_COMP_LOOP_and_134_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[4:0]==5'b01011);
      COMP_LOOP_COMP_LOOP_and_10_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[0]) & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11)
          & (~((COMP_LOOP_acc_psp_sva_mx0w0[1]) | (VEC_LOOP_j_10_0_sva_9_0[2])));
      COMP_LOOP_COMP_LOOP_and_136_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[4:0]==5'b01101);
      COMP_LOOP_COMP_LOOP_and_12_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[0]) & (VEC_LOOP_j_10_0_sva_9_0[2])
          & (VEC_LOOP_j_10_0_sva_9_0[0]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[1]) |
          (VEC_LOOP_j_10_0_sva_9_0[1])));
      COMP_LOOP_COMP_LOOP_and_13_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[0]) & (VEC_LOOP_j_10_0_sva_9_0[2:1]==2'b11)
          & (~((COMP_LOOP_acc_psp_sva_mx0w0[1]) | (VEC_LOOP_j_10_0_sva_9_0[0])));
      COMP_LOOP_COMP_LOOP_and_14_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[0]) & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111)
          & (~ (COMP_LOOP_acc_psp_sva_mx0w0[1]));
      COMP_LOOP_COMP_LOOP_and_140_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[4:0]==5'b10001);
      COMP_LOOP_COMP_LOOP_and_141_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[4:0]==5'b10010);
      COMP_LOOP_COMP_LOOP_and_142_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[4:0]==5'b10011);
      COMP_LOOP_COMP_LOOP_and_18_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1]) & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11)
          & (~((COMP_LOOP_acc_psp_sva_mx0w0[0]) | (VEC_LOOP_j_10_0_sva_9_0[2])));
      COMP_LOOP_COMP_LOOP_and_144_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[4:0]==5'b10101);
      COMP_LOOP_COMP_LOOP_and_20_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1]) & (VEC_LOOP_j_10_0_sva_9_0[2])
          & (VEC_LOOP_j_10_0_sva_9_0[0]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[0]) |
          (VEC_LOOP_j_10_0_sva_9_0[1])));
      COMP_LOOP_COMP_LOOP_and_21_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1]) & (VEC_LOOP_j_10_0_sva_9_0[2:1]==2'b11)
          & (~((COMP_LOOP_acc_psp_sva_mx0w0[0]) | (VEC_LOOP_j_10_0_sva_9_0[0])));
      COMP_LOOP_COMP_LOOP_and_22_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1]) & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111)
          & (~ (COMP_LOOP_acc_psp_sva_mx0w0[0]));
      COMP_LOOP_COMP_LOOP_and_23_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b000);
      COMP_LOOP_COMP_LOOP_and_24_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b001);
      COMP_LOOP_COMP_LOOP_and_25_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b010);
      COMP_LOOP_COMP_LOOP_and_26_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b011);
      COMP_LOOP_COMP_LOOP_and_27_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b100);
      COMP_LOOP_COMP_LOOP_and_28_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b101);
      COMP_LOOP_COMP_LOOP_and_29_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b110);
      COMP_LOOP_COMP_LOOP_and_30_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_6_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_tmp_1459, mux_1492_nl, fsm_output[5]) ) begin
      COMP_LOOP_acc_1_cse_6_sva <= COMP_LOOP_acc_1_cse_6_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_4_sva <= 10'b0000000000;
    end
    else if ( mux_1497_nl | (fsm_output[7]) ) begin
      COMP_LOOP_acc_1_cse_4_sva <= COMP_LOOP_acc_1_cse_4_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_2_sva <= 10'b0000000000;
    end
    else if ( ~(mux_1499_nl & nor_1025_cse) ) begin
      COMP_LOOP_acc_1_cse_2_sva <= COMP_LOOP_acc_1_cse_2_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_2_sva <= 10'b0000000000;
    end
    else if ( ~(mux_1500_nl & nor_1025_cse) ) begin
      COMP_LOOP_acc_10_cse_10_1_2_sva <= COMP_LOOP_2_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( ~(mux_1502_nl & nor_1025_cse) ) begin
      COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_3_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_5_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_nor_5_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[4:0]!=5'b00000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_126_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_nor_126_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[4:1]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_127_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_nor_127_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[4]) | (COMP_LOOP_2_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[2]) | (COMP_LOOP_2_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_157_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_157_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b00011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_129_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_nor_129_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[4]) | (COMP_LOOP_2_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[1]) | (COMP_LOOP_2_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_159_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_159_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b00101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_160_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_160_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b00110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_161_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_161_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b00111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_133_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_nor_133_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[4]) | (COMP_LOOP_2_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[1]) | (COMP_LOOP_2_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_163_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_163_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b01001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_164_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_164_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b01010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_165_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_165_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b01011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_166_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_166_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b01100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_167_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_167_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b01101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_168_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_168_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b01110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_169_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_169_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b01111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_140_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_nor_140_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_171_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_171_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b10001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_172_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_172_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b10010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_173_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_173_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b10011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_174_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_174_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b10100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_175_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_175_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b10101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_176_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_176_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b10110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_177_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_177_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b10111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_178_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_178_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b11000);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_179_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_179_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b11001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_180_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_180_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b11010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_181_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_181_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b11011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_182_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_182_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b11100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_183_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_183_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b11101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_184_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_184_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b11110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_185_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_252 ) begin
      COMP_LOOP_COMP_LOOP_and_185_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[4:0]==5'b11111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_11_psp_sva <= 9'b000000000;
    end
    else if ( mux_1505_nl | (fsm_output[7]) ) begin
      COMP_LOOP_acc_11_psp_sva <= nl_COMP_LOOP_acc_11_psp_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_3_sva <= 10'b0000000000;
    end
    else if ( mux_1507_nl | (fsm_output[7]) ) begin
      COMP_LOOP_acc_10_cse_10_1_3_sva <= COMP_LOOP_3_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( mux_1509_nl | (fsm_output[7]) ) begin
      COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm <= readslicef_9_1_8(COMP_LOOP_acc_12_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_9_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_nor_9_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[4:0]!=5'b00000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_226_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_nor_226_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[4:1]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_227_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_nor_227_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[4]) | (COMP_LOOP_3_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_3_acc_10_itm_10_1_1[2]) | (COMP_LOOP_3_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_281_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_281_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b00011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_229_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_nor_229_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[4]) | (COMP_LOOP_3_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_3_acc_10_itm_10_1_1[1]) | (COMP_LOOP_3_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_283_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_283_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b00101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_284_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_284_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b00110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_285_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_285_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b00111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_233_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_nor_233_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[4]) | (COMP_LOOP_3_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_3_acc_10_itm_10_1_1[1]) | (COMP_LOOP_3_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_287_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_287_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b01001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_288_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_288_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b01010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_289_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_289_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b01011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_290_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_290_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b01100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_291_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_291_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b01101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_292_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_292_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b01110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_293_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_293_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b01111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_240_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_nor_240_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_295_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_295_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b10001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_296_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_296_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b10010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_297_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_297_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b10011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_298_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_298_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b10100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_299_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_299_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b10101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_300_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_300_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b10110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_301_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_301_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b10111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_302_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_302_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b11000);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_303_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_303_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b11001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_304_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_304_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b11010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_305_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_305_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b11011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_306_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_306_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b11100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_307_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_307_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b11101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_308_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_308_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b11110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_309_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_256 ) begin
      COMP_LOOP_COMP_LOOP_and_309_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[4:0]==5'b11111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_4_sva <= 10'b0000000000;
    end
    else if ( mux_1511_nl | (fsm_output[7]) ) begin
      COMP_LOOP_acc_10_cse_10_1_4_sva <= COMP_LOOP_4_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( mux_1513_nl | (fsm_output[7]) ) begin
      COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_5_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_13_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_nor_13_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[4:0]!=5'b00000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_326_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_nor_326_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[4:1]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_327_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_nor_327_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[4]) | (COMP_LOOP_4_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_4_acc_10_itm_10_1_1[2]) | (COMP_LOOP_4_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_405_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_405_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b00011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_329_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_nor_329_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[4]) | (COMP_LOOP_4_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_4_acc_10_itm_10_1_1[1]) | (COMP_LOOP_4_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_407_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_407_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b00101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_408_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_408_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b00110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_409_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_409_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b00111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_333_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_nor_333_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[4]) | (COMP_LOOP_4_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_4_acc_10_itm_10_1_1[1]) | (COMP_LOOP_4_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_411_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_411_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b01001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_412_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_412_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b01010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_413_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_413_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b01011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_414_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_414_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b01100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_415_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_415_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b01101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_416_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_416_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b01110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_417_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_417_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b01111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_340_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_nor_340_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_419_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_419_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b10001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_420_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_420_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b10010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_421_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_421_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b10011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_422_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_422_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b10100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_423_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_423_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b10101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_424_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_424_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b10110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_425_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_425_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b10111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_426_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_426_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b11000);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_427_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_427_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b11001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_428_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_428_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b11010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_429_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_429_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b11011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_430_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_430_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b11100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_431_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_431_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b11101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_432_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_432_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b11110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_433_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_259 ) begin
      COMP_LOOP_COMP_LOOP_and_433_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[4:0]==5'b11111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_13_psp_sva <= 8'b00000000;
    end
    else if ( MUX_s_1_2_2(mux_1518_nl, (fsm_output[7]), fsm_output[5]) ) begin
      COMP_LOOP_acc_13_psp_sva <= nl_COMP_LOOP_acc_13_psp_sva[7:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_5_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_1520_nl, (fsm_output[7]), fsm_output[5]) ) begin
      COMP_LOOP_acc_10_cse_10_1_5_sva <= COMP_LOOP_5_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_1523_nl, (fsm_output[7]), fsm_output[5]) ) begin
      COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_6_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_17_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_nor_17_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[4:0]!=5'b00000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_426_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_nor_426_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[4:1]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_427_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_nor_427_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[4]) | (COMP_LOOP_5_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[2]) | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_529_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_529_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b00011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_429_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_nor_429_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[4]) | (COMP_LOOP_5_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[1]) | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_531_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_531_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b00101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_532_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_532_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b00110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_533_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_533_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b00111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_433_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_nor_433_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[4]) | (COMP_LOOP_5_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[1]) | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_535_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_535_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b01001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_536_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_536_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b01010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_537_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_537_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b01011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_538_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_538_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b01100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_539_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_539_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b01101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_540_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_540_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b01110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_541_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_541_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b01111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_440_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_nor_440_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_543_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_543_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b10001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_544_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_544_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b10010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_545_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_545_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b10011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_546_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_546_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b10100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_547_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_547_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b10101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_548_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_548_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b10110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_549_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_549_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b10111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_550_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_550_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b11000);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_551_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_551_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b11001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_552_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_552_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b11010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_553_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_553_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b11011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_554_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_554_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b11100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_555_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_555_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b11101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_556_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_556_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b11110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_557_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_260 ) begin
      COMP_LOOP_COMP_LOOP_and_557_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[4:0]==5'b11111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_84 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_82_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_84 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_82_itm <= (z_out_7[2:0]==3'b011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_84_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_84 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_84_itm <= (z_out_7[2:0]==3'b101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_85_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_84 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_85_itm <= (z_out_7[2:0]==3'b110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_86_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_84 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_86_itm <= (z_out_7[2:0]==3'b111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_6_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_tmp_1459, and_491_cse, fsm_output[5]) ) begin
      COMP_LOOP_acc_10_cse_10_1_6_sva <= COMP_LOOP_6_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_tmp_1459, mux_1528_nl, fsm_output[5]) ) begin
      COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_7_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_21_itm <= 1'b0;
      COMP_LOOP_nor_526_itm <= 1'b0;
      COMP_LOOP_nor_527_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_653_itm <= 1'b0;
      COMP_LOOP_nor_529_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_655_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_656_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_657_itm <= 1'b0;
      COMP_LOOP_nor_533_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_659_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_660_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_661_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_662_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_663_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_664_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_665_itm <= 1'b0;
      COMP_LOOP_nor_540_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_667_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_668_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_669_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_670_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_671_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_672_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_673_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_674_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_675_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_676_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_677_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_678_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_679_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_680_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_681_itm <= 1'b0;
    end
    else if ( mux_1531_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_21_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[4:0]!=5'b00000));
      COMP_LOOP_nor_526_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[4:1]!=4'b0000));
      COMP_LOOP_nor_527_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[4]) | (COMP_LOOP_6_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[2]) | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_653_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b00011);
      COMP_LOOP_nor_529_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[4]) | (COMP_LOOP_6_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[1]) | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_655_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b00101);
      COMP_LOOP_COMP_LOOP_and_656_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b00110);
      COMP_LOOP_COMP_LOOP_and_657_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b00111);
      COMP_LOOP_nor_533_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[4]) | (COMP_LOOP_6_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[1]) | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_659_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b01001);
      COMP_LOOP_COMP_LOOP_and_660_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b01010);
      COMP_LOOP_COMP_LOOP_and_661_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b01011);
      COMP_LOOP_COMP_LOOP_and_662_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b01100);
      COMP_LOOP_COMP_LOOP_and_663_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b01101);
      COMP_LOOP_COMP_LOOP_and_664_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b01110);
      COMP_LOOP_COMP_LOOP_and_665_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b01111);
      COMP_LOOP_nor_540_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[3:0]!=4'b0000));
      COMP_LOOP_COMP_LOOP_and_667_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b10001);
      COMP_LOOP_COMP_LOOP_and_668_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b10010);
      COMP_LOOP_COMP_LOOP_and_669_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b10011);
      COMP_LOOP_COMP_LOOP_and_670_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b10100);
      COMP_LOOP_COMP_LOOP_and_671_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b10101);
      COMP_LOOP_COMP_LOOP_and_672_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b10110);
      COMP_LOOP_COMP_LOOP_and_673_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b10111);
      COMP_LOOP_COMP_LOOP_and_674_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b11000);
      COMP_LOOP_COMP_LOOP_and_675_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b11001);
      COMP_LOOP_COMP_LOOP_and_676_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b11010);
      COMP_LOOP_COMP_LOOP_and_677_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b11011);
      COMP_LOOP_COMP_LOOP_and_678_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b11100);
      COMP_LOOP_COMP_LOOP_and_679_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b11101);
      COMP_LOOP_COMP_LOOP_and_680_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b11110);
      COMP_LOOP_COMP_LOOP_and_681_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[4:0]==5'b11111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_14_psp_sva <= 9'b000000000;
    end
    else if ( MUX_s_1_2_2(mux_1532_nl, and_464_cse, fsm_output[5]) ) begin
      COMP_LOOP_acc_14_psp_sva <= nl_COMP_LOOP_acc_14_psp_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_7_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2((~ or_tmp_2048), and_464_cse, or_162_nl) ) begin
      COMP_LOOP_acc_10_cse_10_1_7_sva <= COMP_LOOP_7_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( mux_1536_itm ) begin
      COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm <= readslicef_8_1_7(COMP_LOOP_acc_15_nl);
      reg_COMP_LOOP_k_10_3_ftd <= z_out_2[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_25_itm <= 1'b0;
      COMP_LOOP_nor_626_itm <= 1'b0;
      COMP_LOOP_nor_627_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_777_itm <= 1'b0;
      COMP_LOOP_nor_629_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_779_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_780_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_781_itm <= 1'b0;
      COMP_LOOP_nor_633_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_783_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_784_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_785_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_786_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_787_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_788_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_789_itm <= 1'b0;
      COMP_LOOP_nor_640_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_791_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_792_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_793_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_794_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_795_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_796_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_797_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_798_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_799_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_800_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_801_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_802_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_803_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_804_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_805_itm <= 1'b0;
    end
    else if ( mux_1538_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_25_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[4:0]!=5'b00000));
      COMP_LOOP_nor_626_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[4:1]!=4'b0000));
      COMP_LOOP_nor_627_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[4]) | (COMP_LOOP_7_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[2]) | (COMP_LOOP_7_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_777_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b00011);
      COMP_LOOP_nor_629_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[4]) | (COMP_LOOP_7_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[1]) | (COMP_LOOP_7_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_779_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b00101);
      COMP_LOOP_COMP_LOOP_and_780_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b00110);
      COMP_LOOP_COMP_LOOP_and_781_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b00111);
      COMP_LOOP_nor_633_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[4]) | (COMP_LOOP_7_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[1]) | (COMP_LOOP_7_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_783_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b01001);
      COMP_LOOP_COMP_LOOP_and_784_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b01010);
      COMP_LOOP_COMP_LOOP_and_785_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b01011);
      COMP_LOOP_COMP_LOOP_and_786_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b01100);
      COMP_LOOP_COMP_LOOP_and_787_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b01101);
      COMP_LOOP_COMP_LOOP_and_788_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b01110);
      COMP_LOOP_COMP_LOOP_and_789_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b01111);
      COMP_LOOP_nor_640_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[3:0]!=4'b0000));
      COMP_LOOP_COMP_LOOP_and_791_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b10001);
      COMP_LOOP_COMP_LOOP_and_792_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b10010);
      COMP_LOOP_COMP_LOOP_and_793_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b10011);
      COMP_LOOP_COMP_LOOP_and_794_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b10100);
      COMP_LOOP_COMP_LOOP_and_795_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b10101);
      COMP_LOOP_COMP_LOOP_and_796_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b10110);
      COMP_LOOP_COMP_LOOP_and_797_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b10111);
      COMP_LOOP_COMP_LOOP_and_798_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b11000);
      COMP_LOOP_COMP_LOOP_and_799_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b11001);
      COMP_LOOP_COMP_LOOP_and_800_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b11010);
      COMP_LOOP_COMP_LOOP_and_801_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b11011);
      COMP_LOOP_COMP_LOOP_and_802_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b11100);
      COMP_LOOP_COMP_LOOP_and_803_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b11101);
      COMP_LOOP_COMP_LOOP_and_804_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b11110);
      COMP_LOOP_COMP_LOOP_and_805_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[4:0]==5'b11111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_717, and_305_nl, fsm_output[5]) ) begin
      COMP_LOOP_acc_1_cse_sva <= nl_COMP_LOOP_acc_1_cse_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_717, and_464_cse, fsm_output[5]) ) begin
      COMP_LOOP_acc_10_cse_10_1_sva <= COMP_LOOP_8_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(not_tmp_717, and_304_nl, fsm_output[5]) ) begin
      COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_1_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_29_itm <= 1'b0;
      COMP_LOOP_nor_726_itm <= 1'b0;
      COMP_LOOP_nor_727_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_901_itm <= 1'b0;
      COMP_LOOP_nor_729_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_903_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_904_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_905_itm <= 1'b0;
      COMP_LOOP_nor_733_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_907_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_908_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_909_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_910_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_911_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_912_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_913_itm <= 1'b0;
      COMP_LOOP_nor_740_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_915_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_916_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_917_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_918_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_919_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_920_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_921_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_922_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_923_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_924_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_925_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_926_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_927_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_928_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_929_itm <= 1'b0;
    end
    else if ( mux_1543_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_29_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[4:0]!=5'b00000));
      COMP_LOOP_nor_726_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[4:1]!=4'b0000));
      COMP_LOOP_nor_727_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[4]) | (COMP_LOOP_8_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[2]) | (COMP_LOOP_8_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_901_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b00011);
      COMP_LOOP_nor_729_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[4]) | (COMP_LOOP_8_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[1]) | (COMP_LOOP_8_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_903_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b00101);
      COMP_LOOP_COMP_LOOP_and_904_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b00110);
      COMP_LOOP_COMP_LOOP_and_905_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b00111);
      COMP_LOOP_nor_733_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[4]) | (COMP_LOOP_8_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[1]) | (COMP_LOOP_8_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_907_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b01001);
      COMP_LOOP_COMP_LOOP_and_908_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b01010);
      COMP_LOOP_COMP_LOOP_and_909_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b01011);
      COMP_LOOP_COMP_LOOP_and_910_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b01100);
      COMP_LOOP_COMP_LOOP_and_911_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b01101);
      COMP_LOOP_COMP_LOOP_and_912_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b01110);
      COMP_LOOP_COMP_LOOP_and_913_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b01111);
      COMP_LOOP_nor_740_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[3:0]!=4'b0000));
      COMP_LOOP_COMP_LOOP_and_915_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b10001);
      COMP_LOOP_COMP_LOOP_and_916_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b10010);
      COMP_LOOP_COMP_LOOP_and_917_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b10011);
      COMP_LOOP_COMP_LOOP_and_918_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b10100);
      COMP_LOOP_COMP_LOOP_and_919_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b10101);
      COMP_LOOP_COMP_LOOP_and_920_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b10110);
      COMP_LOOP_COMP_LOOP_and_921_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b10111);
      COMP_LOOP_COMP_LOOP_and_922_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b11000);
      COMP_LOOP_COMP_LOOP_and_923_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b11001);
      COMP_LOOP_COMP_LOOP_and_924_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b11010);
      COMP_LOOP_COMP_LOOP_and_925_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b11011);
      COMP_LOOP_COMP_LOOP_and_926_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b11100);
      COMP_LOOP_COMP_LOOP_and_927_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b11101);
      COMP_LOOP_COMP_LOOP_and_928_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b11110);
      COMP_LOOP_COMP_LOOP_and_929_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[4:0]==5'b11111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm <= 1'b0;
    end
    else if ( COMP_LOOP_tmp_or_cse ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_33_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_36_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse,
          {and_dcpl_46 , and_dcpl_49 , and_dcpl_171 , COMP_LOOP_or_59_cse , and_dcpl_173});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_35_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_38_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_cse,
          {and_dcpl_46 , and_dcpl_49 , and_dcpl_171 , COMP_LOOP_or_59_cse , and_dcpl_173});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_36_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_39_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse,
          {and_dcpl_46 , and_dcpl_49 , and_dcpl_171 , COMP_LOOP_or_59_cse , and_dcpl_173});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_37_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_40_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_cse,
          {and_dcpl_46 , and_dcpl_49 , and_dcpl_171 , COMP_LOOP_or_59_cse , and_dcpl_173});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_39_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_42_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_cse,
          {and_dcpl_46 , and_dcpl_49 , and_dcpl_171 , COMP_LOOP_or_59_cse , and_dcpl_173});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_40_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_43_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_cse,
          {and_dcpl_46 , and_dcpl_49 , and_dcpl_171 , COMP_LOOP_or_59_cse , and_dcpl_173});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_41_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_44_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_cse,
          {and_dcpl_46 , and_dcpl_49 , and_dcpl_171 , COMP_LOOP_or_59_cse , and_dcpl_173});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_42_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_45_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_cse,
          {and_dcpl_46 , and_dcpl_49 , and_dcpl_171 , COMP_LOOP_or_59_cse , and_dcpl_173});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_43_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_46_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_cse,
          {and_dcpl_46 , and_dcpl_49 , and_dcpl_171 , COMP_LOOP_or_59_cse , and_dcpl_173});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_44_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_47_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse,
          {and_dcpl_46 , and_dcpl_49 , and_dcpl_171 , COMP_LOOP_or_59_cse , and_dcpl_173});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_45_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_48_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_cse,
          {and_dcpl_46 , and_dcpl_49 , and_dcpl_171 , COMP_LOOP_or_59_cse , and_dcpl_173});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_47_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_cse,
          {and_dcpl_46 , and_dcpl_49 , and_dcpl_171 , COMP_LOOP_or_59_cse , and_dcpl_173});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm <= 1'b0;
      COMP_LOOP_tmp_nor_1_itm <= 1'b0;
      COMP_LOOP_tmp_nor_14_itm <= 1'b0;
      COMP_LOOP_tmp_nor_3_itm <= 1'b0;
      COMP_LOOP_tmp_nor_42_itm <= 1'b0;
      COMP_LOOP_tmp_nor_49_itm <= 1'b0;
    end
    else if ( COMP_LOOP_tmp_or_12_cse ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_48_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_cse, {and_dcpl_46 , and_dcpl_49 , COMP_LOOP_or_59_cse
          , and_dcpl_173});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_49_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_cse, {and_dcpl_46 , and_dcpl_49 , COMP_LOOP_or_59_cse
          , and_dcpl_173});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_50_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_cse, {and_dcpl_46 , and_dcpl_49 , COMP_LOOP_or_59_cse
          , and_dcpl_173});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_51_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_cse, {and_dcpl_46 , and_dcpl_49 , COMP_LOOP_or_59_cse
          , and_dcpl_173});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_52_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_cse, {and_dcpl_46 , and_dcpl_49 , COMP_LOOP_or_59_cse
          , and_dcpl_173});
      COMP_LOOP_tmp_nor_1_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_26_nl, COMP_LOOP_tmp_nor_1_cse,
          COMP_LOOP_tmp_nor_35_cse, COMP_LOOP_tmp_nor_101_cse, {and_dcpl_46 , and_dcpl_49
          , COMP_LOOP_or_41_cse , and_dcpl_176});
      COMP_LOOP_tmp_nor_14_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_27_nl, COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse,
          COMP_LOOP_tmp_nor_1_cse, COMP_LOOP_tmp_nor_105_cse, {and_dcpl_46 , and_dcpl_49
          , COMP_LOOP_or_41_cse , and_dcpl_176});
      COMP_LOOP_tmp_nor_3_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_nor_29_nl, COMP_LOOP_tmp_nor_101_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse, {and_dcpl_46 , COMP_LOOP_or_39_cse
          , and_dcpl_176});
      COMP_LOOP_tmp_nor_42_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_nor_33_nl, COMP_LOOP_tmp_nor_105_cse,
          COMP_LOOP_tmp_nor_35_cse, {and_dcpl_46 , COMP_LOOP_or_39_cse , and_dcpl_176});
      COMP_LOOP_tmp_nor_49_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_40_nl, COMP_LOOP_tmp_nor_35_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse, COMP_LOOP_tmp_nor_1_cse, {and_dcpl_46
          , and_dcpl_49 , COMP_LOOP_or_41_cse , and_dcpl_176});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_122_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_123_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_124_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_126_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_127_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_128_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_129_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_130_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_131_itm <= 1'b0;
    end
    else if ( COMP_LOOP_tmp_or_17_cse ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_53_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_36_cse, {and_dcpl_46 , and_dcpl_49 , and_dcpl_172
          , and_dcpl_174});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_122_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_54_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_38_cse, {and_dcpl_46 , and_dcpl_49 , and_dcpl_172
          , and_dcpl_174});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_123_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_55_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_39_cse, {and_dcpl_46 , and_dcpl_49 , and_dcpl_172
          , and_dcpl_174});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_124_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_56_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_40_cse, {and_dcpl_46 , and_dcpl_49 , and_dcpl_172
          , and_dcpl_174});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_126_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_57_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_42_cse, {and_dcpl_46 , and_dcpl_49 , and_dcpl_172
          , and_dcpl_174});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_127_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_58_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_43_cse, {and_dcpl_46 , and_dcpl_49 , and_dcpl_172
          , and_dcpl_174});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_128_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_59_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_44_cse, {and_dcpl_46 , and_dcpl_49 , and_dcpl_172
          , and_dcpl_174});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_129_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_60_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_45_cse, {and_dcpl_46 , and_dcpl_49 , and_dcpl_172
          , and_dcpl_174});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_130_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_61_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_46_cse, {and_dcpl_46 , and_dcpl_49 , and_dcpl_172
          , and_dcpl_174});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_131_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_nor_1_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_47_cse,
          {and_dcpl_46 , COMP_LOOP_or_42_cse , and_dcpl_174});
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_mux1h_itm_mx0c0 | COMP_LOOP_tmp_mux1h_itm_mx0c1 | COMP_LOOP_tmp_mux1h_itm_mx0c2
        | COMP_LOOP_tmp_mux1h_itm_mx0c3 ) begin
      COMP_LOOP_tmp_mux1h_itm <= MUX1HOT_v_64_4_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_8_i_q_d,
          twiddle_rsc_0_16_i_q_d, twiddle_rsc_0_24_i_q_d, {COMP_LOOP_tmp_mux1h_itm_mx0c0
          , COMP_LOOP_tmp_mux1h_itm_mx0c1 , COMP_LOOP_tmp_mux1h_itm_mx0c2 , COMP_LOOP_tmp_mux1h_itm_mx0c3});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_2_tmp_mul_idiv_sva <= 10'b0000000000;
    end
    else if ( COMP_LOOP_or_39_cse ) begin
      COMP_LOOP_2_tmp_mul_idiv_sva <= z_out_7;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_2_tmp_lshift_ncse_sva <= 10'b0000000000;
    end
    else if ( and_dcpl_49 | and_dcpl_176 ) begin
      COMP_LOOP_2_tmp_lshift_ncse_sva <= MUX_v_10_2_2(z_out_1, z_out_7, and_dcpl_176);
    end
  end
  always @(posedge clk) begin
    if ( and_dcpl_49 | and_dcpl_171 | and_dcpl_278 | and_dcpl_176 | COMP_LOOP_1_acc_8_itm_mx0c4
        | and_dcpl_54 | and_dcpl_222 | and_dcpl_58 | and_dcpl_226 | and_dcpl_65 |
        and_dcpl_229 | and_dcpl_68 | and_dcpl_232 | and_dcpl_75 | and_dcpl_234 |
        and_dcpl_78 | and_dcpl_236 | and_dcpl_83 | and_dcpl_238 ) begin
      COMP_LOOP_1_acc_8_itm <= MUX1HOT_v_64_36_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d,
          vec_rsc_0_2_i_q_d, vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d,
          vec_rsc_0_6_i_q_d, vec_rsc_0_7_i_q_d, vec_rsc_0_8_i_q_d, vec_rsc_0_9_i_q_d,
          vec_rsc_0_10_i_q_d, vec_rsc_0_11_i_q_d, vec_rsc_0_12_i_q_d, vec_rsc_0_13_i_q_d,
          vec_rsc_0_14_i_q_d, vec_rsc_0_15_i_q_d, vec_rsc_0_16_i_q_d, vec_rsc_0_17_i_q_d,
          vec_rsc_0_18_i_q_d, vec_rsc_0_19_i_q_d, vec_rsc_0_20_i_q_d, vec_rsc_0_21_i_q_d,
          vec_rsc_0_22_i_q_d, vec_rsc_0_23_i_q_d, vec_rsc_0_24_i_q_d, vec_rsc_0_25_i_q_d,
          vec_rsc_0_26_i_q_d, vec_rsc_0_27_i_q_d, vec_rsc_0_28_i_q_d, vec_rsc_0_29_i_q_d,
          vec_rsc_0_30_i_q_d, vec_rsc_0_31_i_q_d, COMP_LOOP_acc_17_nl, twiddle_rsc_0_10_i_q_d,
          twiddle_rsc_0_26_i_q_d, COMP_LOOP_1_modulo_dev_cmp_return_rsc_z, {COMP_LOOP_or_nl
          , COMP_LOOP_or_1_nl , COMP_LOOP_or_2_nl , COMP_LOOP_or_3_nl , COMP_LOOP_or_4_nl
          , COMP_LOOP_or_5_nl , COMP_LOOP_or_6_nl , COMP_LOOP_or_7_nl , COMP_LOOP_or_8_nl
          , COMP_LOOP_or_9_nl , COMP_LOOP_or_10_nl , COMP_LOOP_or_11_nl , COMP_LOOP_or_12_nl
          , COMP_LOOP_or_13_nl , COMP_LOOP_or_14_nl , COMP_LOOP_or_15_nl , COMP_LOOP_or_16_nl
          , COMP_LOOP_or_17_nl , COMP_LOOP_or_18_nl , COMP_LOOP_or_19_nl , COMP_LOOP_or_20_nl
          , COMP_LOOP_or_21_nl , COMP_LOOP_or_22_nl , COMP_LOOP_or_23_nl , COMP_LOOP_or_24_nl
          , COMP_LOOP_or_25_nl , COMP_LOOP_or_26_nl , COMP_LOOP_or_27_nl , COMP_LOOP_or_28_nl
          , COMP_LOOP_or_29_nl , COMP_LOOP_or_30_nl , COMP_LOOP_or_31_nl , COMP_LOOP_or_36_itm
          , and_dcpl_278 , and_dcpl_176 , COMP_LOOP_1_acc_8_itm_mx0c4});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_3_tmp_lshift_ncse_sva <= 9'b000000000;
      COMP_LOOP_tmp_nor_25_itm <= 1'b0;
      COMP_LOOP_tmp_nor_26_itm <= 1'b0;
      COMP_LOOP_tmp_nor_28_itm <= 1'b0;
      COMP_LOOP_tmp_nor_31_itm <= 1'b0;
    end
    else if ( COMP_LOOP_tmp_or_35_cse ) begin
      COMP_LOOP_3_tmp_lshift_ncse_sva <= MUX_v_9_2_2((z_out_1[8:0]), (z_out_7[8:0]),
          and_dcpl_174);
      COMP_LOOP_tmp_nor_25_itm <= COMP_LOOP_tmp_nor_78_cse;
      COMP_LOOP_tmp_nor_26_itm <= COMP_LOOP_tmp_nor_79_cse;
      COMP_LOOP_tmp_nor_28_itm <= COMP_LOOP_tmp_nor_81_cse;
      COMP_LOOP_tmp_nor_31_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse;
    end
  end
  always @(posedge clk) begin
    if ( ~ and_294_tmp ) begin
      COMP_LOOP_tmp_mux1h_1_itm <= MUX1HOT_v_64_32_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_1_i_q_d,
          twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_3_i_q_d, twiddle_rsc_0_4_i_q_d, twiddle_rsc_0_5_i_q_d,
          twiddle_rsc_0_6_i_q_d, twiddle_rsc_0_7_i_q_d, twiddle_rsc_0_8_i_q_d, twiddle_rsc_0_9_i_q_d,
          twiddle_rsc_0_10_i_q_d, twiddle_rsc_0_11_i_q_d, twiddle_rsc_0_12_i_q_d,
          twiddle_rsc_0_13_i_q_d, twiddle_rsc_0_14_i_q_d, twiddle_rsc_0_15_i_q_d,
          twiddle_rsc_0_16_i_q_d, twiddle_rsc_0_17_i_q_d, twiddle_rsc_0_18_i_q_d,
          twiddle_rsc_0_19_i_q_d, twiddle_rsc_0_20_i_q_d, twiddle_rsc_0_21_i_q_d,
          twiddle_rsc_0_22_i_q_d, twiddle_rsc_0_23_i_q_d, twiddle_rsc_0_24_i_q_d,
          twiddle_rsc_0_25_i_q_d, twiddle_rsc_0_26_i_q_d, twiddle_rsc_0_27_i_q_d,
          twiddle_rsc_0_28_i_q_d, twiddle_rsc_0_29_i_q_d, twiddle_rsc_0_30_i_q_d,
          twiddle_rsc_0_31_i_q_d, {COMP_LOOP_tmp_and_127_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl
          , COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_nl , COMP_LOOP_tmp_and_128_nl , COMP_LOOP_tmp_and_129_nl
          , COMP_LOOP_tmp_and_130_nl , COMP_LOOP_tmp_and_131_nl , COMP_LOOP_tmp_and_132_nl
          , COMP_LOOP_tmp_and_133_nl , COMP_LOOP_tmp_and_134_nl , COMP_LOOP_tmp_and_135_nl
          , COMP_LOOP_tmp_and_136_nl , COMP_LOOP_tmp_and_137_nl , COMP_LOOP_tmp_and_138_nl
          , COMP_LOOP_tmp_and_139_nl , COMP_LOOP_tmp_and_140_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_18_nl
          , COMP_LOOP_tmp_and_141_nl , COMP_LOOP_tmp_and_142_nl , COMP_LOOP_tmp_and_143_nl
          , COMP_LOOP_tmp_and_144_nl , COMP_LOOP_tmp_and_145_nl , COMP_LOOP_tmp_and_146_nl
          , COMP_LOOP_tmp_and_147_nl , COMP_LOOP_tmp_and_148_nl , COMP_LOOP_tmp_and_149_nl
          , COMP_LOOP_tmp_and_150_nl , COMP_LOOP_tmp_and_151_nl , COMP_LOOP_tmp_and_152_nl
          , COMP_LOOP_tmp_and_153_nl , COMP_LOOP_tmp_and_154_nl , COMP_LOOP_tmp_and_155_nl});
    end
  end
  always @(posedge clk) begin
    if ( ~ nor_1119_tmp ) begin
      COMP_LOOP_tmp_mux1h_2_itm <= MUX1HOT_v_64_16_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_2_i_q_d,
          twiddle_rsc_0_4_i_q_d, twiddle_rsc_0_6_i_q_d, twiddle_rsc_0_8_i_q_d, twiddle_rsc_0_10_i_q_d,
          twiddle_rsc_0_12_i_q_d, twiddle_rsc_0_14_i_q_d, twiddle_rsc_0_16_i_q_d,
          twiddle_rsc_0_18_i_q_d, twiddle_rsc_0_20_i_q_d, twiddle_rsc_0_22_i_q_d,
          twiddle_rsc_0_24_i_q_d, twiddle_rsc_0_26_i_q_d, twiddle_rsc_0_28_i_q_d,
          twiddle_rsc_0_30_i_q_d, {COMP_LOOP_tmp_and_115_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_34_nl
          , COMP_LOOP_tmp_COMP_LOOP_tmp_and_35_nl , COMP_LOOP_tmp_and_116_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_37_nl
          , COMP_LOOP_tmp_and_117_nl , COMP_LOOP_tmp_and_118_nl , COMP_LOOP_tmp_and_119_nl
          , COMP_LOOP_tmp_COMP_LOOP_tmp_and_41_nl , COMP_LOOP_tmp_and_120_nl , COMP_LOOP_tmp_and_121_nl
          , COMP_LOOP_tmp_and_122_nl , COMP_LOOP_tmp_and_123_nl , COMP_LOOP_tmp_and_124_nl
          , COMP_LOOP_tmp_and_125_nl , COMP_LOOP_tmp_and_126_nl});
    end
  end
  always @(posedge clk) begin
    if ( ~ nor_tmp ) begin
      COMP_LOOP_tmp_mux1h_3_itm <= MUX1HOT_v_64_32_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_1_i_q_d,
          twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_3_i_q_d, twiddle_rsc_0_4_i_q_d, twiddle_rsc_0_5_i_q_d,
          twiddle_rsc_0_6_i_q_d, twiddle_rsc_0_7_i_q_d, twiddle_rsc_0_8_i_q_d, twiddle_rsc_0_9_i_q_d,
          twiddle_rsc_0_10_i_q_d, twiddle_rsc_0_11_i_q_d, twiddle_rsc_0_12_i_q_d,
          twiddle_rsc_0_13_i_q_d, twiddle_rsc_0_14_i_q_d, twiddle_rsc_0_15_i_q_d,
          twiddle_rsc_0_16_i_q_d, twiddle_rsc_0_17_i_q_d, twiddle_rsc_0_18_i_q_d,
          twiddle_rsc_0_19_i_q_d, twiddle_rsc_0_20_i_q_d, twiddle_rsc_0_21_i_q_d,
          twiddle_rsc_0_22_i_q_d, twiddle_rsc_0_23_i_q_d, twiddle_rsc_0_24_i_q_d,
          twiddle_rsc_0_25_i_q_d, twiddle_rsc_0_26_i_q_d, twiddle_rsc_0_27_i_q_d,
          twiddle_rsc_0_28_i_q_d, twiddle_rsc_0_29_i_q_d, twiddle_rsc_0_30_i_q_d,
          twiddle_rsc_0_31_i_q_d, {COMP_LOOP_tmp_and_83_nl , COMP_LOOP_tmp_and_84_nl
          , COMP_LOOP_tmp_and_85_nl , COMP_LOOP_tmp_and_86_nl , COMP_LOOP_tmp_and_87_nl
          , COMP_LOOP_tmp_and_88_nl , COMP_LOOP_tmp_and_89_nl , COMP_LOOP_tmp_and_90_nl
          , COMP_LOOP_tmp_and_91_nl , COMP_LOOP_tmp_and_92_nl , COMP_LOOP_tmp_and_93_nl
          , COMP_LOOP_tmp_and_94_nl , COMP_LOOP_tmp_and_95_nl , COMP_LOOP_tmp_and_96_nl
          , COMP_LOOP_tmp_and_97_nl , COMP_LOOP_tmp_and_98_nl , COMP_LOOP_tmp_and_99_nl
          , COMP_LOOP_tmp_and_100_nl , COMP_LOOP_tmp_and_101_nl , COMP_LOOP_tmp_and_102_nl
          , COMP_LOOP_tmp_and_103_nl , COMP_LOOP_tmp_and_104_nl , COMP_LOOP_tmp_and_105_nl
          , COMP_LOOP_tmp_and_106_nl , COMP_LOOP_tmp_and_107_nl , COMP_LOOP_tmp_and_108_nl
          , COMP_LOOP_tmp_and_109_nl , COMP_LOOP_tmp_and_110_nl , COMP_LOOP_tmp_and_111_nl
          , COMP_LOOP_tmp_and_112_nl , COMP_LOOP_tmp_and_113_nl , COMP_LOOP_tmp_and_114_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm <= 1'b0;
    end
    else if ( COMP_LOOP_tmp_or_40_cse ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_cse;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_cse, and_dcpl_176);
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse, and_dcpl_176);
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_cse, and_dcpl_176);
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_cse, and_dcpl_176);
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_cse, and_dcpl_176);
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_cse, and_dcpl_176);
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_cse, and_dcpl_176);
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_cse, and_dcpl_176);
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_cse, and_dcpl_176);
    end
  end
  always @(posedge clk) begin
    if ( ~ nor_1117_tmp ) begin
      COMP_LOOP_tmp_mux1h_4_itm <= MUX1HOT_v_64_8_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_4_i_q_d,
          twiddle_rsc_0_8_i_q_d, twiddle_rsc_0_12_i_q_d, twiddle_rsc_0_16_i_q_d,
          twiddle_rsc_0_20_i_q_d, twiddle_rsc_0_24_i_q_d, twiddle_rsc_0_28_i_q_d,
          {COMP_LOOP_tmp_and_78_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_80_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_81_nl
          , COMP_LOOP_tmp_and_79_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_83_nl , COMP_LOOP_tmp_and_80_nl
          , COMP_LOOP_tmp_and_81_nl , COMP_LOOP_tmp_and_82_nl});
    end
  end
  always @(posedge clk) begin
    if ( ((~((COMP_LOOP_2_tmp_lshift_ncse_sva[0]) & COMP_LOOP_tmp_nor_42_itm)) |
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_rgt
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_rgt
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_rgt
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_rgt
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm | and_dcpl_278 | and_dcpl_176)
        & mux_1585_nl ) begin
      tmp_21_sva_1 <= MUX1HOT_v_64_33_2(twiddle_rsc_0_1_i_q_d, twiddle_rsc_0_22_i_q_d,
          twiddle_rsc_0_0_i_q_d, tmp_21_sva_2, tmp_21_sva_3, twiddle_rsc_0_4_i_q_d,
          tmp_21_sva_5, tmp_21_sva_6, tmp_21_sva_7, twiddle_rsc_0_8_i_q_d, tmp_21_sva_9,
          COMP_LOOP_1_acc_8_itm, tmp_21_sva_11, twiddle_rsc_0_12_i_q_d, tmp_21_sva_13,
          tmp_21_sva_14, tmp_21_sva_15, twiddle_rsc_0_16_i_q_d, tmp_21_sva_17, tmp_21_sva_18,
          tmp_21_sva_19, twiddle_rsc_0_20_i_q_d, tmp_21_sva_21, tmp_21_sva_22, tmp_21_sva_23,
          twiddle_rsc_0_24_i_q_d, tmp_21_sva_25, tmp_21_sva_26, tmp_21_sva_27, twiddle_rsc_0_28_i_q_d,
          tmp_21_sva_29, tmp_21_sva_30, tmp_21_sva_31, {and_dcpl_278 , and_dcpl_176
          , COMP_LOOP_tmp_and_47_nl , COMP_LOOP_tmp_and_48_nl , COMP_LOOP_tmp_and_49_nl
          , COMP_LOOP_tmp_and_50_nl , COMP_LOOP_tmp_and_51_nl , COMP_LOOP_tmp_and_52_nl
          , COMP_LOOP_tmp_and_53_nl , COMP_LOOP_tmp_and_54_nl , COMP_LOOP_tmp_and_55_nl
          , COMP_LOOP_tmp_and_56_nl , COMP_LOOP_tmp_and_57_nl , COMP_LOOP_tmp_and_58_nl
          , COMP_LOOP_tmp_and_59_nl , COMP_LOOP_tmp_and_60_nl , COMP_LOOP_tmp_and_61_nl
          , COMP_LOOP_tmp_and_62_nl , COMP_LOOP_tmp_and_63_nl , COMP_LOOP_tmp_and_64_nl
          , COMP_LOOP_tmp_and_65_nl , COMP_LOOP_tmp_and_66_nl , COMP_LOOP_tmp_and_67_nl
          , COMP_LOOP_tmp_and_68_nl , COMP_LOOP_tmp_and_69_nl , COMP_LOOP_tmp_and_70_nl
          , COMP_LOOP_tmp_and_71_nl , COMP_LOOP_tmp_and_72_nl , COMP_LOOP_tmp_and_73_nl
          , COMP_LOOP_tmp_and_74_nl , COMP_LOOP_tmp_and_75_nl , COMP_LOOP_tmp_and_76_nl
          , COMP_LOOP_tmp_and_77_nl});
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm
        ) begin
      tmp_21_sva_3 <= twiddle_rsc_0_3_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm
        ) begin
      tmp_21_sva_5 <= twiddle_rsc_0_5_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm
        ) begin
      tmp_21_sva_7 <= twiddle_rsc_0_7_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm
        ) begin
      tmp_21_sva_9 <= twiddle_rsc_0_9_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm
        ) begin
      tmp_21_sva_19 <= twiddle_rsc_0_19_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm
        ) begin
      tmp_21_sva_21 <= twiddle_rsc_0_21_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm
        ) begin
      tmp_21_sva_23 <= twiddle_rsc_0_23_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm
        ) begin
      tmp_21_sva_25 <= twiddle_rsc_0_25_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm
        ) begin
      tmp_21_sva_27 <= twiddle_rsc_0_27_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm
        ) begin
      tmp_21_sva_29 <= twiddle_rsc_0_29_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm
        ) begin
      tmp_21_sva_31 <= twiddle_rsc_0_31_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_109 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_132_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_109 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_132_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_48_cse;
    end
  end
  always @(posedge clk) begin
    if ( mux_1592_tmp ) begin
      COMP_LOOP_tmp_mux1h_5_itm <= MUX1HOT_v_64_32_2(twiddle_rsc_0_0_i_q_d, tmp_21_sva_1,
          tmp_21_sva_2, tmp_21_sva_3, twiddle_rsc_0_4_i_q_d, tmp_21_sva_5, tmp_21_sva_6,
          tmp_21_sva_7, twiddle_rsc_0_8_i_q_d, tmp_21_sva_9, COMP_LOOP_1_acc_8_itm,
          tmp_21_sva_11, twiddle_rsc_0_12_i_q_d, tmp_21_sva_13, tmp_21_sva_14, tmp_21_sva_15,
          twiddle_rsc_0_16_i_q_d, tmp_21_sva_17, tmp_21_sva_18, tmp_21_sva_19, twiddle_rsc_0_20_i_q_d,
          tmp_21_sva_21, tmp_21_sva_22, tmp_21_sva_23, twiddle_rsc_0_24_i_q_d, tmp_21_sva_25,
          tmp_21_sva_26, tmp_21_sva_27, twiddle_rsc_0_28_i_q_d, tmp_21_sva_29, tmp_21_sva_30,
          tmp_21_sva_31, {COMP_LOOP_tmp_and_15_nl , COMP_LOOP_tmp_and_16_nl , COMP_LOOP_tmp_and_17_nl
          , COMP_LOOP_tmp_and_18_nl , COMP_LOOP_tmp_and_19_nl , COMP_LOOP_tmp_and_20_nl
          , COMP_LOOP_tmp_and_21_nl , COMP_LOOP_tmp_and_22_nl , COMP_LOOP_tmp_and_23_nl
          , COMP_LOOP_tmp_and_24_nl , COMP_LOOP_tmp_and_25_nl , COMP_LOOP_tmp_and_26_nl
          , COMP_LOOP_tmp_and_27_nl , COMP_LOOP_tmp_and_28_nl , COMP_LOOP_tmp_and_29_nl
          , COMP_LOOP_tmp_and_30_nl , COMP_LOOP_tmp_and_31_nl , COMP_LOOP_tmp_and_32_nl
          , COMP_LOOP_tmp_and_33_nl , COMP_LOOP_tmp_and_34_nl , COMP_LOOP_tmp_and_35_nl
          , COMP_LOOP_tmp_and_36_nl , COMP_LOOP_tmp_and_37_nl , COMP_LOOP_tmp_and_38_nl
          , COMP_LOOP_tmp_and_39_nl , COMP_LOOP_tmp_and_40_nl , COMP_LOOP_tmp_and_41_nl
          , COMP_LOOP_tmp_and_42_nl , COMP_LOOP_tmp_and_43_nl , COMP_LOOP_tmp_and_44_nl
          , COMP_LOOP_tmp_and_45_nl , COMP_LOOP_tmp_and_46_nl});
    end
  end
  always @(posedge clk) begin
    if ( ((~((COMP_LOOP_3_tmp_lshift_ncse_sva[0]) & COMP_LOOP_tmp_nor_25_itm)) |
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_119_rgt
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_121_rgt
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_122_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_123_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_124_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_125_rgt
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_126_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_127_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_128_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_129_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_130_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_131_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_132_itm | and_dcpl_176) & mux_1597_nl )
        begin
      COMP_LOOP_tmp_mux1h_6_itm <= MUX1HOT_v_64_16_2(twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_0_i_q_d,
          twiddle_rsc_0_4_i_q_d, tmp_21_sva_13, twiddle_rsc_0_8_i_q_d, tmp_21_sva_14,
          twiddle_rsc_0_12_i_q_d, tmp_21_sva_15, twiddle_rsc_0_16_i_q_d, tmp_21_sva_17,
          twiddle_rsc_0_20_i_q_d, tmp_21_sva_1, twiddle_rsc_0_24_i_q_d, COMP_LOOP_1_acc_8_itm,
          twiddle_rsc_0_28_i_q_d, tmp_21_sva_11, {and_dcpl_176 , COMP_LOOP_tmp_and_nl
          , COMP_LOOP_tmp_and_1_nl , COMP_LOOP_tmp_and_2_nl , COMP_LOOP_tmp_and_3_nl
          , COMP_LOOP_tmp_and_4_nl , COMP_LOOP_tmp_and_5_nl , COMP_LOOP_tmp_and_6_nl
          , COMP_LOOP_tmp_and_7_nl , COMP_LOOP_tmp_and_8_nl , COMP_LOOP_tmp_and_9_nl
          , COMP_LOOP_tmp_and_10_nl , COMP_LOOP_tmp_and_11_nl , COMP_LOOP_tmp_and_12_nl
          , COMP_LOOP_tmp_and_13_nl , COMP_LOOP_tmp_and_14_nl});
    end
  end
  assign nor_1019_nl = ~((fsm_output[2]) | (fsm_output[4]) | (fsm_output[3]) | (fsm_output[0])
      | (fsm_output[1]) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_320_nl = MUX_s_1_2_2(and_33_cse, nor_tmp_95, fsm_output[2]);
  assign VEC_LOOP_j_not_1_nl = ~ VEC_LOOP_j_10_0_sva_9_0_mx0c0;
  assign nor_1160_nl = ~((fsm_output[2]) | (fsm_output[4]) | (fsm_output[3]) | (fsm_output[1])
      | (fsm_output[6]) | (fsm_output[7]));
  assign and_nl = or_220_cse & (fsm_output[7:6]==2'b11);
  assign nor_1021_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[7]));
  assign and_451_nl = (fsm_output[1]) & (fsm_output[6]) & (fsm_output[7]);
  assign mux_312_nl = MUX_s_1_2_2(nor_1021_nl, and_451_nl, fsm_output[5]);
  assign nand_nl = ~(mux_312_nl & and_dcpl_244 & nor_1023_cse);
  assign or_2285_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[5]) | (fsm_output[4])
      | (fsm_output[3]);
  assign mux_1604_nl = MUX_s_1_2_2(or_2285_nl, mux_tmp_1564, fsm_output[6]);
  assign or_2284_nl = (fsm_output[7]) | (fsm_output[5]) | (fsm_output[4]) | (fsm_output[3]);
  assign or_nl = (~ (fsm_output[7])) | (fsm_output[5]);
  assign mux_nl = MUX_s_1_2_2(or_tmp_2098, or_nl, fsm_output[2]);
  assign mux_1602_nl = MUX_s_1_2_2(mux_tmp_1564, mux_nl, fsm_output[0]);
  assign mux_1603_nl = MUX_s_1_2_2(or_2284_nl, mux_1602_nl, fsm_output[6]);
  assign mux_1492_nl = MUX_s_1_2_2(mux_tmp_1456, and_491_cse, fsm_output[2]);
  assign mux_1496_nl = MUX_s_1_2_2(and_tmp_11, and_485_cse, fsm_output[2]);
  assign mux_1497_nl = MUX_s_1_2_2(not_tmp_692, mux_1496_nl, fsm_output[5]);
  assign and_260_nl = (fsm_output[4:3]==2'b11) & or_32_cse;
  assign mux_1498_nl = MUX_s_1_2_2(and_260_nl, and_479_cse, fsm_output[2]);
  assign mux_1499_nl = MUX_s_1_2_2(or_tmp_2057, (~ mux_1498_nl), fsm_output[5]);
  assign mux_1500_nl = MUX_s_1_2_2(or_tmp_2057, (~ and_479_cse), fsm_output[5]);
  assign nl_COMP_LOOP_3_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_3_sva_6_0 , 3'b010}) + 11'b00000000001;
  assign COMP_LOOP_3_acc_nl = nl_COMP_LOOP_3_acc_nl[10:0];
  assign and_310_nl = (fsm_output[4]) & (fsm_output[3]) & (fsm_output[1]);
  assign mux_1501_nl = MUX_s_1_2_2(and_310_nl, and_479_cse, fsm_output[2]);
  assign mux_1502_nl = MUX_s_1_2_2(or_tmp_2057, (~ mux_1501_nl), fsm_output[5]);
  assign nl_COMP_LOOP_acc_11_psp_sva  = (VEC_LOOP_j_10_0_sva_9_0[9:1]) + ({COMP_LOOP_k_10_3_sva_6_0
      , 2'b01});
  assign mux_1504_nl = MUX_s_1_2_2(mux_tmp_1468, and_tmp_11, fsm_output[2]);
  assign mux_1505_nl = MUX_s_1_2_2(mux_1504_nl, (fsm_output[6]), fsm_output[5]);
  assign mux_1506_nl = MUX_s_1_2_2(mux_tmp_1468, and_485_cse, fsm_output[2]);
  assign mux_1507_nl = MUX_s_1_2_2(mux_1506_nl, (fsm_output[6]), fsm_output[5]);
  assign nl_COMP_LOOP_acc_12_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:3]))})
      + conv_u2u_8_9({COMP_LOOP_k_10_3_sva_6_0 , 1'b0}) + 9'b000000001;
  assign COMP_LOOP_acc_12_nl = nl_COMP_LOOP_acc_12_nl[8:0];
  assign mux_1508_nl = MUX_s_1_2_2(mux_tmp_1468, and_tmp_13, fsm_output[2]);
  assign mux_1509_nl = MUX_s_1_2_2(mux_1508_nl, (fsm_output[6]), fsm_output[5]);
  assign mux_1511_nl = MUX_s_1_2_2(not_tmp_692, and_485_cse, fsm_output[5]);
  assign nl_COMP_LOOP_5_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_3_sva_6_0 , 3'b100}) + 11'b00000000001;
  assign COMP_LOOP_5_acc_nl = nl_COMP_LOOP_5_acc_nl[10:0];
  assign mux_1512_nl = MUX_s_1_2_2(and_tmp_13, and_485_cse, fsm_output[2]);
  assign mux_1513_nl = MUX_s_1_2_2(not_tmp_692, mux_1512_nl, fsm_output[5]);
  assign nl_COMP_LOOP_acc_13_psp_sva  = (VEC_LOOP_j_10_0_sva_9_0[9:2]) + ({COMP_LOOP_k_10_3_sva_6_0
      , 1'b1});
  assign mux_1518_nl = MUX_s_1_2_2(mux_tmp_1482, mux_tmp_1456, fsm_output[2]);
  assign mux_1520_nl = MUX_s_1_2_2(mux_tmp_1482, and_491_cse, fsm_output[2]);
  assign nl_COMP_LOOP_6_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_3_sva_6_0 , 3'b101}) + 11'b00000000001;
  assign COMP_LOOP_6_acc_nl = nl_COMP_LOOP_6_acc_nl[10:0];
  assign mux_1523_nl = MUX_s_1_2_2(mux_tmp_1482, mux_tmp_1487, fsm_output[2]);
  assign nl_COMP_LOOP_7_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_3_sva_6_0 , 3'b110}) + 11'b00000000001;
  assign COMP_LOOP_7_acc_nl = nl_COMP_LOOP_7_acc_nl[10:0];
  assign mux_1528_nl = MUX_s_1_2_2(mux_tmp_1487, and_491_cse, fsm_output[2]);
  assign nl_COMP_LOOP_acc_14_psp_sva  = (VEC_LOOP_j_10_0_sva_9_0[9:1]) + ({COMP_LOOP_k_10_3_sva_6_0
      , 2'b11});
  assign mux_1532_nl = MUX_s_1_2_2(mux_tmp_1452, nor_tmp_95, fsm_output[2]);
  assign or_162_nl = (fsm_output[5:2]!=4'b0000);
  assign nl_COMP_LOOP_acc_15_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:4]))})
      + conv_u2u_7_8(COMP_LOOP_k_10_3_sva_6_0) + 8'b00000001;
  assign COMP_LOOP_acc_15_nl = nl_COMP_LOOP_acc_15_nl[7:0];
  assign nl_COMP_LOOP_acc_1_cse_sva  = VEC_LOOP_j_10_0_sva_9_0 + ({COMP_LOOP_k_10_3_sva_6_0
      , 3'b111});
  assign and_305_nl = ((fsm_output[4:0]!=5'b00000)) & (fsm_output[7:6]==2'b11);
  assign nl_COMP_LOOP_1_acc_nl = ({z_out_2 , 3'b000}) + ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + 11'b00000000001;
  assign COMP_LOOP_1_acc_nl = nl_COMP_LOOP_1_acc_nl[10:0];
  assign and_304_nl = ((fsm_output[4:1]!=4'b0000)) & (fsm_output[7:6]==2'b11);
  assign COMP_LOOP_COMP_LOOP_and_33_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b00011);
  assign COMP_LOOP_COMP_LOOP_and_35_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b00101);
  assign COMP_LOOP_COMP_LOOP_and_36_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b00110);
  assign COMP_LOOP_COMP_LOOP_and_37_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b00111);
  assign COMP_LOOP_COMP_LOOP_and_39_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b01001);
  assign COMP_LOOP_COMP_LOOP_and_40_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b01010);
  assign COMP_LOOP_COMP_LOOP_and_41_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b01011);
  assign COMP_LOOP_COMP_LOOP_and_42_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b01100);
  assign COMP_LOOP_COMP_LOOP_and_43_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b01101);
  assign COMP_LOOP_COMP_LOOP_and_44_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b01110);
  assign COMP_LOOP_COMP_LOOP_and_45_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b01111);
  assign COMP_LOOP_COMP_LOOP_and_47_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b10001);
  assign COMP_LOOP_COMP_LOOP_and_48_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b10010);
  assign COMP_LOOP_COMP_LOOP_and_49_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b10011);
  assign COMP_LOOP_COMP_LOOP_and_50_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b10100);
  assign COMP_LOOP_COMP_LOOP_and_51_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b10101);
  assign COMP_LOOP_COMP_LOOP_and_52_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b10110);
  assign COMP_LOOP_nor_26_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:1]!=4'b0000));
  assign COMP_LOOP_nor_27_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4]) | (COMP_LOOP_1_acc_10_itm_10_1_1[3])
      | (COMP_LOOP_1_acc_10_itm_10_1_1[2]) | (COMP_LOOP_1_acc_10_itm_10_1_1[0]));
  assign COMP_LOOP_nor_29_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4]) | (COMP_LOOP_1_acc_10_itm_10_1_1[3])
      | (COMP_LOOP_1_acc_10_itm_10_1_1[1]) | (COMP_LOOP_1_acc_10_itm_10_1_1[0]));
  assign COMP_LOOP_nor_33_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4]) | (COMP_LOOP_1_acc_10_itm_10_1_1[2])
      | (COMP_LOOP_1_acc_10_itm_10_1_1[1]) | (COMP_LOOP_1_acc_10_itm_10_1_1[0]));
  assign COMP_LOOP_nor_40_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[3:0]!=4'b0000));
  assign COMP_LOOP_COMP_LOOP_and_53_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b10111);
  assign COMP_LOOP_COMP_LOOP_and_54_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b11000);
  assign COMP_LOOP_COMP_LOOP_and_55_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b11001);
  assign COMP_LOOP_COMP_LOOP_and_56_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b11010);
  assign COMP_LOOP_COMP_LOOP_and_57_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b11011);
  assign COMP_LOOP_COMP_LOOP_and_58_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b11100);
  assign COMP_LOOP_COMP_LOOP_and_59_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b11101);
  assign COMP_LOOP_COMP_LOOP_and_60_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b11110);
  assign COMP_LOOP_COMP_LOOP_and_61_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[4:0]==5'b11111);
  assign COMP_LOOP_COMP_LOOP_nor_1_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b00000));
  assign COMP_LOOP_COMP_LOOP_mux_2_nl = MUX_v_64_2_2(COMP_LOOP_1_acc_8_itm, z_out_9,
      COMP_LOOP_or_33_itm);
  assign nl_COMP_LOOP_acc_17_nl = COMP_LOOP_mux_385_cse + COMP_LOOP_COMP_LOOP_mux_2_nl;
  assign COMP_LOOP_acc_17_nl = nl_COMP_LOOP_acc_17_nl[63:0];
  assign COMP_LOOP_or_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_131_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_30_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_29_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_28_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_27_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_26_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_25_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_24_itm & and_dcpl_83);
  assign COMP_LOOP_or_1_nl = ((COMP_LOOP_acc_10_cse_10_1_1_sva[0]) & COMP_LOOP_tmp_nor_1_itm
      & and_dcpl_49) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_30_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_29_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_28_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_27_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_26_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_25_itm & and_dcpl_83);
  assign COMP_LOOP_or_2_nl = ((COMP_LOOP_acc_10_cse_10_1_1_sva[1]) & COMP_LOOP_tmp_nor_14_itm
      & and_dcpl_49) | (COMP_LOOP_COMP_LOOP_and_625_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_30_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_29_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_28_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_27_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_26_itm & and_dcpl_83);
  assign COMP_LOOP_or_3_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_126_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_625_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_30_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_29_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_28_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_27_itm & and_dcpl_83);
  assign COMP_LOOP_or_4_nl = ((COMP_LOOP_acc_10_cse_10_1_1_sva[2]) & COMP_LOOP_tmp_nor_3_itm
      & and_dcpl_49) | (COMP_LOOP_COMP_LOOP_and_377_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_126_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_625_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_30_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_29_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_28_itm & and_dcpl_83);
  assign COMP_LOOP_or_5_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_128_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_377_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_126_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_625_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_30_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_29_itm & and_dcpl_83);
  assign COMP_LOOP_or_6_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_129_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_128_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_377_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_126_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_625_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_30_itm & and_dcpl_83);
  assign COMP_LOOP_or_7_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_130_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_129_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_128_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_377_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_126_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_625_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_83);
  assign COMP_LOOP_or_8_nl = ((COMP_LOOP_acc_10_cse_10_1_1_sva[3]) & COMP_LOOP_tmp_nor_42_itm
      & and_dcpl_49) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_130_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_129_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_128_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_377_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_126_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_625_itm & and_dcpl_83);
  assign COMP_LOOP_or_9_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_132_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_130_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_129_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_128_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_377_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_126_itm & and_dcpl_83);
  assign COMP_LOOP_or_10_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_133_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_132_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_130_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_129_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_128_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_377_itm & and_dcpl_83);
  assign COMP_LOOP_or_11_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_134_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_133_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_132_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_130_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_129_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_128_itm & and_dcpl_83);
  assign COMP_LOOP_or_12_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_134_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_133_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_132_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_130_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_129_itm & and_dcpl_83);
  assign COMP_LOOP_or_13_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_136_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_134_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_133_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_132_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_130_itm & and_dcpl_83);
  assign COMP_LOOP_or_14_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_136_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_134_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_133_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_132_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_83);
  assign COMP_LOOP_or_15_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_136_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_134_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_133_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_132_itm & and_dcpl_83);
  assign COMP_LOOP_or_16_nl = ((COMP_LOOP_acc_10_cse_10_1_1_sva[4]) & COMP_LOOP_tmp_nor_49_itm
      & and_dcpl_49) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_136_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_134_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_133_itm & and_dcpl_83);
  assign COMP_LOOP_or_17_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_140_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_136_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_134_itm & and_dcpl_83);
  assign COMP_LOOP_or_18_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_141_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_140_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_136_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_83);
  assign COMP_LOOP_or_19_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_142_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_141_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_140_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_136_itm & and_dcpl_83);
  assign COMP_LOOP_or_20_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_18_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_142_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_141_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_140_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_83);
  assign COMP_LOOP_or_21_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_144_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_18_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_142_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_141_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_140_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_83);
  assign COMP_LOOP_or_22_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_20_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_144_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_18_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_142_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_141_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_140_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_83);
  assign COMP_LOOP_or_23_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_21_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_20_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_144_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_18_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_142_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_141_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_140_itm & and_dcpl_83);
  assign COMP_LOOP_or_24_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_122_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_22_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_21_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_20_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_144_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_18_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_142_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_141_itm & and_dcpl_83);
  assign COMP_LOOP_or_25_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_123_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_23_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_22_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_21_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_20_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_144_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_18_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_142_itm & and_dcpl_83);
  assign COMP_LOOP_or_26_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_124_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_24_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_23_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_22_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_21_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_20_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_144_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_18_itm & and_dcpl_83);
  assign COMP_LOOP_or_27_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_126_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_25_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_24_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_23_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_22_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_21_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_20_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_144_itm & and_dcpl_83);
  assign COMP_LOOP_or_28_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_127_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_26_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_25_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_24_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_23_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_22_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_21_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_20_itm & and_dcpl_83);
  assign COMP_LOOP_or_29_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_128_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_27_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_26_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_25_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_24_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_23_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_22_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_21_itm & and_dcpl_83);
  assign COMP_LOOP_or_30_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_129_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_28_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_27_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_26_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_25_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_24_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_23_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_22_itm & and_dcpl_83);
  assign COMP_LOOP_or_31_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_130_itm & and_dcpl_49)
      | (COMP_LOOP_COMP_LOOP_and_29_itm & and_dcpl_54) | (COMP_LOOP_COMP_LOOP_and_28_itm
      & and_dcpl_58) | (COMP_LOOP_COMP_LOOP_and_27_itm & and_dcpl_65) | (COMP_LOOP_COMP_LOOP_and_26_itm
      & and_dcpl_68) | (COMP_LOOP_COMP_LOOP_and_25_itm & and_dcpl_75) | (COMP_LOOP_COMP_LOOP_and_24_itm
      & and_dcpl_78) | (COMP_LOOP_COMP_LOOP_and_23_itm & and_dcpl_83);
  assign COMP_LOOP_tmp_and_127_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_131_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[0])
      & COMP_LOOP_tmp_nor_49_itm & (~ and_294_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[1])
      & COMP_LOOP_tmp_nor_1_itm & (~ and_294_tmp);
  assign COMP_LOOP_tmp_and_128_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_127_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_129_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_169 & (~ and_294_tmp);
  assign COMP_LOOP_tmp_and_130_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_128_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_131_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_129_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_132_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_130_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_133_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_167 & (~ and_294_tmp);
  assign COMP_LOOP_tmp_and_134_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_135_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_136_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_137_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_138_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_139_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_140_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_18_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[4])
      & COMP_LOOP_tmp_nor_14_itm & (~ and_294_tmp);
  assign COMP_LOOP_tmp_and_141_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_142_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_143_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_144_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_145_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_146_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_147_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_148_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_149_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_150_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_151_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_152_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_122_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_153_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_123_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_154_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_124_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_155_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_126_itm & (~
      and_294_tmp);
  assign COMP_LOOP_tmp_and_115_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm & (~
      nor_1119_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_34_nl = (COMP_LOOP_3_tmp_mul_idiv_sva_3_0[0])
      & COMP_LOOP_tmp_nor_25_itm & (~ nor_1119_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_35_nl = (COMP_LOOP_3_tmp_mul_idiv_sva_3_0[1])
      & COMP_LOOP_tmp_nor_26_itm & (~ nor_1119_tmp);
  assign COMP_LOOP_tmp_and_116_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm & (~
      nor_1119_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_37_nl = (COMP_LOOP_3_tmp_mul_idiv_sva_3_0[2])
      & COMP_LOOP_tmp_nor_28_itm & (~ nor_1119_tmp);
  assign COMP_LOOP_tmp_and_117_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm & (~
      nor_1119_tmp);
  assign COMP_LOOP_tmp_and_118_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm & (~
      nor_1119_tmp);
  assign COMP_LOOP_tmp_and_119_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm & (~
      nor_1119_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_41_nl = (COMP_LOOP_3_tmp_mul_idiv_sva_3_0[3])
      & COMP_LOOP_tmp_nor_31_itm & (~ nor_1119_tmp);
  assign COMP_LOOP_tmp_and_120_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm & (~
      nor_1119_tmp);
  assign COMP_LOOP_tmp_and_121_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm & (~
      nor_1119_tmp);
  assign COMP_LOOP_tmp_and_122_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm & (~
      nor_1119_tmp);
  assign COMP_LOOP_tmp_and_123_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm & (~
      nor_1119_tmp);
  assign COMP_LOOP_tmp_and_124_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm & (~
      nor_1119_tmp);
  assign COMP_LOOP_tmp_and_125_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm & (~
      nor_1119_tmp);
  assign COMP_LOOP_tmp_and_126_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm & (~
      nor_1119_tmp);
  assign COMP_LOOP_tmp_and_83_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_131_itm & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_84_nl = and_1_cse & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_85_nl = and_4_cse & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_86_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_87_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_169 & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_88_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_89_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_90_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_91_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_167 & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_92_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_93_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_94_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_95_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_96_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_97_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_98_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_99_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_165 & (~ nor_tmp);
  assign COMP_LOOP_tmp_and_100_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm & (~
      nor_tmp);
  assign COMP_LOOP_tmp_and_101_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm & (~
      nor_tmp);
  assign COMP_LOOP_tmp_and_102_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm & (~
      nor_tmp);
  assign COMP_LOOP_tmp_and_103_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm & (~
      nor_tmp);
  assign COMP_LOOP_tmp_and_104_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm & (~
      nor_tmp);
  assign COMP_LOOP_tmp_and_105_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm & (~
      nor_tmp);
  assign COMP_LOOP_tmp_and_106_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_itm & (~
      nor_tmp);
  assign COMP_LOOP_tmp_and_107_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_122_itm & (~
      nor_tmp);
  assign COMP_LOOP_tmp_and_108_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_123_itm & (~
      nor_tmp);
  assign COMP_LOOP_tmp_and_109_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_124_itm & (~
      nor_tmp);
  assign COMP_LOOP_tmp_and_110_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_126_itm & (~
      nor_tmp);
  assign COMP_LOOP_tmp_and_111_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_127_itm & (~
      nor_tmp);
  assign COMP_LOOP_tmp_and_112_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_128_itm & (~
      nor_tmp);
  assign COMP_LOOP_tmp_and_113_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_129_itm & (~
      nor_tmp);
  assign COMP_LOOP_tmp_and_114_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_130_itm & (~
      nor_tmp);
  assign COMP_LOOP_tmp_and_78_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_itm & (~ nor_1117_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_80_nl = (COMP_LOOP_5_tmp_mul_idiv_sva[2:0]==3'b001)
      & (~ nor_1117_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_81_nl = (COMP_LOOP_5_tmp_mul_idiv_sva[2:0]==3'b010)
      & (~ nor_1117_tmp);
  assign COMP_LOOP_tmp_and_79_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_82_itm & (~ nor_1117_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_83_nl = (COMP_LOOP_5_tmp_mul_idiv_sva[2:0]==3'b100)
      & (~ nor_1117_tmp);
  assign COMP_LOOP_tmp_and_80_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_84_itm & (~ nor_1117_tmp);
  assign COMP_LOOP_tmp_and_81_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_85_itm & (~ nor_1117_tmp);
  assign COMP_LOOP_tmp_and_82_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_86_itm & (~ nor_1117_tmp);
  assign COMP_LOOP_tmp_and_47_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_48_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_rgt & and_298_m1c;
  assign COMP_LOOP_tmp_and_49_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_50_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_rgt & and_298_m1c;
  assign COMP_LOOP_tmp_and_51_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_52_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_53_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_54_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_rgt & and_298_m1c;
  assign COMP_LOOP_tmp_and_55_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_56_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_57_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_58_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_59_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_60_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_61_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_62_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_rgt & and_298_m1c;
  assign COMP_LOOP_tmp_and_63_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_64_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_65_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_66_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_67_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_68_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_69_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_70_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_71_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_72_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_73_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_74_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_75_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_76_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm & and_298_m1c;
  assign COMP_LOOP_tmp_and_77_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm & and_298_m1c;
  assign nor_337_nl = ~(((fsm_output[3]) & (fsm_output[0]) & (fsm_output[1])) | (fsm_output[7:6]!=2'b00));
  assign mux_1583_nl = MUX_s_1_2_2(nor_337_nl, and_449_cse, fsm_output[4]);
  assign mux_1582_nl = MUX_s_1_2_2((~ or_tmp_2075), and_464_cse, fsm_output[4]);
  assign mux_1584_nl = MUX_s_1_2_2(mux_1583_nl, mux_1582_nl, fsm_output[2]);
  assign mux_1585_nl = MUX_s_1_2_2(mux_1584_nl, and_464_cse, fsm_output[5]);
  assign COMP_LOOP_tmp_and_15_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_16_nl = and_1_cse & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_17_nl = and_4_cse & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_18_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_19_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_169 & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_20_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_21_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_22_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_23_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_167 & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_24_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_25_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_26_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_27_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_28_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_29_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_30_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_31_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_165 & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_32_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_33_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_34_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_35_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_36_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_37_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_38_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_39_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_40_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_41_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_42_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_43_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_44_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_45_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_46_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm & mux_1592_tmp;
  assign COMP_LOOP_tmp_and_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm & and_dcpl_177;
  assign COMP_LOOP_tmp_and_1_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_119_rgt & and_dcpl_177;
  assign COMP_LOOP_tmp_and_2_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_itm & and_dcpl_177;
  assign COMP_LOOP_tmp_and_3_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_121_rgt & and_dcpl_177;
  assign COMP_LOOP_tmp_and_4_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_122_itm & and_dcpl_177;
  assign COMP_LOOP_tmp_and_5_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_123_itm & and_dcpl_177;
  assign COMP_LOOP_tmp_and_6_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_124_itm & and_dcpl_177;
  assign COMP_LOOP_tmp_and_7_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_125_rgt & and_dcpl_177;
  assign COMP_LOOP_tmp_and_8_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_126_itm & and_dcpl_177;
  assign COMP_LOOP_tmp_and_9_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_127_itm & and_dcpl_177;
  assign COMP_LOOP_tmp_and_10_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_128_itm & and_dcpl_177;
  assign COMP_LOOP_tmp_and_11_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_129_itm & and_dcpl_177;
  assign COMP_LOOP_tmp_and_12_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_130_itm & and_dcpl_177;
  assign COMP_LOOP_tmp_and_13_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_131_itm & and_dcpl_177;
  assign COMP_LOOP_tmp_and_14_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_132_itm & and_dcpl_177;
  assign mux_1594_nl = MUX_s_1_2_2(mux_189_cse, and_464_cse, and_496_cse);
  assign mux_1595_nl = MUX_s_1_2_2(mux_1594_nl, and_464_cse, fsm_output[4]);
  assign mux_217_nl = MUX_s_1_2_2(mux_189_cse, and_464_cse, or_212_cse);
  assign mux_1596_nl = MUX_s_1_2_2(mux_1595_nl, mux_217_nl, fsm_output[2]);
  assign and_478_nl = (and_479_cse | (fsm_output[6])) & (fsm_output[7]);
  assign mux_1597_nl = MUX_s_1_2_2(mux_1596_nl, and_478_nl, fsm_output[5]);
  assign and_755_nl = (fsm_output[7:6]==2'b11) & and_dcpl_31 & and_dcpl_29 & (fsm_output[2])
      & (fsm_output[5]);
  assign COMP_LOOP_mux_382_nl = MUX_v_7_2_2(COMP_LOOP_k_10_3_sva_6_0, ({3'b001 ,
      (~ z_out_4)}), and_755_nl);
  assign nl_z_out_2 = conv_u2u_7_8(COMP_LOOP_mux_382_nl) + 8'b00000001;
  assign z_out_2 = nl_z_out_2[7:0];
  assign COMP_LOOP_mux_383_nl = MUX_v_11_2_2(({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))}),
      STAGE_LOOP_lshift_psp_sva, and_dcpl_334);
  assign COMP_LOOP_COMP_LOOP_nand_1_nl = ~(and_dcpl_334 & (~(nor_1025_cse & (fsm_output[1:0]==2'b10)
      & and_dcpl_29 & and_dcpl_28)));
  assign COMP_LOOP_mux_384_nl = MUX_v_10_2_2(({COMP_LOOP_k_10_3_sva_6_0 , 3'b001}),
      VEC_LOOP_j_10_0_sva_9_0, and_dcpl_334);
  assign nl_acc_1_nl = ({COMP_LOOP_mux_383_nl , COMP_LOOP_COMP_LOOP_nand_1_nl}) +
      conv_u2u_11_12({COMP_LOOP_mux_384_nl , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[11:0];
  assign z_out_3 = readslicef_12_11_1(acc_1_nl);
  assign STAGE_LOOP_mux_4_nl = MUX_v_4_2_2(STAGE_LOOP_i_3_0_sva, (~ STAGE_LOOP_i_3_0_sva),
      and_dcpl_347);
  assign nl_z_out_4 = STAGE_LOOP_mux_4_nl + ({1'b1 , (~ and_dcpl_347) , 2'b11});
  assign z_out_4 = nl_z_out_4[3:0];
  assign COMP_LOOP_mux_385_cse = MUX_v_64_2_2(z_out_9, COMP_LOOP_1_acc_8_itm, COMP_LOOP_or_33_itm);
  assign COMP_LOOP_tmp_nor_135_cse = ~(and_dcpl_420 | and_dcpl_435 | and_dcpl_436);
  assign COMP_LOOP_tmp_mux_21_nl = MUX_s_1_2_2((z_out_1[9]), (COMP_LOOP_2_tmp_lshift_ncse_sva[9]),
      COMP_LOOP_tmp_or_54_ssc);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_174_nl = COMP_LOOP_tmp_mux_21_nl & COMP_LOOP_tmp_nor_135_cse;
  assign COMP_LOOP_tmp_or_76_nl = and_dcpl_423 | and_dcpl_435;
  assign COMP_LOOP_tmp_mux1h_94_nl = MUX1HOT_v_9_4_2(({1'b0 , (z_out[7:0])}), (z_out_1[8:0]),
      (COMP_LOOP_2_tmp_lshift_ncse_sva[8:0]), COMP_LOOP_3_tmp_lshift_ncse_sva, {and_dcpl_420
      , COMP_LOOP_tmp_or_76_nl , COMP_LOOP_tmp_or_54_ssc , and_dcpl_436});
  assign COMP_LOOP_tmp_and_161_nl = (COMP_LOOP_k_10_3_sva_6_0[6]) & COMP_LOOP_tmp_nor_135_cse;
  assign COMP_LOOP_tmp_or_77_nl = and_dcpl_423 | and_dcpl_428 | and_dcpl_429 | and_dcpl_434;
  assign COMP_LOOP_tmp_mux1h_95_nl = MUX1HOT_v_6_3_2(({1'b0 , (COMP_LOOP_k_10_3_sva_6_0[6:2])}),
      (COMP_LOOP_k_10_3_sva_6_0[5:0]), (COMP_LOOP_k_10_3_sva_6_0[6:1]), {and_dcpl_420
      , COMP_LOOP_tmp_or_77_nl , COMP_LOOP_tmp_or_71_itm});
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_mux_18_nl = MUX_s_1_2_2((COMP_LOOP_k_10_3_sva_6_0[1]),
      (COMP_LOOP_k_10_3_sva_6_0[0]), COMP_LOOP_tmp_or_71_itm);
  assign COMP_LOOP_tmp_or_78_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_mux_18_nl & (~(and_dcpl_423
      | and_dcpl_428))) | and_dcpl_429 | and_dcpl_434;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_or_1_nl = ((COMP_LOOP_k_10_3_sva_6_0[0]) & (~(and_dcpl_423
      | and_dcpl_429 | and_dcpl_435))) | and_dcpl_428 | and_dcpl_434 | and_dcpl_436;
  assign nl_z_out_7 = ({COMP_LOOP_tmp_COMP_LOOP_tmp_and_174_nl , COMP_LOOP_tmp_mux1h_94_nl})
      * ({COMP_LOOP_tmp_and_161_nl , COMP_LOOP_tmp_mux1h_95_nl , COMP_LOOP_tmp_or_78_nl
      , COMP_LOOP_tmp_COMP_LOOP_tmp_or_1_nl , 1'b1});
  assign z_out_7 = nl_z_out_7[9:0];
  assign and_756_nl = nor_1025_cse & (fsm_output[1:0]==2'b10) & and_dcpl_30;
  assign COMP_LOOP_tmp_mux1h_96_nl = MUX1HOT_v_64_9_2(({57'b000000000000000000000000000000000000000000000000000000000
      , (z_out_1[6:0])}), COMP_LOOP_tmp_mux1h_itm, COMP_LOOP_tmp_mux1h_1_itm, COMP_LOOP_tmp_mux1h_2_itm,
      COMP_LOOP_tmp_mux1h_3_itm, COMP_LOOP_tmp_mux1h_4_itm, COMP_LOOP_tmp_mux1h_5_itm,
      COMP_LOOP_tmp_mux1h_6_itm, tmp_21_sva_1, {and_756_nl , and_dcpl_448 , and_dcpl_452
      , and_dcpl_456 , and_dcpl_458 , and_dcpl_461 , and_dcpl_465 , and_dcpl_468
      , and_dcpl_472});
  assign COMP_LOOP_tmp_or_79_nl = and_dcpl_448 | and_dcpl_452 | and_dcpl_456 | and_dcpl_458
      | and_dcpl_461 | and_dcpl_465 | and_dcpl_468 | and_dcpl_472;
  assign COMP_LOOP_tmp_mux_22_nl = MUX_v_64_2_2(({57'b000000000000000000000000000000000000000000000000000000000
      , COMP_LOOP_k_10_3_sva_6_0}), COMP_LOOP_1_modulo_dev_cmp_return_rsc_z, COMP_LOOP_tmp_or_79_nl);
  assign nl_z_out_8 = COMP_LOOP_tmp_mux1h_96_nl * COMP_LOOP_tmp_mux_22_nl;
  assign z_out_8 = nl_z_out_8[63:0];
  assign COMP_LOOP_mux1h_657_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_nor_itm, COMP_LOOP_COMP_LOOP_nor_5_itm,
      COMP_LOOP_COMP_LOOP_nor_9_itm, COMP_LOOP_COMP_LOOP_nor_13_itm, COMP_LOOP_COMP_LOOP_nor_17_itm,
      COMP_LOOP_COMP_LOOP_nor_21_itm, COMP_LOOP_COMP_LOOP_nor_25_itm, COMP_LOOP_COMP_LOOP_nor_29_itm,
      {and_dcpl_479 , and_605_cse , and_609_cse , and_614_cse , and_617_cse , and_621_cse
      , and_624_cse , and_628_cse});
  assign COMP_LOOP_COMP_LOOP_and_930_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[0]) &
      COMP_LOOP_nor_126_itm;
  assign COMP_LOOP_COMP_LOOP_and_931_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[0]) &
      COMP_LOOP_nor_226_itm;
  assign COMP_LOOP_COMP_LOOP_and_932_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[0]) &
      COMP_LOOP_nor_326_itm;
  assign COMP_LOOP_COMP_LOOP_and_933_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[0]) &
      COMP_LOOP_nor_426_itm;
  assign COMP_LOOP_COMP_LOOP_and_934_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[0]) &
      COMP_LOOP_nor_526_itm;
  assign COMP_LOOP_COMP_LOOP_and_935_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) &
      COMP_LOOP_nor_626_itm;
  assign COMP_LOOP_COMP_LOOP_and_936_nl = (COMP_LOOP_acc_10_cse_10_1_sva[0]) & COMP_LOOP_nor_726_itm;
  assign COMP_LOOP_mux1h_658_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_625_itm,
      COMP_LOOP_COMP_LOOP_and_930_nl, COMP_LOOP_COMP_LOOP_and_931_nl, COMP_LOOP_COMP_LOOP_and_932_nl,
      COMP_LOOP_COMP_LOOP_and_933_nl, COMP_LOOP_COMP_LOOP_and_934_nl, COMP_LOOP_COMP_LOOP_and_935_nl,
      COMP_LOOP_COMP_LOOP_and_936_nl, {and_dcpl_479 , and_605_cse , and_609_cse ,
      and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_COMP_LOOP_and_937_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[1]) &
      COMP_LOOP_nor_127_itm;
  assign COMP_LOOP_COMP_LOOP_and_938_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[1]) &
      COMP_LOOP_nor_227_itm;
  assign COMP_LOOP_COMP_LOOP_and_939_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[1]) &
      COMP_LOOP_nor_327_itm;
  assign COMP_LOOP_COMP_LOOP_and_940_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[1]) &
      COMP_LOOP_nor_427_itm;
  assign COMP_LOOP_COMP_LOOP_and_941_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[1]) &
      COMP_LOOP_nor_527_itm;
  assign COMP_LOOP_COMP_LOOP_and_942_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[1]) &
      COMP_LOOP_nor_627_itm;
  assign COMP_LOOP_COMP_LOOP_and_943_nl = (COMP_LOOP_acc_10_cse_10_1_sva[1]) & COMP_LOOP_nor_727_itm;
  assign COMP_LOOP_mux1h_659_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_126_itm,
      COMP_LOOP_COMP_LOOP_and_937_nl, COMP_LOOP_COMP_LOOP_and_938_nl, COMP_LOOP_COMP_LOOP_and_939_nl,
      COMP_LOOP_COMP_LOOP_and_940_nl, COMP_LOOP_COMP_LOOP_and_941_nl, COMP_LOOP_COMP_LOOP_and_942_nl,
      COMP_LOOP_COMP_LOOP_and_943_nl, {and_dcpl_479 , and_605_cse , and_609_cse ,
      and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_660_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_377_itm,
      COMP_LOOP_COMP_LOOP_and_157_itm, COMP_LOOP_COMP_LOOP_and_281_itm, COMP_LOOP_COMP_LOOP_and_405_itm,
      COMP_LOOP_COMP_LOOP_and_529_itm, COMP_LOOP_COMP_LOOP_and_653_itm, COMP_LOOP_COMP_LOOP_and_777_itm,
      COMP_LOOP_COMP_LOOP_and_901_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_COMP_LOOP_and_944_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[2]) &
      COMP_LOOP_nor_129_itm;
  assign COMP_LOOP_COMP_LOOP_and_945_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[2]) &
      COMP_LOOP_nor_229_itm;
  assign COMP_LOOP_COMP_LOOP_and_946_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[2]) &
      COMP_LOOP_nor_329_itm;
  assign COMP_LOOP_COMP_LOOP_and_947_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[2]) &
      COMP_LOOP_nor_429_itm;
  assign COMP_LOOP_COMP_LOOP_and_948_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[2]) &
      COMP_LOOP_nor_529_itm;
  assign COMP_LOOP_COMP_LOOP_and_949_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[2]) &
      COMP_LOOP_nor_629_itm;
  assign COMP_LOOP_COMP_LOOP_and_950_nl = (COMP_LOOP_acc_10_cse_10_1_sva[2]) & COMP_LOOP_nor_729_itm;
  assign COMP_LOOP_mux1h_661_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_128_itm,
      COMP_LOOP_COMP_LOOP_and_944_nl, COMP_LOOP_COMP_LOOP_and_945_nl, COMP_LOOP_COMP_LOOP_and_946_nl,
      COMP_LOOP_COMP_LOOP_and_947_nl, COMP_LOOP_COMP_LOOP_and_948_nl, COMP_LOOP_COMP_LOOP_and_949_nl,
      COMP_LOOP_COMP_LOOP_and_950_nl, {and_dcpl_479 , and_605_cse , and_609_cse ,
      and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_662_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_129_itm,
      COMP_LOOP_COMP_LOOP_and_159_itm, COMP_LOOP_COMP_LOOP_and_283_itm, COMP_LOOP_COMP_LOOP_and_407_itm,
      COMP_LOOP_COMP_LOOP_and_531_itm, COMP_LOOP_COMP_LOOP_and_655_itm, COMP_LOOP_COMP_LOOP_and_779_itm,
      COMP_LOOP_COMP_LOOP_and_903_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_663_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_130_itm,
      COMP_LOOP_COMP_LOOP_and_160_itm, COMP_LOOP_COMP_LOOP_and_284_itm, COMP_LOOP_COMP_LOOP_and_408_itm,
      COMP_LOOP_COMP_LOOP_and_532_itm, COMP_LOOP_COMP_LOOP_and_656_itm, COMP_LOOP_COMP_LOOP_and_780_itm,
      COMP_LOOP_COMP_LOOP_and_904_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_664_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_6_itm,
      COMP_LOOP_COMP_LOOP_and_161_itm, COMP_LOOP_COMP_LOOP_and_285_itm, COMP_LOOP_COMP_LOOP_and_409_itm,
      COMP_LOOP_COMP_LOOP_and_533_itm, COMP_LOOP_COMP_LOOP_and_657_itm, COMP_LOOP_COMP_LOOP_and_781_itm,
      COMP_LOOP_COMP_LOOP_and_905_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_COMP_LOOP_and_951_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[3]) &
      COMP_LOOP_nor_133_itm;
  assign COMP_LOOP_COMP_LOOP_and_952_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[3]) &
      COMP_LOOP_nor_233_itm;
  assign COMP_LOOP_COMP_LOOP_and_953_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[3]) &
      COMP_LOOP_nor_333_itm;
  assign COMP_LOOP_COMP_LOOP_and_954_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[3]) &
      COMP_LOOP_nor_433_itm;
  assign COMP_LOOP_COMP_LOOP_and_955_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3]) &
      COMP_LOOP_nor_533_itm;
  assign COMP_LOOP_COMP_LOOP_and_956_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3]) &
      COMP_LOOP_nor_633_itm;
  assign COMP_LOOP_COMP_LOOP_and_957_nl = (COMP_LOOP_acc_10_cse_10_1_sva[3]) & COMP_LOOP_nor_733_itm;
  assign COMP_LOOP_mux1h_665_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_132_itm,
      COMP_LOOP_COMP_LOOP_and_951_nl, COMP_LOOP_COMP_LOOP_and_952_nl, COMP_LOOP_COMP_LOOP_and_953_nl,
      COMP_LOOP_COMP_LOOP_and_954_nl, COMP_LOOP_COMP_LOOP_and_955_nl, COMP_LOOP_COMP_LOOP_and_956_nl,
      COMP_LOOP_COMP_LOOP_and_957_nl, {and_dcpl_479 , and_605_cse , and_609_cse ,
      and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_666_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_133_itm,
      COMP_LOOP_COMP_LOOP_and_163_itm, COMP_LOOP_COMP_LOOP_and_287_itm, COMP_LOOP_COMP_LOOP_and_411_itm,
      COMP_LOOP_COMP_LOOP_and_535_itm, COMP_LOOP_COMP_LOOP_and_659_itm, COMP_LOOP_COMP_LOOP_and_783_itm,
      COMP_LOOP_COMP_LOOP_and_907_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_667_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_134_itm,
      COMP_LOOP_COMP_LOOP_and_164_itm, COMP_LOOP_COMP_LOOP_and_288_itm, COMP_LOOP_COMP_LOOP_and_412_itm,
      COMP_LOOP_COMP_LOOP_and_536_itm, COMP_LOOP_COMP_LOOP_and_660_itm, COMP_LOOP_COMP_LOOP_and_784_itm,
      COMP_LOOP_COMP_LOOP_and_908_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_668_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_10_itm,
      COMP_LOOP_COMP_LOOP_and_165_itm, COMP_LOOP_COMP_LOOP_and_289_itm, COMP_LOOP_COMP_LOOP_and_413_itm,
      COMP_LOOP_COMP_LOOP_and_537_itm, COMP_LOOP_COMP_LOOP_and_661_itm, COMP_LOOP_COMP_LOOP_and_785_itm,
      COMP_LOOP_COMP_LOOP_and_909_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_669_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_136_itm,
      COMP_LOOP_COMP_LOOP_and_166_itm, COMP_LOOP_COMP_LOOP_and_290_itm, COMP_LOOP_COMP_LOOP_and_414_itm,
      COMP_LOOP_COMP_LOOP_and_538_itm, COMP_LOOP_COMP_LOOP_and_662_itm, COMP_LOOP_COMP_LOOP_and_786_itm,
      COMP_LOOP_COMP_LOOP_and_910_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_670_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_12_itm,
      COMP_LOOP_COMP_LOOP_and_167_itm, COMP_LOOP_COMP_LOOP_and_291_itm, COMP_LOOP_COMP_LOOP_and_415_itm,
      COMP_LOOP_COMP_LOOP_and_539_itm, COMP_LOOP_COMP_LOOP_and_663_itm, COMP_LOOP_COMP_LOOP_and_787_itm,
      COMP_LOOP_COMP_LOOP_and_911_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_671_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_13_itm,
      COMP_LOOP_COMP_LOOP_and_168_itm, COMP_LOOP_COMP_LOOP_and_292_itm, COMP_LOOP_COMP_LOOP_and_416_itm,
      COMP_LOOP_COMP_LOOP_and_540_itm, COMP_LOOP_COMP_LOOP_and_664_itm, COMP_LOOP_COMP_LOOP_and_788_itm,
      COMP_LOOP_COMP_LOOP_and_912_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_672_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_14_itm,
      COMP_LOOP_COMP_LOOP_and_169_itm, COMP_LOOP_COMP_LOOP_and_293_itm, COMP_LOOP_COMP_LOOP_and_417_itm,
      COMP_LOOP_COMP_LOOP_and_541_itm, COMP_LOOP_COMP_LOOP_and_665_itm, COMP_LOOP_COMP_LOOP_and_789_itm,
      COMP_LOOP_COMP_LOOP_and_913_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_COMP_LOOP_and_958_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4]) &
      COMP_LOOP_nor_140_itm;
  assign COMP_LOOP_COMP_LOOP_and_959_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[4]) &
      COMP_LOOP_nor_240_itm;
  assign COMP_LOOP_COMP_LOOP_and_960_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4]) &
      COMP_LOOP_nor_340_itm;
  assign COMP_LOOP_COMP_LOOP_and_961_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4]) &
      COMP_LOOP_nor_440_itm;
  assign COMP_LOOP_COMP_LOOP_and_962_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4]) &
      COMP_LOOP_nor_540_itm;
  assign COMP_LOOP_COMP_LOOP_and_963_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[4]) &
      COMP_LOOP_nor_640_itm;
  assign COMP_LOOP_COMP_LOOP_and_964_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4]) & COMP_LOOP_nor_740_itm;
  assign COMP_LOOP_mux1h_673_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_140_itm,
      COMP_LOOP_COMP_LOOP_and_958_nl, COMP_LOOP_COMP_LOOP_and_959_nl, COMP_LOOP_COMP_LOOP_and_960_nl,
      COMP_LOOP_COMP_LOOP_and_961_nl, COMP_LOOP_COMP_LOOP_and_962_nl, COMP_LOOP_COMP_LOOP_and_963_nl,
      COMP_LOOP_COMP_LOOP_and_964_nl, {and_dcpl_479 , and_605_cse , and_609_cse ,
      and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_674_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_141_itm,
      COMP_LOOP_COMP_LOOP_and_171_itm, COMP_LOOP_COMP_LOOP_and_295_itm, COMP_LOOP_COMP_LOOP_and_419_itm,
      COMP_LOOP_COMP_LOOP_and_543_itm, COMP_LOOP_COMP_LOOP_and_667_itm, COMP_LOOP_COMP_LOOP_and_791_itm,
      COMP_LOOP_COMP_LOOP_and_915_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_675_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_142_itm,
      COMP_LOOP_COMP_LOOP_and_172_itm, COMP_LOOP_COMP_LOOP_and_296_itm, COMP_LOOP_COMP_LOOP_and_420_itm,
      COMP_LOOP_COMP_LOOP_and_544_itm, COMP_LOOP_COMP_LOOP_and_668_itm, COMP_LOOP_COMP_LOOP_and_792_itm,
      COMP_LOOP_COMP_LOOP_and_916_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_676_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_18_itm,
      COMP_LOOP_COMP_LOOP_and_173_itm, COMP_LOOP_COMP_LOOP_and_297_itm, COMP_LOOP_COMP_LOOP_and_421_itm,
      COMP_LOOP_COMP_LOOP_and_545_itm, COMP_LOOP_COMP_LOOP_and_669_itm, COMP_LOOP_COMP_LOOP_and_793_itm,
      COMP_LOOP_COMP_LOOP_and_917_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_677_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_144_itm,
      COMP_LOOP_COMP_LOOP_and_174_itm, COMP_LOOP_COMP_LOOP_and_298_itm, COMP_LOOP_COMP_LOOP_and_422_itm,
      COMP_LOOP_COMP_LOOP_and_546_itm, COMP_LOOP_COMP_LOOP_and_670_itm, COMP_LOOP_COMP_LOOP_and_794_itm,
      COMP_LOOP_COMP_LOOP_and_918_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_678_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_20_itm,
      COMP_LOOP_COMP_LOOP_and_175_itm, COMP_LOOP_COMP_LOOP_and_299_itm, COMP_LOOP_COMP_LOOP_and_423_itm,
      COMP_LOOP_COMP_LOOP_and_547_itm, COMP_LOOP_COMP_LOOP_and_671_itm, COMP_LOOP_COMP_LOOP_and_795_itm,
      COMP_LOOP_COMP_LOOP_and_919_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_679_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_21_itm,
      COMP_LOOP_COMP_LOOP_and_176_itm, COMP_LOOP_COMP_LOOP_and_300_itm, COMP_LOOP_COMP_LOOP_and_424_itm,
      COMP_LOOP_COMP_LOOP_and_548_itm, COMP_LOOP_COMP_LOOP_and_672_itm, COMP_LOOP_COMP_LOOP_and_796_itm,
      COMP_LOOP_COMP_LOOP_and_920_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_680_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_22_itm,
      COMP_LOOP_COMP_LOOP_and_177_itm, COMP_LOOP_COMP_LOOP_and_301_itm, COMP_LOOP_COMP_LOOP_and_425_itm,
      COMP_LOOP_COMP_LOOP_and_549_itm, COMP_LOOP_COMP_LOOP_and_673_itm, COMP_LOOP_COMP_LOOP_and_797_itm,
      COMP_LOOP_COMP_LOOP_and_921_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_681_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_23_itm,
      COMP_LOOP_COMP_LOOP_and_178_itm, COMP_LOOP_COMP_LOOP_and_302_itm, COMP_LOOP_COMP_LOOP_and_426_itm,
      COMP_LOOP_COMP_LOOP_and_550_itm, COMP_LOOP_COMP_LOOP_and_674_itm, COMP_LOOP_COMP_LOOP_and_798_itm,
      COMP_LOOP_COMP_LOOP_and_922_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_682_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_24_itm,
      COMP_LOOP_COMP_LOOP_and_179_itm, COMP_LOOP_COMP_LOOP_and_303_itm, COMP_LOOP_COMP_LOOP_and_427_itm,
      COMP_LOOP_COMP_LOOP_and_551_itm, COMP_LOOP_COMP_LOOP_and_675_itm, COMP_LOOP_COMP_LOOP_and_799_itm,
      COMP_LOOP_COMP_LOOP_and_923_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_683_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_25_itm,
      COMP_LOOP_COMP_LOOP_and_180_itm, COMP_LOOP_COMP_LOOP_and_304_itm, COMP_LOOP_COMP_LOOP_and_428_itm,
      COMP_LOOP_COMP_LOOP_and_552_itm, COMP_LOOP_COMP_LOOP_and_676_itm, COMP_LOOP_COMP_LOOP_and_800_itm,
      COMP_LOOP_COMP_LOOP_and_924_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_684_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_26_itm,
      COMP_LOOP_COMP_LOOP_and_181_itm, COMP_LOOP_COMP_LOOP_and_305_itm, COMP_LOOP_COMP_LOOP_and_429_itm,
      COMP_LOOP_COMP_LOOP_and_553_itm, COMP_LOOP_COMP_LOOP_and_677_itm, COMP_LOOP_COMP_LOOP_and_801_itm,
      COMP_LOOP_COMP_LOOP_and_925_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_685_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_27_itm,
      COMP_LOOP_COMP_LOOP_and_182_itm, COMP_LOOP_COMP_LOOP_and_306_itm, COMP_LOOP_COMP_LOOP_and_430_itm,
      COMP_LOOP_COMP_LOOP_and_554_itm, COMP_LOOP_COMP_LOOP_and_678_itm, COMP_LOOP_COMP_LOOP_and_802_itm,
      COMP_LOOP_COMP_LOOP_and_926_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_686_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_28_itm,
      COMP_LOOP_COMP_LOOP_and_183_itm, COMP_LOOP_COMP_LOOP_and_307_itm, COMP_LOOP_COMP_LOOP_and_431_itm,
      COMP_LOOP_COMP_LOOP_and_555_itm, COMP_LOOP_COMP_LOOP_and_679_itm, COMP_LOOP_COMP_LOOP_and_803_itm,
      COMP_LOOP_COMP_LOOP_and_927_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_687_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_29_itm,
      COMP_LOOP_COMP_LOOP_and_184_itm, COMP_LOOP_COMP_LOOP_and_308_itm, COMP_LOOP_COMP_LOOP_and_432_itm,
      COMP_LOOP_COMP_LOOP_and_556_itm, COMP_LOOP_COMP_LOOP_and_680_itm, COMP_LOOP_COMP_LOOP_and_804_itm,
      COMP_LOOP_COMP_LOOP_and_928_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign COMP_LOOP_mux1h_688_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_30_itm,
      COMP_LOOP_COMP_LOOP_and_185_itm, COMP_LOOP_COMP_LOOP_and_309_itm, COMP_LOOP_COMP_LOOP_and_433_itm,
      COMP_LOOP_COMP_LOOP_and_557_itm, COMP_LOOP_COMP_LOOP_and_681_itm, COMP_LOOP_COMP_LOOP_and_805_itm,
      COMP_LOOP_COMP_LOOP_and_929_itm, {and_dcpl_479 , and_605_cse , and_609_cse
      , and_614_cse , and_617_cse , and_621_cse , and_624_cse , and_628_cse});
  assign z_out_9 = MUX1HOT_v_64_32_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d, vec_rsc_0_2_i_q_d,
      vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d, vec_rsc_0_6_i_q_d,
      vec_rsc_0_7_i_q_d, vec_rsc_0_8_i_q_d, vec_rsc_0_9_i_q_d, vec_rsc_0_10_i_q_d,
      vec_rsc_0_11_i_q_d, vec_rsc_0_12_i_q_d, vec_rsc_0_13_i_q_d, vec_rsc_0_14_i_q_d,
      vec_rsc_0_15_i_q_d, vec_rsc_0_16_i_q_d, vec_rsc_0_17_i_q_d, vec_rsc_0_18_i_q_d,
      vec_rsc_0_19_i_q_d, vec_rsc_0_20_i_q_d, vec_rsc_0_21_i_q_d, vec_rsc_0_22_i_q_d,
      vec_rsc_0_23_i_q_d, vec_rsc_0_24_i_q_d, vec_rsc_0_25_i_q_d, vec_rsc_0_26_i_q_d,
      vec_rsc_0_27_i_q_d, vec_rsc_0_28_i_q_d, vec_rsc_0_29_i_q_d, vec_rsc_0_30_i_q_d,
      vec_rsc_0_31_i_q_d, {COMP_LOOP_mux1h_657_nl , COMP_LOOP_mux1h_658_nl , COMP_LOOP_mux1h_659_nl
      , COMP_LOOP_mux1h_660_nl , COMP_LOOP_mux1h_661_nl , COMP_LOOP_mux1h_662_nl
      , COMP_LOOP_mux1h_663_nl , COMP_LOOP_mux1h_664_nl , COMP_LOOP_mux1h_665_nl
      , COMP_LOOP_mux1h_666_nl , COMP_LOOP_mux1h_667_nl , COMP_LOOP_mux1h_668_nl
      , COMP_LOOP_mux1h_669_nl , COMP_LOOP_mux1h_670_nl , COMP_LOOP_mux1h_671_nl
      , COMP_LOOP_mux1h_672_nl , COMP_LOOP_mux1h_673_nl , COMP_LOOP_mux1h_674_nl
      , COMP_LOOP_mux1h_675_nl , COMP_LOOP_mux1h_676_nl , COMP_LOOP_mux1h_677_nl
      , COMP_LOOP_mux1h_678_nl , COMP_LOOP_mux1h_679_nl , COMP_LOOP_mux1h_680_nl
      , COMP_LOOP_mux1h_681_nl , COMP_LOOP_mux1h_682_nl , COMP_LOOP_mux1h_683_nl
      , COMP_LOOP_mux1h_684_nl , COMP_LOOP_mux1h_685_nl , COMP_LOOP_mux1h_686_nl
      , COMP_LOOP_mux1h_687_nl , COMP_LOOP_mux1h_688_nl});

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_5_2;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [4:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_8_2;
    input [0:0] input_7;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [7:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    result = result | ( input_7 & {1{sel[7]}});
    MUX1HOT_s_1_8_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_16_2;
    input [4:0] input_15;
    input [4:0] input_14;
    input [4:0] input_13;
    input [4:0] input_12;
    input [4:0] input_11;
    input [4:0] input_10;
    input [4:0] input_9;
    input [4:0] input_8;
    input [4:0] input_7;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [15:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    result = result | ( input_3 & {5{sel[3]}});
    result = result | ( input_4 & {5{sel[4]}});
    result = result | ( input_5 & {5{sel[5]}});
    result = result | ( input_6 & {5{sel[6]}});
    result = result | ( input_7 & {5{sel[7]}});
    result = result | ( input_8 & {5{sel[8]}});
    result = result | ( input_9 & {5{sel[9]}});
    result = result | ( input_10 & {5{sel[10]}});
    result = result | ( input_11 & {5{sel[11]}});
    result = result | ( input_12 & {5{sel[12]}});
    result = result | ( input_13 & {5{sel[13]}});
    result = result | ( input_14 & {5{sel[14]}});
    result = result | ( input_15 & {5{sel[15]}});
    MUX1HOT_v_5_16_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_6_2;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [5:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    result = result | ( input_3 & {5{sel[3]}});
    result = result | ( input_4 & {5{sel[4]}});
    result = result | ( input_5 & {5{sel[5]}});
    MUX1HOT_v_5_6_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_7_2;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [6:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    result = result | ( input_3 & {5{sel[3]}});
    result = result | ( input_4 & {5{sel[4]}});
    result = result | ( input_5 & {5{sel[5]}});
    result = result | ( input_6 & {5{sel[6]}});
    MUX1HOT_v_5_7_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_16_2;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [15:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    MUX1HOT_v_64_16_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_32_2;
    input [63:0] input_31;
    input [63:0] input_30;
    input [63:0] input_29;
    input [63:0] input_28;
    input [63:0] input_27;
    input [63:0] input_26;
    input [63:0] input_25;
    input [63:0] input_24;
    input [63:0] input_23;
    input [63:0] input_22;
    input [63:0] input_21;
    input [63:0] input_20;
    input [63:0] input_19;
    input [63:0] input_18;
    input [63:0] input_17;
    input [63:0] input_16;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [31:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    result = result | ( input_16 & {64{sel[16]}});
    result = result | ( input_17 & {64{sel[17]}});
    result = result | ( input_18 & {64{sel[18]}});
    result = result | ( input_19 & {64{sel[19]}});
    result = result | ( input_20 & {64{sel[20]}});
    result = result | ( input_21 & {64{sel[21]}});
    result = result | ( input_22 & {64{sel[22]}});
    result = result | ( input_23 & {64{sel[23]}});
    result = result | ( input_24 & {64{sel[24]}});
    result = result | ( input_25 & {64{sel[25]}});
    result = result | ( input_26 & {64{sel[26]}});
    result = result | ( input_27 & {64{sel[27]}});
    result = result | ( input_28 & {64{sel[28]}});
    result = result | ( input_29 & {64{sel[29]}});
    result = result | ( input_30 & {64{sel[30]}});
    result = result | ( input_31 & {64{sel[31]}});
    MUX1HOT_v_64_32_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_33_2;
    input [63:0] input_32;
    input [63:0] input_31;
    input [63:0] input_30;
    input [63:0] input_29;
    input [63:0] input_28;
    input [63:0] input_27;
    input [63:0] input_26;
    input [63:0] input_25;
    input [63:0] input_24;
    input [63:0] input_23;
    input [63:0] input_22;
    input [63:0] input_21;
    input [63:0] input_20;
    input [63:0] input_19;
    input [63:0] input_18;
    input [63:0] input_17;
    input [63:0] input_16;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [32:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    result = result | ( input_16 & {64{sel[16]}});
    result = result | ( input_17 & {64{sel[17]}});
    result = result | ( input_18 & {64{sel[18]}});
    result = result | ( input_19 & {64{sel[19]}});
    result = result | ( input_20 & {64{sel[20]}});
    result = result | ( input_21 & {64{sel[21]}});
    result = result | ( input_22 & {64{sel[22]}});
    result = result | ( input_23 & {64{sel[23]}});
    result = result | ( input_24 & {64{sel[24]}});
    result = result | ( input_25 & {64{sel[25]}});
    result = result | ( input_26 & {64{sel[26]}});
    result = result | ( input_27 & {64{sel[27]}});
    result = result | ( input_28 & {64{sel[28]}});
    result = result | ( input_29 & {64{sel[29]}});
    result = result | ( input_30 & {64{sel[30]}});
    result = result | ( input_31 & {64{sel[31]}});
    result = result | ( input_32 & {64{sel[32]}});
    MUX1HOT_v_64_33_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_36_2;
    input [63:0] input_35;
    input [63:0] input_34;
    input [63:0] input_33;
    input [63:0] input_32;
    input [63:0] input_31;
    input [63:0] input_30;
    input [63:0] input_29;
    input [63:0] input_28;
    input [63:0] input_27;
    input [63:0] input_26;
    input [63:0] input_25;
    input [63:0] input_24;
    input [63:0] input_23;
    input [63:0] input_22;
    input [63:0] input_21;
    input [63:0] input_20;
    input [63:0] input_19;
    input [63:0] input_18;
    input [63:0] input_17;
    input [63:0] input_16;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [35:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    result = result | ( input_16 & {64{sel[16]}});
    result = result | ( input_17 & {64{sel[17]}});
    result = result | ( input_18 & {64{sel[18]}});
    result = result | ( input_19 & {64{sel[19]}});
    result = result | ( input_20 & {64{sel[20]}});
    result = result | ( input_21 & {64{sel[21]}});
    result = result | ( input_22 & {64{sel[22]}});
    result = result | ( input_23 & {64{sel[23]}});
    result = result | ( input_24 & {64{sel[24]}});
    result = result | ( input_25 & {64{sel[25]}});
    result = result | ( input_26 & {64{sel[26]}});
    result = result | ( input_27 & {64{sel[27]}});
    result = result | ( input_28 & {64{sel[28]}});
    result = result | ( input_29 & {64{sel[29]}});
    result = result | ( input_30 & {64{sel[30]}});
    result = result | ( input_31 & {64{sel[31]}});
    result = result | ( input_32 & {64{sel[32]}});
    result = result | ( input_33 & {64{sel[33]}});
    result = result | ( input_34 & {64{sel[34]}});
    result = result | ( input_35 & {64{sel[35]}});
    MUX1HOT_v_64_36_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_4_2;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [3:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    MUX1HOT_v_64_4_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_8_2;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [7:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    MUX1HOT_v_64_8_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_9_2;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [8:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    MUX1HOT_v_64_9_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_4_2;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [3:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    result = result | ( input_3 & {9{sel[3]}});
    MUX1HOT_v_9_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [9:0] readslicef_11_10_1;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_11_10_1 = tmp[9:0];
  end
  endfunction


  function automatic [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function automatic [10:0] readslicef_12_11_1;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_12_11_1 = tmp[10:0];
  end
  endfunction


  function automatic [63:0] readslicef_65_64_1;
    input [64:0] vector;
    reg [64:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_65_64_1 = tmp[63:0];
  end
  endfunction


  function automatic [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_12 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF
// ------------------------------------------------------------------


module inPlaceNTT_DIF (
  clk, rst, vec_rsc_0_0_wadr, vec_rsc_0_0_d, vec_rsc_0_0_we, vec_rsc_0_0_radr, vec_rsc_0_0_q,
      vec_rsc_triosy_0_0_lz, vec_rsc_0_1_wadr, vec_rsc_0_1_d, vec_rsc_0_1_we, vec_rsc_0_1_radr,
      vec_rsc_0_1_q, vec_rsc_triosy_0_1_lz, vec_rsc_0_2_wadr, vec_rsc_0_2_d, vec_rsc_0_2_we,
      vec_rsc_0_2_radr, vec_rsc_0_2_q, vec_rsc_triosy_0_2_lz, vec_rsc_0_3_wadr, vec_rsc_0_3_d,
      vec_rsc_0_3_we, vec_rsc_0_3_radr, vec_rsc_0_3_q, vec_rsc_triosy_0_3_lz, vec_rsc_0_4_wadr,
      vec_rsc_0_4_d, vec_rsc_0_4_we, vec_rsc_0_4_radr, vec_rsc_0_4_q, vec_rsc_triosy_0_4_lz,
      vec_rsc_0_5_wadr, vec_rsc_0_5_d, vec_rsc_0_5_we, vec_rsc_0_5_radr, vec_rsc_0_5_q,
      vec_rsc_triosy_0_5_lz, vec_rsc_0_6_wadr, vec_rsc_0_6_d, vec_rsc_0_6_we, vec_rsc_0_6_radr,
      vec_rsc_0_6_q, vec_rsc_triosy_0_6_lz, vec_rsc_0_7_wadr, vec_rsc_0_7_d, vec_rsc_0_7_we,
      vec_rsc_0_7_radr, vec_rsc_0_7_q, vec_rsc_triosy_0_7_lz, vec_rsc_0_8_wadr, vec_rsc_0_8_d,
      vec_rsc_0_8_we, vec_rsc_0_8_radr, vec_rsc_0_8_q, vec_rsc_triosy_0_8_lz, vec_rsc_0_9_wadr,
      vec_rsc_0_9_d, vec_rsc_0_9_we, vec_rsc_0_9_radr, vec_rsc_0_9_q, vec_rsc_triosy_0_9_lz,
      vec_rsc_0_10_wadr, vec_rsc_0_10_d, vec_rsc_0_10_we, vec_rsc_0_10_radr, vec_rsc_0_10_q,
      vec_rsc_triosy_0_10_lz, vec_rsc_0_11_wadr, vec_rsc_0_11_d, vec_rsc_0_11_we,
      vec_rsc_0_11_radr, vec_rsc_0_11_q, vec_rsc_triosy_0_11_lz, vec_rsc_0_12_wadr,
      vec_rsc_0_12_d, vec_rsc_0_12_we, vec_rsc_0_12_radr, vec_rsc_0_12_q, vec_rsc_triosy_0_12_lz,
      vec_rsc_0_13_wadr, vec_rsc_0_13_d, vec_rsc_0_13_we, vec_rsc_0_13_radr, vec_rsc_0_13_q,
      vec_rsc_triosy_0_13_lz, vec_rsc_0_14_wadr, vec_rsc_0_14_d, vec_rsc_0_14_we,
      vec_rsc_0_14_radr, vec_rsc_0_14_q, vec_rsc_triosy_0_14_lz, vec_rsc_0_15_wadr,
      vec_rsc_0_15_d, vec_rsc_0_15_we, vec_rsc_0_15_radr, vec_rsc_0_15_q, vec_rsc_triosy_0_15_lz,
      vec_rsc_0_16_wadr, vec_rsc_0_16_d, vec_rsc_0_16_we, vec_rsc_0_16_radr, vec_rsc_0_16_q,
      vec_rsc_triosy_0_16_lz, vec_rsc_0_17_wadr, vec_rsc_0_17_d, vec_rsc_0_17_we,
      vec_rsc_0_17_radr, vec_rsc_0_17_q, vec_rsc_triosy_0_17_lz, vec_rsc_0_18_wadr,
      vec_rsc_0_18_d, vec_rsc_0_18_we, vec_rsc_0_18_radr, vec_rsc_0_18_q, vec_rsc_triosy_0_18_lz,
      vec_rsc_0_19_wadr, vec_rsc_0_19_d, vec_rsc_0_19_we, vec_rsc_0_19_radr, vec_rsc_0_19_q,
      vec_rsc_triosy_0_19_lz, vec_rsc_0_20_wadr, vec_rsc_0_20_d, vec_rsc_0_20_we,
      vec_rsc_0_20_radr, vec_rsc_0_20_q, vec_rsc_triosy_0_20_lz, vec_rsc_0_21_wadr,
      vec_rsc_0_21_d, vec_rsc_0_21_we, vec_rsc_0_21_radr, vec_rsc_0_21_q, vec_rsc_triosy_0_21_lz,
      vec_rsc_0_22_wadr, vec_rsc_0_22_d, vec_rsc_0_22_we, vec_rsc_0_22_radr, vec_rsc_0_22_q,
      vec_rsc_triosy_0_22_lz, vec_rsc_0_23_wadr, vec_rsc_0_23_d, vec_rsc_0_23_we,
      vec_rsc_0_23_radr, vec_rsc_0_23_q, vec_rsc_triosy_0_23_lz, vec_rsc_0_24_wadr,
      vec_rsc_0_24_d, vec_rsc_0_24_we, vec_rsc_0_24_radr, vec_rsc_0_24_q, vec_rsc_triosy_0_24_lz,
      vec_rsc_0_25_wadr, vec_rsc_0_25_d, vec_rsc_0_25_we, vec_rsc_0_25_radr, vec_rsc_0_25_q,
      vec_rsc_triosy_0_25_lz, vec_rsc_0_26_wadr, vec_rsc_0_26_d, vec_rsc_0_26_we,
      vec_rsc_0_26_radr, vec_rsc_0_26_q, vec_rsc_triosy_0_26_lz, vec_rsc_0_27_wadr,
      vec_rsc_0_27_d, vec_rsc_0_27_we, vec_rsc_0_27_radr, vec_rsc_0_27_q, vec_rsc_triosy_0_27_lz,
      vec_rsc_0_28_wadr, vec_rsc_0_28_d, vec_rsc_0_28_we, vec_rsc_0_28_radr, vec_rsc_0_28_q,
      vec_rsc_triosy_0_28_lz, vec_rsc_0_29_wadr, vec_rsc_0_29_d, vec_rsc_0_29_we,
      vec_rsc_0_29_radr, vec_rsc_0_29_q, vec_rsc_triosy_0_29_lz, vec_rsc_0_30_wadr,
      vec_rsc_0_30_d, vec_rsc_0_30_we, vec_rsc_0_30_radr, vec_rsc_0_30_q, vec_rsc_triosy_0_30_lz,
      vec_rsc_0_31_wadr, vec_rsc_0_31_d, vec_rsc_0_31_we, vec_rsc_0_31_radr, vec_rsc_0_31_q,
      vec_rsc_triosy_0_31_lz, p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz,
      twiddle_rsc_0_0_radr, twiddle_rsc_0_0_q, twiddle_rsc_triosy_0_0_lz, twiddle_rsc_0_1_radr,
      twiddle_rsc_0_1_q, twiddle_rsc_triosy_0_1_lz, twiddle_rsc_0_2_radr, twiddle_rsc_0_2_q,
      twiddle_rsc_triosy_0_2_lz, twiddle_rsc_0_3_radr, twiddle_rsc_0_3_q, twiddle_rsc_triosy_0_3_lz,
      twiddle_rsc_0_4_radr, twiddle_rsc_0_4_q, twiddle_rsc_triosy_0_4_lz, twiddle_rsc_0_5_radr,
      twiddle_rsc_0_5_q, twiddle_rsc_triosy_0_5_lz, twiddle_rsc_0_6_radr, twiddle_rsc_0_6_q,
      twiddle_rsc_triosy_0_6_lz, twiddle_rsc_0_7_radr, twiddle_rsc_0_7_q, twiddle_rsc_triosy_0_7_lz,
      twiddle_rsc_0_8_radr, twiddle_rsc_0_8_q, twiddle_rsc_triosy_0_8_lz, twiddle_rsc_0_9_radr,
      twiddle_rsc_0_9_q, twiddle_rsc_triosy_0_9_lz, twiddle_rsc_0_10_radr, twiddle_rsc_0_10_q,
      twiddle_rsc_triosy_0_10_lz, twiddle_rsc_0_11_radr, twiddle_rsc_0_11_q, twiddle_rsc_triosy_0_11_lz,
      twiddle_rsc_0_12_radr, twiddle_rsc_0_12_q, twiddle_rsc_triosy_0_12_lz, twiddle_rsc_0_13_radr,
      twiddle_rsc_0_13_q, twiddle_rsc_triosy_0_13_lz, twiddle_rsc_0_14_radr, twiddle_rsc_0_14_q,
      twiddle_rsc_triosy_0_14_lz, twiddle_rsc_0_15_radr, twiddle_rsc_0_15_q, twiddle_rsc_triosy_0_15_lz,
      twiddle_rsc_0_16_radr, twiddle_rsc_0_16_q, twiddle_rsc_triosy_0_16_lz, twiddle_rsc_0_17_radr,
      twiddle_rsc_0_17_q, twiddle_rsc_triosy_0_17_lz, twiddle_rsc_0_18_radr, twiddle_rsc_0_18_q,
      twiddle_rsc_triosy_0_18_lz, twiddle_rsc_0_19_radr, twiddle_rsc_0_19_q, twiddle_rsc_triosy_0_19_lz,
      twiddle_rsc_0_20_radr, twiddle_rsc_0_20_q, twiddle_rsc_triosy_0_20_lz, twiddle_rsc_0_21_radr,
      twiddle_rsc_0_21_q, twiddle_rsc_triosy_0_21_lz, twiddle_rsc_0_22_radr, twiddle_rsc_0_22_q,
      twiddle_rsc_triosy_0_22_lz, twiddle_rsc_0_23_radr, twiddle_rsc_0_23_q, twiddle_rsc_triosy_0_23_lz,
      twiddle_rsc_0_24_radr, twiddle_rsc_0_24_q, twiddle_rsc_triosy_0_24_lz, twiddle_rsc_0_25_radr,
      twiddle_rsc_0_25_q, twiddle_rsc_triosy_0_25_lz, twiddle_rsc_0_26_radr, twiddle_rsc_0_26_q,
      twiddle_rsc_triosy_0_26_lz, twiddle_rsc_0_27_radr, twiddle_rsc_0_27_q, twiddle_rsc_triosy_0_27_lz,
      twiddle_rsc_0_28_radr, twiddle_rsc_0_28_q, twiddle_rsc_triosy_0_28_lz, twiddle_rsc_0_29_radr,
      twiddle_rsc_0_29_q, twiddle_rsc_triosy_0_29_lz, twiddle_rsc_0_30_radr, twiddle_rsc_0_30_q,
      twiddle_rsc_triosy_0_30_lz, twiddle_rsc_0_31_radr, twiddle_rsc_0_31_q, twiddle_rsc_triosy_0_31_lz
);
  input clk;
  input rst;
  output [4:0] vec_rsc_0_0_wadr;
  output [63:0] vec_rsc_0_0_d;
  output vec_rsc_0_0_we;
  output [4:0] vec_rsc_0_0_radr;
  input [63:0] vec_rsc_0_0_q;
  output vec_rsc_triosy_0_0_lz;
  output [4:0] vec_rsc_0_1_wadr;
  output [63:0] vec_rsc_0_1_d;
  output vec_rsc_0_1_we;
  output [4:0] vec_rsc_0_1_radr;
  input [63:0] vec_rsc_0_1_q;
  output vec_rsc_triosy_0_1_lz;
  output [4:0] vec_rsc_0_2_wadr;
  output [63:0] vec_rsc_0_2_d;
  output vec_rsc_0_2_we;
  output [4:0] vec_rsc_0_2_radr;
  input [63:0] vec_rsc_0_2_q;
  output vec_rsc_triosy_0_2_lz;
  output [4:0] vec_rsc_0_3_wadr;
  output [63:0] vec_rsc_0_3_d;
  output vec_rsc_0_3_we;
  output [4:0] vec_rsc_0_3_radr;
  input [63:0] vec_rsc_0_3_q;
  output vec_rsc_triosy_0_3_lz;
  output [4:0] vec_rsc_0_4_wadr;
  output [63:0] vec_rsc_0_4_d;
  output vec_rsc_0_4_we;
  output [4:0] vec_rsc_0_4_radr;
  input [63:0] vec_rsc_0_4_q;
  output vec_rsc_triosy_0_4_lz;
  output [4:0] vec_rsc_0_5_wadr;
  output [63:0] vec_rsc_0_5_d;
  output vec_rsc_0_5_we;
  output [4:0] vec_rsc_0_5_radr;
  input [63:0] vec_rsc_0_5_q;
  output vec_rsc_triosy_0_5_lz;
  output [4:0] vec_rsc_0_6_wadr;
  output [63:0] vec_rsc_0_6_d;
  output vec_rsc_0_6_we;
  output [4:0] vec_rsc_0_6_radr;
  input [63:0] vec_rsc_0_6_q;
  output vec_rsc_triosy_0_6_lz;
  output [4:0] vec_rsc_0_7_wadr;
  output [63:0] vec_rsc_0_7_d;
  output vec_rsc_0_7_we;
  output [4:0] vec_rsc_0_7_radr;
  input [63:0] vec_rsc_0_7_q;
  output vec_rsc_triosy_0_7_lz;
  output [4:0] vec_rsc_0_8_wadr;
  output [63:0] vec_rsc_0_8_d;
  output vec_rsc_0_8_we;
  output [4:0] vec_rsc_0_8_radr;
  input [63:0] vec_rsc_0_8_q;
  output vec_rsc_triosy_0_8_lz;
  output [4:0] vec_rsc_0_9_wadr;
  output [63:0] vec_rsc_0_9_d;
  output vec_rsc_0_9_we;
  output [4:0] vec_rsc_0_9_radr;
  input [63:0] vec_rsc_0_9_q;
  output vec_rsc_triosy_0_9_lz;
  output [4:0] vec_rsc_0_10_wadr;
  output [63:0] vec_rsc_0_10_d;
  output vec_rsc_0_10_we;
  output [4:0] vec_rsc_0_10_radr;
  input [63:0] vec_rsc_0_10_q;
  output vec_rsc_triosy_0_10_lz;
  output [4:0] vec_rsc_0_11_wadr;
  output [63:0] vec_rsc_0_11_d;
  output vec_rsc_0_11_we;
  output [4:0] vec_rsc_0_11_radr;
  input [63:0] vec_rsc_0_11_q;
  output vec_rsc_triosy_0_11_lz;
  output [4:0] vec_rsc_0_12_wadr;
  output [63:0] vec_rsc_0_12_d;
  output vec_rsc_0_12_we;
  output [4:0] vec_rsc_0_12_radr;
  input [63:0] vec_rsc_0_12_q;
  output vec_rsc_triosy_0_12_lz;
  output [4:0] vec_rsc_0_13_wadr;
  output [63:0] vec_rsc_0_13_d;
  output vec_rsc_0_13_we;
  output [4:0] vec_rsc_0_13_radr;
  input [63:0] vec_rsc_0_13_q;
  output vec_rsc_triosy_0_13_lz;
  output [4:0] vec_rsc_0_14_wadr;
  output [63:0] vec_rsc_0_14_d;
  output vec_rsc_0_14_we;
  output [4:0] vec_rsc_0_14_radr;
  input [63:0] vec_rsc_0_14_q;
  output vec_rsc_triosy_0_14_lz;
  output [4:0] vec_rsc_0_15_wadr;
  output [63:0] vec_rsc_0_15_d;
  output vec_rsc_0_15_we;
  output [4:0] vec_rsc_0_15_radr;
  input [63:0] vec_rsc_0_15_q;
  output vec_rsc_triosy_0_15_lz;
  output [4:0] vec_rsc_0_16_wadr;
  output [63:0] vec_rsc_0_16_d;
  output vec_rsc_0_16_we;
  output [4:0] vec_rsc_0_16_radr;
  input [63:0] vec_rsc_0_16_q;
  output vec_rsc_triosy_0_16_lz;
  output [4:0] vec_rsc_0_17_wadr;
  output [63:0] vec_rsc_0_17_d;
  output vec_rsc_0_17_we;
  output [4:0] vec_rsc_0_17_radr;
  input [63:0] vec_rsc_0_17_q;
  output vec_rsc_triosy_0_17_lz;
  output [4:0] vec_rsc_0_18_wadr;
  output [63:0] vec_rsc_0_18_d;
  output vec_rsc_0_18_we;
  output [4:0] vec_rsc_0_18_radr;
  input [63:0] vec_rsc_0_18_q;
  output vec_rsc_triosy_0_18_lz;
  output [4:0] vec_rsc_0_19_wadr;
  output [63:0] vec_rsc_0_19_d;
  output vec_rsc_0_19_we;
  output [4:0] vec_rsc_0_19_radr;
  input [63:0] vec_rsc_0_19_q;
  output vec_rsc_triosy_0_19_lz;
  output [4:0] vec_rsc_0_20_wadr;
  output [63:0] vec_rsc_0_20_d;
  output vec_rsc_0_20_we;
  output [4:0] vec_rsc_0_20_radr;
  input [63:0] vec_rsc_0_20_q;
  output vec_rsc_triosy_0_20_lz;
  output [4:0] vec_rsc_0_21_wadr;
  output [63:0] vec_rsc_0_21_d;
  output vec_rsc_0_21_we;
  output [4:0] vec_rsc_0_21_radr;
  input [63:0] vec_rsc_0_21_q;
  output vec_rsc_triosy_0_21_lz;
  output [4:0] vec_rsc_0_22_wadr;
  output [63:0] vec_rsc_0_22_d;
  output vec_rsc_0_22_we;
  output [4:0] vec_rsc_0_22_radr;
  input [63:0] vec_rsc_0_22_q;
  output vec_rsc_triosy_0_22_lz;
  output [4:0] vec_rsc_0_23_wadr;
  output [63:0] vec_rsc_0_23_d;
  output vec_rsc_0_23_we;
  output [4:0] vec_rsc_0_23_radr;
  input [63:0] vec_rsc_0_23_q;
  output vec_rsc_triosy_0_23_lz;
  output [4:0] vec_rsc_0_24_wadr;
  output [63:0] vec_rsc_0_24_d;
  output vec_rsc_0_24_we;
  output [4:0] vec_rsc_0_24_radr;
  input [63:0] vec_rsc_0_24_q;
  output vec_rsc_triosy_0_24_lz;
  output [4:0] vec_rsc_0_25_wadr;
  output [63:0] vec_rsc_0_25_d;
  output vec_rsc_0_25_we;
  output [4:0] vec_rsc_0_25_radr;
  input [63:0] vec_rsc_0_25_q;
  output vec_rsc_triosy_0_25_lz;
  output [4:0] vec_rsc_0_26_wadr;
  output [63:0] vec_rsc_0_26_d;
  output vec_rsc_0_26_we;
  output [4:0] vec_rsc_0_26_radr;
  input [63:0] vec_rsc_0_26_q;
  output vec_rsc_triosy_0_26_lz;
  output [4:0] vec_rsc_0_27_wadr;
  output [63:0] vec_rsc_0_27_d;
  output vec_rsc_0_27_we;
  output [4:0] vec_rsc_0_27_radr;
  input [63:0] vec_rsc_0_27_q;
  output vec_rsc_triosy_0_27_lz;
  output [4:0] vec_rsc_0_28_wadr;
  output [63:0] vec_rsc_0_28_d;
  output vec_rsc_0_28_we;
  output [4:0] vec_rsc_0_28_radr;
  input [63:0] vec_rsc_0_28_q;
  output vec_rsc_triosy_0_28_lz;
  output [4:0] vec_rsc_0_29_wadr;
  output [63:0] vec_rsc_0_29_d;
  output vec_rsc_0_29_we;
  output [4:0] vec_rsc_0_29_radr;
  input [63:0] vec_rsc_0_29_q;
  output vec_rsc_triosy_0_29_lz;
  output [4:0] vec_rsc_0_30_wadr;
  output [63:0] vec_rsc_0_30_d;
  output vec_rsc_0_30_we;
  output [4:0] vec_rsc_0_30_radr;
  input [63:0] vec_rsc_0_30_q;
  output vec_rsc_triosy_0_30_lz;
  output [4:0] vec_rsc_0_31_wadr;
  output [63:0] vec_rsc_0_31_d;
  output vec_rsc_0_31_we;
  output [4:0] vec_rsc_0_31_radr;
  input [63:0] vec_rsc_0_31_q;
  output vec_rsc_triosy_0_31_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  output [4:0] twiddle_rsc_0_0_radr;
  input [63:0] twiddle_rsc_0_0_q;
  output twiddle_rsc_triosy_0_0_lz;
  output [4:0] twiddle_rsc_0_1_radr;
  input [63:0] twiddle_rsc_0_1_q;
  output twiddle_rsc_triosy_0_1_lz;
  output [4:0] twiddle_rsc_0_2_radr;
  input [63:0] twiddle_rsc_0_2_q;
  output twiddle_rsc_triosy_0_2_lz;
  output [4:0] twiddle_rsc_0_3_radr;
  input [63:0] twiddle_rsc_0_3_q;
  output twiddle_rsc_triosy_0_3_lz;
  output [4:0] twiddle_rsc_0_4_radr;
  input [63:0] twiddle_rsc_0_4_q;
  output twiddle_rsc_triosy_0_4_lz;
  output [4:0] twiddle_rsc_0_5_radr;
  input [63:0] twiddle_rsc_0_5_q;
  output twiddle_rsc_triosy_0_5_lz;
  output [4:0] twiddle_rsc_0_6_radr;
  input [63:0] twiddle_rsc_0_6_q;
  output twiddle_rsc_triosy_0_6_lz;
  output [4:0] twiddle_rsc_0_7_radr;
  input [63:0] twiddle_rsc_0_7_q;
  output twiddle_rsc_triosy_0_7_lz;
  output [4:0] twiddle_rsc_0_8_radr;
  input [63:0] twiddle_rsc_0_8_q;
  output twiddle_rsc_triosy_0_8_lz;
  output [4:0] twiddle_rsc_0_9_radr;
  input [63:0] twiddle_rsc_0_9_q;
  output twiddle_rsc_triosy_0_9_lz;
  output [4:0] twiddle_rsc_0_10_radr;
  input [63:0] twiddle_rsc_0_10_q;
  output twiddle_rsc_triosy_0_10_lz;
  output [4:0] twiddle_rsc_0_11_radr;
  input [63:0] twiddle_rsc_0_11_q;
  output twiddle_rsc_triosy_0_11_lz;
  output [4:0] twiddle_rsc_0_12_radr;
  input [63:0] twiddle_rsc_0_12_q;
  output twiddle_rsc_triosy_0_12_lz;
  output [4:0] twiddle_rsc_0_13_radr;
  input [63:0] twiddle_rsc_0_13_q;
  output twiddle_rsc_triosy_0_13_lz;
  output [4:0] twiddle_rsc_0_14_radr;
  input [63:0] twiddle_rsc_0_14_q;
  output twiddle_rsc_triosy_0_14_lz;
  output [4:0] twiddle_rsc_0_15_radr;
  input [63:0] twiddle_rsc_0_15_q;
  output twiddle_rsc_triosy_0_15_lz;
  output [4:0] twiddle_rsc_0_16_radr;
  input [63:0] twiddle_rsc_0_16_q;
  output twiddle_rsc_triosy_0_16_lz;
  output [4:0] twiddle_rsc_0_17_radr;
  input [63:0] twiddle_rsc_0_17_q;
  output twiddle_rsc_triosy_0_17_lz;
  output [4:0] twiddle_rsc_0_18_radr;
  input [63:0] twiddle_rsc_0_18_q;
  output twiddle_rsc_triosy_0_18_lz;
  output [4:0] twiddle_rsc_0_19_radr;
  input [63:0] twiddle_rsc_0_19_q;
  output twiddle_rsc_triosy_0_19_lz;
  output [4:0] twiddle_rsc_0_20_radr;
  input [63:0] twiddle_rsc_0_20_q;
  output twiddle_rsc_triosy_0_20_lz;
  output [4:0] twiddle_rsc_0_21_radr;
  input [63:0] twiddle_rsc_0_21_q;
  output twiddle_rsc_triosy_0_21_lz;
  output [4:0] twiddle_rsc_0_22_radr;
  input [63:0] twiddle_rsc_0_22_q;
  output twiddle_rsc_triosy_0_22_lz;
  output [4:0] twiddle_rsc_0_23_radr;
  input [63:0] twiddle_rsc_0_23_q;
  output twiddle_rsc_triosy_0_23_lz;
  output [4:0] twiddle_rsc_0_24_radr;
  input [63:0] twiddle_rsc_0_24_q;
  output twiddle_rsc_triosy_0_24_lz;
  output [4:0] twiddle_rsc_0_25_radr;
  input [63:0] twiddle_rsc_0_25_q;
  output twiddle_rsc_triosy_0_25_lz;
  output [4:0] twiddle_rsc_0_26_radr;
  input [63:0] twiddle_rsc_0_26_q;
  output twiddle_rsc_triosy_0_26_lz;
  output [4:0] twiddle_rsc_0_27_radr;
  input [63:0] twiddle_rsc_0_27_q;
  output twiddle_rsc_triosy_0_27_lz;
  output [4:0] twiddle_rsc_0_28_radr;
  input [63:0] twiddle_rsc_0_28_q;
  output twiddle_rsc_triosy_0_28_lz;
  output [4:0] twiddle_rsc_0_29_radr;
  input [63:0] twiddle_rsc_0_29_q;
  output twiddle_rsc_triosy_0_29_lz;
  output [4:0] twiddle_rsc_0_30_radr;
  input [63:0] twiddle_rsc_0_30_q;
  output twiddle_rsc_triosy_0_30_lz;
  output [4:0] twiddle_rsc_0_31_radr;
  input [63:0] twiddle_rsc_0_31_q;
  output twiddle_rsc_triosy_0_31_lz;


  // Interconnect Declarations
  wire [63:0] vec_rsc_0_0_i_q_d;
  wire vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_1_i_q_d;
  wire vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_2_i_q_d;
  wire vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_3_i_q_d;
  wire vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_4_i_q_d;
  wire vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_5_i_q_d;
  wire vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_6_i_q_d;
  wire vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_7_i_q_d;
  wire vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_8_i_q_d;
  wire vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_9_i_q_d;
  wire vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_10_i_q_d;
  wire vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_11_i_q_d;
  wire vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_12_i_q_d;
  wire vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_13_i_q_d;
  wire vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_14_i_q_d;
  wire vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_15_i_q_d;
  wire vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_16_i_q_d;
  wire vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_17_i_q_d;
  wire vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_18_i_q_d;
  wire vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_19_i_q_d;
  wire vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_20_i_q_d;
  wire vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_21_i_q_d;
  wire vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_22_i_q_d;
  wire vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_23_i_q_d;
  wire vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_24_i_q_d;
  wire vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_25_i_q_d;
  wire vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_26_i_q_d;
  wire vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_27_i_q_d;
  wire vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_28_i_q_d;
  wire vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_29_i_q_d;
  wire vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_30_i_q_d;
  wire vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_31_i_q_d;
  wire vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_0_i_q_d;
  wire twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_1_i_q_d;
  wire twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_2_i_q_d;
  wire twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_3_i_q_d;
  wire twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_4_i_q_d;
  wire twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_5_i_q_d;
  wire twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_6_i_q_d;
  wire twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_7_i_q_d;
  wire twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_8_i_q_d;
  wire twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_9_i_q_d;
  wire twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_10_i_q_d;
  wire twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_11_i_q_d;
  wire twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_12_i_q_d;
  wire twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_13_i_q_d;
  wire twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_14_i_q_d;
  wire twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_15_i_q_d;
  wire twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_16_i_q_d;
  wire twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_17_i_q_d;
  wire twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_18_i_q_d;
  wire twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_19_i_q_d;
  wire twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_20_i_q_d;
  wire twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_21_i_q_d;
  wire twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_22_i_q_d;
  wire twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_23_i_q_d;
  wire twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_24_i_q_d;
  wire twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_25_i_q_d;
  wire twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_26_i_q_d;
  wire twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_27_i_q_d;
  wire twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_28_i_q_d;
  wire twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_29_i_q_d;
  wire twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_30_i_q_d;
  wire twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_31_i_q_d;
  wire twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_0_i_d_d_iff;
  wire [4:0] vec_rsc_0_0_i_radr_d_iff;
  wire [4:0] vec_rsc_0_0_i_wadr_d_iff;
  wire vec_rsc_0_0_i_we_d_iff;
  wire vec_rsc_0_1_i_we_d_iff;
  wire vec_rsc_0_2_i_we_d_iff;
  wire vec_rsc_0_3_i_we_d_iff;
  wire vec_rsc_0_4_i_we_d_iff;
  wire vec_rsc_0_5_i_we_d_iff;
  wire vec_rsc_0_6_i_we_d_iff;
  wire vec_rsc_0_7_i_we_d_iff;
  wire vec_rsc_0_8_i_we_d_iff;
  wire vec_rsc_0_9_i_we_d_iff;
  wire vec_rsc_0_10_i_we_d_iff;
  wire vec_rsc_0_11_i_we_d_iff;
  wire vec_rsc_0_12_i_we_d_iff;
  wire vec_rsc_0_13_i_we_d_iff;
  wire vec_rsc_0_14_i_we_d_iff;
  wire vec_rsc_0_15_i_we_d_iff;
  wire vec_rsc_0_16_i_we_d_iff;
  wire vec_rsc_0_17_i_we_d_iff;
  wire vec_rsc_0_18_i_we_d_iff;
  wire vec_rsc_0_19_i_we_d_iff;
  wire vec_rsc_0_20_i_we_d_iff;
  wire vec_rsc_0_21_i_we_d_iff;
  wire vec_rsc_0_22_i_we_d_iff;
  wire vec_rsc_0_23_i_we_d_iff;
  wire vec_rsc_0_24_i_we_d_iff;
  wire vec_rsc_0_25_i_we_d_iff;
  wire vec_rsc_0_26_i_we_d_iff;
  wire vec_rsc_0_27_i_we_d_iff;
  wire vec_rsc_0_28_i_we_d_iff;
  wire vec_rsc_0_29_i_we_d_iff;
  wire vec_rsc_0_30_i_we_d_iff;
  wire vec_rsc_0_31_i_we_d_iff;
  wire [4:0] twiddle_rsc_0_0_i_radr_d_iff;
  wire [4:0] twiddle_rsc_0_1_i_radr_d_iff;
  wire [4:0] twiddle_rsc_0_2_i_radr_d_iff;
  wire [4:0] twiddle_rsc_0_4_i_radr_d_iff;


  // Interconnect Declarations for Component Instantiations 
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_5_64_32_32_64_1_gen vec_rsc_0_0_i
      (
      .q(vec_rsc_0_0_q),
      .radr(vec_rsc_0_0_radr),
      .we(vec_rsc_0_0_we),
      .d(vec_rsc_0_0_d),
      .wadr(vec_rsc_0_0_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_0_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_5_64_32_32_64_1_gen vec_rsc_0_1_i
      (
      .q(vec_rsc_0_1_q),
      .radr(vec_rsc_0_1_radr),
      .we(vec_rsc_0_1_we),
      .d(vec_rsc_0_1_d),
      .wadr(vec_rsc_0_1_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_1_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_1_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_1_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_5_64_32_32_64_1_gen vec_rsc_0_2_i
      (
      .q(vec_rsc_0_2_q),
      .radr(vec_rsc_0_2_radr),
      .we(vec_rsc_0_2_we),
      .d(vec_rsc_0_2_d),
      .wadr(vec_rsc_0_2_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_2_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_2_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_2_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_5_64_32_32_64_1_gen vec_rsc_0_3_i
      (
      .q(vec_rsc_0_3_q),
      .radr(vec_rsc_0_3_radr),
      .we(vec_rsc_0_3_we),
      .d(vec_rsc_0_3_d),
      .wadr(vec_rsc_0_3_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_3_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_3_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_3_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_5_64_32_32_64_1_gen vec_rsc_0_4_i
      (
      .q(vec_rsc_0_4_q),
      .radr(vec_rsc_0_4_radr),
      .we(vec_rsc_0_4_we),
      .d(vec_rsc_0_4_d),
      .wadr(vec_rsc_0_4_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_4_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_4_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_4_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_5_64_32_32_64_1_gen vec_rsc_0_5_i
      (
      .q(vec_rsc_0_5_q),
      .radr(vec_rsc_0_5_radr),
      .we(vec_rsc_0_5_we),
      .d(vec_rsc_0_5_d),
      .wadr(vec_rsc_0_5_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_5_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_5_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_5_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_5_64_32_32_64_1_gen vec_rsc_0_6_i
      (
      .q(vec_rsc_0_6_q),
      .radr(vec_rsc_0_6_radr),
      .we(vec_rsc_0_6_we),
      .d(vec_rsc_0_6_d),
      .wadr(vec_rsc_0_6_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_6_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_6_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_6_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_5_64_32_32_64_1_gen vec_rsc_0_7_i
      (
      .q(vec_rsc_0_7_q),
      .radr(vec_rsc_0_7_radr),
      .we(vec_rsc_0_7_we),
      .d(vec_rsc_0_7_d),
      .wadr(vec_rsc_0_7_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_7_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_7_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_7_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_5_64_32_32_64_1_gen vec_rsc_0_8_i
      (
      .q(vec_rsc_0_8_q),
      .radr(vec_rsc_0_8_radr),
      .we(vec_rsc_0_8_we),
      .d(vec_rsc_0_8_d),
      .wadr(vec_rsc_0_8_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_8_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_8_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_8_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_5_64_32_32_64_1_gen vec_rsc_0_9_i
      (
      .q(vec_rsc_0_9_q),
      .radr(vec_rsc_0_9_radr),
      .we(vec_rsc_0_9_we),
      .d(vec_rsc_0_9_d),
      .wadr(vec_rsc_0_9_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_9_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_9_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_9_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_5_64_32_32_64_1_gen vec_rsc_0_10_i
      (
      .q(vec_rsc_0_10_q),
      .radr(vec_rsc_0_10_radr),
      .we(vec_rsc_0_10_we),
      .d(vec_rsc_0_10_d),
      .wadr(vec_rsc_0_10_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_10_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_10_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_10_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_5_64_32_32_64_1_gen vec_rsc_0_11_i
      (
      .q(vec_rsc_0_11_q),
      .radr(vec_rsc_0_11_radr),
      .we(vec_rsc_0_11_we),
      .d(vec_rsc_0_11_d),
      .wadr(vec_rsc_0_11_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_11_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_11_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_11_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_5_64_32_32_64_1_gen vec_rsc_0_12_i
      (
      .q(vec_rsc_0_12_q),
      .radr(vec_rsc_0_12_radr),
      .we(vec_rsc_0_12_we),
      .d(vec_rsc_0_12_d),
      .wadr(vec_rsc_0_12_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_12_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_12_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_12_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_5_64_32_32_64_1_gen vec_rsc_0_13_i
      (
      .q(vec_rsc_0_13_q),
      .radr(vec_rsc_0_13_radr),
      .we(vec_rsc_0_13_we),
      .d(vec_rsc_0_13_d),
      .wadr(vec_rsc_0_13_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_13_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_13_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_13_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_5_64_32_32_64_1_gen vec_rsc_0_14_i
      (
      .q(vec_rsc_0_14_q),
      .radr(vec_rsc_0_14_radr),
      .we(vec_rsc_0_14_we),
      .d(vec_rsc_0_14_d),
      .wadr(vec_rsc_0_14_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_14_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_14_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_14_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_5_64_32_32_64_1_gen vec_rsc_0_15_i
      (
      .q(vec_rsc_0_15_q),
      .radr(vec_rsc_0_15_radr),
      .we(vec_rsc_0_15_we),
      .d(vec_rsc_0_15_d),
      .wadr(vec_rsc_0_15_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_15_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_15_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_15_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_5_64_32_32_64_1_gen vec_rsc_0_16_i
      (
      .q(vec_rsc_0_16_q),
      .radr(vec_rsc_0_16_radr),
      .we(vec_rsc_0_16_we),
      .d(vec_rsc_0_16_d),
      .wadr(vec_rsc_0_16_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_16_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_5_64_32_32_64_1_gen vec_rsc_0_17_i
      (
      .q(vec_rsc_0_17_q),
      .radr(vec_rsc_0_17_radr),
      .we(vec_rsc_0_17_we),
      .d(vec_rsc_0_17_d),
      .wadr(vec_rsc_0_17_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_17_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_17_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_17_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_5_64_32_32_64_1_gen vec_rsc_0_18_i
      (
      .q(vec_rsc_0_18_q),
      .radr(vec_rsc_0_18_radr),
      .we(vec_rsc_0_18_we),
      .d(vec_rsc_0_18_d),
      .wadr(vec_rsc_0_18_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_18_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_18_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_18_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_5_64_32_32_64_1_gen vec_rsc_0_19_i
      (
      .q(vec_rsc_0_19_q),
      .radr(vec_rsc_0_19_radr),
      .we(vec_rsc_0_19_we),
      .d(vec_rsc_0_19_d),
      .wadr(vec_rsc_0_19_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_19_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_19_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_19_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_5_64_32_32_64_1_gen vec_rsc_0_20_i
      (
      .q(vec_rsc_0_20_q),
      .radr(vec_rsc_0_20_radr),
      .we(vec_rsc_0_20_we),
      .d(vec_rsc_0_20_d),
      .wadr(vec_rsc_0_20_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_20_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_20_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_20_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_5_64_32_32_64_1_gen vec_rsc_0_21_i
      (
      .q(vec_rsc_0_21_q),
      .radr(vec_rsc_0_21_radr),
      .we(vec_rsc_0_21_we),
      .d(vec_rsc_0_21_d),
      .wadr(vec_rsc_0_21_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_21_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_21_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_21_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_5_64_32_32_64_1_gen vec_rsc_0_22_i
      (
      .q(vec_rsc_0_22_q),
      .radr(vec_rsc_0_22_radr),
      .we(vec_rsc_0_22_we),
      .d(vec_rsc_0_22_d),
      .wadr(vec_rsc_0_22_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_22_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_22_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_22_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_5_64_32_32_64_1_gen vec_rsc_0_23_i
      (
      .q(vec_rsc_0_23_q),
      .radr(vec_rsc_0_23_radr),
      .we(vec_rsc_0_23_we),
      .d(vec_rsc_0_23_d),
      .wadr(vec_rsc_0_23_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_23_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_23_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_23_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_5_64_32_32_64_1_gen vec_rsc_0_24_i
      (
      .q(vec_rsc_0_24_q),
      .radr(vec_rsc_0_24_radr),
      .we(vec_rsc_0_24_we),
      .d(vec_rsc_0_24_d),
      .wadr(vec_rsc_0_24_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_24_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_24_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_24_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_5_64_32_32_64_1_gen vec_rsc_0_25_i
      (
      .q(vec_rsc_0_25_q),
      .radr(vec_rsc_0_25_radr),
      .we(vec_rsc_0_25_we),
      .d(vec_rsc_0_25_d),
      .wadr(vec_rsc_0_25_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_25_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_25_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_25_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_5_64_32_32_64_1_gen vec_rsc_0_26_i
      (
      .q(vec_rsc_0_26_q),
      .radr(vec_rsc_0_26_radr),
      .we(vec_rsc_0_26_we),
      .d(vec_rsc_0_26_d),
      .wadr(vec_rsc_0_26_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_26_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_26_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_26_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_5_64_32_32_64_1_gen vec_rsc_0_27_i
      (
      .q(vec_rsc_0_27_q),
      .radr(vec_rsc_0_27_radr),
      .we(vec_rsc_0_27_we),
      .d(vec_rsc_0_27_d),
      .wadr(vec_rsc_0_27_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_27_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_27_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_27_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_5_64_32_32_64_1_gen vec_rsc_0_28_i
      (
      .q(vec_rsc_0_28_q),
      .radr(vec_rsc_0_28_radr),
      .we(vec_rsc_0_28_we),
      .d(vec_rsc_0_28_d),
      .wadr(vec_rsc_0_28_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_28_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_28_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_28_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_5_64_32_32_64_1_gen vec_rsc_0_29_i
      (
      .q(vec_rsc_0_29_q),
      .radr(vec_rsc_0_29_radr),
      .we(vec_rsc_0_29_we),
      .d(vec_rsc_0_29_d),
      .wadr(vec_rsc_0_29_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_29_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_29_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_29_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_5_64_32_32_64_1_gen vec_rsc_0_30_i
      (
      .q(vec_rsc_0_30_q),
      .radr(vec_rsc_0_30_radr),
      .we(vec_rsc_0_30_we),
      .d(vec_rsc_0_30_d),
      .wadr(vec_rsc_0_30_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_30_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_30_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_30_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_5_64_32_32_64_1_gen vec_rsc_0_31_i
      (
      .q(vec_rsc_0_31_q),
      .radr(vec_rsc_0_31_radr),
      .we(vec_rsc_0_31_we),
      .d(vec_rsc_0_31_d),
      .wadr(vec_rsc_0_31_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_31_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_31_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_31_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_41_5_64_32_32_64_1_gen twiddle_rsc_0_0_i
      (
      .q(twiddle_rsc_0_0_q),
      .radr(twiddle_rsc_0_0_radr),
      .q_d(twiddle_rsc_0_0_i_q_d),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_42_5_64_32_32_64_1_gen twiddle_rsc_0_1_i
      (
      .q(twiddle_rsc_0_1_q),
      .radr(twiddle_rsc_0_1_radr),
      .q_d(twiddle_rsc_0_1_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_43_5_64_32_32_64_1_gen twiddle_rsc_0_2_i
      (
      .q(twiddle_rsc_0_2_q),
      .radr(twiddle_rsc_0_2_radr),
      .q_d(twiddle_rsc_0_2_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_44_5_64_32_32_64_1_gen twiddle_rsc_0_3_i
      (
      .q(twiddle_rsc_0_3_q),
      .radr(twiddle_rsc_0_3_radr),
      .q_d(twiddle_rsc_0_3_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_45_5_64_32_32_64_1_gen twiddle_rsc_0_4_i
      (
      .q(twiddle_rsc_0_4_q),
      .radr(twiddle_rsc_0_4_radr),
      .q_d(twiddle_rsc_0_4_i_q_d),
      .radr_d(twiddle_rsc_0_4_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_46_5_64_32_32_64_1_gen twiddle_rsc_0_5_i
      (
      .q(twiddle_rsc_0_5_q),
      .radr(twiddle_rsc_0_5_radr),
      .q_d(twiddle_rsc_0_5_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_47_5_64_32_32_64_1_gen twiddle_rsc_0_6_i
      (
      .q(twiddle_rsc_0_6_q),
      .radr(twiddle_rsc_0_6_radr),
      .q_d(twiddle_rsc_0_6_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_48_5_64_32_32_64_1_gen twiddle_rsc_0_7_i
      (
      .q(twiddle_rsc_0_7_q),
      .radr(twiddle_rsc_0_7_radr),
      .q_d(twiddle_rsc_0_7_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_49_5_64_32_32_64_1_gen twiddle_rsc_0_8_i
      (
      .q(twiddle_rsc_0_8_q),
      .radr(twiddle_rsc_0_8_radr),
      .q_d(twiddle_rsc_0_8_i_q_d),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_50_5_64_32_32_64_1_gen twiddle_rsc_0_9_i
      (
      .q(twiddle_rsc_0_9_q),
      .radr(twiddle_rsc_0_9_radr),
      .q_d(twiddle_rsc_0_9_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_51_5_64_32_32_64_1_gen twiddle_rsc_0_10_i
      (
      .q(twiddle_rsc_0_10_q),
      .radr(twiddle_rsc_0_10_radr),
      .q_d(twiddle_rsc_0_10_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_52_5_64_32_32_64_1_gen twiddle_rsc_0_11_i
      (
      .q(twiddle_rsc_0_11_q),
      .radr(twiddle_rsc_0_11_radr),
      .q_d(twiddle_rsc_0_11_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_53_5_64_32_32_64_1_gen twiddle_rsc_0_12_i
      (
      .q(twiddle_rsc_0_12_q),
      .radr(twiddle_rsc_0_12_radr),
      .q_d(twiddle_rsc_0_12_i_q_d),
      .radr_d(twiddle_rsc_0_4_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_54_5_64_32_32_64_1_gen twiddle_rsc_0_13_i
      (
      .q(twiddle_rsc_0_13_q),
      .radr(twiddle_rsc_0_13_radr),
      .q_d(twiddle_rsc_0_13_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_55_5_64_32_32_64_1_gen twiddle_rsc_0_14_i
      (
      .q(twiddle_rsc_0_14_q),
      .radr(twiddle_rsc_0_14_radr),
      .q_d(twiddle_rsc_0_14_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_56_5_64_32_32_64_1_gen twiddle_rsc_0_15_i
      (
      .q(twiddle_rsc_0_15_q),
      .radr(twiddle_rsc_0_15_radr),
      .q_d(twiddle_rsc_0_15_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_57_5_64_32_32_64_1_gen twiddle_rsc_0_16_i
      (
      .q(twiddle_rsc_0_16_q),
      .radr(twiddle_rsc_0_16_radr),
      .q_d(twiddle_rsc_0_16_i_q_d),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_58_5_64_32_32_64_1_gen twiddle_rsc_0_17_i
      (
      .q(twiddle_rsc_0_17_q),
      .radr(twiddle_rsc_0_17_radr),
      .q_d(twiddle_rsc_0_17_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_59_5_64_32_32_64_1_gen twiddle_rsc_0_18_i
      (
      .q(twiddle_rsc_0_18_q),
      .radr(twiddle_rsc_0_18_radr),
      .q_d(twiddle_rsc_0_18_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_60_5_64_32_32_64_1_gen twiddle_rsc_0_19_i
      (
      .q(twiddle_rsc_0_19_q),
      .radr(twiddle_rsc_0_19_radr),
      .q_d(twiddle_rsc_0_19_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_61_5_64_32_32_64_1_gen twiddle_rsc_0_20_i
      (
      .q(twiddle_rsc_0_20_q),
      .radr(twiddle_rsc_0_20_radr),
      .q_d(twiddle_rsc_0_20_i_q_d),
      .radr_d(twiddle_rsc_0_4_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_62_5_64_32_32_64_1_gen twiddle_rsc_0_21_i
      (
      .q(twiddle_rsc_0_21_q),
      .radr(twiddle_rsc_0_21_radr),
      .q_d(twiddle_rsc_0_21_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_63_5_64_32_32_64_1_gen twiddle_rsc_0_22_i
      (
      .q(twiddle_rsc_0_22_q),
      .radr(twiddle_rsc_0_22_radr),
      .q_d(twiddle_rsc_0_22_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_64_5_64_32_32_64_1_gen twiddle_rsc_0_23_i
      (
      .q(twiddle_rsc_0_23_q),
      .radr(twiddle_rsc_0_23_radr),
      .q_d(twiddle_rsc_0_23_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_65_5_64_32_32_64_1_gen twiddle_rsc_0_24_i
      (
      .q(twiddle_rsc_0_24_q),
      .radr(twiddle_rsc_0_24_radr),
      .q_d(twiddle_rsc_0_24_i_q_d),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_66_5_64_32_32_64_1_gen twiddle_rsc_0_25_i
      (
      .q(twiddle_rsc_0_25_q),
      .radr(twiddle_rsc_0_25_radr),
      .q_d(twiddle_rsc_0_25_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_67_5_64_32_32_64_1_gen twiddle_rsc_0_26_i
      (
      .q(twiddle_rsc_0_26_q),
      .radr(twiddle_rsc_0_26_radr),
      .q_d(twiddle_rsc_0_26_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_68_5_64_32_32_64_1_gen twiddle_rsc_0_27_i
      (
      .q(twiddle_rsc_0_27_q),
      .radr(twiddle_rsc_0_27_radr),
      .q_d(twiddle_rsc_0_27_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_69_5_64_32_32_64_1_gen twiddle_rsc_0_28_i
      (
      .q(twiddle_rsc_0_28_q),
      .radr(twiddle_rsc_0_28_radr),
      .q_d(twiddle_rsc_0_28_i_q_d),
      .radr_d(twiddle_rsc_0_4_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_70_5_64_32_32_64_1_gen twiddle_rsc_0_29_i
      (
      .q(twiddle_rsc_0_29_q),
      .radr(twiddle_rsc_0_29_radr),
      .q_d(twiddle_rsc_0_29_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_71_5_64_32_32_64_1_gen twiddle_rsc_0_30_i
      (
      .q(twiddle_rsc_0_30_q),
      .radr(twiddle_rsc_0_30_radr),
      .q_d(twiddle_rsc_0_30_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_72_5_64_32_32_64_1_gen twiddle_rsc_0_31_i
      (
      .q(twiddle_rsc_0_31_q),
      .radr(twiddle_rsc_0_31_radr),
      .q_d(twiddle_rsc_0_31_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_core inPlaceNTT_DIF_core_inst (
      .clk(clk),
      .rst(rst),
      .vec_rsc_triosy_0_0_lz(vec_rsc_triosy_0_0_lz),
      .vec_rsc_triosy_0_1_lz(vec_rsc_triosy_0_1_lz),
      .vec_rsc_triosy_0_2_lz(vec_rsc_triosy_0_2_lz),
      .vec_rsc_triosy_0_3_lz(vec_rsc_triosy_0_3_lz),
      .vec_rsc_triosy_0_4_lz(vec_rsc_triosy_0_4_lz),
      .vec_rsc_triosy_0_5_lz(vec_rsc_triosy_0_5_lz),
      .vec_rsc_triosy_0_6_lz(vec_rsc_triosy_0_6_lz),
      .vec_rsc_triosy_0_7_lz(vec_rsc_triosy_0_7_lz),
      .vec_rsc_triosy_0_8_lz(vec_rsc_triosy_0_8_lz),
      .vec_rsc_triosy_0_9_lz(vec_rsc_triosy_0_9_lz),
      .vec_rsc_triosy_0_10_lz(vec_rsc_triosy_0_10_lz),
      .vec_rsc_triosy_0_11_lz(vec_rsc_triosy_0_11_lz),
      .vec_rsc_triosy_0_12_lz(vec_rsc_triosy_0_12_lz),
      .vec_rsc_triosy_0_13_lz(vec_rsc_triosy_0_13_lz),
      .vec_rsc_triosy_0_14_lz(vec_rsc_triosy_0_14_lz),
      .vec_rsc_triosy_0_15_lz(vec_rsc_triosy_0_15_lz),
      .vec_rsc_triosy_0_16_lz(vec_rsc_triosy_0_16_lz),
      .vec_rsc_triosy_0_17_lz(vec_rsc_triosy_0_17_lz),
      .vec_rsc_triosy_0_18_lz(vec_rsc_triosy_0_18_lz),
      .vec_rsc_triosy_0_19_lz(vec_rsc_triosy_0_19_lz),
      .vec_rsc_triosy_0_20_lz(vec_rsc_triosy_0_20_lz),
      .vec_rsc_triosy_0_21_lz(vec_rsc_triosy_0_21_lz),
      .vec_rsc_triosy_0_22_lz(vec_rsc_triosy_0_22_lz),
      .vec_rsc_triosy_0_23_lz(vec_rsc_triosy_0_23_lz),
      .vec_rsc_triosy_0_24_lz(vec_rsc_triosy_0_24_lz),
      .vec_rsc_triosy_0_25_lz(vec_rsc_triosy_0_25_lz),
      .vec_rsc_triosy_0_26_lz(vec_rsc_triosy_0_26_lz),
      .vec_rsc_triosy_0_27_lz(vec_rsc_triosy_0_27_lz),
      .vec_rsc_triosy_0_28_lz(vec_rsc_triosy_0_28_lz),
      .vec_rsc_triosy_0_29_lz(vec_rsc_triosy_0_29_lz),
      .vec_rsc_triosy_0_30_lz(vec_rsc_triosy_0_30_lz),
      .vec_rsc_triosy_0_31_lz(vec_rsc_triosy_0_31_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .twiddle_rsc_triosy_0_0_lz(twiddle_rsc_triosy_0_0_lz),
      .twiddle_rsc_triosy_0_1_lz(twiddle_rsc_triosy_0_1_lz),
      .twiddle_rsc_triosy_0_2_lz(twiddle_rsc_triosy_0_2_lz),
      .twiddle_rsc_triosy_0_3_lz(twiddle_rsc_triosy_0_3_lz),
      .twiddle_rsc_triosy_0_4_lz(twiddle_rsc_triosy_0_4_lz),
      .twiddle_rsc_triosy_0_5_lz(twiddle_rsc_triosy_0_5_lz),
      .twiddle_rsc_triosy_0_6_lz(twiddle_rsc_triosy_0_6_lz),
      .twiddle_rsc_triosy_0_7_lz(twiddle_rsc_triosy_0_7_lz),
      .twiddle_rsc_triosy_0_8_lz(twiddle_rsc_triosy_0_8_lz),
      .twiddle_rsc_triosy_0_9_lz(twiddle_rsc_triosy_0_9_lz),
      .twiddle_rsc_triosy_0_10_lz(twiddle_rsc_triosy_0_10_lz),
      .twiddle_rsc_triosy_0_11_lz(twiddle_rsc_triosy_0_11_lz),
      .twiddle_rsc_triosy_0_12_lz(twiddle_rsc_triosy_0_12_lz),
      .twiddle_rsc_triosy_0_13_lz(twiddle_rsc_triosy_0_13_lz),
      .twiddle_rsc_triosy_0_14_lz(twiddle_rsc_triosy_0_14_lz),
      .twiddle_rsc_triosy_0_15_lz(twiddle_rsc_triosy_0_15_lz),
      .twiddle_rsc_triosy_0_16_lz(twiddle_rsc_triosy_0_16_lz),
      .twiddle_rsc_triosy_0_17_lz(twiddle_rsc_triosy_0_17_lz),
      .twiddle_rsc_triosy_0_18_lz(twiddle_rsc_triosy_0_18_lz),
      .twiddle_rsc_triosy_0_19_lz(twiddle_rsc_triosy_0_19_lz),
      .twiddle_rsc_triosy_0_20_lz(twiddle_rsc_triosy_0_20_lz),
      .twiddle_rsc_triosy_0_21_lz(twiddle_rsc_triosy_0_21_lz),
      .twiddle_rsc_triosy_0_22_lz(twiddle_rsc_triosy_0_22_lz),
      .twiddle_rsc_triosy_0_23_lz(twiddle_rsc_triosy_0_23_lz),
      .twiddle_rsc_triosy_0_24_lz(twiddle_rsc_triosy_0_24_lz),
      .twiddle_rsc_triosy_0_25_lz(twiddle_rsc_triosy_0_25_lz),
      .twiddle_rsc_triosy_0_26_lz(twiddle_rsc_triosy_0_26_lz),
      .twiddle_rsc_triosy_0_27_lz(twiddle_rsc_triosy_0_27_lz),
      .twiddle_rsc_triosy_0_28_lz(twiddle_rsc_triosy_0_28_lz),
      .twiddle_rsc_triosy_0_29_lz(twiddle_rsc_triosy_0_29_lz),
      .twiddle_rsc_triosy_0_30_lz(twiddle_rsc_triosy_0_30_lz),
      .twiddle_rsc_triosy_0_31_lz(twiddle_rsc_triosy_0_31_lz),
      .vec_rsc_0_0_i_q_d(vec_rsc_0_0_i_q_d),
      .vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_1_i_q_d(vec_rsc_0_1_i_q_d),
      .vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_2_i_q_d(vec_rsc_0_2_i_q_d),
      .vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_3_i_q_d(vec_rsc_0_3_i_q_d),
      .vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_4_i_q_d(vec_rsc_0_4_i_q_d),
      .vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_5_i_q_d(vec_rsc_0_5_i_q_d),
      .vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_6_i_q_d(vec_rsc_0_6_i_q_d),
      .vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_7_i_q_d(vec_rsc_0_7_i_q_d),
      .vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_8_i_q_d(vec_rsc_0_8_i_q_d),
      .vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_9_i_q_d(vec_rsc_0_9_i_q_d),
      .vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_10_i_q_d(vec_rsc_0_10_i_q_d),
      .vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_11_i_q_d(vec_rsc_0_11_i_q_d),
      .vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_12_i_q_d(vec_rsc_0_12_i_q_d),
      .vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_13_i_q_d(vec_rsc_0_13_i_q_d),
      .vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_14_i_q_d(vec_rsc_0_14_i_q_d),
      .vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_15_i_q_d(vec_rsc_0_15_i_q_d),
      .vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_16_i_q_d(vec_rsc_0_16_i_q_d),
      .vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_17_i_q_d(vec_rsc_0_17_i_q_d),
      .vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_18_i_q_d(vec_rsc_0_18_i_q_d),
      .vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_19_i_q_d(vec_rsc_0_19_i_q_d),
      .vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_20_i_q_d(vec_rsc_0_20_i_q_d),
      .vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_21_i_q_d(vec_rsc_0_21_i_q_d),
      .vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_22_i_q_d(vec_rsc_0_22_i_q_d),
      .vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_23_i_q_d(vec_rsc_0_23_i_q_d),
      .vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_24_i_q_d(vec_rsc_0_24_i_q_d),
      .vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_25_i_q_d(vec_rsc_0_25_i_q_d),
      .vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_26_i_q_d(vec_rsc_0_26_i_q_d),
      .vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_27_i_q_d(vec_rsc_0_27_i_q_d),
      .vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_28_i_q_d(vec_rsc_0_28_i_q_d),
      .vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_29_i_q_d(vec_rsc_0_29_i_q_d),
      .vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_30_i_q_d(vec_rsc_0_30_i_q_d),
      .vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_31_i_q_d(vec_rsc_0_31_i_q_d),
      .vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_0_i_q_d(twiddle_rsc_0_0_i_q_d),
      .twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_1_i_q_d(twiddle_rsc_0_1_i_q_d),
      .twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_2_i_q_d(twiddle_rsc_0_2_i_q_d),
      .twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_3_i_q_d(twiddle_rsc_0_3_i_q_d),
      .twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_4_i_q_d(twiddle_rsc_0_4_i_q_d),
      .twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_5_i_q_d(twiddle_rsc_0_5_i_q_d),
      .twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_6_i_q_d(twiddle_rsc_0_6_i_q_d),
      .twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_7_i_q_d(twiddle_rsc_0_7_i_q_d),
      .twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_8_i_q_d(twiddle_rsc_0_8_i_q_d),
      .twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_9_i_q_d(twiddle_rsc_0_9_i_q_d),
      .twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_10_i_q_d(twiddle_rsc_0_10_i_q_d),
      .twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_11_i_q_d(twiddle_rsc_0_11_i_q_d),
      .twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_12_i_q_d(twiddle_rsc_0_12_i_q_d),
      .twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_13_i_q_d(twiddle_rsc_0_13_i_q_d),
      .twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_14_i_q_d(twiddle_rsc_0_14_i_q_d),
      .twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_15_i_q_d(twiddle_rsc_0_15_i_q_d),
      .twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_16_i_q_d(twiddle_rsc_0_16_i_q_d),
      .twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_17_i_q_d(twiddle_rsc_0_17_i_q_d),
      .twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_18_i_q_d(twiddle_rsc_0_18_i_q_d),
      .twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_19_i_q_d(twiddle_rsc_0_19_i_q_d),
      .twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_20_i_q_d(twiddle_rsc_0_20_i_q_d),
      .twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_21_i_q_d(twiddle_rsc_0_21_i_q_d),
      .twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_22_i_q_d(twiddle_rsc_0_22_i_q_d),
      .twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_23_i_q_d(twiddle_rsc_0_23_i_q_d),
      .twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_24_i_q_d(twiddle_rsc_0_24_i_q_d),
      .twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_25_i_q_d(twiddle_rsc_0_25_i_q_d),
      .twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_26_i_q_d(twiddle_rsc_0_26_i_q_d),
      .twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_27_i_q_d(twiddle_rsc_0_27_i_q_d),
      .twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_28_i_q_d(twiddle_rsc_0_28_i_q_d),
      .twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_29_i_q_d(twiddle_rsc_0_29_i_q_d),
      .twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_30_i_q_d(twiddle_rsc_0_30_i_q_d),
      .twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_31_i_q_d(twiddle_rsc_0_31_i_q_d),
      .twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_0_i_d_d_pff(vec_rsc_0_0_i_d_d_iff),
      .vec_rsc_0_0_i_radr_d_pff(vec_rsc_0_0_i_radr_d_iff),
      .vec_rsc_0_0_i_wadr_d_pff(vec_rsc_0_0_i_wadr_d_iff),
      .vec_rsc_0_0_i_we_d_pff(vec_rsc_0_0_i_we_d_iff),
      .vec_rsc_0_1_i_we_d_pff(vec_rsc_0_1_i_we_d_iff),
      .vec_rsc_0_2_i_we_d_pff(vec_rsc_0_2_i_we_d_iff),
      .vec_rsc_0_3_i_we_d_pff(vec_rsc_0_3_i_we_d_iff),
      .vec_rsc_0_4_i_we_d_pff(vec_rsc_0_4_i_we_d_iff),
      .vec_rsc_0_5_i_we_d_pff(vec_rsc_0_5_i_we_d_iff),
      .vec_rsc_0_6_i_we_d_pff(vec_rsc_0_6_i_we_d_iff),
      .vec_rsc_0_7_i_we_d_pff(vec_rsc_0_7_i_we_d_iff),
      .vec_rsc_0_8_i_we_d_pff(vec_rsc_0_8_i_we_d_iff),
      .vec_rsc_0_9_i_we_d_pff(vec_rsc_0_9_i_we_d_iff),
      .vec_rsc_0_10_i_we_d_pff(vec_rsc_0_10_i_we_d_iff),
      .vec_rsc_0_11_i_we_d_pff(vec_rsc_0_11_i_we_d_iff),
      .vec_rsc_0_12_i_we_d_pff(vec_rsc_0_12_i_we_d_iff),
      .vec_rsc_0_13_i_we_d_pff(vec_rsc_0_13_i_we_d_iff),
      .vec_rsc_0_14_i_we_d_pff(vec_rsc_0_14_i_we_d_iff),
      .vec_rsc_0_15_i_we_d_pff(vec_rsc_0_15_i_we_d_iff),
      .vec_rsc_0_16_i_we_d_pff(vec_rsc_0_16_i_we_d_iff),
      .vec_rsc_0_17_i_we_d_pff(vec_rsc_0_17_i_we_d_iff),
      .vec_rsc_0_18_i_we_d_pff(vec_rsc_0_18_i_we_d_iff),
      .vec_rsc_0_19_i_we_d_pff(vec_rsc_0_19_i_we_d_iff),
      .vec_rsc_0_20_i_we_d_pff(vec_rsc_0_20_i_we_d_iff),
      .vec_rsc_0_21_i_we_d_pff(vec_rsc_0_21_i_we_d_iff),
      .vec_rsc_0_22_i_we_d_pff(vec_rsc_0_22_i_we_d_iff),
      .vec_rsc_0_23_i_we_d_pff(vec_rsc_0_23_i_we_d_iff),
      .vec_rsc_0_24_i_we_d_pff(vec_rsc_0_24_i_we_d_iff),
      .vec_rsc_0_25_i_we_d_pff(vec_rsc_0_25_i_we_d_iff),
      .vec_rsc_0_26_i_we_d_pff(vec_rsc_0_26_i_we_d_iff),
      .vec_rsc_0_27_i_we_d_pff(vec_rsc_0_27_i_we_d_iff),
      .vec_rsc_0_28_i_we_d_pff(vec_rsc_0_28_i_we_d_iff),
      .vec_rsc_0_29_i_we_d_pff(vec_rsc_0_29_i_we_d_iff),
      .vec_rsc_0_30_i_we_d_pff(vec_rsc_0_30_i_we_d_iff),
      .vec_rsc_0_31_i_we_d_pff(vec_rsc_0_31_i_we_d_iff),
      .twiddle_rsc_0_0_i_radr_d_pff(twiddle_rsc_0_0_i_radr_d_iff),
      .twiddle_rsc_0_1_i_radr_d_pff(twiddle_rsc_0_1_i_radr_d_iff),
      .twiddle_rsc_0_2_i_radr_d_pff(twiddle_rsc_0_2_i_radr_d_iff),
      .twiddle_rsc_0_4_i_radr_d_pff(twiddle_rsc_0_4_i_radr_d_iff)
    );
endmodule



