
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.v 
module mgc_rem(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_b-1:0] z;  
   reg  [width_b-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  rem_s(a,b,z);
	else
          rem_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.v 
module mgc_div(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_a-1:0] z;  
   reg  [width_a-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  div_s(a,b,z);
	else
          div_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Wed Jun 30 21:42:36 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_9_64_512_512_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_9_64_512_512_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [8:0] adra;
  input [8:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_9_64_512_512_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_9_64_512_512_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [8:0] adra;
  input [8:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_9_64_512_512_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_9_64_512_512_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [8:0] adra;
  input [8:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_9_64_512_512_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_9_64_512_512_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [8:0] adra;
  input [8:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_9_64_512_512_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_9_64_512_512_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [8:0] adra;
  input [8:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_9_64_512_512_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_9_64_512_512_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [8:0] adra;
  input [8:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_9_64_512_512_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_9_64_512_512_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [8:0] adra;
  input [8:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_9_64_512_512_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_9_64_512_512_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [8:0] adra;
  input [8:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core_core_fsm (
  clk, rst, fsm_output, STAGE_LOOP_C_8_tr0, modExp_while_C_38_tr0, COMP_LOOP_C_1_tr0,
      COMP_LOOP_1_modExp_1_while_C_38_tr0, COMP_LOOP_C_62_tr0, COMP_LOOP_2_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_124_tr0, COMP_LOOP_3_modExp_1_while_C_38_tr0, COMP_LOOP_C_186_tr0,
      COMP_LOOP_4_modExp_1_while_C_38_tr0, COMP_LOOP_C_248_tr0, COMP_LOOP_5_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_310_tr0, COMP_LOOP_6_modExp_1_while_C_38_tr0, COMP_LOOP_C_372_tr0,
      COMP_LOOP_7_modExp_1_while_C_38_tr0, COMP_LOOP_C_434_tr0, COMP_LOOP_8_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_496_tr0, VEC_LOOP_C_0_tr0, STAGE_LOOP_C_9_tr0
);
  input clk;
  input rst;
  output [9:0] fsm_output;
  reg [9:0] fsm_output;
  input STAGE_LOOP_C_8_tr0;
  input modExp_while_C_38_tr0;
  input COMP_LOOP_C_1_tr0;
  input COMP_LOOP_1_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_62_tr0;
  input COMP_LOOP_2_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_124_tr0;
  input COMP_LOOP_3_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_186_tr0;
  input COMP_LOOP_4_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_248_tr0;
  input COMP_LOOP_5_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_310_tr0;
  input COMP_LOOP_6_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_372_tr0;
  input COMP_LOOP_7_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_434_tr0;
  input COMP_LOOP_8_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_496_tr0;
  input VEC_LOOP_C_0_tr0;
  input STAGE_LOOP_C_9_tr0;


  // FSM State Type Declaration for inPlaceNTT_DIT_core_core_fsm_1
  parameter
    main_C_0 = 10'd0,
    STAGE_LOOP_C_0 = 10'd1,
    STAGE_LOOP_C_1 = 10'd2,
    STAGE_LOOP_C_2 = 10'd3,
    STAGE_LOOP_C_3 = 10'd4,
    STAGE_LOOP_C_4 = 10'd5,
    STAGE_LOOP_C_5 = 10'd6,
    STAGE_LOOP_C_6 = 10'd7,
    STAGE_LOOP_C_7 = 10'd8,
    STAGE_LOOP_C_8 = 10'd9,
    modExp_while_C_0 = 10'd10,
    modExp_while_C_1 = 10'd11,
    modExp_while_C_2 = 10'd12,
    modExp_while_C_3 = 10'd13,
    modExp_while_C_4 = 10'd14,
    modExp_while_C_5 = 10'd15,
    modExp_while_C_6 = 10'd16,
    modExp_while_C_7 = 10'd17,
    modExp_while_C_8 = 10'd18,
    modExp_while_C_9 = 10'd19,
    modExp_while_C_10 = 10'd20,
    modExp_while_C_11 = 10'd21,
    modExp_while_C_12 = 10'd22,
    modExp_while_C_13 = 10'd23,
    modExp_while_C_14 = 10'd24,
    modExp_while_C_15 = 10'd25,
    modExp_while_C_16 = 10'd26,
    modExp_while_C_17 = 10'd27,
    modExp_while_C_18 = 10'd28,
    modExp_while_C_19 = 10'd29,
    modExp_while_C_20 = 10'd30,
    modExp_while_C_21 = 10'd31,
    modExp_while_C_22 = 10'd32,
    modExp_while_C_23 = 10'd33,
    modExp_while_C_24 = 10'd34,
    modExp_while_C_25 = 10'd35,
    modExp_while_C_26 = 10'd36,
    modExp_while_C_27 = 10'd37,
    modExp_while_C_28 = 10'd38,
    modExp_while_C_29 = 10'd39,
    modExp_while_C_30 = 10'd40,
    modExp_while_C_31 = 10'd41,
    modExp_while_C_32 = 10'd42,
    modExp_while_C_33 = 10'd43,
    modExp_while_C_34 = 10'd44,
    modExp_while_C_35 = 10'd45,
    modExp_while_C_36 = 10'd46,
    modExp_while_C_37 = 10'd47,
    modExp_while_C_38 = 10'd48,
    COMP_LOOP_C_0 = 10'd49,
    COMP_LOOP_C_1 = 10'd50,
    COMP_LOOP_1_modExp_1_while_C_0 = 10'd51,
    COMP_LOOP_1_modExp_1_while_C_1 = 10'd52,
    COMP_LOOP_1_modExp_1_while_C_2 = 10'd53,
    COMP_LOOP_1_modExp_1_while_C_3 = 10'd54,
    COMP_LOOP_1_modExp_1_while_C_4 = 10'd55,
    COMP_LOOP_1_modExp_1_while_C_5 = 10'd56,
    COMP_LOOP_1_modExp_1_while_C_6 = 10'd57,
    COMP_LOOP_1_modExp_1_while_C_7 = 10'd58,
    COMP_LOOP_1_modExp_1_while_C_8 = 10'd59,
    COMP_LOOP_1_modExp_1_while_C_9 = 10'd60,
    COMP_LOOP_1_modExp_1_while_C_10 = 10'd61,
    COMP_LOOP_1_modExp_1_while_C_11 = 10'd62,
    COMP_LOOP_1_modExp_1_while_C_12 = 10'd63,
    COMP_LOOP_1_modExp_1_while_C_13 = 10'd64,
    COMP_LOOP_1_modExp_1_while_C_14 = 10'd65,
    COMP_LOOP_1_modExp_1_while_C_15 = 10'd66,
    COMP_LOOP_1_modExp_1_while_C_16 = 10'd67,
    COMP_LOOP_1_modExp_1_while_C_17 = 10'd68,
    COMP_LOOP_1_modExp_1_while_C_18 = 10'd69,
    COMP_LOOP_1_modExp_1_while_C_19 = 10'd70,
    COMP_LOOP_1_modExp_1_while_C_20 = 10'd71,
    COMP_LOOP_1_modExp_1_while_C_21 = 10'd72,
    COMP_LOOP_1_modExp_1_while_C_22 = 10'd73,
    COMP_LOOP_1_modExp_1_while_C_23 = 10'd74,
    COMP_LOOP_1_modExp_1_while_C_24 = 10'd75,
    COMP_LOOP_1_modExp_1_while_C_25 = 10'd76,
    COMP_LOOP_1_modExp_1_while_C_26 = 10'd77,
    COMP_LOOP_1_modExp_1_while_C_27 = 10'd78,
    COMP_LOOP_1_modExp_1_while_C_28 = 10'd79,
    COMP_LOOP_1_modExp_1_while_C_29 = 10'd80,
    COMP_LOOP_1_modExp_1_while_C_30 = 10'd81,
    COMP_LOOP_1_modExp_1_while_C_31 = 10'd82,
    COMP_LOOP_1_modExp_1_while_C_32 = 10'd83,
    COMP_LOOP_1_modExp_1_while_C_33 = 10'd84,
    COMP_LOOP_1_modExp_1_while_C_34 = 10'd85,
    COMP_LOOP_1_modExp_1_while_C_35 = 10'd86,
    COMP_LOOP_1_modExp_1_while_C_36 = 10'd87,
    COMP_LOOP_1_modExp_1_while_C_37 = 10'd88,
    COMP_LOOP_1_modExp_1_while_C_38 = 10'd89,
    COMP_LOOP_C_2 = 10'd90,
    COMP_LOOP_C_3 = 10'd91,
    COMP_LOOP_C_4 = 10'd92,
    COMP_LOOP_C_5 = 10'd93,
    COMP_LOOP_C_6 = 10'd94,
    COMP_LOOP_C_7 = 10'd95,
    COMP_LOOP_C_8 = 10'd96,
    COMP_LOOP_C_9 = 10'd97,
    COMP_LOOP_C_10 = 10'd98,
    COMP_LOOP_C_11 = 10'd99,
    COMP_LOOP_C_12 = 10'd100,
    COMP_LOOP_C_13 = 10'd101,
    COMP_LOOP_C_14 = 10'd102,
    COMP_LOOP_C_15 = 10'd103,
    COMP_LOOP_C_16 = 10'd104,
    COMP_LOOP_C_17 = 10'd105,
    COMP_LOOP_C_18 = 10'd106,
    COMP_LOOP_C_19 = 10'd107,
    COMP_LOOP_C_20 = 10'd108,
    COMP_LOOP_C_21 = 10'd109,
    COMP_LOOP_C_22 = 10'd110,
    COMP_LOOP_C_23 = 10'd111,
    COMP_LOOP_C_24 = 10'd112,
    COMP_LOOP_C_25 = 10'd113,
    COMP_LOOP_C_26 = 10'd114,
    COMP_LOOP_C_27 = 10'd115,
    COMP_LOOP_C_28 = 10'd116,
    COMP_LOOP_C_29 = 10'd117,
    COMP_LOOP_C_30 = 10'd118,
    COMP_LOOP_C_31 = 10'd119,
    COMP_LOOP_C_32 = 10'd120,
    COMP_LOOP_C_33 = 10'd121,
    COMP_LOOP_C_34 = 10'd122,
    COMP_LOOP_C_35 = 10'd123,
    COMP_LOOP_C_36 = 10'd124,
    COMP_LOOP_C_37 = 10'd125,
    COMP_LOOP_C_38 = 10'd126,
    COMP_LOOP_C_39 = 10'd127,
    COMP_LOOP_C_40 = 10'd128,
    COMP_LOOP_C_41 = 10'd129,
    COMP_LOOP_C_42 = 10'd130,
    COMP_LOOP_C_43 = 10'd131,
    COMP_LOOP_C_44 = 10'd132,
    COMP_LOOP_C_45 = 10'd133,
    COMP_LOOP_C_46 = 10'd134,
    COMP_LOOP_C_47 = 10'd135,
    COMP_LOOP_C_48 = 10'd136,
    COMP_LOOP_C_49 = 10'd137,
    COMP_LOOP_C_50 = 10'd138,
    COMP_LOOP_C_51 = 10'd139,
    COMP_LOOP_C_52 = 10'd140,
    COMP_LOOP_C_53 = 10'd141,
    COMP_LOOP_C_54 = 10'd142,
    COMP_LOOP_C_55 = 10'd143,
    COMP_LOOP_C_56 = 10'd144,
    COMP_LOOP_C_57 = 10'd145,
    COMP_LOOP_C_58 = 10'd146,
    COMP_LOOP_C_59 = 10'd147,
    COMP_LOOP_C_60 = 10'd148,
    COMP_LOOP_C_61 = 10'd149,
    COMP_LOOP_C_62 = 10'd150,
    COMP_LOOP_C_63 = 10'd151,
    COMP_LOOP_2_modExp_1_while_C_0 = 10'd152,
    COMP_LOOP_2_modExp_1_while_C_1 = 10'd153,
    COMP_LOOP_2_modExp_1_while_C_2 = 10'd154,
    COMP_LOOP_2_modExp_1_while_C_3 = 10'd155,
    COMP_LOOP_2_modExp_1_while_C_4 = 10'd156,
    COMP_LOOP_2_modExp_1_while_C_5 = 10'd157,
    COMP_LOOP_2_modExp_1_while_C_6 = 10'd158,
    COMP_LOOP_2_modExp_1_while_C_7 = 10'd159,
    COMP_LOOP_2_modExp_1_while_C_8 = 10'd160,
    COMP_LOOP_2_modExp_1_while_C_9 = 10'd161,
    COMP_LOOP_2_modExp_1_while_C_10 = 10'd162,
    COMP_LOOP_2_modExp_1_while_C_11 = 10'd163,
    COMP_LOOP_2_modExp_1_while_C_12 = 10'd164,
    COMP_LOOP_2_modExp_1_while_C_13 = 10'd165,
    COMP_LOOP_2_modExp_1_while_C_14 = 10'd166,
    COMP_LOOP_2_modExp_1_while_C_15 = 10'd167,
    COMP_LOOP_2_modExp_1_while_C_16 = 10'd168,
    COMP_LOOP_2_modExp_1_while_C_17 = 10'd169,
    COMP_LOOP_2_modExp_1_while_C_18 = 10'd170,
    COMP_LOOP_2_modExp_1_while_C_19 = 10'd171,
    COMP_LOOP_2_modExp_1_while_C_20 = 10'd172,
    COMP_LOOP_2_modExp_1_while_C_21 = 10'd173,
    COMP_LOOP_2_modExp_1_while_C_22 = 10'd174,
    COMP_LOOP_2_modExp_1_while_C_23 = 10'd175,
    COMP_LOOP_2_modExp_1_while_C_24 = 10'd176,
    COMP_LOOP_2_modExp_1_while_C_25 = 10'd177,
    COMP_LOOP_2_modExp_1_while_C_26 = 10'd178,
    COMP_LOOP_2_modExp_1_while_C_27 = 10'd179,
    COMP_LOOP_2_modExp_1_while_C_28 = 10'd180,
    COMP_LOOP_2_modExp_1_while_C_29 = 10'd181,
    COMP_LOOP_2_modExp_1_while_C_30 = 10'd182,
    COMP_LOOP_2_modExp_1_while_C_31 = 10'd183,
    COMP_LOOP_2_modExp_1_while_C_32 = 10'd184,
    COMP_LOOP_2_modExp_1_while_C_33 = 10'd185,
    COMP_LOOP_2_modExp_1_while_C_34 = 10'd186,
    COMP_LOOP_2_modExp_1_while_C_35 = 10'd187,
    COMP_LOOP_2_modExp_1_while_C_36 = 10'd188,
    COMP_LOOP_2_modExp_1_while_C_37 = 10'd189,
    COMP_LOOP_2_modExp_1_while_C_38 = 10'd190,
    COMP_LOOP_C_64 = 10'd191,
    COMP_LOOP_C_65 = 10'd192,
    COMP_LOOP_C_66 = 10'd193,
    COMP_LOOP_C_67 = 10'd194,
    COMP_LOOP_C_68 = 10'd195,
    COMP_LOOP_C_69 = 10'd196,
    COMP_LOOP_C_70 = 10'd197,
    COMP_LOOP_C_71 = 10'd198,
    COMP_LOOP_C_72 = 10'd199,
    COMP_LOOP_C_73 = 10'd200,
    COMP_LOOP_C_74 = 10'd201,
    COMP_LOOP_C_75 = 10'd202,
    COMP_LOOP_C_76 = 10'd203,
    COMP_LOOP_C_77 = 10'd204,
    COMP_LOOP_C_78 = 10'd205,
    COMP_LOOP_C_79 = 10'd206,
    COMP_LOOP_C_80 = 10'd207,
    COMP_LOOP_C_81 = 10'd208,
    COMP_LOOP_C_82 = 10'd209,
    COMP_LOOP_C_83 = 10'd210,
    COMP_LOOP_C_84 = 10'd211,
    COMP_LOOP_C_85 = 10'd212,
    COMP_LOOP_C_86 = 10'd213,
    COMP_LOOP_C_87 = 10'd214,
    COMP_LOOP_C_88 = 10'd215,
    COMP_LOOP_C_89 = 10'd216,
    COMP_LOOP_C_90 = 10'd217,
    COMP_LOOP_C_91 = 10'd218,
    COMP_LOOP_C_92 = 10'd219,
    COMP_LOOP_C_93 = 10'd220,
    COMP_LOOP_C_94 = 10'd221,
    COMP_LOOP_C_95 = 10'd222,
    COMP_LOOP_C_96 = 10'd223,
    COMP_LOOP_C_97 = 10'd224,
    COMP_LOOP_C_98 = 10'd225,
    COMP_LOOP_C_99 = 10'd226,
    COMP_LOOP_C_100 = 10'd227,
    COMP_LOOP_C_101 = 10'd228,
    COMP_LOOP_C_102 = 10'd229,
    COMP_LOOP_C_103 = 10'd230,
    COMP_LOOP_C_104 = 10'd231,
    COMP_LOOP_C_105 = 10'd232,
    COMP_LOOP_C_106 = 10'd233,
    COMP_LOOP_C_107 = 10'd234,
    COMP_LOOP_C_108 = 10'd235,
    COMP_LOOP_C_109 = 10'd236,
    COMP_LOOP_C_110 = 10'd237,
    COMP_LOOP_C_111 = 10'd238,
    COMP_LOOP_C_112 = 10'd239,
    COMP_LOOP_C_113 = 10'd240,
    COMP_LOOP_C_114 = 10'd241,
    COMP_LOOP_C_115 = 10'd242,
    COMP_LOOP_C_116 = 10'd243,
    COMP_LOOP_C_117 = 10'd244,
    COMP_LOOP_C_118 = 10'd245,
    COMP_LOOP_C_119 = 10'd246,
    COMP_LOOP_C_120 = 10'd247,
    COMP_LOOP_C_121 = 10'd248,
    COMP_LOOP_C_122 = 10'd249,
    COMP_LOOP_C_123 = 10'd250,
    COMP_LOOP_C_124 = 10'd251,
    COMP_LOOP_C_125 = 10'd252,
    COMP_LOOP_3_modExp_1_while_C_0 = 10'd253,
    COMP_LOOP_3_modExp_1_while_C_1 = 10'd254,
    COMP_LOOP_3_modExp_1_while_C_2 = 10'd255,
    COMP_LOOP_3_modExp_1_while_C_3 = 10'd256,
    COMP_LOOP_3_modExp_1_while_C_4 = 10'd257,
    COMP_LOOP_3_modExp_1_while_C_5 = 10'd258,
    COMP_LOOP_3_modExp_1_while_C_6 = 10'd259,
    COMP_LOOP_3_modExp_1_while_C_7 = 10'd260,
    COMP_LOOP_3_modExp_1_while_C_8 = 10'd261,
    COMP_LOOP_3_modExp_1_while_C_9 = 10'd262,
    COMP_LOOP_3_modExp_1_while_C_10 = 10'd263,
    COMP_LOOP_3_modExp_1_while_C_11 = 10'd264,
    COMP_LOOP_3_modExp_1_while_C_12 = 10'd265,
    COMP_LOOP_3_modExp_1_while_C_13 = 10'd266,
    COMP_LOOP_3_modExp_1_while_C_14 = 10'd267,
    COMP_LOOP_3_modExp_1_while_C_15 = 10'd268,
    COMP_LOOP_3_modExp_1_while_C_16 = 10'd269,
    COMP_LOOP_3_modExp_1_while_C_17 = 10'd270,
    COMP_LOOP_3_modExp_1_while_C_18 = 10'd271,
    COMP_LOOP_3_modExp_1_while_C_19 = 10'd272,
    COMP_LOOP_3_modExp_1_while_C_20 = 10'd273,
    COMP_LOOP_3_modExp_1_while_C_21 = 10'd274,
    COMP_LOOP_3_modExp_1_while_C_22 = 10'd275,
    COMP_LOOP_3_modExp_1_while_C_23 = 10'd276,
    COMP_LOOP_3_modExp_1_while_C_24 = 10'd277,
    COMP_LOOP_3_modExp_1_while_C_25 = 10'd278,
    COMP_LOOP_3_modExp_1_while_C_26 = 10'd279,
    COMP_LOOP_3_modExp_1_while_C_27 = 10'd280,
    COMP_LOOP_3_modExp_1_while_C_28 = 10'd281,
    COMP_LOOP_3_modExp_1_while_C_29 = 10'd282,
    COMP_LOOP_3_modExp_1_while_C_30 = 10'd283,
    COMP_LOOP_3_modExp_1_while_C_31 = 10'd284,
    COMP_LOOP_3_modExp_1_while_C_32 = 10'd285,
    COMP_LOOP_3_modExp_1_while_C_33 = 10'd286,
    COMP_LOOP_3_modExp_1_while_C_34 = 10'd287,
    COMP_LOOP_3_modExp_1_while_C_35 = 10'd288,
    COMP_LOOP_3_modExp_1_while_C_36 = 10'd289,
    COMP_LOOP_3_modExp_1_while_C_37 = 10'd290,
    COMP_LOOP_3_modExp_1_while_C_38 = 10'd291,
    COMP_LOOP_C_126 = 10'd292,
    COMP_LOOP_C_127 = 10'd293,
    COMP_LOOP_C_128 = 10'd294,
    COMP_LOOP_C_129 = 10'd295,
    COMP_LOOP_C_130 = 10'd296,
    COMP_LOOP_C_131 = 10'd297,
    COMP_LOOP_C_132 = 10'd298,
    COMP_LOOP_C_133 = 10'd299,
    COMP_LOOP_C_134 = 10'd300,
    COMP_LOOP_C_135 = 10'd301,
    COMP_LOOP_C_136 = 10'd302,
    COMP_LOOP_C_137 = 10'd303,
    COMP_LOOP_C_138 = 10'd304,
    COMP_LOOP_C_139 = 10'd305,
    COMP_LOOP_C_140 = 10'd306,
    COMP_LOOP_C_141 = 10'd307,
    COMP_LOOP_C_142 = 10'd308,
    COMP_LOOP_C_143 = 10'd309,
    COMP_LOOP_C_144 = 10'd310,
    COMP_LOOP_C_145 = 10'd311,
    COMP_LOOP_C_146 = 10'd312,
    COMP_LOOP_C_147 = 10'd313,
    COMP_LOOP_C_148 = 10'd314,
    COMP_LOOP_C_149 = 10'd315,
    COMP_LOOP_C_150 = 10'd316,
    COMP_LOOP_C_151 = 10'd317,
    COMP_LOOP_C_152 = 10'd318,
    COMP_LOOP_C_153 = 10'd319,
    COMP_LOOP_C_154 = 10'd320,
    COMP_LOOP_C_155 = 10'd321,
    COMP_LOOP_C_156 = 10'd322,
    COMP_LOOP_C_157 = 10'd323,
    COMP_LOOP_C_158 = 10'd324,
    COMP_LOOP_C_159 = 10'd325,
    COMP_LOOP_C_160 = 10'd326,
    COMP_LOOP_C_161 = 10'd327,
    COMP_LOOP_C_162 = 10'd328,
    COMP_LOOP_C_163 = 10'd329,
    COMP_LOOP_C_164 = 10'd330,
    COMP_LOOP_C_165 = 10'd331,
    COMP_LOOP_C_166 = 10'd332,
    COMP_LOOP_C_167 = 10'd333,
    COMP_LOOP_C_168 = 10'd334,
    COMP_LOOP_C_169 = 10'd335,
    COMP_LOOP_C_170 = 10'd336,
    COMP_LOOP_C_171 = 10'd337,
    COMP_LOOP_C_172 = 10'd338,
    COMP_LOOP_C_173 = 10'd339,
    COMP_LOOP_C_174 = 10'd340,
    COMP_LOOP_C_175 = 10'd341,
    COMP_LOOP_C_176 = 10'd342,
    COMP_LOOP_C_177 = 10'd343,
    COMP_LOOP_C_178 = 10'd344,
    COMP_LOOP_C_179 = 10'd345,
    COMP_LOOP_C_180 = 10'd346,
    COMP_LOOP_C_181 = 10'd347,
    COMP_LOOP_C_182 = 10'd348,
    COMP_LOOP_C_183 = 10'd349,
    COMP_LOOP_C_184 = 10'd350,
    COMP_LOOP_C_185 = 10'd351,
    COMP_LOOP_C_186 = 10'd352,
    COMP_LOOP_C_187 = 10'd353,
    COMP_LOOP_4_modExp_1_while_C_0 = 10'd354,
    COMP_LOOP_4_modExp_1_while_C_1 = 10'd355,
    COMP_LOOP_4_modExp_1_while_C_2 = 10'd356,
    COMP_LOOP_4_modExp_1_while_C_3 = 10'd357,
    COMP_LOOP_4_modExp_1_while_C_4 = 10'd358,
    COMP_LOOP_4_modExp_1_while_C_5 = 10'd359,
    COMP_LOOP_4_modExp_1_while_C_6 = 10'd360,
    COMP_LOOP_4_modExp_1_while_C_7 = 10'd361,
    COMP_LOOP_4_modExp_1_while_C_8 = 10'd362,
    COMP_LOOP_4_modExp_1_while_C_9 = 10'd363,
    COMP_LOOP_4_modExp_1_while_C_10 = 10'd364,
    COMP_LOOP_4_modExp_1_while_C_11 = 10'd365,
    COMP_LOOP_4_modExp_1_while_C_12 = 10'd366,
    COMP_LOOP_4_modExp_1_while_C_13 = 10'd367,
    COMP_LOOP_4_modExp_1_while_C_14 = 10'd368,
    COMP_LOOP_4_modExp_1_while_C_15 = 10'd369,
    COMP_LOOP_4_modExp_1_while_C_16 = 10'd370,
    COMP_LOOP_4_modExp_1_while_C_17 = 10'd371,
    COMP_LOOP_4_modExp_1_while_C_18 = 10'd372,
    COMP_LOOP_4_modExp_1_while_C_19 = 10'd373,
    COMP_LOOP_4_modExp_1_while_C_20 = 10'd374,
    COMP_LOOP_4_modExp_1_while_C_21 = 10'd375,
    COMP_LOOP_4_modExp_1_while_C_22 = 10'd376,
    COMP_LOOP_4_modExp_1_while_C_23 = 10'd377,
    COMP_LOOP_4_modExp_1_while_C_24 = 10'd378,
    COMP_LOOP_4_modExp_1_while_C_25 = 10'd379,
    COMP_LOOP_4_modExp_1_while_C_26 = 10'd380,
    COMP_LOOP_4_modExp_1_while_C_27 = 10'd381,
    COMP_LOOP_4_modExp_1_while_C_28 = 10'd382,
    COMP_LOOP_4_modExp_1_while_C_29 = 10'd383,
    COMP_LOOP_4_modExp_1_while_C_30 = 10'd384,
    COMP_LOOP_4_modExp_1_while_C_31 = 10'd385,
    COMP_LOOP_4_modExp_1_while_C_32 = 10'd386,
    COMP_LOOP_4_modExp_1_while_C_33 = 10'd387,
    COMP_LOOP_4_modExp_1_while_C_34 = 10'd388,
    COMP_LOOP_4_modExp_1_while_C_35 = 10'd389,
    COMP_LOOP_4_modExp_1_while_C_36 = 10'd390,
    COMP_LOOP_4_modExp_1_while_C_37 = 10'd391,
    COMP_LOOP_4_modExp_1_while_C_38 = 10'd392,
    COMP_LOOP_C_188 = 10'd393,
    COMP_LOOP_C_189 = 10'd394,
    COMP_LOOP_C_190 = 10'd395,
    COMP_LOOP_C_191 = 10'd396,
    COMP_LOOP_C_192 = 10'd397,
    COMP_LOOP_C_193 = 10'd398,
    COMP_LOOP_C_194 = 10'd399,
    COMP_LOOP_C_195 = 10'd400,
    COMP_LOOP_C_196 = 10'd401,
    COMP_LOOP_C_197 = 10'd402,
    COMP_LOOP_C_198 = 10'd403,
    COMP_LOOP_C_199 = 10'd404,
    COMP_LOOP_C_200 = 10'd405,
    COMP_LOOP_C_201 = 10'd406,
    COMP_LOOP_C_202 = 10'd407,
    COMP_LOOP_C_203 = 10'd408,
    COMP_LOOP_C_204 = 10'd409,
    COMP_LOOP_C_205 = 10'd410,
    COMP_LOOP_C_206 = 10'd411,
    COMP_LOOP_C_207 = 10'd412,
    COMP_LOOP_C_208 = 10'd413,
    COMP_LOOP_C_209 = 10'd414,
    COMP_LOOP_C_210 = 10'd415,
    COMP_LOOP_C_211 = 10'd416,
    COMP_LOOP_C_212 = 10'd417,
    COMP_LOOP_C_213 = 10'd418,
    COMP_LOOP_C_214 = 10'd419,
    COMP_LOOP_C_215 = 10'd420,
    COMP_LOOP_C_216 = 10'd421,
    COMP_LOOP_C_217 = 10'd422,
    COMP_LOOP_C_218 = 10'd423,
    COMP_LOOP_C_219 = 10'd424,
    COMP_LOOP_C_220 = 10'd425,
    COMP_LOOP_C_221 = 10'd426,
    COMP_LOOP_C_222 = 10'd427,
    COMP_LOOP_C_223 = 10'd428,
    COMP_LOOP_C_224 = 10'd429,
    COMP_LOOP_C_225 = 10'd430,
    COMP_LOOP_C_226 = 10'd431,
    COMP_LOOP_C_227 = 10'd432,
    COMP_LOOP_C_228 = 10'd433,
    COMP_LOOP_C_229 = 10'd434,
    COMP_LOOP_C_230 = 10'd435,
    COMP_LOOP_C_231 = 10'd436,
    COMP_LOOP_C_232 = 10'd437,
    COMP_LOOP_C_233 = 10'd438,
    COMP_LOOP_C_234 = 10'd439,
    COMP_LOOP_C_235 = 10'd440,
    COMP_LOOP_C_236 = 10'd441,
    COMP_LOOP_C_237 = 10'd442,
    COMP_LOOP_C_238 = 10'd443,
    COMP_LOOP_C_239 = 10'd444,
    COMP_LOOP_C_240 = 10'd445,
    COMP_LOOP_C_241 = 10'd446,
    COMP_LOOP_C_242 = 10'd447,
    COMP_LOOP_C_243 = 10'd448,
    COMP_LOOP_C_244 = 10'd449,
    COMP_LOOP_C_245 = 10'd450,
    COMP_LOOP_C_246 = 10'd451,
    COMP_LOOP_C_247 = 10'd452,
    COMP_LOOP_C_248 = 10'd453,
    COMP_LOOP_C_249 = 10'd454,
    COMP_LOOP_5_modExp_1_while_C_0 = 10'd455,
    COMP_LOOP_5_modExp_1_while_C_1 = 10'd456,
    COMP_LOOP_5_modExp_1_while_C_2 = 10'd457,
    COMP_LOOP_5_modExp_1_while_C_3 = 10'd458,
    COMP_LOOP_5_modExp_1_while_C_4 = 10'd459,
    COMP_LOOP_5_modExp_1_while_C_5 = 10'd460,
    COMP_LOOP_5_modExp_1_while_C_6 = 10'd461,
    COMP_LOOP_5_modExp_1_while_C_7 = 10'd462,
    COMP_LOOP_5_modExp_1_while_C_8 = 10'd463,
    COMP_LOOP_5_modExp_1_while_C_9 = 10'd464,
    COMP_LOOP_5_modExp_1_while_C_10 = 10'd465,
    COMP_LOOP_5_modExp_1_while_C_11 = 10'd466,
    COMP_LOOP_5_modExp_1_while_C_12 = 10'd467,
    COMP_LOOP_5_modExp_1_while_C_13 = 10'd468,
    COMP_LOOP_5_modExp_1_while_C_14 = 10'd469,
    COMP_LOOP_5_modExp_1_while_C_15 = 10'd470,
    COMP_LOOP_5_modExp_1_while_C_16 = 10'd471,
    COMP_LOOP_5_modExp_1_while_C_17 = 10'd472,
    COMP_LOOP_5_modExp_1_while_C_18 = 10'd473,
    COMP_LOOP_5_modExp_1_while_C_19 = 10'd474,
    COMP_LOOP_5_modExp_1_while_C_20 = 10'd475,
    COMP_LOOP_5_modExp_1_while_C_21 = 10'd476,
    COMP_LOOP_5_modExp_1_while_C_22 = 10'd477,
    COMP_LOOP_5_modExp_1_while_C_23 = 10'd478,
    COMP_LOOP_5_modExp_1_while_C_24 = 10'd479,
    COMP_LOOP_5_modExp_1_while_C_25 = 10'd480,
    COMP_LOOP_5_modExp_1_while_C_26 = 10'd481,
    COMP_LOOP_5_modExp_1_while_C_27 = 10'd482,
    COMP_LOOP_5_modExp_1_while_C_28 = 10'd483,
    COMP_LOOP_5_modExp_1_while_C_29 = 10'd484,
    COMP_LOOP_5_modExp_1_while_C_30 = 10'd485,
    COMP_LOOP_5_modExp_1_while_C_31 = 10'd486,
    COMP_LOOP_5_modExp_1_while_C_32 = 10'd487,
    COMP_LOOP_5_modExp_1_while_C_33 = 10'd488,
    COMP_LOOP_5_modExp_1_while_C_34 = 10'd489,
    COMP_LOOP_5_modExp_1_while_C_35 = 10'd490,
    COMP_LOOP_5_modExp_1_while_C_36 = 10'd491,
    COMP_LOOP_5_modExp_1_while_C_37 = 10'd492,
    COMP_LOOP_5_modExp_1_while_C_38 = 10'd493,
    COMP_LOOP_C_250 = 10'd494,
    COMP_LOOP_C_251 = 10'd495,
    COMP_LOOP_C_252 = 10'd496,
    COMP_LOOP_C_253 = 10'd497,
    COMP_LOOP_C_254 = 10'd498,
    COMP_LOOP_C_255 = 10'd499,
    COMP_LOOP_C_256 = 10'd500,
    COMP_LOOP_C_257 = 10'd501,
    COMP_LOOP_C_258 = 10'd502,
    COMP_LOOP_C_259 = 10'd503,
    COMP_LOOP_C_260 = 10'd504,
    COMP_LOOP_C_261 = 10'd505,
    COMP_LOOP_C_262 = 10'd506,
    COMP_LOOP_C_263 = 10'd507,
    COMP_LOOP_C_264 = 10'd508,
    COMP_LOOP_C_265 = 10'd509,
    COMP_LOOP_C_266 = 10'd510,
    COMP_LOOP_C_267 = 10'd511,
    COMP_LOOP_C_268 = 10'd512,
    COMP_LOOP_C_269 = 10'd513,
    COMP_LOOP_C_270 = 10'd514,
    COMP_LOOP_C_271 = 10'd515,
    COMP_LOOP_C_272 = 10'd516,
    COMP_LOOP_C_273 = 10'd517,
    COMP_LOOP_C_274 = 10'd518,
    COMP_LOOP_C_275 = 10'd519,
    COMP_LOOP_C_276 = 10'd520,
    COMP_LOOP_C_277 = 10'd521,
    COMP_LOOP_C_278 = 10'd522,
    COMP_LOOP_C_279 = 10'd523,
    COMP_LOOP_C_280 = 10'd524,
    COMP_LOOP_C_281 = 10'd525,
    COMP_LOOP_C_282 = 10'd526,
    COMP_LOOP_C_283 = 10'd527,
    COMP_LOOP_C_284 = 10'd528,
    COMP_LOOP_C_285 = 10'd529,
    COMP_LOOP_C_286 = 10'd530,
    COMP_LOOP_C_287 = 10'd531,
    COMP_LOOP_C_288 = 10'd532,
    COMP_LOOP_C_289 = 10'd533,
    COMP_LOOP_C_290 = 10'd534,
    COMP_LOOP_C_291 = 10'd535,
    COMP_LOOP_C_292 = 10'd536,
    COMP_LOOP_C_293 = 10'd537,
    COMP_LOOP_C_294 = 10'd538,
    COMP_LOOP_C_295 = 10'd539,
    COMP_LOOP_C_296 = 10'd540,
    COMP_LOOP_C_297 = 10'd541,
    COMP_LOOP_C_298 = 10'd542,
    COMP_LOOP_C_299 = 10'd543,
    COMP_LOOP_C_300 = 10'd544,
    COMP_LOOP_C_301 = 10'd545,
    COMP_LOOP_C_302 = 10'd546,
    COMP_LOOP_C_303 = 10'd547,
    COMP_LOOP_C_304 = 10'd548,
    COMP_LOOP_C_305 = 10'd549,
    COMP_LOOP_C_306 = 10'd550,
    COMP_LOOP_C_307 = 10'd551,
    COMP_LOOP_C_308 = 10'd552,
    COMP_LOOP_C_309 = 10'd553,
    COMP_LOOP_C_310 = 10'd554,
    COMP_LOOP_C_311 = 10'd555,
    COMP_LOOP_6_modExp_1_while_C_0 = 10'd556,
    COMP_LOOP_6_modExp_1_while_C_1 = 10'd557,
    COMP_LOOP_6_modExp_1_while_C_2 = 10'd558,
    COMP_LOOP_6_modExp_1_while_C_3 = 10'd559,
    COMP_LOOP_6_modExp_1_while_C_4 = 10'd560,
    COMP_LOOP_6_modExp_1_while_C_5 = 10'd561,
    COMP_LOOP_6_modExp_1_while_C_6 = 10'd562,
    COMP_LOOP_6_modExp_1_while_C_7 = 10'd563,
    COMP_LOOP_6_modExp_1_while_C_8 = 10'd564,
    COMP_LOOP_6_modExp_1_while_C_9 = 10'd565,
    COMP_LOOP_6_modExp_1_while_C_10 = 10'd566,
    COMP_LOOP_6_modExp_1_while_C_11 = 10'd567,
    COMP_LOOP_6_modExp_1_while_C_12 = 10'd568,
    COMP_LOOP_6_modExp_1_while_C_13 = 10'd569,
    COMP_LOOP_6_modExp_1_while_C_14 = 10'd570,
    COMP_LOOP_6_modExp_1_while_C_15 = 10'd571,
    COMP_LOOP_6_modExp_1_while_C_16 = 10'd572,
    COMP_LOOP_6_modExp_1_while_C_17 = 10'd573,
    COMP_LOOP_6_modExp_1_while_C_18 = 10'd574,
    COMP_LOOP_6_modExp_1_while_C_19 = 10'd575,
    COMP_LOOP_6_modExp_1_while_C_20 = 10'd576,
    COMP_LOOP_6_modExp_1_while_C_21 = 10'd577,
    COMP_LOOP_6_modExp_1_while_C_22 = 10'd578,
    COMP_LOOP_6_modExp_1_while_C_23 = 10'd579,
    COMP_LOOP_6_modExp_1_while_C_24 = 10'd580,
    COMP_LOOP_6_modExp_1_while_C_25 = 10'd581,
    COMP_LOOP_6_modExp_1_while_C_26 = 10'd582,
    COMP_LOOP_6_modExp_1_while_C_27 = 10'd583,
    COMP_LOOP_6_modExp_1_while_C_28 = 10'd584,
    COMP_LOOP_6_modExp_1_while_C_29 = 10'd585,
    COMP_LOOP_6_modExp_1_while_C_30 = 10'd586,
    COMP_LOOP_6_modExp_1_while_C_31 = 10'd587,
    COMP_LOOP_6_modExp_1_while_C_32 = 10'd588,
    COMP_LOOP_6_modExp_1_while_C_33 = 10'd589,
    COMP_LOOP_6_modExp_1_while_C_34 = 10'd590,
    COMP_LOOP_6_modExp_1_while_C_35 = 10'd591,
    COMP_LOOP_6_modExp_1_while_C_36 = 10'd592,
    COMP_LOOP_6_modExp_1_while_C_37 = 10'd593,
    COMP_LOOP_6_modExp_1_while_C_38 = 10'd594,
    COMP_LOOP_C_312 = 10'd595,
    COMP_LOOP_C_313 = 10'd596,
    COMP_LOOP_C_314 = 10'd597,
    COMP_LOOP_C_315 = 10'd598,
    COMP_LOOP_C_316 = 10'd599,
    COMP_LOOP_C_317 = 10'd600,
    COMP_LOOP_C_318 = 10'd601,
    COMP_LOOP_C_319 = 10'd602,
    COMP_LOOP_C_320 = 10'd603,
    COMP_LOOP_C_321 = 10'd604,
    COMP_LOOP_C_322 = 10'd605,
    COMP_LOOP_C_323 = 10'd606,
    COMP_LOOP_C_324 = 10'd607,
    COMP_LOOP_C_325 = 10'd608,
    COMP_LOOP_C_326 = 10'd609,
    COMP_LOOP_C_327 = 10'd610,
    COMP_LOOP_C_328 = 10'd611,
    COMP_LOOP_C_329 = 10'd612,
    COMP_LOOP_C_330 = 10'd613,
    COMP_LOOP_C_331 = 10'd614,
    COMP_LOOP_C_332 = 10'd615,
    COMP_LOOP_C_333 = 10'd616,
    COMP_LOOP_C_334 = 10'd617,
    COMP_LOOP_C_335 = 10'd618,
    COMP_LOOP_C_336 = 10'd619,
    COMP_LOOP_C_337 = 10'd620,
    COMP_LOOP_C_338 = 10'd621,
    COMP_LOOP_C_339 = 10'd622,
    COMP_LOOP_C_340 = 10'd623,
    COMP_LOOP_C_341 = 10'd624,
    COMP_LOOP_C_342 = 10'd625,
    COMP_LOOP_C_343 = 10'd626,
    COMP_LOOP_C_344 = 10'd627,
    COMP_LOOP_C_345 = 10'd628,
    COMP_LOOP_C_346 = 10'd629,
    COMP_LOOP_C_347 = 10'd630,
    COMP_LOOP_C_348 = 10'd631,
    COMP_LOOP_C_349 = 10'd632,
    COMP_LOOP_C_350 = 10'd633,
    COMP_LOOP_C_351 = 10'd634,
    COMP_LOOP_C_352 = 10'd635,
    COMP_LOOP_C_353 = 10'd636,
    COMP_LOOP_C_354 = 10'd637,
    COMP_LOOP_C_355 = 10'd638,
    COMP_LOOP_C_356 = 10'd639,
    COMP_LOOP_C_357 = 10'd640,
    COMP_LOOP_C_358 = 10'd641,
    COMP_LOOP_C_359 = 10'd642,
    COMP_LOOP_C_360 = 10'd643,
    COMP_LOOP_C_361 = 10'd644,
    COMP_LOOP_C_362 = 10'd645,
    COMP_LOOP_C_363 = 10'd646,
    COMP_LOOP_C_364 = 10'd647,
    COMP_LOOP_C_365 = 10'd648,
    COMP_LOOP_C_366 = 10'd649,
    COMP_LOOP_C_367 = 10'd650,
    COMP_LOOP_C_368 = 10'd651,
    COMP_LOOP_C_369 = 10'd652,
    COMP_LOOP_C_370 = 10'd653,
    COMP_LOOP_C_371 = 10'd654,
    COMP_LOOP_C_372 = 10'd655,
    COMP_LOOP_C_373 = 10'd656,
    COMP_LOOP_7_modExp_1_while_C_0 = 10'd657,
    COMP_LOOP_7_modExp_1_while_C_1 = 10'd658,
    COMP_LOOP_7_modExp_1_while_C_2 = 10'd659,
    COMP_LOOP_7_modExp_1_while_C_3 = 10'd660,
    COMP_LOOP_7_modExp_1_while_C_4 = 10'd661,
    COMP_LOOP_7_modExp_1_while_C_5 = 10'd662,
    COMP_LOOP_7_modExp_1_while_C_6 = 10'd663,
    COMP_LOOP_7_modExp_1_while_C_7 = 10'd664,
    COMP_LOOP_7_modExp_1_while_C_8 = 10'd665,
    COMP_LOOP_7_modExp_1_while_C_9 = 10'd666,
    COMP_LOOP_7_modExp_1_while_C_10 = 10'd667,
    COMP_LOOP_7_modExp_1_while_C_11 = 10'd668,
    COMP_LOOP_7_modExp_1_while_C_12 = 10'd669,
    COMP_LOOP_7_modExp_1_while_C_13 = 10'd670,
    COMP_LOOP_7_modExp_1_while_C_14 = 10'd671,
    COMP_LOOP_7_modExp_1_while_C_15 = 10'd672,
    COMP_LOOP_7_modExp_1_while_C_16 = 10'd673,
    COMP_LOOP_7_modExp_1_while_C_17 = 10'd674,
    COMP_LOOP_7_modExp_1_while_C_18 = 10'd675,
    COMP_LOOP_7_modExp_1_while_C_19 = 10'd676,
    COMP_LOOP_7_modExp_1_while_C_20 = 10'd677,
    COMP_LOOP_7_modExp_1_while_C_21 = 10'd678,
    COMP_LOOP_7_modExp_1_while_C_22 = 10'd679,
    COMP_LOOP_7_modExp_1_while_C_23 = 10'd680,
    COMP_LOOP_7_modExp_1_while_C_24 = 10'd681,
    COMP_LOOP_7_modExp_1_while_C_25 = 10'd682,
    COMP_LOOP_7_modExp_1_while_C_26 = 10'd683,
    COMP_LOOP_7_modExp_1_while_C_27 = 10'd684,
    COMP_LOOP_7_modExp_1_while_C_28 = 10'd685,
    COMP_LOOP_7_modExp_1_while_C_29 = 10'd686,
    COMP_LOOP_7_modExp_1_while_C_30 = 10'd687,
    COMP_LOOP_7_modExp_1_while_C_31 = 10'd688,
    COMP_LOOP_7_modExp_1_while_C_32 = 10'd689,
    COMP_LOOP_7_modExp_1_while_C_33 = 10'd690,
    COMP_LOOP_7_modExp_1_while_C_34 = 10'd691,
    COMP_LOOP_7_modExp_1_while_C_35 = 10'd692,
    COMP_LOOP_7_modExp_1_while_C_36 = 10'd693,
    COMP_LOOP_7_modExp_1_while_C_37 = 10'd694,
    COMP_LOOP_7_modExp_1_while_C_38 = 10'd695,
    COMP_LOOP_C_374 = 10'd696,
    COMP_LOOP_C_375 = 10'd697,
    COMP_LOOP_C_376 = 10'd698,
    COMP_LOOP_C_377 = 10'd699,
    COMP_LOOP_C_378 = 10'd700,
    COMP_LOOP_C_379 = 10'd701,
    COMP_LOOP_C_380 = 10'd702,
    COMP_LOOP_C_381 = 10'd703,
    COMP_LOOP_C_382 = 10'd704,
    COMP_LOOP_C_383 = 10'd705,
    COMP_LOOP_C_384 = 10'd706,
    COMP_LOOP_C_385 = 10'd707,
    COMP_LOOP_C_386 = 10'd708,
    COMP_LOOP_C_387 = 10'd709,
    COMP_LOOP_C_388 = 10'd710,
    COMP_LOOP_C_389 = 10'd711,
    COMP_LOOP_C_390 = 10'd712,
    COMP_LOOP_C_391 = 10'd713,
    COMP_LOOP_C_392 = 10'd714,
    COMP_LOOP_C_393 = 10'd715,
    COMP_LOOP_C_394 = 10'd716,
    COMP_LOOP_C_395 = 10'd717,
    COMP_LOOP_C_396 = 10'd718,
    COMP_LOOP_C_397 = 10'd719,
    COMP_LOOP_C_398 = 10'd720,
    COMP_LOOP_C_399 = 10'd721,
    COMP_LOOP_C_400 = 10'd722,
    COMP_LOOP_C_401 = 10'd723,
    COMP_LOOP_C_402 = 10'd724,
    COMP_LOOP_C_403 = 10'd725,
    COMP_LOOP_C_404 = 10'd726,
    COMP_LOOP_C_405 = 10'd727,
    COMP_LOOP_C_406 = 10'd728,
    COMP_LOOP_C_407 = 10'd729,
    COMP_LOOP_C_408 = 10'd730,
    COMP_LOOP_C_409 = 10'd731,
    COMP_LOOP_C_410 = 10'd732,
    COMP_LOOP_C_411 = 10'd733,
    COMP_LOOP_C_412 = 10'd734,
    COMP_LOOP_C_413 = 10'd735,
    COMP_LOOP_C_414 = 10'd736,
    COMP_LOOP_C_415 = 10'd737,
    COMP_LOOP_C_416 = 10'd738,
    COMP_LOOP_C_417 = 10'd739,
    COMP_LOOP_C_418 = 10'd740,
    COMP_LOOP_C_419 = 10'd741,
    COMP_LOOP_C_420 = 10'd742,
    COMP_LOOP_C_421 = 10'd743,
    COMP_LOOP_C_422 = 10'd744,
    COMP_LOOP_C_423 = 10'd745,
    COMP_LOOP_C_424 = 10'd746,
    COMP_LOOP_C_425 = 10'd747,
    COMP_LOOP_C_426 = 10'd748,
    COMP_LOOP_C_427 = 10'd749,
    COMP_LOOP_C_428 = 10'd750,
    COMP_LOOP_C_429 = 10'd751,
    COMP_LOOP_C_430 = 10'd752,
    COMP_LOOP_C_431 = 10'd753,
    COMP_LOOP_C_432 = 10'd754,
    COMP_LOOP_C_433 = 10'd755,
    COMP_LOOP_C_434 = 10'd756,
    COMP_LOOP_C_435 = 10'd757,
    COMP_LOOP_8_modExp_1_while_C_0 = 10'd758,
    COMP_LOOP_8_modExp_1_while_C_1 = 10'd759,
    COMP_LOOP_8_modExp_1_while_C_2 = 10'd760,
    COMP_LOOP_8_modExp_1_while_C_3 = 10'd761,
    COMP_LOOP_8_modExp_1_while_C_4 = 10'd762,
    COMP_LOOP_8_modExp_1_while_C_5 = 10'd763,
    COMP_LOOP_8_modExp_1_while_C_6 = 10'd764,
    COMP_LOOP_8_modExp_1_while_C_7 = 10'd765,
    COMP_LOOP_8_modExp_1_while_C_8 = 10'd766,
    COMP_LOOP_8_modExp_1_while_C_9 = 10'd767,
    COMP_LOOP_8_modExp_1_while_C_10 = 10'd768,
    COMP_LOOP_8_modExp_1_while_C_11 = 10'd769,
    COMP_LOOP_8_modExp_1_while_C_12 = 10'd770,
    COMP_LOOP_8_modExp_1_while_C_13 = 10'd771,
    COMP_LOOP_8_modExp_1_while_C_14 = 10'd772,
    COMP_LOOP_8_modExp_1_while_C_15 = 10'd773,
    COMP_LOOP_8_modExp_1_while_C_16 = 10'd774,
    COMP_LOOP_8_modExp_1_while_C_17 = 10'd775,
    COMP_LOOP_8_modExp_1_while_C_18 = 10'd776,
    COMP_LOOP_8_modExp_1_while_C_19 = 10'd777,
    COMP_LOOP_8_modExp_1_while_C_20 = 10'd778,
    COMP_LOOP_8_modExp_1_while_C_21 = 10'd779,
    COMP_LOOP_8_modExp_1_while_C_22 = 10'd780,
    COMP_LOOP_8_modExp_1_while_C_23 = 10'd781,
    COMP_LOOP_8_modExp_1_while_C_24 = 10'd782,
    COMP_LOOP_8_modExp_1_while_C_25 = 10'd783,
    COMP_LOOP_8_modExp_1_while_C_26 = 10'd784,
    COMP_LOOP_8_modExp_1_while_C_27 = 10'd785,
    COMP_LOOP_8_modExp_1_while_C_28 = 10'd786,
    COMP_LOOP_8_modExp_1_while_C_29 = 10'd787,
    COMP_LOOP_8_modExp_1_while_C_30 = 10'd788,
    COMP_LOOP_8_modExp_1_while_C_31 = 10'd789,
    COMP_LOOP_8_modExp_1_while_C_32 = 10'd790,
    COMP_LOOP_8_modExp_1_while_C_33 = 10'd791,
    COMP_LOOP_8_modExp_1_while_C_34 = 10'd792,
    COMP_LOOP_8_modExp_1_while_C_35 = 10'd793,
    COMP_LOOP_8_modExp_1_while_C_36 = 10'd794,
    COMP_LOOP_8_modExp_1_while_C_37 = 10'd795,
    COMP_LOOP_8_modExp_1_while_C_38 = 10'd796,
    COMP_LOOP_C_436 = 10'd797,
    COMP_LOOP_C_437 = 10'd798,
    COMP_LOOP_C_438 = 10'd799,
    COMP_LOOP_C_439 = 10'd800,
    COMP_LOOP_C_440 = 10'd801,
    COMP_LOOP_C_441 = 10'd802,
    COMP_LOOP_C_442 = 10'd803,
    COMP_LOOP_C_443 = 10'd804,
    COMP_LOOP_C_444 = 10'd805,
    COMP_LOOP_C_445 = 10'd806,
    COMP_LOOP_C_446 = 10'd807,
    COMP_LOOP_C_447 = 10'd808,
    COMP_LOOP_C_448 = 10'd809,
    COMP_LOOP_C_449 = 10'd810,
    COMP_LOOP_C_450 = 10'd811,
    COMP_LOOP_C_451 = 10'd812,
    COMP_LOOP_C_452 = 10'd813,
    COMP_LOOP_C_453 = 10'd814,
    COMP_LOOP_C_454 = 10'd815,
    COMP_LOOP_C_455 = 10'd816,
    COMP_LOOP_C_456 = 10'd817,
    COMP_LOOP_C_457 = 10'd818,
    COMP_LOOP_C_458 = 10'd819,
    COMP_LOOP_C_459 = 10'd820,
    COMP_LOOP_C_460 = 10'd821,
    COMP_LOOP_C_461 = 10'd822,
    COMP_LOOP_C_462 = 10'd823,
    COMP_LOOP_C_463 = 10'd824,
    COMP_LOOP_C_464 = 10'd825,
    COMP_LOOP_C_465 = 10'd826,
    COMP_LOOP_C_466 = 10'd827,
    COMP_LOOP_C_467 = 10'd828,
    COMP_LOOP_C_468 = 10'd829,
    COMP_LOOP_C_469 = 10'd830,
    COMP_LOOP_C_470 = 10'd831,
    COMP_LOOP_C_471 = 10'd832,
    COMP_LOOP_C_472 = 10'd833,
    COMP_LOOP_C_473 = 10'd834,
    COMP_LOOP_C_474 = 10'd835,
    COMP_LOOP_C_475 = 10'd836,
    COMP_LOOP_C_476 = 10'd837,
    COMP_LOOP_C_477 = 10'd838,
    COMP_LOOP_C_478 = 10'd839,
    COMP_LOOP_C_479 = 10'd840,
    COMP_LOOP_C_480 = 10'd841,
    COMP_LOOP_C_481 = 10'd842,
    COMP_LOOP_C_482 = 10'd843,
    COMP_LOOP_C_483 = 10'd844,
    COMP_LOOP_C_484 = 10'd845,
    COMP_LOOP_C_485 = 10'd846,
    COMP_LOOP_C_486 = 10'd847,
    COMP_LOOP_C_487 = 10'd848,
    COMP_LOOP_C_488 = 10'd849,
    COMP_LOOP_C_489 = 10'd850,
    COMP_LOOP_C_490 = 10'd851,
    COMP_LOOP_C_491 = 10'd852,
    COMP_LOOP_C_492 = 10'd853,
    COMP_LOOP_C_493 = 10'd854,
    COMP_LOOP_C_494 = 10'd855,
    COMP_LOOP_C_495 = 10'd856,
    COMP_LOOP_C_496 = 10'd857,
    VEC_LOOP_C_0 = 10'd858,
    STAGE_LOOP_C_9 = 10'd859,
    main_C_1 = 10'd860;

  reg [9:0] state_var;
  reg [9:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : inPlaceNTT_DIT_core_core_fsm_1
    case (state_var)
      STAGE_LOOP_C_0 : begin
        fsm_output = 10'b0000000001;
        state_var_NS = STAGE_LOOP_C_1;
      end
      STAGE_LOOP_C_1 : begin
        fsm_output = 10'b0000000010;
        state_var_NS = STAGE_LOOP_C_2;
      end
      STAGE_LOOP_C_2 : begin
        fsm_output = 10'b0000000011;
        state_var_NS = STAGE_LOOP_C_3;
      end
      STAGE_LOOP_C_3 : begin
        fsm_output = 10'b0000000100;
        state_var_NS = STAGE_LOOP_C_4;
      end
      STAGE_LOOP_C_4 : begin
        fsm_output = 10'b0000000101;
        state_var_NS = STAGE_LOOP_C_5;
      end
      STAGE_LOOP_C_5 : begin
        fsm_output = 10'b0000000110;
        state_var_NS = STAGE_LOOP_C_6;
      end
      STAGE_LOOP_C_6 : begin
        fsm_output = 10'b0000000111;
        state_var_NS = STAGE_LOOP_C_7;
      end
      STAGE_LOOP_C_7 : begin
        fsm_output = 10'b0000001000;
        state_var_NS = STAGE_LOOP_C_8;
      end
      STAGE_LOOP_C_8 : begin
        fsm_output = 10'b0000001001;
        if ( STAGE_LOOP_C_8_tr0 ) begin
          state_var_NS = COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_while_C_0;
        end
      end
      modExp_while_C_0 : begin
        fsm_output = 10'b0000001010;
        state_var_NS = modExp_while_C_1;
      end
      modExp_while_C_1 : begin
        fsm_output = 10'b0000001011;
        state_var_NS = modExp_while_C_2;
      end
      modExp_while_C_2 : begin
        fsm_output = 10'b0000001100;
        state_var_NS = modExp_while_C_3;
      end
      modExp_while_C_3 : begin
        fsm_output = 10'b0000001101;
        state_var_NS = modExp_while_C_4;
      end
      modExp_while_C_4 : begin
        fsm_output = 10'b0000001110;
        state_var_NS = modExp_while_C_5;
      end
      modExp_while_C_5 : begin
        fsm_output = 10'b0000001111;
        state_var_NS = modExp_while_C_6;
      end
      modExp_while_C_6 : begin
        fsm_output = 10'b0000010000;
        state_var_NS = modExp_while_C_7;
      end
      modExp_while_C_7 : begin
        fsm_output = 10'b0000010001;
        state_var_NS = modExp_while_C_8;
      end
      modExp_while_C_8 : begin
        fsm_output = 10'b0000010010;
        state_var_NS = modExp_while_C_9;
      end
      modExp_while_C_9 : begin
        fsm_output = 10'b0000010011;
        state_var_NS = modExp_while_C_10;
      end
      modExp_while_C_10 : begin
        fsm_output = 10'b0000010100;
        state_var_NS = modExp_while_C_11;
      end
      modExp_while_C_11 : begin
        fsm_output = 10'b0000010101;
        state_var_NS = modExp_while_C_12;
      end
      modExp_while_C_12 : begin
        fsm_output = 10'b0000010110;
        state_var_NS = modExp_while_C_13;
      end
      modExp_while_C_13 : begin
        fsm_output = 10'b0000010111;
        state_var_NS = modExp_while_C_14;
      end
      modExp_while_C_14 : begin
        fsm_output = 10'b0000011000;
        state_var_NS = modExp_while_C_15;
      end
      modExp_while_C_15 : begin
        fsm_output = 10'b0000011001;
        state_var_NS = modExp_while_C_16;
      end
      modExp_while_C_16 : begin
        fsm_output = 10'b0000011010;
        state_var_NS = modExp_while_C_17;
      end
      modExp_while_C_17 : begin
        fsm_output = 10'b0000011011;
        state_var_NS = modExp_while_C_18;
      end
      modExp_while_C_18 : begin
        fsm_output = 10'b0000011100;
        state_var_NS = modExp_while_C_19;
      end
      modExp_while_C_19 : begin
        fsm_output = 10'b0000011101;
        state_var_NS = modExp_while_C_20;
      end
      modExp_while_C_20 : begin
        fsm_output = 10'b0000011110;
        state_var_NS = modExp_while_C_21;
      end
      modExp_while_C_21 : begin
        fsm_output = 10'b0000011111;
        state_var_NS = modExp_while_C_22;
      end
      modExp_while_C_22 : begin
        fsm_output = 10'b0000100000;
        state_var_NS = modExp_while_C_23;
      end
      modExp_while_C_23 : begin
        fsm_output = 10'b0000100001;
        state_var_NS = modExp_while_C_24;
      end
      modExp_while_C_24 : begin
        fsm_output = 10'b0000100010;
        state_var_NS = modExp_while_C_25;
      end
      modExp_while_C_25 : begin
        fsm_output = 10'b0000100011;
        state_var_NS = modExp_while_C_26;
      end
      modExp_while_C_26 : begin
        fsm_output = 10'b0000100100;
        state_var_NS = modExp_while_C_27;
      end
      modExp_while_C_27 : begin
        fsm_output = 10'b0000100101;
        state_var_NS = modExp_while_C_28;
      end
      modExp_while_C_28 : begin
        fsm_output = 10'b0000100110;
        state_var_NS = modExp_while_C_29;
      end
      modExp_while_C_29 : begin
        fsm_output = 10'b0000100111;
        state_var_NS = modExp_while_C_30;
      end
      modExp_while_C_30 : begin
        fsm_output = 10'b0000101000;
        state_var_NS = modExp_while_C_31;
      end
      modExp_while_C_31 : begin
        fsm_output = 10'b0000101001;
        state_var_NS = modExp_while_C_32;
      end
      modExp_while_C_32 : begin
        fsm_output = 10'b0000101010;
        state_var_NS = modExp_while_C_33;
      end
      modExp_while_C_33 : begin
        fsm_output = 10'b0000101011;
        state_var_NS = modExp_while_C_34;
      end
      modExp_while_C_34 : begin
        fsm_output = 10'b0000101100;
        state_var_NS = modExp_while_C_35;
      end
      modExp_while_C_35 : begin
        fsm_output = 10'b0000101101;
        state_var_NS = modExp_while_C_36;
      end
      modExp_while_C_36 : begin
        fsm_output = 10'b0000101110;
        state_var_NS = modExp_while_C_37;
      end
      modExp_while_C_37 : begin
        fsm_output = 10'b0000101111;
        state_var_NS = modExp_while_C_38;
      end
      modExp_while_C_38 : begin
        fsm_output = 10'b0000110000;
        if ( modExp_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_while_C_0;
        end
      end
      COMP_LOOP_C_0 : begin
        fsm_output = 10'b0000110001;
        state_var_NS = COMP_LOOP_C_1;
      end
      COMP_LOOP_C_1 : begin
        fsm_output = 10'b0000110010;
        if ( COMP_LOOP_C_1_tr0 ) begin
          state_var_NS = COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_1_modExp_1_while_C_0 : begin
        fsm_output = 10'b0000110011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_1;
      end
      COMP_LOOP_1_modExp_1_while_C_1 : begin
        fsm_output = 10'b0000110100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_2;
      end
      COMP_LOOP_1_modExp_1_while_C_2 : begin
        fsm_output = 10'b0000110101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_3;
      end
      COMP_LOOP_1_modExp_1_while_C_3 : begin
        fsm_output = 10'b0000110110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_4;
      end
      COMP_LOOP_1_modExp_1_while_C_4 : begin
        fsm_output = 10'b0000110111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_5;
      end
      COMP_LOOP_1_modExp_1_while_C_5 : begin
        fsm_output = 10'b0000111000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_6;
      end
      COMP_LOOP_1_modExp_1_while_C_6 : begin
        fsm_output = 10'b0000111001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_7;
      end
      COMP_LOOP_1_modExp_1_while_C_7 : begin
        fsm_output = 10'b0000111010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_8;
      end
      COMP_LOOP_1_modExp_1_while_C_8 : begin
        fsm_output = 10'b0000111011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_9;
      end
      COMP_LOOP_1_modExp_1_while_C_9 : begin
        fsm_output = 10'b0000111100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_10;
      end
      COMP_LOOP_1_modExp_1_while_C_10 : begin
        fsm_output = 10'b0000111101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_11;
      end
      COMP_LOOP_1_modExp_1_while_C_11 : begin
        fsm_output = 10'b0000111110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_12;
      end
      COMP_LOOP_1_modExp_1_while_C_12 : begin
        fsm_output = 10'b0000111111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_13;
      end
      COMP_LOOP_1_modExp_1_while_C_13 : begin
        fsm_output = 10'b0001000000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_14;
      end
      COMP_LOOP_1_modExp_1_while_C_14 : begin
        fsm_output = 10'b0001000001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_15;
      end
      COMP_LOOP_1_modExp_1_while_C_15 : begin
        fsm_output = 10'b0001000010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_16;
      end
      COMP_LOOP_1_modExp_1_while_C_16 : begin
        fsm_output = 10'b0001000011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_17;
      end
      COMP_LOOP_1_modExp_1_while_C_17 : begin
        fsm_output = 10'b0001000100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_18;
      end
      COMP_LOOP_1_modExp_1_while_C_18 : begin
        fsm_output = 10'b0001000101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_19;
      end
      COMP_LOOP_1_modExp_1_while_C_19 : begin
        fsm_output = 10'b0001000110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_20;
      end
      COMP_LOOP_1_modExp_1_while_C_20 : begin
        fsm_output = 10'b0001000111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_21;
      end
      COMP_LOOP_1_modExp_1_while_C_21 : begin
        fsm_output = 10'b0001001000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_22;
      end
      COMP_LOOP_1_modExp_1_while_C_22 : begin
        fsm_output = 10'b0001001001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_23;
      end
      COMP_LOOP_1_modExp_1_while_C_23 : begin
        fsm_output = 10'b0001001010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_24;
      end
      COMP_LOOP_1_modExp_1_while_C_24 : begin
        fsm_output = 10'b0001001011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_25;
      end
      COMP_LOOP_1_modExp_1_while_C_25 : begin
        fsm_output = 10'b0001001100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_26;
      end
      COMP_LOOP_1_modExp_1_while_C_26 : begin
        fsm_output = 10'b0001001101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_27;
      end
      COMP_LOOP_1_modExp_1_while_C_27 : begin
        fsm_output = 10'b0001001110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_28;
      end
      COMP_LOOP_1_modExp_1_while_C_28 : begin
        fsm_output = 10'b0001001111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_29;
      end
      COMP_LOOP_1_modExp_1_while_C_29 : begin
        fsm_output = 10'b0001010000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_30;
      end
      COMP_LOOP_1_modExp_1_while_C_30 : begin
        fsm_output = 10'b0001010001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_31;
      end
      COMP_LOOP_1_modExp_1_while_C_31 : begin
        fsm_output = 10'b0001010010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_32;
      end
      COMP_LOOP_1_modExp_1_while_C_32 : begin
        fsm_output = 10'b0001010011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_33;
      end
      COMP_LOOP_1_modExp_1_while_C_33 : begin
        fsm_output = 10'b0001010100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_34;
      end
      COMP_LOOP_1_modExp_1_while_C_34 : begin
        fsm_output = 10'b0001010101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_35;
      end
      COMP_LOOP_1_modExp_1_while_C_35 : begin
        fsm_output = 10'b0001010110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_36;
      end
      COMP_LOOP_1_modExp_1_while_C_36 : begin
        fsm_output = 10'b0001010111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_37;
      end
      COMP_LOOP_1_modExp_1_while_C_37 : begin
        fsm_output = 10'b0001011000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_38;
      end
      COMP_LOOP_1_modExp_1_while_C_38 : begin
        fsm_output = 10'b0001011001;
        if ( COMP_LOOP_1_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_2 : begin
        fsm_output = 10'b0001011010;
        state_var_NS = COMP_LOOP_C_3;
      end
      COMP_LOOP_C_3 : begin
        fsm_output = 10'b0001011011;
        state_var_NS = COMP_LOOP_C_4;
      end
      COMP_LOOP_C_4 : begin
        fsm_output = 10'b0001011100;
        state_var_NS = COMP_LOOP_C_5;
      end
      COMP_LOOP_C_5 : begin
        fsm_output = 10'b0001011101;
        state_var_NS = COMP_LOOP_C_6;
      end
      COMP_LOOP_C_6 : begin
        fsm_output = 10'b0001011110;
        state_var_NS = COMP_LOOP_C_7;
      end
      COMP_LOOP_C_7 : begin
        fsm_output = 10'b0001011111;
        state_var_NS = COMP_LOOP_C_8;
      end
      COMP_LOOP_C_8 : begin
        fsm_output = 10'b0001100000;
        state_var_NS = COMP_LOOP_C_9;
      end
      COMP_LOOP_C_9 : begin
        fsm_output = 10'b0001100001;
        state_var_NS = COMP_LOOP_C_10;
      end
      COMP_LOOP_C_10 : begin
        fsm_output = 10'b0001100010;
        state_var_NS = COMP_LOOP_C_11;
      end
      COMP_LOOP_C_11 : begin
        fsm_output = 10'b0001100011;
        state_var_NS = COMP_LOOP_C_12;
      end
      COMP_LOOP_C_12 : begin
        fsm_output = 10'b0001100100;
        state_var_NS = COMP_LOOP_C_13;
      end
      COMP_LOOP_C_13 : begin
        fsm_output = 10'b0001100101;
        state_var_NS = COMP_LOOP_C_14;
      end
      COMP_LOOP_C_14 : begin
        fsm_output = 10'b0001100110;
        state_var_NS = COMP_LOOP_C_15;
      end
      COMP_LOOP_C_15 : begin
        fsm_output = 10'b0001100111;
        state_var_NS = COMP_LOOP_C_16;
      end
      COMP_LOOP_C_16 : begin
        fsm_output = 10'b0001101000;
        state_var_NS = COMP_LOOP_C_17;
      end
      COMP_LOOP_C_17 : begin
        fsm_output = 10'b0001101001;
        state_var_NS = COMP_LOOP_C_18;
      end
      COMP_LOOP_C_18 : begin
        fsm_output = 10'b0001101010;
        state_var_NS = COMP_LOOP_C_19;
      end
      COMP_LOOP_C_19 : begin
        fsm_output = 10'b0001101011;
        state_var_NS = COMP_LOOP_C_20;
      end
      COMP_LOOP_C_20 : begin
        fsm_output = 10'b0001101100;
        state_var_NS = COMP_LOOP_C_21;
      end
      COMP_LOOP_C_21 : begin
        fsm_output = 10'b0001101101;
        state_var_NS = COMP_LOOP_C_22;
      end
      COMP_LOOP_C_22 : begin
        fsm_output = 10'b0001101110;
        state_var_NS = COMP_LOOP_C_23;
      end
      COMP_LOOP_C_23 : begin
        fsm_output = 10'b0001101111;
        state_var_NS = COMP_LOOP_C_24;
      end
      COMP_LOOP_C_24 : begin
        fsm_output = 10'b0001110000;
        state_var_NS = COMP_LOOP_C_25;
      end
      COMP_LOOP_C_25 : begin
        fsm_output = 10'b0001110001;
        state_var_NS = COMP_LOOP_C_26;
      end
      COMP_LOOP_C_26 : begin
        fsm_output = 10'b0001110010;
        state_var_NS = COMP_LOOP_C_27;
      end
      COMP_LOOP_C_27 : begin
        fsm_output = 10'b0001110011;
        state_var_NS = COMP_LOOP_C_28;
      end
      COMP_LOOP_C_28 : begin
        fsm_output = 10'b0001110100;
        state_var_NS = COMP_LOOP_C_29;
      end
      COMP_LOOP_C_29 : begin
        fsm_output = 10'b0001110101;
        state_var_NS = COMP_LOOP_C_30;
      end
      COMP_LOOP_C_30 : begin
        fsm_output = 10'b0001110110;
        state_var_NS = COMP_LOOP_C_31;
      end
      COMP_LOOP_C_31 : begin
        fsm_output = 10'b0001110111;
        state_var_NS = COMP_LOOP_C_32;
      end
      COMP_LOOP_C_32 : begin
        fsm_output = 10'b0001111000;
        state_var_NS = COMP_LOOP_C_33;
      end
      COMP_LOOP_C_33 : begin
        fsm_output = 10'b0001111001;
        state_var_NS = COMP_LOOP_C_34;
      end
      COMP_LOOP_C_34 : begin
        fsm_output = 10'b0001111010;
        state_var_NS = COMP_LOOP_C_35;
      end
      COMP_LOOP_C_35 : begin
        fsm_output = 10'b0001111011;
        state_var_NS = COMP_LOOP_C_36;
      end
      COMP_LOOP_C_36 : begin
        fsm_output = 10'b0001111100;
        state_var_NS = COMP_LOOP_C_37;
      end
      COMP_LOOP_C_37 : begin
        fsm_output = 10'b0001111101;
        state_var_NS = COMP_LOOP_C_38;
      end
      COMP_LOOP_C_38 : begin
        fsm_output = 10'b0001111110;
        state_var_NS = COMP_LOOP_C_39;
      end
      COMP_LOOP_C_39 : begin
        fsm_output = 10'b0001111111;
        state_var_NS = COMP_LOOP_C_40;
      end
      COMP_LOOP_C_40 : begin
        fsm_output = 10'b0010000000;
        state_var_NS = COMP_LOOP_C_41;
      end
      COMP_LOOP_C_41 : begin
        fsm_output = 10'b0010000001;
        state_var_NS = COMP_LOOP_C_42;
      end
      COMP_LOOP_C_42 : begin
        fsm_output = 10'b0010000010;
        state_var_NS = COMP_LOOP_C_43;
      end
      COMP_LOOP_C_43 : begin
        fsm_output = 10'b0010000011;
        state_var_NS = COMP_LOOP_C_44;
      end
      COMP_LOOP_C_44 : begin
        fsm_output = 10'b0010000100;
        state_var_NS = COMP_LOOP_C_45;
      end
      COMP_LOOP_C_45 : begin
        fsm_output = 10'b0010000101;
        state_var_NS = COMP_LOOP_C_46;
      end
      COMP_LOOP_C_46 : begin
        fsm_output = 10'b0010000110;
        state_var_NS = COMP_LOOP_C_47;
      end
      COMP_LOOP_C_47 : begin
        fsm_output = 10'b0010000111;
        state_var_NS = COMP_LOOP_C_48;
      end
      COMP_LOOP_C_48 : begin
        fsm_output = 10'b0010001000;
        state_var_NS = COMP_LOOP_C_49;
      end
      COMP_LOOP_C_49 : begin
        fsm_output = 10'b0010001001;
        state_var_NS = COMP_LOOP_C_50;
      end
      COMP_LOOP_C_50 : begin
        fsm_output = 10'b0010001010;
        state_var_NS = COMP_LOOP_C_51;
      end
      COMP_LOOP_C_51 : begin
        fsm_output = 10'b0010001011;
        state_var_NS = COMP_LOOP_C_52;
      end
      COMP_LOOP_C_52 : begin
        fsm_output = 10'b0010001100;
        state_var_NS = COMP_LOOP_C_53;
      end
      COMP_LOOP_C_53 : begin
        fsm_output = 10'b0010001101;
        state_var_NS = COMP_LOOP_C_54;
      end
      COMP_LOOP_C_54 : begin
        fsm_output = 10'b0010001110;
        state_var_NS = COMP_LOOP_C_55;
      end
      COMP_LOOP_C_55 : begin
        fsm_output = 10'b0010001111;
        state_var_NS = COMP_LOOP_C_56;
      end
      COMP_LOOP_C_56 : begin
        fsm_output = 10'b0010010000;
        state_var_NS = COMP_LOOP_C_57;
      end
      COMP_LOOP_C_57 : begin
        fsm_output = 10'b0010010001;
        state_var_NS = COMP_LOOP_C_58;
      end
      COMP_LOOP_C_58 : begin
        fsm_output = 10'b0010010010;
        state_var_NS = COMP_LOOP_C_59;
      end
      COMP_LOOP_C_59 : begin
        fsm_output = 10'b0010010011;
        state_var_NS = COMP_LOOP_C_60;
      end
      COMP_LOOP_C_60 : begin
        fsm_output = 10'b0010010100;
        state_var_NS = COMP_LOOP_C_61;
      end
      COMP_LOOP_C_61 : begin
        fsm_output = 10'b0010010101;
        state_var_NS = COMP_LOOP_C_62;
      end
      COMP_LOOP_C_62 : begin
        fsm_output = 10'b0010010110;
        if ( COMP_LOOP_C_62_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_63;
        end
      end
      COMP_LOOP_C_63 : begin
        fsm_output = 10'b0010010111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_0;
      end
      COMP_LOOP_2_modExp_1_while_C_0 : begin
        fsm_output = 10'b0010011000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_1;
      end
      COMP_LOOP_2_modExp_1_while_C_1 : begin
        fsm_output = 10'b0010011001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_2;
      end
      COMP_LOOP_2_modExp_1_while_C_2 : begin
        fsm_output = 10'b0010011010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_3;
      end
      COMP_LOOP_2_modExp_1_while_C_3 : begin
        fsm_output = 10'b0010011011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_4;
      end
      COMP_LOOP_2_modExp_1_while_C_4 : begin
        fsm_output = 10'b0010011100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_5;
      end
      COMP_LOOP_2_modExp_1_while_C_5 : begin
        fsm_output = 10'b0010011101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_6;
      end
      COMP_LOOP_2_modExp_1_while_C_6 : begin
        fsm_output = 10'b0010011110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_7;
      end
      COMP_LOOP_2_modExp_1_while_C_7 : begin
        fsm_output = 10'b0010011111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_8;
      end
      COMP_LOOP_2_modExp_1_while_C_8 : begin
        fsm_output = 10'b0010100000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_9;
      end
      COMP_LOOP_2_modExp_1_while_C_9 : begin
        fsm_output = 10'b0010100001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_10;
      end
      COMP_LOOP_2_modExp_1_while_C_10 : begin
        fsm_output = 10'b0010100010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_11;
      end
      COMP_LOOP_2_modExp_1_while_C_11 : begin
        fsm_output = 10'b0010100011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_12;
      end
      COMP_LOOP_2_modExp_1_while_C_12 : begin
        fsm_output = 10'b0010100100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_13;
      end
      COMP_LOOP_2_modExp_1_while_C_13 : begin
        fsm_output = 10'b0010100101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_14;
      end
      COMP_LOOP_2_modExp_1_while_C_14 : begin
        fsm_output = 10'b0010100110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_15;
      end
      COMP_LOOP_2_modExp_1_while_C_15 : begin
        fsm_output = 10'b0010100111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_16;
      end
      COMP_LOOP_2_modExp_1_while_C_16 : begin
        fsm_output = 10'b0010101000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_17;
      end
      COMP_LOOP_2_modExp_1_while_C_17 : begin
        fsm_output = 10'b0010101001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_18;
      end
      COMP_LOOP_2_modExp_1_while_C_18 : begin
        fsm_output = 10'b0010101010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_19;
      end
      COMP_LOOP_2_modExp_1_while_C_19 : begin
        fsm_output = 10'b0010101011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_20;
      end
      COMP_LOOP_2_modExp_1_while_C_20 : begin
        fsm_output = 10'b0010101100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_21;
      end
      COMP_LOOP_2_modExp_1_while_C_21 : begin
        fsm_output = 10'b0010101101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_22;
      end
      COMP_LOOP_2_modExp_1_while_C_22 : begin
        fsm_output = 10'b0010101110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_23;
      end
      COMP_LOOP_2_modExp_1_while_C_23 : begin
        fsm_output = 10'b0010101111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_24;
      end
      COMP_LOOP_2_modExp_1_while_C_24 : begin
        fsm_output = 10'b0010110000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_25;
      end
      COMP_LOOP_2_modExp_1_while_C_25 : begin
        fsm_output = 10'b0010110001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_26;
      end
      COMP_LOOP_2_modExp_1_while_C_26 : begin
        fsm_output = 10'b0010110010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_27;
      end
      COMP_LOOP_2_modExp_1_while_C_27 : begin
        fsm_output = 10'b0010110011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_28;
      end
      COMP_LOOP_2_modExp_1_while_C_28 : begin
        fsm_output = 10'b0010110100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_29;
      end
      COMP_LOOP_2_modExp_1_while_C_29 : begin
        fsm_output = 10'b0010110101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_30;
      end
      COMP_LOOP_2_modExp_1_while_C_30 : begin
        fsm_output = 10'b0010110110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_31;
      end
      COMP_LOOP_2_modExp_1_while_C_31 : begin
        fsm_output = 10'b0010110111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_32;
      end
      COMP_LOOP_2_modExp_1_while_C_32 : begin
        fsm_output = 10'b0010111000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_33;
      end
      COMP_LOOP_2_modExp_1_while_C_33 : begin
        fsm_output = 10'b0010111001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_34;
      end
      COMP_LOOP_2_modExp_1_while_C_34 : begin
        fsm_output = 10'b0010111010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_35;
      end
      COMP_LOOP_2_modExp_1_while_C_35 : begin
        fsm_output = 10'b0010111011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_36;
      end
      COMP_LOOP_2_modExp_1_while_C_36 : begin
        fsm_output = 10'b0010111100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_37;
      end
      COMP_LOOP_2_modExp_1_while_C_37 : begin
        fsm_output = 10'b0010111101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_38;
      end
      COMP_LOOP_2_modExp_1_while_C_38 : begin
        fsm_output = 10'b0010111110;
        if ( COMP_LOOP_2_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_64;
        end
        else begin
          state_var_NS = COMP_LOOP_2_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_64 : begin
        fsm_output = 10'b0010111111;
        state_var_NS = COMP_LOOP_C_65;
      end
      COMP_LOOP_C_65 : begin
        fsm_output = 10'b0011000000;
        state_var_NS = COMP_LOOP_C_66;
      end
      COMP_LOOP_C_66 : begin
        fsm_output = 10'b0011000001;
        state_var_NS = COMP_LOOP_C_67;
      end
      COMP_LOOP_C_67 : begin
        fsm_output = 10'b0011000010;
        state_var_NS = COMP_LOOP_C_68;
      end
      COMP_LOOP_C_68 : begin
        fsm_output = 10'b0011000011;
        state_var_NS = COMP_LOOP_C_69;
      end
      COMP_LOOP_C_69 : begin
        fsm_output = 10'b0011000100;
        state_var_NS = COMP_LOOP_C_70;
      end
      COMP_LOOP_C_70 : begin
        fsm_output = 10'b0011000101;
        state_var_NS = COMP_LOOP_C_71;
      end
      COMP_LOOP_C_71 : begin
        fsm_output = 10'b0011000110;
        state_var_NS = COMP_LOOP_C_72;
      end
      COMP_LOOP_C_72 : begin
        fsm_output = 10'b0011000111;
        state_var_NS = COMP_LOOP_C_73;
      end
      COMP_LOOP_C_73 : begin
        fsm_output = 10'b0011001000;
        state_var_NS = COMP_LOOP_C_74;
      end
      COMP_LOOP_C_74 : begin
        fsm_output = 10'b0011001001;
        state_var_NS = COMP_LOOP_C_75;
      end
      COMP_LOOP_C_75 : begin
        fsm_output = 10'b0011001010;
        state_var_NS = COMP_LOOP_C_76;
      end
      COMP_LOOP_C_76 : begin
        fsm_output = 10'b0011001011;
        state_var_NS = COMP_LOOP_C_77;
      end
      COMP_LOOP_C_77 : begin
        fsm_output = 10'b0011001100;
        state_var_NS = COMP_LOOP_C_78;
      end
      COMP_LOOP_C_78 : begin
        fsm_output = 10'b0011001101;
        state_var_NS = COMP_LOOP_C_79;
      end
      COMP_LOOP_C_79 : begin
        fsm_output = 10'b0011001110;
        state_var_NS = COMP_LOOP_C_80;
      end
      COMP_LOOP_C_80 : begin
        fsm_output = 10'b0011001111;
        state_var_NS = COMP_LOOP_C_81;
      end
      COMP_LOOP_C_81 : begin
        fsm_output = 10'b0011010000;
        state_var_NS = COMP_LOOP_C_82;
      end
      COMP_LOOP_C_82 : begin
        fsm_output = 10'b0011010001;
        state_var_NS = COMP_LOOP_C_83;
      end
      COMP_LOOP_C_83 : begin
        fsm_output = 10'b0011010010;
        state_var_NS = COMP_LOOP_C_84;
      end
      COMP_LOOP_C_84 : begin
        fsm_output = 10'b0011010011;
        state_var_NS = COMP_LOOP_C_85;
      end
      COMP_LOOP_C_85 : begin
        fsm_output = 10'b0011010100;
        state_var_NS = COMP_LOOP_C_86;
      end
      COMP_LOOP_C_86 : begin
        fsm_output = 10'b0011010101;
        state_var_NS = COMP_LOOP_C_87;
      end
      COMP_LOOP_C_87 : begin
        fsm_output = 10'b0011010110;
        state_var_NS = COMP_LOOP_C_88;
      end
      COMP_LOOP_C_88 : begin
        fsm_output = 10'b0011010111;
        state_var_NS = COMP_LOOP_C_89;
      end
      COMP_LOOP_C_89 : begin
        fsm_output = 10'b0011011000;
        state_var_NS = COMP_LOOP_C_90;
      end
      COMP_LOOP_C_90 : begin
        fsm_output = 10'b0011011001;
        state_var_NS = COMP_LOOP_C_91;
      end
      COMP_LOOP_C_91 : begin
        fsm_output = 10'b0011011010;
        state_var_NS = COMP_LOOP_C_92;
      end
      COMP_LOOP_C_92 : begin
        fsm_output = 10'b0011011011;
        state_var_NS = COMP_LOOP_C_93;
      end
      COMP_LOOP_C_93 : begin
        fsm_output = 10'b0011011100;
        state_var_NS = COMP_LOOP_C_94;
      end
      COMP_LOOP_C_94 : begin
        fsm_output = 10'b0011011101;
        state_var_NS = COMP_LOOP_C_95;
      end
      COMP_LOOP_C_95 : begin
        fsm_output = 10'b0011011110;
        state_var_NS = COMP_LOOP_C_96;
      end
      COMP_LOOP_C_96 : begin
        fsm_output = 10'b0011011111;
        state_var_NS = COMP_LOOP_C_97;
      end
      COMP_LOOP_C_97 : begin
        fsm_output = 10'b0011100000;
        state_var_NS = COMP_LOOP_C_98;
      end
      COMP_LOOP_C_98 : begin
        fsm_output = 10'b0011100001;
        state_var_NS = COMP_LOOP_C_99;
      end
      COMP_LOOP_C_99 : begin
        fsm_output = 10'b0011100010;
        state_var_NS = COMP_LOOP_C_100;
      end
      COMP_LOOP_C_100 : begin
        fsm_output = 10'b0011100011;
        state_var_NS = COMP_LOOP_C_101;
      end
      COMP_LOOP_C_101 : begin
        fsm_output = 10'b0011100100;
        state_var_NS = COMP_LOOP_C_102;
      end
      COMP_LOOP_C_102 : begin
        fsm_output = 10'b0011100101;
        state_var_NS = COMP_LOOP_C_103;
      end
      COMP_LOOP_C_103 : begin
        fsm_output = 10'b0011100110;
        state_var_NS = COMP_LOOP_C_104;
      end
      COMP_LOOP_C_104 : begin
        fsm_output = 10'b0011100111;
        state_var_NS = COMP_LOOP_C_105;
      end
      COMP_LOOP_C_105 : begin
        fsm_output = 10'b0011101000;
        state_var_NS = COMP_LOOP_C_106;
      end
      COMP_LOOP_C_106 : begin
        fsm_output = 10'b0011101001;
        state_var_NS = COMP_LOOP_C_107;
      end
      COMP_LOOP_C_107 : begin
        fsm_output = 10'b0011101010;
        state_var_NS = COMP_LOOP_C_108;
      end
      COMP_LOOP_C_108 : begin
        fsm_output = 10'b0011101011;
        state_var_NS = COMP_LOOP_C_109;
      end
      COMP_LOOP_C_109 : begin
        fsm_output = 10'b0011101100;
        state_var_NS = COMP_LOOP_C_110;
      end
      COMP_LOOP_C_110 : begin
        fsm_output = 10'b0011101101;
        state_var_NS = COMP_LOOP_C_111;
      end
      COMP_LOOP_C_111 : begin
        fsm_output = 10'b0011101110;
        state_var_NS = COMP_LOOP_C_112;
      end
      COMP_LOOP_C_112 : begin
        fsm_output = 10'b0011101111;
        state_var_NS = COMP_LOOP_C_113;
      end
      COMP_LOOP_C_113 : begin
        fsm_output = 10'b0011110000;
        state_var_NS = COMP_LOOP_C_114;
      end
      COMP_LOOP_C_114 : begin
        fsm_output = 10'b0011110001;
        state_var_NS = COMP_LOOP_C_115;
      end
      COMP_LOOP_C_115 : begin
        fsm_output = 10'b0011110010;
        state_var_NS = COMP_LOOP_C_116;
      end
      COMP_LOOP_C_116 : begin
        fsm_output = 10'b0011110011;
        state_var_NS = COMP_LOOP_C_117;
      end
      COMP_LOOP_C_117 : begin
        fsm_output = 10'b0011110100;
        state_var_NS = COMP_LOOP_C_118;
      end
      COMP_LOOP_C_118 : begin
        fsm_output = 10'b0011110101;
        state_var_NS = COMP_LOOP_C_119;
      end
      COMP_LOOP_C_119 : begin
        fsm_output = 10'b0011110110;
        state_var_NS = COMP_LOOP_C_120;
      end
      COMP_LOOP_C_120 : begin
        fsm_output = 10'b0011110111;
        state_var_NS = COMP_LOOP_C_121;
      end
      COMP_LOOP_C_121 : begin
        fsm_output = 10'b0011111000;
        state_var_NS = COMP_LOOP_C_122;
      end
      COMP_LOOP_C_122 : begin
        fsm_output = 10'b0011111001;
        state_var_NS = COMP_LOOP_C_123;
      end
      COMP_LOOP_C_123 : begin
        fsm_output = 10'b0011111010;
        state_var_NS = COMP_LOOP_C_124;
      end
      COMP_LOOP_C_124 : begin
        fsm_output = 10'b0011111011;
        if ( COMP_LOOP_C_124_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_125;
        end
      end
      COMP_LOOP_C_125 : begin
        fsm_output = 10'b0011111100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_0;
      end
      COMP_LOOP_3_modExp_1_while_C_0 : begin
        fsm_output = 10'b0011111101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_1;
      end
      COMP_LOOP_3_modExp_1_while_C_1 : begin
        fsm_output = 10'b0011111110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_2;
      end
      COMP_LOOP_3_modExp_1_while_C_2 : begin
        fsm_output = 10'b0011111111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_3;
      end
      COMP_LOOP_3_modExp_1_while_C_3 : begin
        fsm_output = 10'b0100000000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_4;
      end
      COMP_LOOP_3_modExp_1_while_C_4 : begin
        fsm_output = 10'b0100000001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_5;
      end
      COMP_LOOP_3_modExp_1_while_C_5 : begin
        fsm_output = 10'b0100000010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_6;
      end
      COMP_LOOP_3_modExp_1_while_C_6 : begin
        fsm_output = 10'b0100000011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_7;
      end
      COMP_LOOP_3_modExp_1_while_C_7 : begin
        fsm_output = 10'b0100000100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_8;
      end
      COMP_LOOP_3_modExp_1_while_C_8 : begin
        fsm_output = 10'b0100000101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_9;
      end
      COMP_LOOP_3_modExp_1_while_C_9 : begin
        fsm_output = 10'b0100000110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_10;
      end
      COMP_LOOP_3_modExp_1_while_C_10 : begin
        fsm_output = 10'b0100000111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_11;
      end
      COMP_LOOP_3_modExp_1_while_C_11 : begin
        fsm_output = 10'b0100001000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_12;
      end
      COMP_LOOP_3_modExp_1_while_C_12 : begin
        fsm_output = 10'b0100001001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_13;
      end
      COMP_LOOP_3_modExp_1_while_C_13 : begin
        fsm_output = 10'b0100001010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_14;
      end
      COMP_LOOP_3_modExp_1_while_C_14 : begin
        fsm_output = 10'b0100001011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_15;
      end
      COMP_LOOP_3_modExp_1_while_C_15 : begin
        fsm_output = 10'b0100001100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_16;
      end
      COMP_LOOP_3_modExp_1_while_C_16 : begin
        fsm_output = 10'b0100001101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_17;
      end
      COMP_LOOP_3_modExp_1_while_C_17 : begin
        fsm_output = 10'b0100001110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_18;
      end
      COMP_LOOP_3_modExp_1_while_C_18 : begin
        fsm_output = 10'b0100001111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_19;
      end
      COMP_LOOP_3_modExp_1_while_C_19 : begin
        fsm_output = 10'b0100010000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_20;
      end
      COMP_LOOP_3_modExp_1_while_C_20 : begin
        fsm_output = 10'b0100010001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_21;
      end
      COMP_LOOP_3_modExp_1_while_C_21 : begin
        fsm_output = 10'b0100010010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_22;
      end
      COMP_LOOP_3_modExp_1_while_C_22 : begin
        fsm_output = 10'b0100010011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_23;
      end
      COMP_LOOP_3_modExp_1_while_C_23 : begin
        fsm_output = 10'b0100010100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_24;
      end
      COMP_LOOP_3_modExp_1_while_C_24 : begin
        fsm_output = 10'b0100010101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_25;
      end
      COMP_LOOP_3_modExp_1_while_C_25 : begin
        fsm_output = 10'b0100010110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_26;
      end
      COMP_LOOP_3_modExp_1_while_C_26 : begin
        fsm_output = 10'b0100010111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_27;
      end
      COMP_LOOP_3_modExp_1_while_C_27 : begin
        fsm_output = 10'b0100011000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_28;
      end
      COMP_LOOP_3_modExp_1_while_C_28 : begin
        fsm_output = 10'b0100011001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_29;
      end
      COMP_LOOP_3_modExp_1_while_C_29 : begin
        fsm_output = 10'b0100011010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_30;
      end
      COMP_LOOP_3_modExp_1_while_C_30 : begin
        fsm_output = 10'b0100011011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_31;
      end
      COMP_LOOP_3_modExp_1_while_C_31 : begin
        fsm_output = 10'b0100011100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_32;
      end
      COMP_LOOP_3_modExp_1_while_C_32 : begin
        fsm_output = 10'b0100011101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_33;
      end
      COMP_LOOP_3_modExp_1_while_C_33 : begin
        fsm_output = 10'b0100011110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_34;
      end
      COMP_LOOP_3_modExp_1_while_C_34 : begin
        fsm_output = 10'b0100011111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_35;
      end
      COMP_LOOP_3_modExp_1_while_C_35 : begin
        fsm_output = 10'b0100100000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_36;
      end
      COMP_LOOP_3_modExp_1_while_C_36 : begin
        fsm_output = 10'b0100100001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_37;
      end
      COMP_LOOP_3_modExp_1_while_C_37 : begin
        fsm_output = 10'b0100100010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_38;
      end
      COMP_LOOP_3_modExp_1_while_C_38 : begin
        fsm_output = 10'b0100100011;
        if ( COMP_LOOP_3_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_126;
        end
        else begin
          state_var_NS = COMP_LOOP_3_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_126 : begin
        fsm_output = 10'b0100100100;
        state_var_NS = COMP_LOOP_C_127;
      end
      COMP_LOOP_C_127 : begin
        fsm_output = 10'b0100100101;
        state_var_NS = COMP_LOOP_C_128;
      end
      COMP_LOOP_C_128 : begin
        fsm_output = 10'b0100100110;
        state_var_NS = COMP_LOOP_C_129;
      end
      COMP_LOOP_C_129 : begin
        fsm_output = 10'b0100100111;
        state_var_NS = COMP_LOOP_C_130;
      end
      COMP_LOOP_C_130 : begin
        fsm_output = 10'b0100101000;
        state_var_NS = COMP_LOOP_C_131;
      end
      COMP_LOOP_C_131 : begin
        fsm_output = 10'b0100101001;
        state_var_NS = COMP_LOOP_C_132;
      end
      COMP_LOOP_C_132 : begin
        fsm_output = 10'b0100101010;
        state_var_NS = COMP_LOOP_C_133;
      end
      COMP_LOOP_C_133 : begin
        fsm_output = 10'b0100101011;
        state_var_NS = COMP_LOOP_C_134;
      end
      COMP_LOOP_C_134 : begin
        fsm_output = 10'b0100101100;
        state_var_NS = COMP_LOOP_C_135;
      end
      COMP_LOOP_C_135 : begin
        fsm_output = 10'b0100101101;
        state_var_NS = COMP_LOOP_C_136;
      end
      COMP_LOOP_C_136 : begin
        fsm_output = 10'b0100101110;
        state_var_NS = COMP_LOOP_C_137;
      end
      COMP_LOOP_C_137 : begin
        fsm_output = 10'b0100101111;
        state_var_NS = COMP_LOOP_C_138;
      end
      COMP_LOOP_C_138 : begin
        fsm_output = 10'b0100110000;
        state_var_NS = COMP_LOOP_C_139;
      end
      COMP_LOOP_C_139 : begin
        fsm_output = 10'b0100110001;
        state_var_NS = COMP_LOOP_C_140;
      end
      COMP_LOOP_C_140 : begin
        fsm_output = 10'b0100110010;
        state_var_NS = COMP_LOOP_C_141;
      end
      COMP_LOOP_C_141 : begin
        fsm_output = 10'b0100110011;
        state_var_NS = COMP_LOOP_C_142;
      end
      COMP_LOOP_C_142 : begin
        fsm_output = 10'b0100110100;
        state_var_NS = COMP_LOOP_C_143;
      end
      COMP_LOOP_C_143 : begin
        fsm_output = 10'b0100110101;
        state_var_NS = COMP_LOOP_C_144;
      end
      COMP_LOOP_C_144 : begin
        fsm_output = 10'b0100110110;
        state_var_NS = COMP_LOOP_C_145;
      end
      COMP_LOOP_C_145 : begin
        fsm_output = 10'b0100110111;
        state_var_NS = COMP_LOOP_C_146;
      end
      COMP_LOOP_C_146 : begin
        fsm_output = 10'b0100111000;
        state_var_NS = COMP_LOOP_C_147;
      end
      COMP_LOOP_C_147 : begin
        fsm_output = 10'b0100111001;
        state_var_NS = COMP_LOOP_C_148;
      end
      COMP_LOOP_C_148 : begin
        fsm_output = 10'b0100111010;
        state_var_NS = COMP_LOOP_C_149;
      end
      COMP_LOOP_C_149 : begin
        fsm_output = 10'b0100111011;
        state_var_NS = COMP_LOOP_C_150;
      end
      COMP_LOOP_C_150 : begin
        fsm_output = 10'b0100111100;
        state_var_NS = COMP_LOOP_C_151;
      end
      COMP_LOOP_C_151 : begin
        fsm_output = 10'b0100111101;
        state_var_NS = COMP_LOOP_C_152;
      end
      COMP_LOOP_C_152 : begin
        fsm_output = 10'b0100111110;
        state_var_NS = COMP_LOOP_C_153;
      end
      COMP_LOOP_C_153 : begin
        fsm_output = 10'b0100111111;
        state_var_NS = COMP_LOOP_C_154;
      end
      COMP_LOOP_C_154 : begin
        fsm_output = 10'b0101000000;
        state_var_NS = COMP_LOOP_C_155;
      end
      COMP_LOOP_C_155 : begin
        fsm_output = 10'b0101000001;
        state_var_NS = COMP_LOOP_C_156;
      end
      COMP_LOOP_C_156 : begin
        fsm_output = 10'b0101000010;
        state_var_NS = COMP_LOOP_C_157;
      end
      COMP_LOOP_C_157 : begin
        fsm_output = 10'b0101000011;
        state_var_NS = COMP_LOOP_C_158;
      end
      COMP_LOOP_C_158 : begin
        fsm_output = 10'b0101000100;
        state_var_NS = COMP_LOOP_C_159;
      end
      COMP_LOOP_C_159 : begin
        fsm_output = 10'b0101000101;
        state_var_NS = COMP_LOOP_C_160;
      end
      COMP_LOOP_C_160 : begin
        fsm_output = 10'b0101000110;
        state_var_NS = COMP_LOOP_C_161;
      end
      COMP_LOOP_C_161 : begin
        fsm_output = 10'b0101000111;
        state_var_NS = COMP_LOOP_C_162;
      end
      COMP_LOOP_C_162 : begin
        fsm_output = 10'b0101001000;
        state_var_NS = COMP_LOOP_C_163;
      end
      COMP_LOOP_C_163 : begin
        fsm_output = 10'b0101001001;
        state_var_NS = COMP_LOOP_C_164;
      end
      COMP_LOOP_C_164 : begin
        fsm_output = 10'b0101001010;
        state_var_NS = COMP_LOOP_C_165;
      end
      COMP_LOOP_C_165 : begin
        fsm_output = 10'b0101001011;
        state_var_NS = COMP_LOOP_C_166;
      end
      COMP_LOOP_C_166 : begin
        fsm_output = 10'b0101001100;
        state_var_NS = COMP_LOOP_C_167;
      end
      COMP_LOOP_C_167 : begin
        fsm_output = 10'b0101001101;
        state_var_NS = COMP_LOOP_C_168;
      end
      COMP_LOOP_C_168 : begin
        fsm_output = 10'b0101001110;
        state_var_NS = COMP_LOOP_C_169;
      end
      COMP_LOOP_C_169 : begin
        fsm_output = 10'b0101001111;
        state_var_NS = COMP_LOOP_C_170;
      end
      COMP_LOOP_C_170 : begin
        fsm_output = 10'b0101010000;
        state_var_NS = COMP_LOOP_C_171;
      end
      COMP_LOOP_C_171 : begin
        fsm_output = 10'b0101010001;
        state_var_NS = COMP_LOOP_C_172;
      end
      COMP_LOOP_C_172 : begin
        fsm_output = 10'b0101010010;
        state_var_NS = COMP_LOOP_C_173;
      end
      COMP_LOOP_C_173 : begin
        fsm_output = 10'b0101010011;
        state_var_NS = COMP_LOOP_C_174;
      end
      COMP_LOOP_C_174 : begin
        fsm_output = 10'b0101010100;
        state_var_NS = COMP_LOOP_C_175;
      end
      COMP_LOOP_C_175 : begin
        fsm_output = 10'b0101010101;
        state_var_NS = COMP_LOOP_C_176;
      end
      COMP_LOOP_C_176 : begin
        fsm_output = 10'b0101010110;
        state_var_NS = COMP_LOOP_C_177;
      end
      COMP_LOOP_C_177 : begin
        fsm_output = 10'b0101010111;
        state_var_NS = COMP_LOOP_C_178;
      end
      COMP_LOOP_C_178 : begin
        fsm_output = 10'b0101011000;
        state_var_NS = COMP_LOOP_C_179;
      end
      COMP_LOOP_C_179 : begin
        fsm_output = 10'b0101011001;
        state_var_NS = COMP_LOOP_C_180;
      end
      COMP_LOOP_C_180 : begin
        fsm_output = 10'b0101011010;
        state_var_NS = COMP_LOOP_C_181;
      end
      COMP_LOOP_C_181 : begin
        fsm_output = 10'b0101011011;
        state_var_NS = COMP_LOOP_C_182;
      end
      COMP_LOOP_C_182 : begin
        fsm_output = 10'b0101011100;
        state_var_NS = COMP_LOOP_C_183;
      end
      COMP_LOOP_C_183 : begin
        fsm_output = 10'b0101011101;
        state_var_NS = COMP_LOOP_C_184;
      end
      COMP_LOOP_C_184 : begin
        fsm_output = 10'b0101011110;
        state_var_NS = COMP_LOOP_C_185;
      end
      COMP_LOOP_C_185 : begin
        fsm_output = 10'b0101011111;
        state_var_NS = COMP_LOOP_C_186;
      end
      COMP_LOOP_C_186 : begin
        fsm_output = 10'b0101100000;
        if ( COMP_LOOP_C_186_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_187;
        end
      end
      COMP_LOOP_C_187 : begin
        fsm_output = 10'b0101100001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_0;
      end
      COMP_LOOP_4_modExp_1_while_C_0 : begin
        fsm_output = 10'b0101100010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_1;
      end
      COMP_LOOP_4_modExp_1_while_C_1 : begin
        fsm_output = 10'b0101100011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_2;
      end
      COMP_LOOP_4_modExp_1_while_C_2 : begin
        fsm_output = 10'b0101100100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_3;
      end
      COMP_LOOP_4_modExp_1_while_C_3 : begin
        fsm_output = 10'b0101100101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_4;
      end
      COMP_LOOP_4_modExp_1_while_C_4 : begin
        fsm_output = 10'b0101100110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_5;
      end
      COMP_LOOP_4_modExp_1_while_C_5 : begin
        fsm_output = 10'b0101100111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_6;
      end
      COMP_LOOP_4_modExp_1_while_C_6 : begin
        fsm_output = 10'b0101101000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_7;
      end
      COMP_LOOP_4_modExp_1_while_C_7 : begin
        fsm_output = 10'b0101101001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_8;
      end
      COMP_LOOP_4_modExp_1_while_C_8 : begin
        fsm_output = 10'b0101101010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_9;
      end
      COMP_LOOP_4_modExp_1_while_C_9 : begin
        fsm_output = 10'b0101101011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_10;
      end
      COMP_LOOP_4_modExp_1_while_C_10 : begin
        fsm_output = 10'b0101101100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_11;
      end
      COMP_LOOP_4_modExp_1_while_C_11 : begin
        fsm_output = 10'b0101101101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_12;
      end
      COMP_LOOP_4_modExp_1_while_C_12 : begin
        fsm_output = 10'b0101101110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_13;
      end
      COMP_LOOP_4_modExp_1_while_C_13 : begin
        fsm_output = 10'b0101101111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_14;
      end
      COMP_LOOP_4_modExp_1_while_C_14 : begin
        fsm_output = 10'b0101110000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_15;
      end
      COMP_LOOP_4_modExp_1_while_C_15 : begin
        fsm_output = 10'b0101110001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_16;
      end
      COMP_LOOP_4_modExp_1_while_C_16 : begin
        fsm_output = 10'b0101110010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_17;
      end
      COMP_LOOP_4_modExp_1_while_C_17 : begin
        fsm_output = 10'b0101110011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_18;
      end
      COMP_LOOP_4_modExp_1_while_C_18 : begin
        fsm_output = 10'b0101110100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_19;
      end
      COMP_LOOP_4_modExp_1_while_C_19 : begin
        fsm_output = 10'b0101110101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_20;
      end
      COMP_LOOP_4_modExp_1_while_C_20 : begin
        fsm_output = 10'b0101110110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_21;
      end
      COMP_LOOP_4_modExp_1_while_C_21 : begin
        fsm_output = 10'b0101110111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_22;
      end
      COMP_LOOP_4_modExp_1_while_C_22 : begin
        fsm_output = 10'b0101111000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_23;
      end
      COMP_LOOP_4_modExp_1_while_C_23 : begin
        fsm_output = 10'b0101111001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_24;
      end
      COMP_LOOP_4_modExp_1_while_C_24 : begin
        fsm_output = 10'b0101111010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_25;
      end
      COMP_LOOP_4_modExp_1_while_C_25 : begin
        fsm_output = 10'b0101111011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_26;
      end
      COMP_LOOP_4_modExp_1_while_C_26 : begin
        fsm_output = 10'b0101111100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_27;
      end
      COMP_LOOP_4_modExp_1_while_C_27 : begin
        fsm_output = 10'b0101111101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_28;
      end
      COMP_LOOP_4_modExp_1_while_C_28 : begin
        fsm_output = 10'b0101111110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_29;
      end
      COMP_LOOP_4_modExp_1_while_C_29 : begin
        fsm_output = 10'b0101111111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_30;
      end
      COMP_LOOP_4_modExp_1_while_C_30 : begin
        fsm_output = 10'b0110000000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_31;
      end
      COMP_LOOP_4_modExp_1_while_C_31 : begin
        fsm_output = 10'b0110000001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_32;
      end
      COMP_LOOP_4_modExp_1_while_C_32 : begin
        fsm_output = 10'b0110000010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_33;
      end
      COMP_LOOP_4_modExp_1_while_C_33 : begin
        fsm_output = 10'b0110000011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_34;
      end
      COMP_LOOP_4_modExp_1_while_C_34 : begin
        fsm_output = 10'b0110000100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_35;
      end
      COMP_LOOP_4_modExp_1_while_C_35 : begin
        fsm_output = 10'b0110000101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_36;
      end
      COMP_LOOP_4_modExp_1_while_C_36 : begin
        fsm_output = 10'b0110000110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_37;
      end
      COMP_LOOP_4_modExp_1_while_C_37 : begin
        fsm_output = 10'b0110000111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_38;
      end
      COMP_LOOP_4_modExp_1_while_C_38 : begin
        fsm_output = 10'b0110001000;
        if ( COMP_LOOP_4_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_188;
        end
        else begin
          state_var_NS = COMP_LOOP_4_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_188 : begin
        fsm_output = 10'b0110001001;
        state_var_NS = COMP_LOOP_C_189;
      end
      COMP_LOOP_C_189 : begin
        fsm_output = 10'b0110001010;
        state_var_NS = COMP_LOOP_C_190;
      end
      COMP_LOOP_C_190 : begin
        fsm_output = 10'b0110001011;
        state_var_NS = COMP_LOOP_C_191;
      end
      COMP_LOOP_C_191 : begin
        fsm_output = 10'b0110001100;
        state_var_NS = COMP_LOOP_C_192;
      end
      COMP_LOOP_C_192 : begin
        fsm_output = 10'b0110001101;
        state_var_NS = COMP_LOOP_C_193;
      end
      COMP_LOOP_C_193 : begin
        fsm_output = 10'b0110001110;
        state_var_NS = COMP_LOOP_C_194;
      end
      COMP_LOOP_C_194 : begin
        fsm_output = 10'b0110001111;
        state_var_NS = COMP_LOOP_C_195;
      end
      COMP_LOOP_C_195 : begin
        fsm_output = 10'b0110010000;
        state_var_NS = COMP_LOOP_C_196;
      end
      COMP_LOOP_C_196 : begin
        fsm_output = 10'b0110010001;
        state_var_NS = COMP_LOOP_C_197;
      end
      COMP_LOOP_C_197 : begin
        fsm_output = 10'b0110010010;
        state_var_NS = COMP_LOOP_C_198;
      end
      COMP_LOOP_C_198 : begin
        fsm_output = 10'b0110010011;
        state_var_NS = COMP_LOOP_C_199;
      end
      COMP_LOOP_C_199 : begin
        fsm_output = 10'b0110010100;
        state_var_NS = COMP_LOOP_C_200;
      end
      COMP_LOOP_C_200 : begin
        fsm_output = 10'b0110010101;
        state_var_NS = COMP_LOOP_C_201;
      end
      COMP_LOOP_C_201 : begin
        fsm_output = 10'b0110010110;
        state_var_NS = COMP_LOOP_C_202;
      end
      COMP_LOOP_C_202 : begin
        fsm_output = 10'b0110010111;
        state_var_NS = COMP_LOOP_C_203;
      end
      COMP_LOOP_C_203 : begin
        fsm_output = 10'b0110011000;
        state_var_NS = COMP_LOOP_C_204;
      end
      COMP_LOOP_C_204 : begin
        fsm_output = 10'b0110011001;
        state_var_NS = COMP_LOOP_C_205;
      end
      COMP_LOOP_C_205 : begin
        fsm_output = 10'b0110011010;
        state_var_NS = COMP_LOOP_C_206;
      end
      COMP_LOOP_C_206 : begin
        fsm_output = 10'b0110011011;
        state_var_NS = COMP_LOOP_C_207;
      end
      COMP_LOOP_C_207 : begin
        fsm_output = 10'b0110011100;
        state_var_NS = COMP_LOOP_C_208;
      end
      COMP_LOOP_C_208 : begin
        fsm_output = 10'b0110011101;
        state_var_NS = COMP_LOOP_C_209;
      end
      COMP_LOOP_C_209 : begin
        fsm_output = 10'b0110011110;
        state_var_NS = COMP_LOOP_C_210;
      end
      COMP_LOOP_C_210 : begin
        fsm_output = 10'b0110011111;
        state_var_NS = COMP_LOOP_C_211;
      end
      COMP_LOOP_C_211 : begin
        fsm_output = 10'b0110100000;
        state_var_NS = COMP_LOOP_C_212;
      end
      COMP_LOOP_C_212 : begin
        fsm_output = 10'b0110100001;
        state_var_NS = COMP_LOOP_C_213;
      end
      COMP_LOOP_C_213 : begin
        fsm_output = 10'b0110100010;
        state_var_NS = COMP_LOOP_C_214;
      end
      COMP_LOOP_C_214 : begin
        fsm_output = 10'b0110100011;
        state_var_NS = COMP_LOOP_C_215;
      end
      COMP_LOOP_C_215 : begin
        fsm_output = 10'b0110100100;
        state_var_NS = COMP_LOOP_C_216;
      end
      COMP_LOOP_C_216 : begin
        fsm_output = 10'b0110100101;
        state_var_NS = COMP_LOOP_C_217;
      end
      COMP_LOOP_C_217 : begin
        fsm_output = 10'b0110100110;
        state_var_NS = COMP_LOOP_C_218;
      end
      COMP_LOOP_C_218 : begin
        fsm_output = 10'b0110100111;
        state_var_NS = COMP_LOOP_C_219;
      end
      COMP_LOOP_C_219 : begin
        fsm_output = 10'b0110101000;
        state_var_NS = COMP_LOOP_C_220;
      end
      COMP_LOOP_C_220 : begin
        fsm_output = 10'b0110101001;
        state_var_NS = COMP_LOOP_C_221;
      end
      COMP_LOOP_C_221 : begin
        fsm_output = 10'b0110101010;
        state_var_NS = COMP_LOOP_C_222;
      end
      COMP_LOOP_C_222 : begin
        fsm_output = 10'b0110101011;
        state_var_NS = COMP_LOOP_C_223;
      end
      COMP_LOOP_C_223 : begin
        fsm_output = 10'b0110101100;
        state_var_NS = COMP_LOOP_C_224;
      end
      COMP_LOOP_C_224 : begin
        fsm_output = 10'b0110101101;
        state_var_NS = COMP_LOOP_C_225;
      end
      COMP_LOOP_C_225 : begin
        fsm_output = 10'b0110101110;
        state_var_NS = COMP_LOOP_C_226;
      end
      COMP_LOOP_C_226 : begin
        fsm_output = 10'b0110101111;
        state_var_NS = COMP_LOOP_C_227;
      end
      COMP_LOOP_C_227 : begin
        fsm_output = 10'b0110110000;
        state_var_NS = COMP_LOOP_C_228;
      end
      COMP_LOOP_C_228 : begin
        fsm_output = 10'b0110110001;
        state_var_NS = COMP_LOOP_C_229;
      end
      COMP_LOOP_C_229 : begin
        fsm_output = 10'b0110110010;
        state_var_NS = COMP_LOOP_C_230;
      end
      COMP_LOOP_C_230 : begin
        fsm_output = 10'b0110110011;
        state_var_NS = COMP_LOOP_C_231;
      end
      COMP_LOOP_C_231 : begin
        fsm_output = 10'b0110110100;
        state_var_NS = COMP_LOOP_C_232;
      end
      COMP_LOOP_C_232 : begin
        fsm_output = 10'b0110110101;
        state_var_NS = COMP_LOOP_C_233;
      end
      COMP_LOOP_C_233 : begin
        fsm_output = 10'b0110110110;
        state_var_NS = COMP_LOOP_C_234;
      end
      COMP_LOOP_C_234 : begin
        fsm_output = 10'b0110110111;
        state_var_NS = COMP_LOOP_C_235;
      end
      COMP_LOOP_C_235 : begin
        fsm_output = 10'b0110111000;
        state_var_NS = COMP_LOOP_C_236;
      end
      COMP_LOOP_C_236 : begin
        fsm_output = 10'b0110111001;
        state_var_NS = COMP_LOOP_C_237;
      end
      COMP_LOOP_C_237 : begin
        fsm_output = 10'b0110111010;
        state_var_NS = COMP_LOOP_C_238;
      end
      COMP_LOOP_C_238 : begin
        fsm_output = 10'b0110111011;
        state_var_NS = COMP_LOOP_C_239;
      end
      COMP_LOOP_C_239 : begin
        fsm_output = 10'b0110111100;
        state_var_NS = COMP_LOOP_C_240;
      end
      COMP_LOOP_C_240 : begin
        fsm_output = 10'b0110111101;
        state_var_NS = COMP_LOOP_C_241;
      end
      COMP_LOOP_C_241 : begin
        fsm_output = 10'b0110111110;
        state_var_NS = COMP_LOOP_C_242;
      end
      COMP_LOOP_C_242 : begin
        fsm_output = 10'b0110111111;
        state_var_NS = COMP_LOOP_C_243;
      end
      COMP_LOOP_C_243 : begin
        fsm_output = 10'b0111000000;
        state_var_NS = COMP_LOOP_C_244;
      end
      COMP_LOOP_C_244 : begin
        fsm_output = 10'b0111000001;
        state_var_NS = COMP_LOOP_C_245;
      end
      COMP_LOOP_C_245 : begin
        fsm_output = 10'b0111000010;
        state_var_NS = COMP_LOOP_C_246;
      end
      COMP_LOOP_C_246 : begin
        fsm_output = 10'b0111000011;
        state_var_NS = COMP_LOOP_C_247;
      end
      COMP_LOOP_C_247 : begin
        fsm_output = 10'b0111000100;
        state_var_NS = COMP_LOOP_C_248;
      end
      COMP_LOOP_C_248 : begin
        fsm_output = 10'b0111000101;
        if ( COMP_LOOP_C_248_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_249;
        end
      end
      COMP_LOOP_C_249 : begin
        fsm_output = 10'b0111000110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_0;
      end
      COMP_LOOP_5_modExp_1_while_C_0 : begin
        fsm_output = 10'b0111000111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_1;
      end
      COMP_LOOP_5_modExp_1_while_C_1 : begin
        fsm_output = 10'b0111001000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_2;
      end
      COMP_LOOP_5_modExp_1_while_C_2 : begin
        fsm_output = 10'b0111001001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_3;
      end
      COMP_LOOP_5_modExp_1_while_C_3 : begin
        fsm_output = 10'b0111001010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_4;
      end
      COMP_LOOP_5_modExp_1_while_C_4 : begin
        fsm_output = 10'b0111001011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_5;
      end
      COMP_LOOP_5_modExp_1_while_C_5 : begin
        fsm_output = 10'b0111001100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_6;
      end
      COMP_LOOP_5_modExp_1_while_C_6 : begin
        fsm_output = 10'b0111001101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_7;
      end
      COMP_LOOP_5_modExp_1_while_C_7 : begin
        fsm_output = 10'b0111001110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_8;
      end
      COMP_LOOP_5_modExp_1_while_C_8 : begin
        fsm_output = 10'b0111001111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_9;
      end
      COMP_LOOP_5_modExp_1_while_C_9 : begin
        fsm_output = 10'b0111010000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_10;
      end
      COMP_LOOP_5_modExp_1_while_C_10 : begin
        fsm_output = 10'b0111010001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_11;
      end
      COMP_LOOP_5_modExp_1_while_C_11 : begin
        fsm_output = 10'b0111010010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_12;
      end
      COMP_LOOP_5_modExp_1_while_C_12 : begin
        fsm_output = 10'b0111010011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_13;
      end
      COMP_LOOP_5_modExp_1_while_C_13 : begin
        fsm_output = 10'b0111010100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_14;
      end
      COMP_LOOP_5_modExp_1_while_C_14 : begin
        fsm_output = 10'b0111010101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_15;
      end
      COMP_LOOP_5_modExp_1_while_C_15 : begin
        fsm_output = 10'b0111010110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_16;
      end
      COMP_LOOP_5_modExp_1_while_C_16 : begin
        fsm_output = 10'b0111010111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_17;
      end
      COMP_LOOP_5_modExp_1_while_C_17 : begin
        fsm_output = 10'b0111011000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_18;
      end
      COMP_LOOP_5_modExp_1_while_C_18 : begin
        fsm_output = 10'b0111011001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_19;
      end
      COMP_LOOP_5_modExp_1_while_C_19 : begin
        fsm_output = 10'b0111011010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_20;
      end
      COMP_LOOP_5_modExp_1_while_C_20 : begin
        fsm_output = 10'b0111011011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_21;
      end
      COMP_LOOP_5_modExp_1_while_C_21 : begin
        fsm_output = 10'b0111011100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_22;
      end
      COMP_LOOP_5_modExp_1_while_C_22 : begin
        fsm_output = 10'b0111011101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_23;
      end
      COMP_LOOP_5_modExp_1_while_C_23 : begin
        fsm_output = 10'b0111011110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_24;
      end
      COMP_LOOP_5_modExp_1_while_C_24 : begin
        fsm_output = 10'b0111011111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_25;
      end
      COMP_LOOP_5_modExp_1_while_C_25 : begin
        fsm_output = 10'b0111100000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_26;
      end
      COMP_LOOP_5_modExp_1_while_C_26 : begin
        fsm_output = 10'b0111100001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_27;
      end
      COMP_LOOP_5_modExp_1_while_C_27 : begin
        fsm_output = 10'b0111100010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_28;
      end
      COMP_LOOP_5_modExp_1_while_C_28 : begin
        fsm_output = 10'b0111100011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_29;
      end
      COMP_LOOP_5_modExp_1_while_C_29 : begin
        fsm_output = 10'b0111100100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_30;
      end
      COMP_LOOP_5_modExp_1_while_C_30 : begin
        fsm_output = 10'b0111100101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_31;
      end
      COMP_LOOP_5_modExp_1_while_C_31 : begin
        fsm_output = 10'b0111100110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_32;
      end
      COMP_LOOP_5_modExp_1_while_C_32 : begin
        fsm_output = 10'b0111100111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_33;
      end
      COMP_LOOP_5_modExp_1_while_C_33 : begin
        fsm_output = 10'b0111101000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_34;
      end
      COMP_LOOP_5_modExp_1_while_C_34 : begin
        fsm_output = 10'b0111101001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_35;
      end
      COMP_LOOP_5_modExp_1_while_C_35 : begin
        fsm_output = 10'b0111101010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_36;
      end
      COMP_LOOP_5_modExp_1_while_C_36 : begin
        fsm_output = 10'b0111101011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_37;
      end
      COMP_LOOP_5_modExp_1_while_C_37 : begin
        fsm_output = 10'b0111101100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_38;
      end
      COMP_LOOP_5_modExp_1_while_C_38 : begin
        fsm_output = 10'b0111101101;
        if ( COMP_LOOP_5_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_250;
        end
        else begin
          state_var_NS = COMP_LOOP_5_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_250 : begin
        fsm_output = 10'b0111101110;
        state_var_NS = COMP_LOOP_C_251;
      end
      COMP_LOOP_C_251 : begin
        fsm_output = 10'b0111101111;
        state_var_NS = COMP_LOOP_C_252;
      end
      COMP_LOOP_C_252 : begin
        fsm_output = 10'b0111110000;
        state_var_NS = COMP_LOOP_C_253;
      end
      COMP_LOOP_C_253 : begin
        fsm_output = 10'b0111110001;
        state_var_NS = COMP_LOOP_C_254;
      end
      COMP_LOOP_C_254 : begin
        fsm_output = 10'b0111110010;
        state_var_NS = COMP_LOOP_C_255;
      end
      COMP_LOOP_C_255 : begin
        fsm_output = 10'b0111110011;
        state_var_NS = COMP_LOOP_C_256;
      end
      COMP_LOOP_C_256 : begin
        fsm_output = 10'b0111110100;
        state_var_NS = COMP_LOOP_C_257;
      end
      COMP_LOOP_C_257 : begin
        fsm_output = 10'b0111110101;
        state_var_NS = COMP_LOOP_C_258;
      end
      COMP_LOOP_C_258 : begin
        fsm_output = 10'b0111110110;
        state_var_NS = COMP_LOOP_C_259;
      end
      COMP_LOOP_C_259 : begin
        fsm_output = 10'b0111110111;
        state_var_NS = COMP_LOOP_C_260;
      end
      COMP_LOOP_C_260 : begin
        fsm_output = 10'b0111111000;
        state_var_NS = COMP_LOOP_C_261;
      end
      COMP_LOOP_C_261 : begin
        fsm_output = 10'b0111111001;
        state_var_NS = COMP_LOOP_C_262;
      end
      COMP_LOOP_C_262 : begin
        fsm_output = 10'b0111111010;
        state_var_NS = COMP_LOOP_C_263;
      end
      COMP_LOOP_C_263 : begin
        fsm_output = 10'b0111111011;
        state_var_NS = COMP_LOOP_C_264;
      end
      COMP_LOOP_C_264 : begin
        fsm_output = 10'b0111111100;
        state_var_NS = COMP_LOOP_C_265;
      end
      COMP_LOOP_C_265 : begin
        fsm_output = 10'b0111111101;
        state_var_NS = COMP_LOOP_C_266;
      end
      COMP_LOOP_C_266 : begin
        fsm_output = 10'b0111111110;
        state_var_NS = COMP_LOOP_C_267;
      end
      COMP_LOOP_C_267 : begin
        fsm_output = 10'b0111111111;
        state_var_NS = COMP_LOOP_C_268;
      end
      COMP_LOOP_C_268 : begin
        fsm_output = 10'b1000000000;
        state_var_NS = COMP_LOOP_C_269;
      end
      COMP_LOOP_C_269 : begin
        fsm_output = 10'b1000000001;
        state_var_NS = COMP_LOOP_C_270;
      end
      COMP_LOOP_C_270 : begin
        fsm_output = 10'b1000000010;
        state_var_NS = COMP_LOOP_C_271;
      end
      COMP_LOOP_C_271 : begin
        fsm_output = 10'b1000000011;
        state_var_NS = COMP_LOOP_C_272;
      end
      COMP_LOOP_C_272 : begin
        fsm_output = 10'b1000000100;
        state_var_NS = COMP_LOOP_C_273;
      end
      COMP_LOOP_C_273 : begin
        fsm_output = 10'b1000000101;
        state_var_NS = COMP_LOOP_C_274;
      end
      COMP_LOOP_C_274 : begin
        fsm_output = 10'b1000000110;
        state_var_NS = COMP_LOOP_C_275;
      end
      COMP_LOOP_C_275 : begin
        fsm_output = 10'b1000000111;
        state_var_NS = COMP_LOOP_C_276;
      end
      COMP_LOOP_C_276 : begin
        fsm_output = 10'b1000001000;
        state_var_NS = COMP_LOOP_C_277;
      end
      COMP_LOOP_C_277 : begin
        fsm_output = 10'b1000001001;
        state_var_NS = COMP_LOOP_C_278;
      end
      COMP_LOOP_C_278 : begin
        fsm_output = 10'b1000001010;
        state_var_NS = COMP_LOOP_C_279;
      end
      COMP_LOOP_C_279 : begin
        fsm_output = 10'b1000001011;
        state_var_NS = COMP_LOOP_C_280;
      end
      COMP_LOOP_C_280 : begin
        fsm_output = 10'b1000001100;
        state_var_NS = COMP_LOOP_C_281;
      end
      COMP_LOOP_C_281 : begin
        fsm_output = 10'b1000001101;
        state_var_NS = COMP_LOOP_C_282;
      end
      COMP_LOOP_C_282 : begin
        fsm_output = 10'b1000001110;
        state_var_NS = COMP_LOOP_C_283;
      end
      COMP_LOOP_C_283 : begin
        fsm_output = 10'b1000001111;
        state_var_NS = COMP_LOOP_C_284;
      end
      COMP_LOOP_C_284 : begin
        fsm_output = 10'b1000010000;
        state_var_NS = COMP_LOOP_C_285;
      end
      COMP_LOOP_C_285 : begin
        fsm_output = 10'b1000010001;
        state_var_NS = COMP_LOOP_C_286;
      end
      COMP_LOOP_C_286 : begin
        fsm_output = 10'b1000010010;
        state_var_NS = COMP_LOOP_C_287;
      end
      COMP_LOOP_C_287 : begin
        fsm_output = 10'b1000010011;
        state_var_NS = COMP_LOOP_C_288;
      end
      COMP_LOOP_C_288 : begin
        fsm_output = 10'b1000010100;
        state_var_NS = COMP_LOOP_C_289;
      end
      COMP_LOOP_C_289 : begin
        fsm_output = 10'b1000010101;
        state_var_NS = COMP_LOOP_C_290;
      end
      COMP_LOOP_C_290 : begin
        fsm_output = 10'b1000010110;
        state_var_NS = COMP_LOOP_C_291;
      end
      COMP_LOOP_C_291 : begin
        fsm_output = 10'b1000010111;
        state_var_NS = COMP_LOOP_C_292;
      end
      COMP_LOOP_C_292 : begin
        fsm_output = 10'b1000011000;
        state_var_NS = COMP_LOOP_C_293;
      end
      COMP_LOOP_C_293 : begin
        fsm_output = 10'b1000011001;
        state_var_NS = COMP_LOOP_C_294;
      end
      COMP_LOOP_C_294 : begin
        fsm_output = 10'b1000011010;
        state_var_NS = COMP_LOOP_C_295;
      end
      COMP_LOOP_C_295 : begin
        fsm_output = 10'b1000011011;
        state_var_NS = COMP_LOOP_C_296;
      end
      COMP_LOOP_C_296 : begin
        fsm_output = 10'b1000011100;
        state_var_NS = COMP_LOOP_C_297;
      end
      COMP_LOOP_C_297 : begin
        fsm_output = 10'b1000011101;
        state_var_NS = COMP_LOOP_C_298;
      end
      COMP_LOOP_C_298 : begin
        fsm_output = 10'b1000011110;
        state_var_NS = COMP_LOOP_C_299;
      end
      COMP_LOOP_C_299 : begin
        fsm_output = 10'b1000011111;
        state_var_NS = COMP_LOOP_C_300;
      end
      COMP_LOOP_C_300 : begin
        fsm_output = 10'b1000100000;
        state_var_NS = COMP_LOOP_C_301;
      end
      COMP_LOOP_C_301 : begin
        fsm_output = 10'b1000100001;
        state_var_NS = COMP_LOOP_C_302;
      end
      COMP_LOOP_C_302 : begin
        fsm_output = 10'b1000100010;
        state_var_NS = COMP_LOOP_C_303;
      end
      COMP_LOOP_C_303 : begin
        fsm_output = 10'b1000100011;
        state_var_NS = COMP_LOOP_C_304;
      end
      COMP_LOOP_C_304 : begin
        fsm_output = 10'b1000100100;
        state_var_NS = COMP_LOOP_C_305;
      end
      COMP_LOOP_C_305 : begin
        fsm_output = 10'b1000100101;
        state_var_NS = COMP_LOOP_C_306;
      end
      COMP_LOOP_C_306 : begin
        fsm_output = 10'b1000100110;
        state_var_NS = COMP_LOOP_C_307;
      end
      COMP_LOOP_C_307 : begin
        fsm_output = 10'b1000100111;
        state_var_NS = COMP_LOOP_C_308;
      end
      COMP_LOOP_C_308 : begin
        fsm_output = 10'b1000101000;
        state_var_NS = COMP_LOOP_C_309;
      end
      COMP_LOOP_C_309 : begin
        fsm_output = 10'b1000101001;
        state_var_NS = COMP_LOOP_C_310;
      end
      COMP_LOOP_C_310 : begin
        fsm_output = 10'b1000101010;
        if ( COMP_LOOP_C_310_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_311;
        end
      end
      COMP_LOOP_C_311 : begin
        fsm_output = 10'b1000101011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_0;
      end
      COMP_LOOP_6_modExp_1_while_C_0 : begin
        fsm_output = 10'b1000101100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_1;
      end
      COMP_LOOP_6_modExp_1_while_C_1 : begin
        fsm_output = 10'b1000101101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_2;
      end
      COMP_LOOP_6_modExp_1_while_C_2 : begin
        fsm_output = 10'b1000101110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_3;
      end
      COMP_LOOP_6_modExp_1_while_C_3 : begin
        fsm_output = 10'b1000101111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_4;
      end
      COMP_LOOP_6_modExp_1_while_C_4 : begin
        fsm_output = 10'b1000110000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_5;
      end
      COMP_LOOP_6_modExp_1_while_C_5 : begin
        fsm_output = 10'b1000110001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_6;
      end
      COMP_LOOP_6_modExp_1_while_C_6 : begin
        fsm_output = 10'b1000110010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_7;
      end
      COMP_LOOP_6_modExp_1_while_C_7 : begin
        fsm_output = 10'b1000110011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_8;
      end
      COMP_LOOP_6_modExp_1_while_C_8 : begin
        fsm_output = 10'b1000110100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_9;
      end
      COMP_LOOP_6_modExp_1_while_C_9 : begin
        fsm_output = 10'b1000110101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_10;
      end
      COMP_LOOP_6_modExp_1_while_C_10 : begin
        fsm_output = 10'b1000110110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_11;
      end
      COMP_LOOP_6_modExp_1_while_C_11 : begin
        fsm_output = 10'b1000110111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_12;
      end
      COMP_LOOP_6_modExp_1_while_C_12 : begin
        fsm_output = 10'b1000111000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_13;
      end
      COMP_LOOP_6_modExp_1_while_C_13 : begin
        fsm_output = 10'b1000111001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_14;
      end
      COMP_LOOP_6_modExp_1_while_C_14 : begin
        fsm_output = 10'b1000111010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_15;
      end
      COMP_LOOP_6_modExp_1_while_C_15 : begin
        fsm_output = 10'b1000111011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_16;
      end
      COMP_LOOP_6_modExp_1_while_C_16 : begin
        fsm_output = 10'b1000111100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_17;
      end
      COMP_LOOP_6_modExp_1_while_C_17 : begin
        fsm_output = 10'b1000111101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_18;
      end
      COMP_LOOP_6_modExp_1_while_C_18 : begin
        fsm_output = 10'b1000111110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_19;
      end
      COMP_LOOP_6_modExp_1_while_C_19 : begin
        fsm_output = 10'b1000111111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_20;
      end
      COMP_LOOP_6_modExp_1_while_C_20 : begin
        fsm_output = 10'b1001000000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_21;
      end
      COMP_LOOP_6_modExp_1_while_C_21 : begin
        fsm_output = 10'b1001000001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_22;
      end
      COMP_LOOP_6_modExp_1_while_C_22 : begin
        fsm_output = 10'b1001000010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_23;
      end
      COMP_LOOP_6_modExp_1_while_C_23 : begin
        fsm_output = 10'b1001000011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_24;
      end
      COMP_LOOP_6_modExp_1_while_C_24 : begin
        fsm_output = 10'b1001000100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_25;
      end
      COMP_LOOP_6_modExp_1_while_C_25 : begin
        fsm_output = 10'b1001000101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_26;
      end
      COMP_LOOP_6_modExp_1_while_C_26 : begin
        fsm_output = 10'b1001000110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_27;
      end
      COMP_LOOP_6_modExp_1_while_C_27 : begin
        fsm_output = 10'b1001000111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_28;
      end
      COMP_LOOP_6_modExp_1_while_C_28 : begin
        fsm_output = 10'b1001001000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_29;
      end
      COMP_LOOP_6_modExp_1_while_C_29 : begin
        fsm_output = 10'b1001001001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_30;
      end
      COMP_LOOP_6_modExp_1_while_C_30 : begin
        fsm_output = 10'b1001001010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_31;
      end
      COMP_LOOP_6_modExp_1_while_C_31 : begin
        fsm_output = 10'b1001001011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_32;
      end
      COMP_LOOP_6_modExp_1_while_C_32 : begin
        fsm_output = 10'b1001001100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_33;
      end
      COMP_LOOP_6_modExp_1_while_C_33 : begin
        fsm_output = 10'b1001001101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_34;
      end
      COMP_LOOP_6_modExp_1_while_C_34 : begin
        fsm_output = 10'b1001001110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_35;
      end
      COMP_LOOP_6_modExp_1_while_C_35 : begin
        fsm_output = 10'b1001001111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_36;
      end
      COMP_LOOP_6_modExp_1_while_C_36 : begin
        fsm_output = 10'b1001010000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_37;
      end
      COMP_LOOP_6_modExp_1_while_C_37 : begin
        fsm_output = 10'b1001010001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_38;
      end
      COMP_LOOP_6_modExp_1_while_C_38 : begin
        fsm_output = 10'b1001010010;
        if ( COMP_LOOP_6_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_312;
        end
        else begin
          state_var_NS = COMP_LOOP_6_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_312 : begin
        fsm_output = 10'b1001010011;
        state_var_NS = COMP_LOOP_C_313;
      end
      COMP_LOOP_C_313 : begin
        fsm_output = 10'b1001010100;
        state_var_NS = COMP_LOOP_C_314;
      end
      COMP_LOOP_C_314 : begin
        fsm_output = 10'b1001010101;
        state_var_NS = COMP_LOOP_C_315;
      end
      COMP_LOOP_C_315 : begin
        fsm_output = 10'b1001010110;
        state_var_NS = COMP_LOOP_C_316;
      end
      COMP_LOOP_C_316 : begin
        fsm_output = 10'b1001010111;
        state_var_NS = COMP_LOOP_C_317;
      end
      COMP_LOOP_C_317 : begin
        fsm_output = 10'b1001011000;
        state_var_NS = COMP_LOOP_C_318;
      end
      COMP_LOOP_C_318 : begin
        fsm_output = 10'b1001011001;
        state_var_NS = COMP_LOOP_C_319;
      end
      COMP_LOOP_C_319 : begin
        fsm_output = 10'b1001011010;
        state_var_NS = COMP_LOOP_C_320;
      end
      COMP_LOOP_C_320 : begin
        fsm_output = 10'b1001011011;
        state_var_NS = COMP_LOOP_C_321;
      end
      COMP_LOOP_C_321 : begin
        fsm_output = 10'b1001011100;
        state_var_NS = COMP_LOOP_C_322;
      end
      COMP_LOOP_C_322 : begin
        fsm_output = 10'b1001011101;
        state_var_NS = COMP_LOOP_C_323;
      end
      COMP_LOOP_C_323 : begin
        fsm_output = 10'b1001011110;
        state_var_NS = COMP_LOOP_C_324;
      end
      COMP_LOOP_C_324 : begin
        fsm_output = 10'b1001011111;
        state_var_NS = COMP_LOOP_C_325;
      end
      COMP_LOOP_C_325 : begin
        fsm_output = 10'b1001100000;
        state_var_NS = COMP_LOOP_C_326;
      end
      COMP_LOOP_C_326 : begin
        fsm_output = 10'b1001100001;
        state_var_NS = COMP_LOOP_C_327;
      end
      COMP_LOOP_C_327 : begin
        fsm_output = 10'b1001100010;
        state_var_NS = COMP_LOOP_C_328;
      end
      COMP_LOOP_C_328 : begin
        fsm_output = 10'b1001100011;
        state_var_NS = COMP_LOOP_C_329;
      end
      COMP_LOOP_C_329 : begin
        fsm_output = 10'b1001100100;
        state_var_NS = COMP_LOOP_C_330;
      end
      COMP_LOOP_C_330 : begin
        fsm_output = 10'b1001100101;
        state_var_NS = COMP_LOOP_C_331;
      end
      COMP_LOOP_C_331 : begin
        fsm_output = 10'b1001100110;
        state_var_NS = COMP_LOOP_C_332;
      end
      COMP_LOOP_C_332 : begin
        fsm_output = 10'b1001100111;
        state_var_NS = COMP_LOOP_C_333;
      end
      COMP_LOOP_C_333 : begin
        fsm_output = 10'b1001101000;
        state_var_NS = COMP_LOOP_C_334;
      end
      COMP_LOOP_C_334 : begin
        fsm_output = 10'b1001101001;
        state_var_NS = COMP_LOOP_C_335;
      end
      COMP_LOOP_C_335 : begin
        fsm_output = 10'b1001101010;
        state_var_NS = COMP_LOOP_C_336;
      end
      COMP_LOOP_C_336 : begin
        fsm_output = 10'b1001101011;
        state_var_NS = COMP_LOOP_C_337;
      end
      COMP_LOOP_C_337 : begin
        fsm_output = 10'b1001101100;
        state_var_NS = COMP_LOOP_C_338;
      end
      COMP_LOOP_C_338 : begin
        fsm_output = 10'b1001101101;
        state_var_NS = COMP_LOOP_C_339;
      end
      COMP_LOOP_C_339 : begin
        fsm_output = 10'b1001101110;
        state_var_NS = COMP_LOOP_C_340;
      end
      COMP_LOOP_C_340 : begin
        fsm_output = 10'b1001101111;
        state_var_NS = COMP_LOOP_C_341;
      end
      COMP_LOOP_C_341 : begin
        fsm_output = 10'b1001110000;
        state_var_NS = COMP_LOOP_C_342;
      end
      COMP_LOOP_C_342 : begin
        fsm_output = 10'b1001110001;
        state_var_NS = COMP_LOOP_C_343;
      end
      COMP_LOOP_C_343 : begin
        fsm_output = 10'b1001110010;
        state_var_NS = COMP_LOOP_C_344;
      end
      COMP_LOOP_C_344 : begin
        fsm_output = 10'b1001110011;
        state_var_NS = COMP_LOOP_C_345;
      end
      COMP_LOOP_C_345 : begin
        fsm_output = 10'b1001110100;
        state_var_NS = COMP_LOOP_C_346;
      end
      COMP_LOOP_C_346 : begin
        fsm_output = 10'b1001110101;
        state_var_NS = COMP_LOOP_C_347;
      end
      COMP_LOOP_C_347 : begin
        fsm_output = 10'b1001110110;
        state_var_NS = COMP_LOOP_C_348;
      end
      COMP_LOOP_C_348 : begin
        fsm_output = 10'b1001110111;
        state_var_NS = COMP_LOOP_C_349;
      end
      COMP_LOOP_C_349 : begin
        fsm_output = 10'b1001111000;
        state_var_NS = COMP_LOOP_C_350;
      end
      COMP_LOOP_C_350 : begin
        fsm_output = 10'b1001111001;
        state_var_NS = COMP_LOOP_C_351;
      end
      COMP_LOOP_C_351 : begin
        fsm_output = 10'b1001111010;
        state_var_NS = COMP_LOOP_C_352;
      end
      COMP_LOOP_C_352 : begin
        fsm_output = 10'b1001111011;
        state_var_NS = COMP_LOOP_C_353;
      end
      COMP_LOOP_C_353 : begin
        fsm_output = 10'b1001111100;
        state_var_NS = COMP_LOOP_C_354;
      end
      COMP_LOOP_C_354 : begin
        fsm_output = 10'b1001111101;
        state_var_NS = COMP_LOOP_C_355;
      end
      COMP_LOOP_C_355 : begin
        fsm_output = 10'b1001111110;
        state_var_NS = COMP_LOOP_C_356;
      end
      COMP_LOOP_C_356 : begin
        fsm_output = 10'b1001111111;
        state_var_NS = COMP_LOOP_C_357;
      end
      COMP_LOOP_C_357 : begin
        fsm_output = 10'b1010000000;
        state_var_NS = COMP_LOOP_C_358;
      end
      COMP_LOOP_C_358 : begin
        fsm_output = 10'b1010000001;
        state_var_NS = COMP_LOOP_C_359;
      end
      COMP_LOOP_C_359 : begin
        fsm_output = 10'b1010000010;
        state_var_NS = COMP_LOOP_C_360;
      end
      COMP_LOOP_C_360 : begin
        fsm_output = 10'b1010000011;
        state_var_NS = COMP_LOOP_C_361;
      end
      COMP_LOOP_C_361 : begin
        fsm_output = 10'b1010000100;
        state_var_NS = COMP_LOOP_C_362;
      end
      COMP_LOOP_C_362 : begin
        fsm_output = 10'b1010000101;
        state_var_NS = COMP_LOOP_C_363;
      end
      COMP_LOOP_C_363 : begin
        fsm_output = 10'b1010000110;
        state_var_NS = COMP_LOOP_C_364;
      end
      COMP_LOOP_C_364 : begin
        fsm_output = 10'b1010000111;
        state_var_NS = COMP_LOOP_C_365;
      end
      COMP_LOOP_C_365 : begin
        fsm_output = 10'b1010001000;
        state_var_NS = COMP_LOOP_C_366;
      end
      COMP_LOOP_C_366 : begin
        fsm_output = 10'b1010001001;
        state_var_NS = COMP_LOOP_C_367;
      end
      COMP_LOOP_C_367 : begin
        fsm_output = 10'b1010001010;
        state_var_NS = COMP_LOOP_C_368;
      end
      COMP_LOOP_C_368 : begin
        fsm_output = 10'b1010001011;
        state_var_NS = COMP_LOOP_C_369;
      end
      COMP_LOOP_C_369 : begin
        fsm_output = 10'b1010001100;
        state_var_NS = COMP_LOOP_C_370;
      end
      COMP_LOOP_C_370 : begin
        fsm_output = 10'b1010001101;
        state_var_NS = COMP_LOOP_C_371;
      end
      COMP_LOOP_C_371 : begin
        fsm_output = 10'b1010001110;
        state_var_NS = COMP_LOOP_C_372;
      end
      COMP_LOOP_C_372 : begin
        fsm_output = 10'b1010001111;
        if ( COMP_LOOP_C_372_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_373;
        end
      end
      COMP_LOOP_C_373 : begin
        fsm_output = 10'b1010010000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_0;
      end
      COMP_LOOP_7_modExp_1_while_C_0 : begin
        fsm_output = 10'b1010010001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_1;
      end
      COMP_LOOP_7_modExp_1_while_C_1 : begin
        fsm_output = 10'b1010010010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_2;
      end
      COMP_LOOP_7_modExp_1_while_C_2 : begin
        fsm_output = 10'b1010010011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_3;
      end
      COMP_LOOP_7_modExp_1_while_C_3 : begin
        fsm_output = 10'b1010010100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_4;
      end
      COMP_LOOP_7_modExp_1_while_C_4 : begin
        fsm_output = 10'b1010010101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_5;
      end
      COMP_LOOP_7_modExp_1_while_C_5 : begin
        fsm_output = 10'b1010010110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_6;
      end
      COMP_LOOP_7_modExp_1_while_C_6 : begin
        fsm_output = 10'b1010010111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_7;
      end
      COMP_LOOP_7_modExp_1_while_C_7 : begin
        fsm_output = 10'b1010011000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_8;
      end
      COMP_LOOP_7_modExp_1_while_C_8 : begin
        fsm_output = 10'b1010011001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_9;
      end
      COMP_LOOP_7_modExp_1_while_C_9 : begin
        fsm_output = 10'b1010011010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_10;
      end
      COMP_LOOP_7_modExp_1_while_C_10 : begin
        fsm_output = 10'b1010011011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_11;
      end
      COMP_LOOP_7_modExp_1_while_C_11 : begin
        fsm_output = 10'b1010011100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_12;
      end
      COMP_LOOP_7_modExp_1_while_C_12 : begin
        fsm_output = 10'b1010011101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_13;
      end
      COMP_LOOP_7_modExp_1_while_C_13 : begin
        fsm_output = 10'b1010011110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_14;
      end
      COMP_LOOP_7_modExp_1_while_C_14 : begin
        fsm_output = 10'b1010011111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_15;
      end
      COMP_LOOP_7_modExp_1_while_C_15 : begin
        fsm_output = 10'b1010100000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_16;
      end
      COMP_LOOP_7_modExp_1_while_C_16 : begin
        fsm_output = 10'b1010100001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_17;
      end
      COMP_LOOP_7_modExp_1_while_C_17 : begin
        fsm_output = 10'b1010100010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_18;
      end
      COMP_LOOP_7_modExp_1_while_C_18 : begin
        fsm_output = 10'b1010100011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_19;
      end
      COMP_LOOP_7_modExp_1_while_C_19 : begin
        fsm_output = 10'b1010100100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_20;
      end
      COMP_LOOP_7_modExp_1_while_C_20 : begin
        fsm_output = 10'b1010100101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_21;
      end
      COMP_LOOP_7_modExp_1_while_C_21 : begin
        fsm_output = 10'b1010100110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_22;
      end
      COMP_LOOP_7_modExp_1_while_C_22 : begin
        fsm_output = 10'b1010100111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_23;
      end
      COMP_LOOP_7_modExp_1_while_C_23 : begin
        fsm_output = 10'b1010101000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_24;
      end
      COMP_LOOP_7_modExp_1_while_C_24 : begin
        fsm_output = 10'b1010101001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_25;
      end
      COMP_LOOP_7_modExp_1_while_C_25 : begin
        fsm_output = 10'b1010101010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_26;
      end
      COMP_LOOP_7_modExp_1_while_C_26 : begin
        fsm_output = 10'b1010101011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_27;
      end
      COMP_LOOP_7_modExp_1_while_C_27 : begin
        fsm_output = 10'b1010101100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_28;
      end
      COMP_LOOP_7_modExp_1_while_C_28 : begin
        fsm_output = 10'b1010101101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_29;
      end
      COMP_LOOP_7_modExp_1_while_C_29 : begin
        fsm_output = 10'b1010101110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_30;
      end
      COMP_LOOP_7_modExp_1_while_C_30 : begin
        fsm_output = 10'b1010101111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_31;
      end
      COMP_LOOP_7_modExp_1_while_C_31 : begin
        fsm_output = 10'b1010110000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_32;
      end
      COMP_LOOP_7_modExp_1_while_C_32 : begin
        fsm_output = 10'b1010110001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_33;
      end
      COMP_LOOP_7_modExp_1_while_C_33 : begin
        fsm_output = 10'b1010110010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_34;
      end
      COMP_LOOP_7_modExp_1_while_C_34 : begin
        fsm_output = 10'b1010110011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_35;
      end
      COMP_LOOP_7_modExp_1_while_C_35 : begin
        fsm_output = 10'b1010110100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_36;
      end
      COMP_LOOP_7_modExp_1_while_C_36 : begin
        fsm_output = 10'b1010110101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_37;
      end
      COMP_LOOP_7_modExp_1_while_C_37 : begin
        fsm_output = 10'b1010110110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_38;
      end
      COMP_LOOP_7_modExp_1_while_C_38 : begin
        fsm_output = 10'b1010110111;
        if ( COMP_LOOP_7_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_374;
        end
        else begin
          state_var_NS = COMP_LOOP_7_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_374 : begin
        fsm_output = 10'b1010111000;
        state_var_NS = COMP_LOOP_C_375;
      end
      COMP_LOOP_C_375 : begin
        fsm_output = 10'b1010111001;
        state_var_NS = COMP_LOOP_C_376;
      end
      COMP_LOOP_C_376 : begin
        fsm_output = 10'b1010111010;
        state_var_NS = COMP_LOOP_C_377;
      end
      COMP_LOOP_C_377 : begin
        fsm_output = 10'b1010111011;
        state_var_NS = COMP_LOOP_C_378;
      end
      COMP_LOOP_C_378 : begin
        fsm_output = 10'b1010111100;
        state_var_NS = COMP_LOOP_C_379;
      end
      COMP_LOOP_C_379 : begin
        fsm_output = 10'b1010111101;
        state_var_NS = COMP_LOOP_C_380;
      end
      COMP_LOOP_C_380 : begin
        fsm_output = 10'b1010111110;
        state_var_NS = COMP_LOOP_C_381;
      end
      COMP_LOOP_C_381 : begin
        fsm_output = 10'b1010111111;
        state_var_NS = COMP_LOOP_C_382;
      end
      COMP_LOOP_C_382 : begin
        fsm_output = 10'b1011000000;
        state_var_NS = COMP_LOOP_C_383;
      end
      COMP_LOOP_C_383 : begin
        fsm_output = 10'b1011000001;
        state_var_NS = COMP_LOOP_C_384;
      end
      COMP_LOOP_C_384 : begin
        fsm_output = 10'b1011000010;
        state_var_NS = COMP_LOOP_C_385;
      end
      COMP_LOOP_C_385 : begin
        fsm_output = 10'b1011000011;
        state_var_NS = COMP_LOOP_C_386;
      end
      COMP_LOOP_C_386 : begin
        fsm_output = 10'b1011000100;
        state_var_NS = COMP_LOOP_C_387;
      end
      COMP_LOOP_C_387 : begin
        fsm_output = 10'b1011000101;
        state_var_NS = COMP_LOOP_C_388;
      end
      COMP_LOOP_C_388 : begin
        fsm_output = 10'b1011000110;
        state_var_NS = COMP_LOOP_C_389;
      end
      COMP_LOOP_C_389 : begin
        fsm_output = 10'b1011000111;
        state_var_NS = COMP_LOOP_C_390;
      end
      COMP_LOOP_C_390 : begin
        fsm_output = 10'b1011001000;
        state_var_NS = COMP_LOOP_C_391;
      end
      COMP_LOOP_C_391 : begin
        fsm_output = 10'b1011001001;
        state_var_NS = COMP_LOOP_C_392;
      end
      COMP_LOOP_C_392 : begin
        fsm_output = 10'b1011001010;
        state_var_NS = COMP_LOOP_C_393;
      end
      COMP_LOOP_C_393 : begin
        fsm_output = 10'b1011001011;
        state_var_NS = COMP_LOOP_C_394;
      end
      COMP_LOOP_C_394 : begin
        fsm_output = 10'b1011001100;
        state_var_NS = COMP_LOOP_C_395;
      end
      COMP_LOOP_C_395 : begin
        fsm_output = 10'b1011001101;
        state_var_NS = COMP_LOOP_C_396;
      end
      COMP_LOOP_C_396 : begin
        fsm_output = 10'b1011001110;
        state_var_NS = COMP_LOOP_C_397;
      end
      COMP_LOOP_C_397 : begin
        fsm_output = 10'b1011001111;
        state_var_NS = COMP_LOOP_C_398;
      end
      COMP_LOOP_C_398 : begin
        fsm_output = 10'b1011010000;
        state_var_NS = COMP_LOOP_C_399;
      end
      COMP_LOOP_C_399 : begin
        fsm_output = 10'b1011010001;
        state_var_NS = COMP_LOOP_C_400;
      end
      COMP_LOOP_C_400 : begin
        fsm_output = 10'b1011010010;
        state_var_NS = COMP_LOOP_C_401;
      end
      COMP_LOOP_C_401 : begin
        fsm_output = 10'b1011010011;
        state_var_NS = COMP_LOOP_C_402;
      end
      COMP_LOOP_C_402 : begin
        fsm_output = 10'b1011010100;
        state_var_NS = COMP_LOOP_C_403;
      end
      COMP_LOOP_C_403 : begin
        fsm_output = 10'b1011010101;
        state_var_NS = COMP_LOOP_C_404;
      end
      COMP_LOOP_C_404 : begin
        fsm_output = 10'b1011010110;
        state_var_NS = COMP_LOOP_C_405;
      end
      COMP_LOOP_C_405 : begin
        fsm_output = 10'b1011010111;
        state_var_NS = COMP_LOOP_C_406;
      end
      COMP_LOOP_C_406 : begin
        fsm_output = 10'b1011011000;
        state_var_NS = COMP_LOOP_C_407;
      end
      COMP_LOOP_C_407 : begin
        fsm_output = 10'b1011011001;
        state_var_NS = COMP_LOOP_C_408;
      end
      COMP_LOOP_C_408 : begin
        fsm_output = 10'b1011011010;
        state_var_NS = COMP_LOOP_C_409;
      end
      COMP_LOOP_C_409 : begin
        fsm_output = 10'b1011011011;
        state_var_NS = COMP_LOOP_C_410;
      end
      COMP_LOOP_C_410 : begin
        fsm_output = 10'b1011011100;
        state_var_NS = COMP_LOOP_C_411;
      end
      COMP_LOOP_C_411 : begin
        fsm_output = 10'b1011011101;
        state_var_NS = COMP_LOOP_C_412;
      end
      COMP_LOOP_C_412 : begin
        fsm_output = 10'b1011011110;
        state_var_NS = COMP_LOOP_C_413;
      end
      COMP_LOOP_C_413 : begin
        fsm_output = 10'b1011011111;
        state_var_NS = COMP_LOOP_C_414;
      end
      COMP_LOOP_C_414 : begin
        fsm_output = 10'b1011100000;
        state_var_NS = COMP_LOOP_C_415;
      end
      COMP_LOOP_C_415 : begin
        fsm_output = 10'b1011100001;
        state_var_NS = COMP_LOOP_C_416;
      end
      COMP_LOOP_C_416 : begin
        fsm_output = 10'b1011100010;
        state_var_NS = COMP_LOOP_C_417;
      end
      COMP_LOOP_C_417 : begin
        fsm_output = 10'b1011100011;
        state_var_NS = COMP_LOOP_C_418;
      end
      COMP_LOOP_C_418 : begin
        fsm_output = 10'b1011100100;
        state_var_NS = COMP_LOOP_C_419;
      end
      COMP_LOOP_C_419 : begin
        fsm_output = 10'b1011100101;
        state_var_NS = COMP_LOOP_C_420;
      end
      COMP_LOOP_C_420 : begin
        fsm_output = 10'b1011100110;
        state_var_NS = COMP_LOOP_C_421;
      end
      COMP_LOOP_C_421 : begin
        fsm_output = 10'b1011100111;
        state_var_NS = COMP_LOOP_C_422;
      end
      COMP_LOOP_C_422 : begin
        fsm_output = 10'b1011101000;
        state_var_NS = COMP_LOOP_C_423;
      end
      COMP_LOOP_C_423 : begin
        fsm_output = 10'b1011101001;
        state_var_NS = COMP_LOOP_C_424;
      end
      COMP_LOOP_C_424 : begin
        fsm_output = 10'b1011101010;
        state_var_NS = COMP_LOOP_C_425;
      end
      COMP_LOOP_C_425 : begin
        fsm_output = 10'b1011101011;
        state_var_NS = COMP_LOOP_C_426;
      end
      COMP_LOOP_C_426 : begin
        fsm_output = 10'b1011101100;
        state_var_NS = COMP_LOOP_C_427;
      end
      COMP_LOOP_C_427 : begin
        fsm_output = 10'b1011101101;
        state_var_NS = COMP_LOOP_C_428;
      end
      COMP_LOOP_C_428 : begin
        fsm_output = 10'b1011101110;
        state_var_NS = COMP_LOOP_C_429;
      end
      COMP_LOOP_C_429 : begin
        fsm_output = 10'b1011101111;
        state_var_NS = COMP_LOOP_C_430;
      end
      COMP_LOOP_C_430 : begin
        fsm_output = 10'b1011110000;
        state_var_NS = COMP_LOOP_C_431;
      end
      COMP_LOOP_C_431 : begin
        fsm_output = 10'b1011110001;
        state_var_NS = COMP_LOOP_C_432;
      end
      COMP_LOOP_C_432 : begin
        fsm_output = 10'b1011110010;
        state_var_NS = COMP_LOOP_C_433;
      end
      COMP_LOOP_C_433 : begin
        fsm_output = 10'b1011110011;
        state_var_NS = COMP_LOOP_C_434;
      end
      COMP_LOOP_C_434 : begin
        fsm_output = 10'b1011110100;
        if ( COMP_LOOP_C_434_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_435;
        end
      end
      COMP_LOOP_C_435 : begin
        fsm_output = 10'b1011110101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_0;
      end
      COMP_LOOP_8_modExp_1_while_C_0 : begin
        fsm_output = 10'b1011110110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_1;
      end
      COMP_LOOP_8_modExp_1_while_C_1 : begin
        fsm_output = 10'b1011110111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_2;
      end
      COMP_LOOP_8_modExp_1_while_C_2 : begin
        fsm_output = 10'b1011111000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_3;
      end
      COMP_LOOP_8_modExp_1_while_C_3 : begin
        fsm_output = 10'b1011111001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_4;
      end
      COMP_LOOP_8_modExp_1_while_C_4 : begin
        fsm_output = 10'b1011111010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_5;
      end
      COMP_LOOP_8_modExp_1_while_C_5 : begin
        fsm_output = 10'b1011111011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_6;
      end
      COMP_LOOP_8_modExp_1_while_C_6 : begin
        fsm_output = 10'b1011111100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_7;
      end
      COMP_LOOP_8_modExp_1_while_C_7 : begin
        fsm_output = 10'b1011111101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_8;
      end
      COMP_LOOP_8_modExp_1_while_C_8 : begin
        fsm_output = 10'b1011111110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_9;
      end
      COMP_LOOP_8_modExp_1_while_C_9 : begin
        fsm_output = 10'b1011111111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_10;
      end
      COMP_LOOP_8_modExp_1_while_C_10 : begin
        fsm_output = 10'b1100000000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_11;
      end
      COMP_LOOP_8_modExp_1_while_C_11 : begin
        fsm_output = 10'b1100000001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_12;
      end
      COMP_LOOP_8_modExp_1_while_C_12 : begin
        fsm_output = 10'b1100000010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_13;
      end
      COMP_LOOP_8_modExp_1_while_C_13 : begin
        fsm_output = 10'b1100000011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_14;
      end
      COMP_LOOP_8_modExp_1_while_C_14 : begin
        fsm_output = 10'b1100000100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_15;
      end
      COMP_LOOP_8_modExp_1_while_C_15 : begin
        fsm_output = 10'b1100000101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_16;
      end
      COMP_LOOP_8_modExp_1_while_C_16 : begin
        fsm_output = 10'b1100000110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_17;
      end
      COMP_LOOP_8_modExp_1_while_C_17 : begin
        fsm_output = 10'b1100000111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_18;
      end
      COMP_LOOP_8_modExp_1_while_C_18 : begin
        fsm_output = 10'b1100001000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_19;
      end
      COMP_LOOP_8_modExp_1_while_C_19 : begin
        fsm_output = 10'b1100001001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_20;
      end
      COMP_LOOP_8_modExp_1_while_C_20 : begin
        fsm_output = 10'b1100001010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_21;
      end
      COMP_LOOP_8_modExp_1_while_C_21 : begin
        fsm_output = 10'b1100001011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_22;
      end
      COMP_LOOP_8_modExp_1_while_C_22 : begin
        fsm_output = 10'b1100001100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_23;
      end
      COMP_LOOP_8_modExp_1_while_C_23 : begin
        fsm_output = 10'b1100001101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_24;
      end
      COMP_LOOP_8_modExp_1_while_C_24 : begin
        fsm_output = 10'b1100001110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_25;
      end
      COMP_LOOP_8_modExp_1_while_C_25 : begin
        fsm_output = 10'b1100001111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_26;
      end
      COMP_LOOP_8_modExp_1_while_C_26 : begin
        fsm_output = 10'b1100010000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_27;
      end
      COMP_LOOP_8_modExp_1_while_C_27 : begin
        fsm_output = 10'b1100010001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_28;
      end
      COMP_LOOP_8_modExp_1_while_C_28 : begin
        fsm_output = 10'b1100010010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_29;
      end
      COMP_LOOP_8_modExp_1_while_C_29 : begin
        fsm_output = 10'b1100010011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_30;
      end
      COMP_LOOP_8_modExp_1_while_C_30 : begin
        fsm_output = 10'b1100010100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_31;
      end
      COMP_LOOP_8_modExp_1_while_C_31 : begin
        fsm_output = 10'b1100010101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_32;
      end
      COMP_LOOP_8_modExp_1_while_C_32 : begin
        fsm_output = 10'b1100010110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_33;
      end
      COMP_LOOP_8_modExp_1_while_C_33 : begin
        fsm_output = 10'b1100010111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_34;
      end
      COMP_LOOP_8_modExp_1_while_C_34 : begin
        fsm_output = 10'b1100011000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_35;
      end
      COMP_LOOP_8_modExp_1_while_C_35 : begin
        fsm_output = 10'b1100011001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_36;
      end
      COMP_LOOP_8_modExp_1_while_C_36 : begin
        fsm_output = 10'b1100011010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_37;
      end
      COMP_LOOP_8_modExp_1_while_C_37 : begin
        fsm_output = 10'b1100011011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_38;
      end
      COMP_LOOP_8_modExp_1_while_C_38 : begin
        fsm_output = 10'b1100011100;
        if ( COMP_LOOP_8_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_436;
        end
        else begin
          state_var_NS = COMP_LOOP_8_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_436 : begin
        fsm_output = 10'b1100011101;
        state_var_NS = COMP_LOOP_C_437;
      end
      COMP_LOOP_C_437 : begin
        fsm_output = 10'b1100011110;
        state_var_NS = COMP_LOOP_C_438;
      end
      COMP_LOOP_C_438 : begin
        fsm_output = 10'b1100011111;
        state_var_NS = COMP_LOOP_C_439;
      end
      COMP_LOOP_C_439 : begin
        fsm_output = 10'b1100100000;
        state_var_NS = COMP_LOOP_C_440;
      end
      COMP_LOOP_C_440 : begin
        fsm_output = 10'b1100100001;
        state_var_NS = COMP_LOOP_C_441;
      end
      COMP_LOOP_C_441 : begin
        fsm_output = 10'b1100100010;
        state_var_NS = COMP_LOOP_C_442;
      end
      COMP_LOOP_C_442 : begin
        fsm_output = 10'b1100100011;
        state_var_NS = COMP_LOOP_C_443;
      end
      COMP_LOOP_C_443 : begin
        fsm_output = 10'b1100100100;
        state_var_NS = COMP_LOOP_C_444;
      end
      COMP_LOOP_C_444 : begin
        fsm_output = 10'b1100100101;
        state_var_NS = COMP_LOOP_C_445;
      end
      COMP_LOOP_C_445 : begin
        fsm_output = 10'b1100100110;
        state_var_NS = COMP_LOOP_C_446;
      end
      COMP_LOOP_C_446 : begin
        fsm_output = 10'b1100100111;
        state_var_NS = COMP_LOOP_C_447;
      end
      COMP_LOOP_C_447 : begin
        fsm_output = 10'b1100101000;
        state_var_NS = COMP_LOOP_C_448;
      end
      COMP_LOOP_C_448 : begin
        fsm_output = 10'b1100101001;
        state_var_NS = COMP_LOOP_C_449;
      end
      COMP_LOOP_C_449 : begin
        fsm_output = 10'b1100101010;
        state_var_NS = COMP_LOOP_C_450;
      end
      COMP_LOOP_C_450 : begin
        fsm_output = 10'b1100101011;
        state_var_NS = COMP_LOOP_C_451;
      end
      COMP_LOOP_C_451 : begin
        fsm_output = 10'b1100101100;
        state_var_NS = COMP_LOOP_C_452;
      end
      COMP_LOOP_C_452 : begin
        fsm_output = 10'b1100101101;
        state_var_NS = COMP_LOOP_C_453;
      end
      COMP_LOOP_C_453 : begin
        fsm_output = 10'b1100101110;
        state_var_NS = COMP_LOOP_C_454;
      end
      COMP_LOOP_C_454 : begin
        fsm_output = 10'b1100101111;
        state_var_NS = COMP_LOOP_C_455;
      end
      COMP_LOOP_C_455 : begin
        fsm_output = 10'b1100110000;
        state_var_NS = COMP_LOOP_C_456;
      end
      COMP_LOOP_C_456 : begin
        fsm_output = 10'b1100110001;
        state_var_NS = COMP_LOOP_C_457;
      end
      COMP_LOOP_C_457 : begin
        fsm_output = 10'b1100110010;
        state_var_NS = COMP_LOOP_C_458;
      end
      COMP_LOOP_C_458 : begin
        fsm_output = 10'b1100110011;
        state_var_NS = COMP_LOOP_C_459;
      end
      COMP_LOOP_C_459 : begin
        fsm_output = 10'b1100110100;
        state_var_NS = COMP_LOOP_C_460;
      end
      COMP_LOOP_C_460 : begin
        fsm_output = 10'b1100110101;
        state_var_NS = COMP_LOOP_C_461;
      end
      COMP_LOOP_C_461 : begin
        fsm_output = 10'b1100110110;
        state_var_NS = COMP_LOOP_C_462;
      end
      COMP_LOOP_C_462 : begin
        fsm_output = 10'b1100110111;
        state_var_NS = COMP_LOOP_C_463;
      end
      COMP_LOOP_C_463 : begin
        fsm_output = 10'b1100111000;
        state_var_NS = COMP_LOOP_C_464;
      end
      COMP_LOOP_C_464 : begin
        fsm_output = 10'b1100111001;
        state_var_NS = COMP_LOOP_C_465;
      end
      COMP_LOOP_C_465 : begin
        fsm_output = 10'b1100111010;
        state_var_NS = COMP_LOOP_C_466;
      end
      COMP_LOOP_C_466 : begin
        fsm_output = 10'b1100111011;
        state_var_NS = COMP_LOOP_C_467;
      end
      COMP_LOOP_C_467 : begin
        fsm_output = 10'b1100111100;
        state_var_NS = COMP_LOOP_C_468;
      end
      COMP_LOOP_C_468 : begin
        fsm_output = 10'b1100111101;
        state_var_NS = COMP_LOOP_C_469;
      end
      COMP_LOOP_C_469 : begin
        fsm_output = 10'b1100111110;
        state_var_NS = COMP_LOOP_C_470;
      end
      COMP_LOOP_C_470 : begin
        fsm_output = 10'b1100111111;
        state_var_NS = COMP_LOOP_C_471;
      end
      COMP_LOOP_C_471 : begin
        fsm_output = 10'b1101000000;
        state_var_NS = COMP_LOOP_C_472;
      end
      COMP_LOOP_C_472 : begin
        fsm_output = 10'b1101000001;
        state_var_NS = COMP_LOOP_C_473;
      end
      COMP_LOOP_C_473 : begin
        fsm_output = 10'b1101000010;
        state_var_NS = COMP_LOOP_C_474;
      end
      COMP_LOOP_C_474 : begin
        fsm_output = 10'b1101000011;
        state_var_NS = COMP_LOOP_C_475;
      end
      COMP_LOOP_C_475 : begin
        fsm_output = 10'b1101000100;
        state_var_NS = COMP_LOOP_C_476;
      end
      COMP_LOOP_C_476 : begin
        fsm_output = 10'b1101000101;
        state_var_NS = COMP_LOOP_C_477;
      end
      COMP_LOOP_C_477 : begin
        fsm_output = 10'b1101000110;
        state_var_NS = COMP_LOOP_C_478;
      end
      COMP_LOOP_C_478 : begin
        fsm_output = 10'b1101000111;
        state_var_NS = COMP_LOOP_C_479;
      end
      COMP_LOOP_C_479 : begin
        fsm_output = 10'b1101001000;
        state_var_NS = COMP_LOOP_C_480;
      end
      COMP_LOOP_C_480 : begin
        fsm_output = 10'b1101001001;
        state_var_NS = COMP_LOOP_C_481;
      end
      COMP_LOOP_C_481 : begin
        fsm_output = 10'b1101001010;
        state_var_NS = COMP_LOOP_C_482;
      end
      COMP_LOOP_C_482 : begin
        fsm_output = 10'b1101001011;
        state_var_NS = COMP_LOOP_C_483;
      end
      COMP_LOOP_C_483 : begin
        fsm_output = 10'b1101001100;
        state_var_NS = COMP_LOOP_C_484;
      end
      COMP_LOOP_C_484 : begin
        fsm_output = 10'b1101001101;
        state_var_NS = COMP_LOOP_C_485;
      end
      COMP_LOOP_C_485 : begin
        fsm_output = 10'b1101001110;
        state_var_NS = COMP_LOOP_C_486;
      end
      COMP_LOOP_C_486 : begin
        fsm_output = 10'b1101001111;
        state_var_NS = COMP_LOOP_C_487;
      end
      COMP_LOOP_C_487 : begin
        fsm_output = 10'b1101010000;
        state_var_NS = COMP_LOOP_C_488;
      end
      COMP_LOOP_C_488 : begin
        fsm_output = 10'b1101010001;
        state_var_NS = COMP_LOOP_C_489;
      end
      COMP_LOOP_C_489 : begin
        fsm_output = 10'b1101010010;
        state_var_NS = COMP_LOOP_C_490;
      end
      COMP_LOOP_C_490 : begin
        fsm_output = 10'b1101010011;
        state_var_NS = COMP_LOOP_C_491;
      end
      COMP_LOOP_C_491 : begin
        fsm_output = 10'b1101010100;
        state_var_NS = COMP_LOOP_C_492;
      end
      COMP_LOOP_C_492 : begin
        fsm_output = 10'b1101010101;
        state_var_NS = COMP_LOOP_C_493;
      end
      COMP_LOOP_C_493 : begin
        fsm_output = 10'b1101010110;
        state_var_NS = COMP_LOOP_C_494;
      end
      COMP_LOOP_C_494 : begin
        fsm_output = 10'b1101010111;
        state_var_NS = COMP_LOOP_C_495;
      end
      COMP_LOOP_C_495 : begin
        fsm_output = 10'b1101011000;
        state_var_NS = COMP_LOOP_C_496;
      end
      COMP_LOOP_C_496 : begin
        fsm_output = 10'b1101011001;
        if ( COMP_LOOP_C_496_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_C_0 : begin
        fsm_output = 10'b1101011010;
        if ( VEC_LOOP_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_9;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      STAGE_LOOP_C_9 : begin
        fsm_output = 10'b1101011011;
        if ( STAGE_LOOP_C_9_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = STAGE_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 10'b1101011100;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 10'b0000000000;
        state_var_NS = STAGE_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core (
  clk, rst, vec_rsc_triosy_0_0_lz, vec_rsc_triosy_0_1_lz, vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz, vec_rsc_triosy_0_4_lz, vec_rsc_triosy_0_5_lz, vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz, p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz,
      vec_rsc_0_0_i_qa_d, vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_1_i_qa_d,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_qa_d, vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_4_i_qa_d,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_qa_d, vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_7_i_qa_d,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_0_i_adra_d_pff, vec_rsc_0_0_i_da_d_pff,
      vec_rsc_0_0_i_wea_d_pff, vec_rsc_0_1_i_wea_d_pff, vec_rsc_0_2_i_wea_d_pff,
      vec_rsc_0_3_i_wea_d_pff, vec_rsc_0_4_i_wea_d_pff, vec_rsc_0_5_i_wea_d_pff,
      vec_rsc_0_6_i_wea_d_pff, vec_rsc_0_7_i_wea_d_pff
);
  input clk;
  input rst;
  output vec_rsc_triosy_0_0_lz;
  output vec_rsc_triosy_0_1_lz;
  output vec_rsc_triosy_0_2_lz;
  output vec_rsc_triosy_0_3_lz;
  output vec_rsc_triosy_0_4_lz;
  output vec_rsc_triosy_0_5_lz;
  output vec_rsc_triosy_0_6_lz;
  output vec_rsc_triosy_0_7_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  input [63:0] vec_rsc_0_0_i_qa_d;
  output vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_1_i_qa_d;
  output vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_2_i_qa_d;
  output vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_3_i_qa_d;
  output vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_4_i_qa_d;
  output vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_5_i_qa_d;
  output vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_6_i_qa_d;
  output vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_7_i_qa_d;
  output vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [8:0] vec_rsc_0_0_i_adra_d_pff;
  output [63:0] vec_rsc_0_0_i_da_d_pff;
  output vec_rsc_0_0_i_wea_d_pff;
  output vec_rsc_0_1_i_wea_d_pff;
  output vec_rsc_0_2_i_wea_d_pff;
  output vec_rsc_0_3_i_wea_d_pff;
  output vec_rsc_0_4_i_wea_d_pff;
  output vec_rsc_0_5_i_wea_d_pff;
  output vec_rsc_0_6_i_wea_d_pff;
  output vec_rsc_0_7_i_wea_d_pff;


  // Interconnect Declarations
  wire [63:0] p_rsci_idat;
  wire [63:0] r_rsci_idat;
  reg [63:0] modulo_result_rem_cmp_a;
  reg [63:0] modulo_result_rem_cmp_b;
  wire [63:0] modulo_result_rem_cmp_z;
  reg [64:0] operator_66_true_div_cmp_a;
  wire [64:0] operator_66_true_div_cmp_z;
  reg [9:0] operator_66_true_div_cmp_b_9_0;
  wire [9:0] fsm_output;
  wire nor_tmp;
  wire or_tmp;
  wire or_tmp_92;
  wire nor_tmp_23;
  wire or_tmp_103;
  wire nor_tmp_27;
  wire mux_tmp_156;
  wire or_tmp_113;
  wire and_dcpl_4;
  wire or_tmp_154;
  wire and_dcpl_11;
  wire and_dcpl_14;
  wire and_dcpl_23;
  wire not_tmp_131;
  wire and_dcpl_46;
  wire and_dcpl_47;
  wire and_dcpl_48;
  wire and_dcpl_50;
  wire and_dcpl_51;
  wire and_dcpl_56;
  wire and_dcpl_57;
  wire and_dcpl_58;
  wire and_dcpl_59;
  wire and_dcpl_60;
  wire and_dcpl_63;
  wire and_dcpl_64;
  wire and_dcpl_65;
  wire and_dcpl_66;
  wire and_dcpl_67;
  wire and_dcpl_68;
  wire and_dcpl_69;
  wire and_dcpl_70;
  wire and_dcpl_73;
  wire and_dcpl_80;
  wire and_dcpl_82;
  wire and_dcpl_84;
  wire and_dcpl_89;
  wire and_dcpl_91;
  wire and_dcpl_93;
  wire and_dcpl_100;
  wire and_dcpl_102;
  wire and_dcpl_103;
  wire and_dcpl_108;
  wire and_dcpl_109;
  wire and_dcpl_110;
  wire and_dcpl_112;
  wire and_dcpl_121;
  wire and_dcpl_122;
  wire and_dcpl_123;
  wire and_dcpl_127;
  wire and_dcpl_128;
  wire and_dcpl_129;
  wire and_dcpl_130;
  wire and_dcpl_137;
  wire and_dcpl_138;
  wire or_tmp_268;
  wire or_tmp_273;
  wire not_tmp_165;
  wire or_tmp_335;
  wire or_tmp_340;
  wire or_tmp_395;
  wire nand_tmp_18;
  wire or_tmp_454;
  wire nand_tmp_21;
  wire or_tmp_525;
  wire or_tmp_535;
  wire or_tmp_590;
  wire or_tmp_600;
  wire or_tmp_655;
  wire nand_tmp_31;
  wire or_tmp_719;
  wire nand_tmp_35;
  wire and_dcpl_140;
  wire and_dcpl_147;
  wire mux_tmp_677;
  wire mux_tmp_688;
  wire mux_tmp_689;
  wire nor_tmp_146;
  wire mux_tmp_705;
  wire or_tmp_788;
  wire mux_tmp_718;
  wire mux_tmp_719;
  wire mux_tmp_722;
  wire or_tmp_792;
  wire nand_tmp_42;
  wire mux_tmp_731;
  wire not_tmp_274;
  wire not_tmp_280;
  wire or_tmp_810;
  wire mux_tmp_776;
  wire not_tmp_297;
  wire not_tmp_309;
  wire not_tmp_312;
  wire not_tmp_315;
  wire and_dcpl_152;
  wire and_dcpl_156;
  wire or_tmp_891;
  wire mux_tmp_845;
  wire not_tmp_347;
  wire and_dcpl_162;
  wire or_tmp_916;
  wire mux_tmp_886;
  wire or_tmp_918;
  wire and_tmp_28;
  wire and_dcpl_164;
  wire and_dcpl_167;
  wire and_dcpl_168;
  wire and_dcpl_171;
  wire and_dcpl_172;
  wire and_dcpl_176;
  wire and_dcpl_180;
  wire and_dcpl_184;
  wire and_dcpl_187;
  wire not_tmp_374;
  wire not_tmp_399;
  wire not_tmp_400;
  wire not_tmp_406;
  wire not_tmp_414;
  wire mux_tmp_997;
  wire mux_tmp_1006;
  wire not_tmp_436;
  wire not_tmp_462;
  wire and_dcpl_219;
  wire not_tmp_480;
  wire nor_tmp_240;
  wire mux_tmp_1159;
  wire nor_tmp_241;
  wire mux_tmp_1160;
  wire and_tmp_44;
  wire mux_tmp_1162;
  wire not_tmp_482;
  wire nor_tmp_244;
  wire mux_tmp_1164;
  wire mux_tmp_1170;
  wire or_tmp_1144;
  wire and_tmp_45;
  wire and_tmp_46;
  wire mux_tmp_1178;
  wire or_tmp_1159;
  wire or_tmp_1165;
  wire mux_tmp_1202;
  wire or_tmp_1174;
  wire or_tmp_1176;
  wire and_dcpl_226;
  wire not_tmp_513;
  wire not_tmp_523;
  wire or_tmp_1261;
  wire mux_tmp_1305;
  reg COMP_LOOP_COMP_LOOP_and_11_itm;
  reg COMP_LOOP_COMP_LOOP_and_145_itm;
  reg COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [11:0] COMP_LOOP_acc_1_cse_6_sva_1;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_6_sva_1;
  reg [11:0] VEC_LOOP_j_sva_11_0;
  reg COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  reg [5:0] COMP_LOOP_k_9_3_sva_5_0;
  wire [6:0] COMP_LOOP_k_9_3_sva_2;
  wire [7:0] nl_COMP_LOOP_k_9_3_sva_2;
  reg [11:0] COMP_LOOP_acc_10_cse_12_1_1_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_6_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_2_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_4_sva;
  reg [10:0] COMP_LOOP_acc_11_psp_sva;
  wire [11:0] nl_COMP_LOOP_acc_11_psp_sva;
  reg [9:0] COMP_LOOP_acc_13_psp_sva;
  reg [10:0] COMP_LOOP_acc_14_psp_sva;
  wire [11:0] nl_COMP_LOOP_acc_14_psp_sva;
  reg [63:0] tmp_10_lpi_4_dfm;
  wire [11:0] COMP_LOOP_acc_1_cse_4_sva_1;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_4_sva_1;
  wire [11:0] COMP_LOOP_acc_1_cse_2_sva_mx0w0;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_2_sva_mx0w0;
  wire and_244_m1c;
  wire mux_984_m1c;
  wire and_224_m1c;
  wire and_226_m1c;
  wire and_229_m1c;
  wire and_230_m1c;
  wire and_233_m1c;
  wire and_235_m1c;
  wire and_237_m1c;
  wire and_187_m1c;
  wire and_416_cse;
  wire nand_190_cse;
  wire nand_168_cse;
  reg reg_vec_rsc_triosy_0_7_obj_ld_cse;
  wire and_389_cse;
  wire or_838_cse;
  wire or_1099_cse;
  wire or_1385_cse;
  wire or_1391_cse;
  wire and_477_cse;
  wire nor_425_cse;
  wire or_247_cse;
  wire and_483_cse;
  wire or_245_cse;
  wire and_314_cse;
  wire nor_393_cse;
  wire nand_100_cse;
  wire or_1189_cse;
  wire and_316_cse;
  wire [63:0] modulo_result_mux_1_cse;
  wire nand_97_cse;
  wire or_81_cse;
  wire or_83_cse;
  wire or_171_cse;
  wire or_216_cse;
  wire or_1202_cse;
  wire and_369_cse;
  wire and_437_cse;
  wire or_329_cse;
  wire or_327_cse;
  wire mux_392_cse;
  wire or_320_cse;
  wire nand_246_cse;
  wire or_314_cse;
  wire or_312_cse;
  wire nand_194_cse;
  wire nand_189_cse;
  wire and_428_cse;
  wire or_817_cse;
  wire or_242_cse;
  wire nor_601_cse;
  wire mux_29_cse;
  wire nand_230_cse;
  wire and_502_cse;
  wire or_816_cse;
  wire or_210_cse;
  wire or_1392_cse;
  wire nand_89_cse;
  wire nor_357_cse;
  wire and_361_cse;
  wire and_462_cse;
  wire and_382_cse;
  wire or_1394_cse;
  wire or_1423_cse;
  wire mux_331_cse;
  wire mux_342_cse;
  wire and_491_cse;
  wire or_115_cse;
  wire and_25_cse;
  wire [8:0] COMP_LOOP_acc_psp_sva_1;
  wire [9:0] nl_COMP_LOOP_acc_psp_sva_1;
  reg [8:0] COMP_LOOP_acc_psp_sva;
  wire mux_696_itm;
  wire mux_1158_itm;
  wire mux_1273_itm;
  wire and_dcpl;
  wire and_dcpl_236;
  wire and_dcpl_238;
  wire and_dcpl_240;
  wire and_dcpl_242;
  wire and_dcpl_243;
  wire and_dcpl_245;
  wire and_dcpl_247;
  wire and_dcpl_255;
  wire and_dcpl_260;
  wire and_dcpl_266;
  wire [9:0] z_out;
  wire and_dcpl_268;
  wire and_dcpl_269;
  wire and_dcpl_276;
  wire and_dcpl_298;
  wire [9:0] z_out_1;
  wire [10:0] nl_z_out_1;
  wire and_dcpl_324;
  wire and_dcpl_340;
  wire and_dcpl_345;
  wire [64:0] z_out_2;
  wire and_dcpl_347;
  wire and_dcpl_349;
  wire and_dcpl_354;
  wire or_tmp_1317;
  wire not_tmp_581;
  wire and_dcpl_357;
  wire and_dcpl_362;
  wire and_dcpl_364;
  wire and_dcpl_367;
  wire and_dcpl_368;
  wire and_dcpl_372;
  wire and_dcpl_379;
  wire and_dcpl_383;
  wire and_dcpl_385;
  wire and_dcpl_388;
  wire and_dcpl_394;
  wire and_dcpl_399;
  wire and_dcpl_404;
  wire and_dcpl_406;
  wire and_dcpl_409;
  wire and_dcpl_411;
  wire [64:0] z_out_3;
  wire [65:0] nl_z_out_3;
  wire or_tmp_1346;
  wire or_tmp_1348;
  wire or_tmp_1349;
  wire not_tmp_600;
  wire [63:0] z_out_4;
  wire signed [128:0] nl_z_out_4;
  reg [63:0] p_sva;
  reg [63:0] r_sva;
  reg [3:0] STAGE_LOOP_i_3_0_sva;
  reg [9:0] STAGE_LOOP_lshift_psp_sva;
  reg [63:0] modExp_result_sva;
  reg modExp_exp_1_7_1_sva;
  reg modExp_exp_1_6_1_sva;
  reg modExp_exp_1_5_1_sva;
  reg modExp_exp_1_4_1_sva;
  reg modExp_exp_1_3_1_sva;
  reg modExp_exp_1_2_1_sva;
  reg modExp_exp_1_1_1_sva;
  reg modExp_exp_1_0_1_sva_1;
  reg [63:0] COMP_LOOP_1_mul_mut;
  reg COMP_LOOP_COMP_LOOP_nor_1_itm;
  reg COMP_LOOP_COMP_LOOP_and_12_itm;
  reg [63:0] COMP_LOOP_1_acc_8_itm;
  reg COMP_LOOP_COMP_LOOP_nor_4_itm;
  reg COMP_LOOP_COMP_LOOP_and_30_itm;
  reg COMP_LOOP_COMP_LOOP_and_32_itm;
  reg COMP_LOOP_COMP_LOOP_and_33_itm;
  reg COMP_LOOP_COMP_LOOP_and_34_itm;
  reg COMP_LOOP_COMP_LOOP_and_86_itm;
  reg COMP_LOOP_COMP_LOOP_and_89_itm;
  reg COMP_LOOP_COMP_LOOP_and_124_itm;
  reg COMP_LOOP_COMP_LOOP_and_125_itm;
  wire STAGE_LOOP_i_3_0_sva_mx0c1;
  wire [3:0] STAGE_LOOP_i_3_0_sva_2;
  wire [4:0] nl_STAGE_LOOP_i_3_0_sva_2;
  wire [63:0] modulo_qr_sva_1_mx0w1;
  wire [64:0] nl_modulo_qr_sva_1_mx0w1;
  wire [63:0] COMP_LOOP_1_acc_5_mut_mx0w5;
  wire [64:0] nl_COMP_LOOP_1_acc_5_mut_mx0w5;
  wire [9:0] STAGE_LOOP_lshift_psp_sva_mx0w0;
  wire VEC_LOOP_j_sva_11_0_mx0c1;
  wire modExp_result_sva_mx0c0;
  wire [62:0] operator_64_false_slc_modExp_exp_63_1_3;
  wire modExp_while_and_3;
  wire modExp_while_and_5;
  wire COMP_LOOP_COMP_LOOP_and_211;
  wire COMP_LOOP_COMP_LOOP_and_213;
  wire COMP_LOOP_COMP_LOOP_and_215;
  wire and_243_m1c;
  wire modExp_result_and_rgt;
  wire modExp_result_and_1_rgt;
  wire COMP_LOOP_COMP_LOOP_and_11_cse;
  wire modExp_while_or_cse;
  wire COMP_LOOP_COMP_LOOP_and_12_cse;
  wire COMP_LOOP_COMP_LOOP_and_37_cse;
  wire COMP_LOOP_COMP_LOOP_and_13_cse;
  wire COMP_LOOP_or_2_cse;
  wire nor_473_cse;
  wire nor_461_cse;
  wire nor_447_cse;
  wire and_494_cse;
  wire operator_64_false_1_or_4_ssc;
  wire operator_64_false_1_or_5_ssc;
  wire and_511_cse;
  wire or_tmp_1365;
  wire mux_tmp;
  wire or_tmp_1367;
  wire nor_tmp_292;
  wire mux_tmp_1374;
  wire mux_tmp_1377;
  wire mux_tmp_1378;
  wire or_tmp_1370;
  wire nor_tmp_296;
  wire or_tmp_1374;
  wire mux_tmp_1399;
  wire or_tmp_1389;
  wire or_tmp_1394;
  wire nor_tmp_301;
  wire or_tmp_1401;
  wire [64:0] operator_64_false_mux1h_2_rgt;
  reg operator_64_false_acc_mut_64;
  reg [63:0] operator_64_false_acc_mut_63_0;
  wire or_136_cse;
  wire and_705_cse;
  wire COMP_LOOP_or_40_itm;
  wire operator_64_false_1_or_1_itm;
  wire STAGE_LOOP_acc_itm_2_1;
  wire or_1440_cse;

  wire[0:0] modulo_result_or_nl;
  wire[0:0] mux_782_nl;
  wire[0:0] and_388_nl;
  wire[0:0] mux_781_nl;
  wire[0:0] mux_780_nl;
  wire[0:0] or_864_nl;
  wire[0:0] or_862_nl;
  wire[0:0] nor_422_nl;
  wire[0:0] mux_779_nl;
  wire[0:0] mux_778_nl;
  wire[0:0] or_859_nl;
  wire[0:0] or_857_nl;
  wire[0:0] mux_777_nl;
  wire[0:0] or_855_nl;
  wire[0:0] mux_728_nl;
  wire[0:0] mux_727_nl;
  wire[0:0] mux_726_nl;
  wire[0:0] mux_725_nl;
  wire[0:0] mux_724_nl;
  wire[0:0] mux_723_nl;
  wire[0:0] mux_721_nl;
  wire[0:0] mux_720_nl;
  wire[0:0] mux_717_nl;
  wire[0:0] mux_716_nl;
  wire[0:0] mux_715_nl;
  wire[0:0] mux_714_nl;
  wire[0:0] mux_713_nl;
  wire[0:0] nand_41_nl;
  wire[0:0] mux_712_nl;
  wire[0:0] mux_711_nl;
  wire[0:0] mux_710_nl;
  wire[0:0] mux_709_nl;
  wire[0:0] mux_708_nl;
  wire[0:0] mux_707_nl;
  wire[0:0] mux_706_nl;
  wire[0:0] mux_704_nl;
  wire[0:0] mux_703_nl;
  wire[0:0] mux_702_nl;
  wire[0:0] mux_701_nl;
  wire[0:0] mux_700_nl;
  wire[0:0] mux_699_nl;
  wire[0:0] mux_698_nl;
  wire[0:0] mux_697_nl;
  wire[0:0] mux_695_nl;
  wire[0:0] mux_694_nl;
  wire[0:0] mux_693_nl;
  wire[0:0] mux_692_nl;
  wire[0:0] mux_691_nl;
  wire[0:0] or_819_nl;
  wire[0:0] mux_690_nl;
  wire[0:0] mux_687_nl;
  wire[0:0] mux_686_nl;
  wire[0:0] mux_685_nl;
  wire[0:0] mux_684_nl;
  wire[0:0] mux_683_nl;
  wire[0:0] nand_40_nl;
  wire[0:0] mux_682_nl;
  wire[0:0] nand_39_nl;
  wire[0:0] or_815_nl;
  wire[0:0] or_813_nl;
  wire[0:0] mux_681_nl;
  wire[0:0] mux_680_nl;
  wire[0:0] mux_679_nl;
  wire[0:0] mux_678_nl;
  wire[0:0] or_808_nl;
  wire[0:0] mux_775_nl;
  wire[0:0] mux_774_nl;
  wire[0:0] mux_773_nl;
  wire[0:0] mux_772_nl;
  wire[0:0] mux_771_nl;
  wire[0:0] mux_770_nl;
  wire[0:0] nand_130_nl;
  wire[0:0] mux_769_nl;
  wire[0:0] nand_44_nl;
  wire[0:0] mux_768_nl;
  wire[0:0] mux_767_nl;
  wire[0:0] nor_423_nl;
  wire[0:0] mux_766_nl;
  wire[0:0] mux_765_nl;
  wire[0:0] mux_764_nl;
  wire[0:0] or_850_nl;
  wire[0:0] mux_763_nl;
  wire[0:0] nor_424_nl;
  wire[0:0] mux_762_nl;
  wire[0:0] mux_761_nl;
  wire[0:0] and_167_nl;
  wire[0:0] mux_760_nl;
  wire[0:0] mux_759_nl;
  wire[0:0] mux_758_nl;
  wire[0:0] mux_757_nl;
  wire[0:0] mux_756_nl;
  wire[0:0] nand_249_nl;
  wire[0:0] or_848_nl;
  wire[0:0] mux_755_nl;
  wire[0:0] mux_754_nl;
  wire[0:0] mux_753_nl;
  wire[0:0] mux_752_nl;
  wire[0:0] mux_751_nl;
  wire[0:0] mux_750_nl;
  wire[0:0] or_847_nl;
  wire[0:0] mux_749_nl;
  wire[0:0] nand_43_nl;
  wire[0:0] mux_748_nl;
  wire[0:0] or_845_nl;
  wire[0:0] mux_747_nl;
  wire[0:0] mux_746_nl;
  wire[0:0] mux_745_nl;
  wire[0:0] mux_744_nl;
  wire[0:0] mux_743_nl;
  wire[0:0] or_843_nl;
  wire[0:0] mux_742_nl;
  wire[0:0] mux_741_nl;
  wire[0:0] or_842_nl;
  wire[0:0] mux_740_nl;
  wire[0:0] and_165_nl;
  wire[0:0] mux_739_nl;
  wire[0:0] mux_738_nl;
  wire[0:0] mux_737_nl;
  wire[0:0] nor_426_nl;
  wire[0:0] mux_736_nl;
  wire[0:0] mux_735_nl;
  wire[0:0] nor_427_nl;
  wire[0:0] mux_734_nl;
  wire[0:0] mux_733_nl;
  wire[0:0] mux_732_nl;
  wire[0:0] mux_730_nl;
  wire[0:0] mux_729_nl;
  wire[0:0] nor_428_nl;
  wire[0:0] nor_429_nl;
  wire[0:0] nor_430_nl;
  wire[0:0] mux_795_nl;
  wire[0:0] mux_794_nl;
  wire[0:0] mux_793_nl;
  wire[0:0] nor_411_nl;
  wire[0:0] mux_792_nl;
  wire[0:0] and_380_nl;
  wire[0:0] nor_412_nl;
  wire[0:0] mux_791_nl;
  wire[0:0] nor_414_nl;
  wire[0:0] mux_790_nl;
  wire[0:0] and_381_nl;
  wire[0:0] or_881_nl;
  wire[0:0] nor_415_nl;
  wire[0:0] mux_789_nl;
  wire[0:0] and_383_nl;
  wire[0:0] or_877_nl;
  wire[0:0] mux_788_nl;
  wire[0:0] nor_416_nl;
  wire[0:0] mux_787_nl;
  wire[0:0] nand_47_nl;
  wire[0:0] mux_786_nl;
  wire[0:0] nand_127_nl;
  wire[0:0] or_872_nl;
  wire[0:0] mux_785_nl;
  wire[0:0] mux_784_nl;
  wire[0:0] nor_417_nl;
  wire[0:0] nor_418_nl;
  wire[0:0] mux_783_nl;
  wire[0:0] nor_419_nl;
  wire[0:0] and_386_nl;
  wire[0:0] nor_659_nl;
  wire[0:0] and_704_nl;
  wire[0:0] mux_812_nl;
  wire[0:0] and_176_nl;
  wire[63:0] modExp_while_if_mux1h_nl;
  wire[0:0] modExp_while_if_or_nl;
  wire[0:0] mux_1122_nl;
  wire[0:0] mux_1121_nl;
  wire[0:0] nor_340_nl;
  wire[0:0] mux_1120_nl;
  wire[0:0] or_1113_nl;
  wire[0:0] mux_1119_nl;
  wire[0:0] or_1111_nl;
  wire[0:0] or_1109_nl;
  wire[0:0] mux_1118_nl;
  wire[0:0] nor_341_nl;
  wire[0:0] and_324_nl;
  wire[0:0] mux_1117_nl;
  wire[0:0] nor_342_nl;
  wire[0:0] and_492_nl;
  wire[0:0] and_325_nl;
  wire[0:0] mux_1116_nl;
  wire[0:0] nor_344_nl;
  wire[0:0] nor_345_nl;
  wire[0:0] modExp_while_if_and_1_nl;
  wire[0:0] modExp_while_if_and_2_nl;
  wire[0:0] and_179_nl;
  wire[0:0] mux_856_nl;
  wire[0:0] mux_855_nl;
  wire[0:0] mux_854_nl;
  wire[0:0] mux_853_nl;
  wire[0:0] mux_852_nl;
  wire[0:0] mux_851_nl;
  wire[0:0] mux_850_nl;
  wire[0:0] mux_849_nl;
  wire[0:0] mux_848_nl;
  wire[0:0] mux_847_nl;
  wire[0:0] or_1388_nl;
  wire[0:0] mux_846_nl;
  wire[0:0] mux_844_nl;
  wire[0:0] or_928_nl;
  wire[0:0] mux_843_nl;
  wire[0:0] mux_842_nl;
  wire[0:0] mux_841_nl;
  wire[0:0] mux_840_nl;
  wire[0:0] and_372_nl;
  wire[0:0] mux_839_nl;
  wire[0:0] mux_838_nl;
  wire[0:0] and_373_nl;
  wire[0:0] nor_397_nl;
  wire[0:0] mux_836_nl;
  wire[0:0] mux_835_nl;
  wire[0:0] or_925_nl;
  wire[0:0] mux_834_nl;
  wire[0:0] mux_833_nl;
  wire[0:0] mux_832_nl;
  wire[0:0] mux_831_nl;
  wire[0:0] mux_830_nl;
  wire[0:0] mux_829_nl;
  wire[0:0] mux_828_nl;
  wire[0:0] mux_826_nl;
  wire[0:0] mux_825_nl;
  wire[0:0] mux_824_nl;
  wire[0:0] mux_823_nl;
  wire[0:0] mux_822_nl;
  wire[0:0] mux_821_nl;
  wire[0:0] mux_820_nl;
  wire[0:0] mux_819_nl;
  wire[0:0] mux_818_nl;
  wire[0:0] or_924_nl;
  wire[0:0] mux_817_nl;
  wire[0:0] mux_816_nl;
  wire[0:0] and_376_nl;
  wire[0:0] or_923_nl;
  wire[0:0] mux_815_nl;
  wire[0:0] mux_1423_nl;
  wire[0:0] mux_1422_nl;
  wire[0:0] mux_1421_nl;
  wire[0:0] mux_1420_nl;
  wire[0:0] mux_1419_nl;
  wire[0:0] or_1550_nl;
  wire[0:0] mux_1418_nl;
  wire[0:0] or_1499_nl;
  wire[0:0] mux_1417_nl;
  wire[0:0] mux_1416_nl;
  wire[0:0] mux_1415_nl;
  wire[0:0] and_707_nl;
  wire[0:0] mux_1414_nl;
  wire[0:0] mux_1413_nl;
  wire[0:0] and_706_nl;
  wire[0:0] or_1497_nl;
  wire[0:0] mux_1412_nl;
  wire[0:0] mux_1411_nl;
  wire[0:0] mux_1410_nl;
  wire[0:0] mux_1409_nl;
  wire[0:0] mux_1408_nl;
  wire[0:0] mux_1407_nl;
  wire[0:0] mux_1406_nl;
  wire[0:0] mux_1405_nl;
  wire[0:0] mux_1404_nl;
  wire[0:0] mux_1403_nl;
  wire[0:0] mux_1402_nl;
  wire[0:0] mux_1401_nl;
  wire[0:0] mux_1399_nl;
  wire[0:0] mux_1398_nl;
  wire[0:0] mux_1397_nl;
  wire[0:0] mux_1396_nl;
  wire[0:0] mux_1395_nl;
  wire[0:0] mux_1394_nl;
  wire[0:0] mux_1393_nl;
  wire[0:0] mux_1392_nl;
  wire[0:0] mux_1391_nl;
  wire[0:0] mux_1390_nl;
  wire[0:0] mux_1389_nl;
  wire[0:0] mux_1388_nl;
  wire[0:0] nand_275_nl;
  wire[0:0] mux_1387_nl;
  wire[0:0] mux_1386_nl;
  wire[0:0] mux_1385_nl;
  wire[0:0] nand_276_nl;
  wire[0:0] and_717_nl;
  wire[0:0] mux_1384_nl;
  wire[0:0] mux_1383_nl;
  wire[0:0] mux_1382_nl;
  wire[0:0] mux_1381_nl;
  wire[0:0] mux_1380_nl;
  wire[0:0] mux_1377_nl;
  wire[0:0] or_1489_nl;
  wire[0:0] mux_1376_nl;
  wire[0:0] mux_1374_nl;
  wire[0:0] and_718_nl;
  wire[0:0] or_1487_nl;
  wire[0:0] mux_1373_nl;
  wire[0:0] nand_266_nl;
  wire[0:0] or_1485_nl;
  wire[0:0] mux_1453_nl;
  wire[0:0] mux_1452_nl;
  wire[0:0] and_710_nl;
  wire[0:0] mux_1451_nl;
  wire[0:0] or_1540_nl;
  wire[0:0] mux_1450_nl;
  wire[0:0] or_1539_nl;
  wire[0:0] mux_1449_nl;
  wire[0:0] mux_1448_nl;
  wire[0:0] or_1537_nl;
  wire[0:0] nor_676_nl;
  wire[0:0] mux_1447_nl;
  wire[0:0] mux_1446_nl;
  wire[0:0] or_1535_nl;
  wire[0:0] or_1534_nl;
  wire[0:0] or_1533_nl;
  wire[0:0] mux_1445_nl;
  wire[0:0] mux_1444_nl;
  wire[0:0] mux_1443_nl;
  wire[0:0] mux_1442_nl;
  wire[0:0] mux_1441_nl;
  wire[0:0] nor_677_nl;
  wire[0:0] nor_678_nl;
  wire[0:0] and_711_nl;
  wire[0:0] nor_679_nl;
  wire[0:0] nor_680_nl;
  wire[0:0] mux_1440_nl;
  wire[0:0] mux_1439_nl;
  wire[0:0] nor_681_nl;
  wire[0:0] nor_682_nl;
  wire[0:0] nor_683_nl;
  wire[0:0] mux_1438_nl;
  wire[0:0] or_1524_nl;
  wire[0:0] mux_1437_nl;
  wire[0:0] mux_1436_nl;
  wire[0:0] mux_1435_nl;
  wire[0:0] nor_684_nl;
  wire[0:0] mux_1434_nl;
  wire[0:0] mux_1433_nl;
  wire[0:0] nor_685_nl;
  wire[0:0] and_712_nl;
  wire[0:0] mux_1432_nl;
  wire[0:0] mux_1431_nl;
  wire[0:0] mux_1430_nl;
  wire[0:0] or_1516_nl;
  wire[0:0] or_1513_nl;
  wire[0:0] mux_1429_nl;
  wire[0:0] and_713_nl;
  wire[0:0] mux_1428_nl;
  wire[0:0] or_1512_nl;
  wire[0:0] mux_1427_nl;
  wire[0:0] nand_278_nl;
  wire[0:0] nor_686_nl;
  wire[0:0] mux_1426_nl;
  wire[0:0] mux_1425_nl;
  wire[0:0] nand_274_nl;
  wire[0:0] or_1505_nl;
  wire[0:0] or_1504_nl;
  wire[0:0] mux_1424_nl;
  wire[0:0] or_1503_nl;
  wire[0:0] or_1501_nl;
  wire[0:0] nand_263_nl;
  wire[0:0] mux_865_nl;
  wire[0:0] nor_630_nl;
  wire[0:0] mux_864_nl;
  wire[0:0] or_940_nl;
  wire[0:0] nor_631_nl;
  wire[0:0] mux_1457_nl;
  wire[0:0] or_1549_nl;
  wire[0:0] mux_1456_nl;
  wire[0:0] or_1547_nl;
  wire[0:0] or_1545_nl;
  wire[0:0] nand_271_nl;
  wire[0:0] mux_1455_nl;
  wire[0:0] nor_674_nl;
  wire[0:0] nor_675_nl;
  wire[0:0] mux_885_nl;
  wire[0:0] mux_884_nl;
  wire[0:0] mux_883_nl;
  wire[0:0] mux_882_nl;
  wire[0:0] nor_389_nl;
  wire[0:0] nor_390_nl;
  wire[0:0] and_185_nl;
  wire[0:0] mux_881_nl;
  wire[0:0] and_360_nl;
  wire[0:0] mux_880_nl;
  wire[0:0] and_184_nl;
  wire[0:0] mux_879_nl;
  wire[0:0] COMP_LOOP_or_15_nl;
  wire[0:0] COMP_LOOP_or_16_nl;
  wire[0:0] COMP_LOOP_or_17_nl;
  wire[0:0] COMP_LOOP_or_18_nl;
  wire[0:0] COMP_LOOP_or_19_nl;
  wire[0:0] COMP_LOOP_or_20_nl;
  wire[0:0] COMP_LOOP_or_21_nl;
  wire[0:0] COMP_LOOP_or_22_nl;
  wire[0:0] mux_913_nl;
  wire[0:0] mux_912_nl;
  wire[0:0] mux_911_nl;
  wire[0:0] mux_910_nl;
  wire[0:0] mux_909_nl;
  wire[0:0] or_964_nl;
  wire[0:0] mux_908_nl;
  wire[0:0] nand_120_nl;
  wire[0:0] mux_907_nl;
  wire[0:0] mux_906_nl;
  wire[0:0] mux_905_nl;
  wire[0:0] mux_904_nl;
  wire[0:0] mux_903_nl;
  wire[0:0] mux_902_nl;
  wire[0:0] mux_901_nl;
  wire[0:0] nand_121_nl;
  wire[0:0] and_192_nl;
  wire[0:0] mux_900_nl;
  wire[0:0] nand_122_nl;
  wire[0:0] mux_899_nl;
  wire[0:0] mux_898_nl;
  wire[0:0] mux_897_nl;
  wire[0:0] nor_388_nl;
  wire[0:0] or_959_nl;
  wire[0:0] mux_896_nl;
  wire[0:0] mux_895_nl;
  wire[0:0] mux_894_nl;
  wire[0:0] mux_893_nl;
  wire[0:0] mux_892_nl;
  wire[0:0] mux_891_nl;
  wire[0:0] mux_890_nl;
  wire[0:0] mux_889_nl;
  wire[0:0] or_958_nl;
  wire[0:0] mux_888_nl;
  wire[0:0] mux_887_nl;
  wire[0:0] mux_34_nl;
  wire[0:0] mux_33_nl;
  wire[0:0] or_42_nl;
  wire[0:0] or_41_nl;
  wire[0:0] or_39_nl;
  wire[0:0] nor_604_nl;
  wire[0:0] nor_605_nl;
  wire[0:0] mux_915_nl;
  wire[0:0] nor_386_nl;
  wire[0:0] nor_387_nl;
  wire[0:0] and_238_nl;
  wire[0:0] COMP_LOOP_or_26_nl;
  wire[0:0] COMP_LOOP_or_27_nl;
  wire[0:0] COMP_LOOP_or_7_nl;
  wire[0:0] COMP_LOOP_or_8_nl;
  wire[0:0] COMP_LOOP_or_9_nl;
  wire[0:0] COMP_LOOP_or_10_nl;
  wire[0:0] COMP_LOOP_or_11_nl;
  wire[0:0] COMP_LOOP_or_12_nl;
  wire[0:0] COMP_LOOP_or_13_nl;
  wire[0:0] COMP_LOOP_or_14_nl;
  wire[0:0] mux_48_nl;
  wire[0:0] and_470_nl;
  wire[0:0] mux_47_nl;
  wire[0:0] mux_46_nl;
  wire[0:0] nor_591_nl;
  wire[0:0] nor_592_nl;
  wire[0:0] mux_45_nl;
  wire[0:0] nor_593_nl;
  wire[0:0] nor_594_nl;
  wire[0:0] nor_595_nl;
  wire[0:0] mux_44_nl;
  wire[0:0] or_62_nl;
  wire[0:0] mux_43_nl;
  wire[0:0] or_61_nl;
  wire[0:0] or_59_nl;
  wire[0:0] mux_42_nl;
  wire[0:0] nand_224_nl;
  wire[0:0] or_56_nl;
  wire[0:0] mux_971_nl;
  wire[0:0] mux_970_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] mux_348_nl;
  wire[0:0] mux_347_nl;
  wire[0:0] or_248_nl;
  wire[0:0] nand_9_nl;
  wire[0:0] mux_346_nl;
  wire[0:0] mux_965_nl;
  wire[0:0] mux_964_nl;
  wire[0:0] mux_963_nl;
  wire[0:0] nor_371_nl;
  wire[0:0] or_246_nl;
  wire[0:0] mux_343_nl;
  wire[0:0] mux_341_nl;
  wire[0:0] mux_960_nl;
  wire[0:0] nand_56_nl;
  wire[0:0] mux_959_nl;
  wire[0:0] or_1009_nl;
  wire[0:0] mux_958_nl;
  wire[0:0] mux_957_nl;
  wire[0:0] mux_956_nl;
  wire[0:0] mux_955_nl;
  wire[0:0] and_246_nl;
  wire[0:0] mux_954_nl;
  wire[0:0] nor_190_nl;
  wire[0:0] mux_333_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] mux_951_nl;
  wire[0:0] mux_950_nl;
  wire[0:0] nor_372_nl;
  wire[0:0] mux_328_nl;
  wire[0:0] mux_948_nl;
  wire[0:0] nor_560_nl;
  wire[0:0] mux_947_nl;
  wire[0:0] mux_334_nl;
  wire[0:0] or_1003_nl;
  wire[0:0] mux_945_nl;
  wire[0:0] mux_944_nl;
  wire[0:0] mux_943_nl;
  wire[0:0] mux_942_nl;
  wire[0:0] or_1002_nl;
  wire[0:0] mux_941_nl;
  wire[0:0] mux_940_nl;
  wire[0:0] or_999_nl;
  wire[0:0] mux_939_nl;
  wire[0:0] mux_938_nl;
  wire[0:0] mux_937_nl;
  wire[0:0] mux_936_nl;
  wire[0:0] or_1383_nl;
  wire[0:0] mux_935_nl;
  wire[0:0] mux_934_nl;
  wire[0:0] nand_117_nl;
  wire[0:0] mux_933_nl;
  wire[0:0] or_996_nl;
  wire[0:0] or_994_nl;
  wire[0:0] mux_932_nl;
  wire[0:0] or_231_nl;
  wire[0:0] mux_313_nl;
  wire[0:0] or_992_nl;
  wire[0:0] mux_930_nl;
  wire[0:0] COMP_LOOP_mux1h_31_nl;
  wire[7:0] COMP_LOOP_acc_12_nl;
  wire[8:0] nl_COMP_LOOP_acc_12_nl;
  wire[0:0] COMP_LOOP_and_76_nl;
  wire[0:0] mux_1032_nl;
  wire[0:0] mux_1031_nl;
  wire[0:0] mux_1030_nl;
  wire[0:0] mux_1029_nl;
  wire[0:0] mux_1028_nl;
  wire[0:0] mux_1027_nl;
  wire[0:0] mux_1026_nl;
  wire[0:0] mux_1025_nl;
  wire[0:0] nor_205_nl;
  wire[0:0] mux_1024_nl;
  wire[0:0] mux_1023_nl;
  wire[0:0] mux_1022_nl;
  wire[0:0] or_1072_nl;
  wire[0:0] mux_1021_nl;
  wire[0:0] mux_1020_nl;
  wire[0:0] mux_1019_nl;
  wire[0:0] and_252_nl;
  wire[0:0] mux_1018_nl;
  wire[0:0] mux_1017_nl;
  wire[0:0] mux_1016_nl;
  wire[0:0] mux_1015_nl;
  wire[0:0] and_340_nl;
  wire[0:0] nor_351_nl;
  wire[0:0] nor_352_nl;
  wire[0:0] mux_1014_nl;
  wire[0:0] mux_1013_nl;
  wire[0:0] and_251_nl;
  wire[0:0] mux_1012_nl;
  wire[0:0] mux_1011_nl;
  wire[0:0] mux_1010_nl;
  wire[0:0] mux_1009_nl;
  wire[0:0] mux_1008_nl;
  wire[0:0] mux_1007_nl;
  wire[0:0] mux_1005_nl;
  wire[0:0] mux_1004_nl;
  wire[0:0] mux_1003_nl;
  wire[0:0] mux_1002_nl;
  wire[0:0] or_1061_nl;
  wire[0:0] mux_1001_nl;
  wire[0:0] mux_1000_nl;
  wire[0:0] mux_999_nl;
  wire[0:0] or_1059_nl;
  wire[0:0] mux_998_nl;
  wire[0:0] mux_996_nl;
  wire[0:0] nor_353_nl;
  wire[0:0] nor_354_nl;
  wire[0:0] mux_995_nl;
  wire[0:0] mux_987_nl;
  wire[0:0] or_1432_nl;
  wire[0:0] or_1433_nl;
  wire[0:0] mux_986_nl;
  wire[0:0] mux_985_nl;
  wire[0:0] or_1040_nl;
  wire[0:0] or_1039_nl;
  wire[0:0] or_1037_nl;
  wire[0:0] mux_1035_nl;
  wire[0:0] nor_347_nl;
  wire[0:0] mux_1034_nl;
  wire[0:0] nand_108_nl;
  wire[0:0] or_1082_nl;
  wire[0:0] nor_348_nl;
  wire[0:0] mux_1033_nl;
  wire[0:0] or_1078_nl;
  wire[0:0] or_1077_nl;
  wire[63:0] COMP_LOOP_1_acc_8_nl;
  wire[64:0] nl_COMP_LOOP_1_acc_8_nl;
  wire[0:0] mux_1139_nl;
  wire[0:0] mux_1138_nl;
  wire[0:0] nor_334_nl;
  wire[0:0] mux_1137_nl;
  wire[0:0] or_1146_nl;
  wire[0:0] or_1145_nl;
  wire[0:0] mux_1136_nl;
  wire[0:0] nor_335_nl;
  wire[0:0] mux_1135_nl;
  wire[0:0] or_1142_nl;
  wire[0:0] or_1141_nl;
  wire[0:0] and_321_nl;
  wire[0:0] mux_1134_nl;
  wire[0:0] nor_336_nl;
  wire[0:0] mux_1133_nl;
  wire[0:0] or_1137_nl;
  wire[0:0] or_1136_nl;
  wire[0:0] and_322_nl;
  wire[0:0] mux_1132_nl;
  wire[0:0] nor_337_nl;
  wire[0:0] nor_338_nl;
  wire[0:0] mux_1156_nl;
  wire[0:0] mux_1155_nl;
  wire[0:0] nand_98_nl;
  wire[0:0] nand_99_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_145_nl;
  wire[9:0] COMP_LOOP_1_acc_nl;
  wire[10:0] nl_COMP_LOOP_1_acc_nl;
  wire[0:0] mux_1174_nl;
  wire[0:0] mux_1173_nl;
  wire[0:0] mux_1172_nl;
  wire[0:0] mux_1171_nl;
  wire[0:0] mux_1169_nl;
  wire[0:0] mux_1168_nl;
  wire[0:0] mux_1167_nl;
  wire[0:0] mux_1166_nl;
  wire[0:0] mux_1165_nl;
  wire[0:0] mux_1163_nl;
  wire[0:0] and_315_nl;
  wire[0:0] mux_1181_nl;
  wire[0:0] mux_1180_nl;
  wire[0:0] mux_1179_nl;
  wire[0:0] mux_1177_nl;
  wire[0:0] and_313_nl;
  wire[0:0] mux_1176_nl;
  wire[0:0] mux_1184_nl;
  wire[0:0] nand_234_nl;
  wire[0:0] mux_1183_nl;
  wire[0:0] or_1193_nl;
  wire[0:0] mux_1186_nl;
  wire[0:0] nor_328_nl;
  wire[0:0] mux_1185_nl;
  wire[0:0] and_272_nl;
  wire[0:0] and_271_nl;
  wire[0:0] or_1200_nl;
  wire[0:0] mux_1187_nl;
  wire[0:0] or_100_nl;
  wire[0:0] or_1197_nl;
  wire[0:0] or_1201_nl;
  wire[0:0] mux_1192_nl;
  wire[0:0] mux_1191_nl;
  wire[0:0] nor_327_nl;
  wire[0:0] mux_1190_nl;
  wire[0:0] and_274_nl;
  wire[0:0] COMP_LOOP_mux_nl;
  wire[0:0] mux_1246_nl;
  wire[0:0] mux_1245_nl;
  wire[0:0] and_306_nl;
  wire[0:0] mux_1244_nl;
  wire[0:0] mux_1243_nl;
  wire[0:0] nor_316_nl;
  wire[0:0] nor_317_nl;
  wire[0:0] nor_318_nl;
  wire[0:0] nor_319_nl;
  wire[0:0] mux_1242_nl;
  wire[0:0] and_307_nl;
  wire[0:0] mux_1241_nl;
  wire[0:0] nor_320_nl;
  wire[0:0] and_493_nl;
  wire[0:0] nor_322_nl;
  wire[0:0] mux_1240_nl;
  wire[0:0] or_1229_nl;
  wire[0:0] nand_95_nl;
  wire[0:0] mux_1196_nl;
  wire[0:0] nor_324_nl;
  wire[0:0] mux_1195_nl;
  wire[0:0] or_1210_nl;
  wire[0:0] nor_325_nl;
  wire[0:0] mux_1194_nl;
  wire[0:0] or_1208_nl;
  wire[0:0] mux_1249_nl;
  wire[0:0] or_1430_nl;
  wire[0:0] or_1431_nl;
  wire[0:0] mux_1248_nl;
  wire[0:0] or_1245_nl;
  wire[0:0] mux_1247_nl;
  wire[0:0] or_1244_nl;
  wire[0:0] or_1243_nl;
  wire[0:0] COMP_LOOP_mux1h_52_nl;
  wire[0:0] mux_1285_nl;
  wire[0:0] mux_1284_nl;
  wire[0:0] nand_259_nl;
  wire[0:0] mux_1283_nl;
  wire[0:0] nor_304_nl;
  wire[0:0] nor_305_nl;
  wire[0:0] nand_260_nl;
  wire[0:0] mux_1282_nl;
  wire[0:0] nand_261_nl;
  wire[0:0] mux_1281_nl;
  wire[0:0] nor_306_nl;
  wire[0:0] nor_307_nl;
  wire[0:0] mux_1280_nl;
  wire[0:0] or_1283_nl;
  wire[0:0] nand_226_nl;
  wire[0:0] or_1483_nl;
  wire[0:0] COMP_LOOP_mux1h_66_nl;
  wire[0:0] COMP_LOOP_mux1h_68_nl;
  wire[0:0] mux_1320_nl;
  wire[0:0] mux_1319_nl;
  wire[0:0] mux_1318_nl;
  wire[0:0] mux_1317_nl;
  wire[0:0] nand_86_nl;
  wire[0:0] or_1323_nl;
  wire[0:0] mux_1316_nl;
  wire[0:0] mux_1315_nl;
  wire[0:0] mux_1314_nl;
  wire[0:0] nand_247_nl;
  wire[0:0] or_1366_nl;
  wire[0:0] or_1367_nl;
  wire[0:0] mux_1313_nl;
  wire[0:0] mux_1312_nl;
  wire[0:0] or_1316_nl;
  wire[0:0] mux_1311_nl;
  wire[0:0] mux_1310_nl;
  wire[0:0] mux_1309_nl;
  wire[0:0] mux_1308_nl;
  wire[0:0] mux_1307_nl;
  wire[0:0] mux_1306_nl;
  wire[0:0] or_1314_nl;
  wire[0:0] mux_1304_nl;
  wire[0:0] mux_1303_nl;
  wire[0:0] mux_1302_nl;
  wire[0:0] mux_1301_nl;
  wire[0:0] mux_1300_nl;
  wire[0:0] mux_1299_nl;
  wire[0:0] mux_1298_nl;
  wire[0:0] mux_1297_nl;
  wire[0:0] mux_1296_nl;
  wire[0:0] mux_1295_nl;
  wire[0:0] or_1311_nl;
  wire[0:0] mux_1294_nl;
  wire[0:0] mux_1293_nl;
  wire[0:0] or_1309_nl;
  wire[0:0] or_1307_nl;
  wire[0:0] mux_1323_nl;
  wire[0:0] or_1434_nl;
  wire[0:0] or_1435_nl;
  wire[0:0] mux_1322_nl;
  wire[0:0] or_1329_nl;
  wire[0:0] mux_1321_nl;
  wire[0:0] or_1328_nl;
  wire[0:0] or_1326_nl;
  wire[0:0] mux_1326_nl;
  wire[0:0] and_282_nl;
  wire[0:0] mux_1325_nl;
  wire[0:0] nor_292_nl;
  wire[0:0] mux_1324_nl;
  wire[0:0] nor_293_nl;
  wire[0:0] and_283_nl;
  wire[0:0] nor_294_nl;
  wire[0:0] nor_295_nl;
  wire[0:0] or_1402_nl;
  wire[0:0] nand_199_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] and_432_nl;
  wire[0:0] mux_381_nl;
  wire[0:0] or_308_nl;
  wire[0:0] or_306_nl;
  wire[0:0] or_325_nl;
  wire[0:0] or_323_nl;
  wire[0:0] mux_418_nl;
  wire[0:0] or_375_nl;
  wire[0:0] or_373_nl;
  wire[0:0] mux_456_nl;
  wire[0:0] nor_512_nl;
  wire[0:0] nor_513_nl;
  wire[0:0] mux_494_nl;
  wire[0:0] nor_496_nl;
  wire[0:0] nor_497_nl;
  wire[0:0] mux_538_nl;
  wire[0:0] or_570_nl;
  wire[0:0] or_568_nl;
  wire[0:0] mux_575_nl;
  wire[0:0] or_635_nl;
  wire[0:0] or_633_nl;
  wire[0:0] mux_612_nl;
  wire[0:0] nor_458_nl;
  wire[0:0] nor_459_nl;
  wire[0:0] mux_649_nl;
  wire[0:0] nor_444_nl;
  wire[0:0] nor_445_nl;
  wire[0:0] or_854_nl;
  wire[0:0] or_853_nl;
  wire[0:0] nor_405_nl;
  wire[0:0] mux_801_nl;
  wire[0:0] mux_800_nl;
  wire[0:0] or_903_nl;
  wire[0:0] or_902_nl;
  wire[0:0] nand_49_nl;
  wire[0:0] mux_799_nl;
  wire[0:0] and_489_nl;
  wire[0:0] nor_407_nl;
  wire[0:0] mux_798_nl;
  wire[0:0] nor_408_nl;
  wire[0:0] mux_797_nl;
  wire[0:0] nor_409_nl;
  wire[0:0] mux_796_nl;
  wire[0:0] or_895_nl;
  wire[0:0] or_893_nl;
  wire[0:0] nor_410_nl;
  wire[0:0] mux_807_nl;
  wire[0:0] nor_400_nl;
  wire[0:0] mux_806_nl;
  wire[0:0] or_1362_nl;
  wire[0:0] or_913_nl;
  wire[0:0] mux_805_nl;
  wire[0:0] nor_401_nl;
  wire[0:0] and_377_nl;
  wire[0:0] mux_804_nl;
  wire[0:0] nor_402_nl;
  wire[0:0] and_378_nl;
  wire[0:0] mux_803_nl;
  wire[0:0] nor_403_nl;
  wire[0:0] nor_404_nl;
  wire[0:0] mux_811_nl;
  wire[0:0] mux_810_nl;
  wire[0:0] mux_809_nl;
  wire[0:0] or_916_nl;
  wire[0:0] mux_814_nl;
  wire[0:0] nor_398_nl;
  wire[0:0] nor_399_nl;
  wire[0:0] or_955_nl;
  wire[0:0] mux_919_nl;
  wire[0:0] mux_918_nl;
  wire[0:0] nor_382_nl;
  wire[0:0] and_474_nl;
  wire[0:0] mux_30_nl;
  wire[0:0] nor_603_nl;
  wire[0:0] and_475_nl;
  wire[0:0] mux_977_nl;
  wire[0:0] nor_366_nl;
  wire[0:0] mux_976_nl;
  wire[0:0] or_1026_nl;
  wire[0:0] or_1024_nl;
  wire[0:0] nor_367_nl;
  wire[0:0] mux_975_nl;
  wire[0:0] and_350_nl;
  wire[0:0] mux_974_nl;
  wire[0:0] nor_368_nl;
  wire[0:0] mux_973_nl;
  wire[0:0] and_351_nl;
  wire[0:0] nor_369_nl;
  wire[0:0] nor_370_nl;
  wire[0:0] mux_993_nl;
  wire[0:0] mux_992_nl;
  wire[0:0] and_344_nl;
  wire[0:0] mux_991_nl;
  wire[0:0] and_345_nl;
  wire[0:0] nor_355_nl;
  wire[0:0] nor_356_nl;
  wire[0:0] mux_990_nl;
  wire[0:0] and_346_nl;
  wire[0:0] mux_989_nl;
  wire[0:0] nor_358_nl;
  wire[0:0] mux_988_nl;
  wire[0:0] nand_111_nl;
  wire[0:0] or_1045_nl;
  wire[0:0] or_1183_nl;
  wire[0:0] mux_1157_nl;
  wire[0:0] and_320_nl;
  wire[0:0] and_263_nl;
  wire[0:0] mux_1161_nl;
  wire[0:0] nor_329_nl;
  wire[0:0] mux_1272_nl;
  wire[0:0] mux_1271_nl;
  wire[0:0] mux_1270_nl;
  wire[0:0] mux_1269_nl;
  wire[0:0] mux_1268_nl;
  wire[0:0] or_1268_nl;
  wire[0:0] mux_1267_nl;
  wire[0:0] or_1267_nl;
  wire[0:0] mux_1266_nl;
  wire[0:0] mux_1265_nl;
  wire[0:0] mux_1264_nl;
  wire[0:0] mux_1263_nl;
  wire[0:0] or_1263_nl;
  wire[0:0] mux_1262_nl;
  wire[0:0] mux_1261_nl;
  wire[0:0] mux_1260_nl;
  wire[0:0] mux_1259_nl;
  wire[0:0] mux_1258_nl;
  wire[0:0] mux_1257_nl;
  wire[0:0] nand_227_nl;
  wire[0:0] or_1258_nl;
  wire[0:0] mux_1256_nl;
  wire[0:0] or_1256_nl;
  wire[0:0] mux_1255_nl;
  wire[0:0] mux_1254_nl;
  wire[0:0] or_1254_nl;
  wire[0:0] mux_1253_nl;
  wire[0:0] mux_1252_nl;
  wire[0:0] mux_1250_nl;
  wire[0:0] or_1249_nl;
  wire[0:0] mux_1276_nl;
  wire[0:0] and_294_nl;
  wire[0:0] mux_1275_nl;
  wire[0:0] nor_310_nl;
  wire[0:0] and_295_nl;
  wire[0:0] mux_1291_nl;
  wire[0:0] mux_1290_nl;
  wire[0:0] nor_300_nl;
  wire[0:0] mux_1289_nl;
  wire[0:0] or_1304_nl;
  wire[0:0] or_1303_nl;
  wire[0:0] nor_628_nl;
  wire[0:0] and_289_nl;
  wire[0:0] mux_1288_nl;
  wire[0:0] nor_303_nl;
  wire[0:0] mux_1287_nl;
  wire[0:0] or_1295_nl;
  wire[0:0] mux_1286_nl;
  wire[0:0] or_1093_nl;
  wire[0:0] or_1292_nl;
  wire[0:0] mux_877_nl;
  wire[0:0] mux_876_nl;
  wire[0:0] mux_875_nl;
  wire[0:0] mux_874_nl;
  wire[0:0] and_363_nl;
  wire[0:0] and_364_nl;
  wire[2:0] STAGE_LOOP_acc_nl;
  wire[3:0] nl_STAGE_LOOP_acc_nl;
  wire[0:0] nor_361_nl;
  wire[0:0] mux_983_nl;
  wire[0:0] mux_982_nl;
  wire[0:0] or_1381_nl;
  wire[0:0] or_1382_nl;
  wire[0:0] nand_113_nl;
  wire[0:0] mux_981_nl;
  wire[0:0] nor_362_nl;
  wire[0:0] and_348_nl;
  wire[0:0] and_349_nl;
  wire[0:0] mux_980_nl;
  wire[0:0] nor_363_nl;
  wire[0:0] mux_979_nl;
  wire[0:0] nor_364_nl;
  wire[0:0] nor_365_nl;
  wire[0:0] and_91_nl;
  wire[0:0] mux_370_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] mux_368_nl;
  wire[0:0] and_419_nl;
  wire[0:0] mux_367_nl;
  wire[0:0] nor_553_nl;
  wire[0:0] nor_554_nl;
  wire[0:0] nor_555_nl;
  wire[0:0] and_420_nl;
  wire[0:0] mux_366_nl;
  wire[0:0] and_421_nl;
  wire[0:0] nor_556_nl;
  wire[0:0] and_422_nl;
  wire[0:0] mux_365_nl;
  wire[0:0] nor_557_nl;
  wire[0:0] nor_558_nl;
  wire[0:0] mux_364_nl;
  wire[0:0] or_269_nl;
  wire[0:0] or_268_nl;
  wire[0:0] and_96_nl;
  wire[0:0] mux_371_nl;
  wire[0:0] nor_551_nl;
  wire[0:0] nor_552_nl;
  wire[0:0] and_104_nl;
  wire[0:0] mux_372_nl;
  wire[0:0] nor_549_nl;
  wire[0:0] nor_550_nl;
  wire[0:0] and_115_nl;
  wire[0:0] mux_373_nl;
  wire[0:0] nor_547_nl;
  wire[0:0] nor_548_nl;
  wire[0:0] and_123_nl;
  wire[0:0] mux_374_nl;
  wire[0:0] nor_545_nl;
  wire[0:0] nor_546_nl;
  wire[0:0] and_136_nl;
  wire[0:0] mux_375_nl;
  wire[0:0] nor_544_nl;
  wire[0:0] and_143_nl;
  wire[0:0] mux_376_nl;
  wire[0:0] nor_542_nl;
  wire[0:0] nor_543_nl;
  wire[0:0] and_152_nl;
  wire[0:0] mux_377_nl;
  wire[0:0] and_500_nl;
  wire[0:0] nor_541_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] mux_398_nl;
  wire[0:0] mux_397_nl;
  wire[0:0] mux_396_nl;
  wire[0:0] mux_395_nl;
  wire[0:0] or_331_nl;
  wire[0:0] mux_394_nl;
  wire[0:0] mux_393_nl;
  wire[0:0] or_326_nl;
  wire[0:0] mux_391_nl;
  wire[0:0] mux_390_nl;
  wire[0:0] mux_389_nl;
  wire[0:0] mux_388_nl;
  wire[0:0] or_321_nl;
  wire[0:0] mux_387_nl;
  wire[0:0] or_316_nl;
  wire[0:0] mux_386_nl;
  wire[0:0] mux_385_nl;
  wire[0:0] or_313_nl;
  wire[0:0] mux_384_nl;
  wire[0:0] mux_383_nl;
  wire[0:0] mux_382_nl;
  wire[0:0] or_311_nl;
  wire[0:0] or_305_nl;
  wire[0:0] mux_380_nl;
  wire[0:0] mux_379_nl;
  wire[0:0] mux_378_nl;
  wire[0:0] or_302_nl;
  wire[0:0] or_301_nl;
  wire[0:0] or_299_nl;
  wire[0:0] or_298_nl;
  wire[0:0] mux_413_nl;
  wire[0:0] nor_528_nl;
  wire[0:0] mux_412_nl;
  wire[0:0] nand_15_nl;
  wire[0:0] mux_411_nl;
  wire[0:0] nor_529_nl;
  wire[0:0] nor_530_nl;
  wire[0:0] or_359_nl;
  wire[0:0] mux_410_nl;
  wire[0:0] or_358_nl;
  wire[0:0] or_357_nl;
  wire[0:0] mux_409_nl;
  wire[0:0] and_417_nl;
  wire[0:0] mux_408_nl;
  wire[0:0] nor_531_nl;
  wire[0:0] nor_532_nl;
  wire[0:0] nor_533_nl;
  wire[0:0] mux_407_nl;
  wire[0:0] mux_406_nl;
  wire[0:0] mux_405_nl;
  wire[0:0] nor_534_nl;
  wire[0:0] nor_535_nl;
  wire[0:0] mux_404_nl;
  wire[0:0] or_347_nl;
  wire[0:0] or_345_nl;
  wire[0:0] nor_536_nl;
  wire[0:0] nor_537_nl;
  wire[0:0] mux_403_nl;
  wire[0:0] mux_402_nl;
  wire[0:0] or_340_nl;
  wire[0:0] mux_401_nl;
  wire[0:0] or_339_nl;
  wire[0:0] or_337_nl;
  wire[0:0] nand_13_nl;
  wire[0:0] mux_400_nl;
  wire[0:0] nor_538_nl;
  wire[0:0] nor_539_nl;
  wire[0:0] or_332_nl;
  wire[0:0] mux_436_nl;
  wire[0:0] mux_435_nl;
  wire[0:0] mux_434_nl;
  wire[0:0] mux_433_nl;
  wire[0:0] mux_432_nl;
  wire[0:0] or_398_nl;
  wire[0:0] mux_431_nl;
  wire[0:0] mux_430_nl;
  wire[0:0] or_393_nl;
  wire[0:0] mux_428_nl;
  wire[0:0] mux_427_nl;
  wire[0:0] mux_426_nl;
  wire[0:0] mux_425_nl;
  wire[0:0] or_388_nl;
  wire[0:0] mux_424_nl;
  wire[0:0] or_383_nl;
  wire[0:0] mux_423_nl;
  wire[0:0] mux_422_nl;
  wire[0:0] or_380_nl;
  wire[0:0] mux_421_nl;
  wire[0:0] mux_420_nl;
  wire[0:0] mux_419_nl;
  wire[0:0] or_378_nl;
  wire[0:0] or_372_nl;
  wire[0:0] mux_417_nl;
  wire[0:0] mux_416_nl;
  wire[0:0] mux_415_nl;
  wire[0:0] or_369_nl;
  wire[0:0] or_368_nl;
  wire[0:0] or_366_nl;
  wire[0:0] or_365_nl;
  wire[0:0] mux_451_nl;
  wire[0:0] mux_450_nl;
  wire[0:0] mux_449_nl;
  wire[0:0] nor_514_nl;
  wire[0:0] mux_448_nl;
  wire[0:0] or_423_nl;
  wire[0:0] or_421_nl;
  wire[0:0] nor_515_nl;
  wire[0:0] nor_516_nl;
  wire[0:0] mux_447_nl;
  wire[0:0] and_414_nl;
  wire[0:0] mux_446_nl;
  wire[0:0] nor_517_nl;
  wire[0:0] nor_518_nl;
  wire[0:0] nor_519_nl;
  wire[0:0] mux_445_nl;
  wire[0:0] or_411_nl;
  wire[0:0] or_410_nl;
  wire[0:0] mux_444_nl;
  wire[0:0] mux_443_nl;
  wire[0:0] nor_520_nl;
  wire[0:0] mux_442_nl;
  wire[0:0] nor_521_nl;
  wire[0:0] nor_522_nl;
  wire[0:0] mux_441_nl;
  wire[0:0] mux_440_nl;
  wire[0:0] mux_439_nl;
  wire[0:0] nor_523_nl;
  wire[0:0] nor_524_nl;
  wire[0:0] and_415_nl;
  wire[0:0] mux_438_nl;
  wire[0:0] mux_437_nl;
  wire[0:0] nor_525_nl;
  wire[0:0] nor_526_nl;
  wire[0:0] or_400_nl;
  wire[0:0] nor_527_nl;
  wire[0:0] mux_474_nl;
  wire[0:0] mux_473_nl;
  wire[0:0] mux_472_nl;
  wire[0:0] mux_471_nl;
  wire[0:0] mux_470_nl;
  wire[0:0] or_457_nl;
  wire[0:0] mux_469_nl;
  wire[0:0] mux_468_nl;
  wire[0:0] or_452_nl;
  wire[0:0] mux_466_nl;
  wire[0:0] mux_465_nl;
  wire[0:0] mux_464_nl;
  wire[0:0] mux_463_nl;
  wire[0:0] or_447_nl;
  wire[0:0] mux_462_nl;
  wire[0:0] or_442_nl;
  wire[0:0] mux_461_nl;
  wire[0:0] mux_460_nl;
  wire[0:0] or_439_nl;
  wire[0:0] mux_459_nl;
  wire[0:0] mux_458_nl;
  wire[0:0] mux_457_nl;
  wire[0:0] or_437_nl;
  wire[0:0] or_432_nl;
  wire[0:0] mux_455_nl;
  wire[0:0] mux_454_nl;
  wire[0:0] mux_453_nl;
  wire[0:0] or_429_nl;
  wire[0:0] or_428_nl;
  wire[0:0] or_426_nl;
  wire[0:0] or_425_nl;
  wire[0:0] mux_489_nl;
  wire[0:0] mux_488_nl;
  wire[0:0] mux_487_nl;
  wire[0:0] nor_498_nl;
  wire[0:0] mux_486_nl;
  wire[0:0] or_482_nl;
  wire[0:0] or_480_nl;
  wire[0:0] nor_499_nl;
  wire[0:0] nor_500_nl;
  wire[0:0] mux_485_nl;
  wire[0:0] and_411_nl;
  wire[0:0] mux_484_nl;
  wire[0:0] nor_501_nl;
  wire[0:0] nor_502_nl;
  wire[0:0] nor_503_nl;
  wire[0:0] mux_483_nl;
  wire[0:0] or_470_nl;
  wire[0:0] or_469_nl;
  wire[0:0] mux_482_nl;
  wire[0:0] mux_481_nl;
  wire[0:0] nor_504_nl;
  wire[0:0] mux_480_nl;
  wire[0:0] nor_505_nl;
  wire[0:0] nor_506_nl;
  wire[0:0] mux_479_nl;
  wire[0:0] mux_478_nl;
  wire[0:0] mux_477_nl;
  wire[0:0] nor_507_nl;
  wire[0:0] nor_508_nl;
  wire[0:0] and_412_nl;
  wire[0:0] mux_476_nl;
  wire[0:0] mux_475_nl;
  wire[0:0] nor_509_nl;
  wire[0:0] nor_510_nl;
  wire[0:0] or_459_nl;
  wire[0:0] nor_511_nl;
  wire[0:0] mux_512_nl;
  wire[0:0] mux_511_nl;
  wire[0:0] mux_510_nl;
  wire[0:0] mux_509_nl;
  wire[0:0] mux_508_nl;
  wire[0:0] or_516_nl;
  wire[0:0] mux_507_nl;
  wire[0:0] mux_506_nl;
  wire[0:0] or_511_nl;
  wire[0:0] mux_504_nl;
  wire[0:0] mux_503_nl;
  wire[0:0] mux_502_nl;
  wire[0:0] mux_501_nl;
  wire[0:0] or_506_nl;
  wire[0:0] mux_500_nl;
  wire[0:0] or_501_nl;
  wire[0:0] mux_499_nl;
  wire[0:0] mux_498_nl;
  wire[0:0] or_498_nl;
  wire[0:0] mux_497_nl;
  wire[0:0] mux_496_nl;
  wire[0:0] mux_495_nl;
  wire[0:0] or_496_nl;
  wire[0:0] or_491_nl;
  wire[0:0] mux_493_nl;
  wire[0:0] mux_492_nl;
  wire[0:0] mux_491_nl;
  wire[0:0] or_488_nl;
  wire[0:0] or_487_nl;
  wire[0:0] or_485_nl;
  wire[0:0] or_484_nl;
  wire[0:0] mux_526_nl;
  wire[0:0] nor_484_nl;
  wire[0:0] mux_525_nl;
  wire[0:0] nand_24_nl;
  wire[0:0] mux_524_nl;
  wire[0:0] nor_485_nl;
  wire[0:0] nor_486_nl;
  wire[0:0] or_544_nl;
  wire[0:0] mux_523_nl;
  wire[0:0] or_543_nl;
  wire[0:0] or_542_nl;
  wire[0:0] mux_522_nl;
  wire[0:0] and_410_nl;
  wire[0:0] mux_521_nl;
  wire[0:0] and_499_nl;
  wire[0:0] nor_488_nl;
  wire[0:0] nor_489_nl;
  wire[0:0] mux_520_nl;
  wire[0:0] mux_519_nl;
  wire[0:0] mux_518_nl;
  wire[0:0] nor_490_nl;
  wire[0:0] nor_491_nl;
  wire[0:0] mux_517_nl;
  wire[0:0] or_532_nl;
  wire[0:0] or_530_nl;
  wire[0:0] nor_492_nl;
  wire[0:0] nor_493_nl;
  wire[0:0] mux_516_nl;
  wire[0:0] mux_515_nl;
  wire[0:0] or_525_nl;
  wire[0:0] mux_514_nl;
  wire[0:0] nand_232_nl;
  wire[0:0] or_522_nl;
  wire[0:0] nand_22_nl;
  wire[0:0] mux_513_nl;
  wire[0:0] nor_494_nl;
  wire[0:0] nor_495_nl;
  wire[0:0] or_517_nl;
  wire[0:0] mux_549_nl;
  wire[0:0] mux_548_nl;
  wire[0:0] mux_547_nl;
  wire[0:0] mux_546_nl;
  wire[0:0] or_582_nl;
  wire[0:0] or_580_nl;
  wire[0:0] mux_545_nl;
  wire[0:0] mux_544_nl;
  wire[0:0] mux_543_nl;
  wire[0:0] or_579_nl;
  wire[0:0] or_578_nl;
  wire[0:0] or_576_nl;
  wire[0:0] mux_542_nl;
  wire[0:0] mux_541_nl;
  wire[0:0] mux_540_nl;
  wire[0:0] mux_539_nl;
  wire[0:0] or_575_nl;
  wire[0:0] mux_537_nl;
  wire[0:0] mux_536_nl;
  wire[0:0] or_566_nl;
  wire[0:0] mux_534_nl;
  wire[0:0] mux_533_nl;
  wire[0:0] mux_532_nl;
  wire[0:0] mux_531_nl;
  wire[0:0] or_559_nl;
  wire[0:0] mux_530_nl;
  wire[0:0] or_554_nl;
  wire[0:0] mux_529_nl;
  wire[0:0] mux_528_nl;
  wire[0:0] or_551_nl;
  wire[0:0] nor_114_nl;
  wire[0:0] mux_563_nl;
  wire[0:0] nor_472_nl;
  wire[0:0] mux_562_nl;
  wire[0:0] nand_27_nl;
  wire[0:0] mux_561_nl;
  wire[0:0] nor_474_nl;
  wire[0:0] or_609_nl;
  wire[0:0] mux_560_nl;
  wire[0:0] or_608_nl;
  wire[0:0] or_607_nl;
  wire[0:0] mux_559_nl;
  wire[0:0] and_409_nl;
  wire[0:0] mux_558_nl;
  wire[0:0] nor_475_nl;
  wire[0:0] nor_476_nl;
  wire[0:0] nor_477_nl;
  wire[0:0] mux_557_nl;
  wire[0:0] mux_556_nl;
  wire[0:0] mux_555_nl;
  wire[0:0] nor_478_nl;
  wire[0:0] nor_479_nl;
  wire[0:0] mux_554_nl;
  wire[0:0] or_598_nl;
  wire[0:0] or_596_nl;
  wire[0:0] nor_480_nl;
  wire[0:0] nor_481_nl;
  wire[0:0] mux_553_nl;
  wire[0:0] mux_552_nl;
  wire[0:0] or_591_nl;
  wire[0:0] mux_551_nl;
  wire[0:0] or_590_nl;
  wire[0:0] or_589_nl;
  wire[0:0] nand_25_nl;
  wire[0:0] mux_550_nl;
  wire[0:0] nor_482_nl;
  wire[0:0] or_583_nl;
  wire[0:0] mux_586_nl;
  wire[0:0] mux_585_nl;
  wire[0:0] mux_584_nl;
  wire[0:0] mux_583_nl;
  wire[0:0] or_647_nl;
  wire[0:0] or_645_nl;
  wire[0:0] mux_582_nl;
  wire[0:0] mux_581_nl;
  wire[0:0] mux_580_nl;
  wire[0:0] or_644_nl;
  wire[0:0] or_643_nl;
  wire[0:0] or_641_nl;
  wire[0:0] mux_579_nl;
  wire[0:0] mux_578_nl;
  wire[0:0] mux_577_nl;
  wire[0:0] mux_576_nl;
  wire[0:0] or_640_nl;
  wire[0:0] mux_574_nl;
  wire[0:0] mux_573_nl;
  wire[0:0] or_631_nl;
  wire[0:0] mux_571_nl;
  wire[0:0] mux_570_nl;
  wire[0:0] mux_569_nl;
  wire[0:0] mux_568_nl;
  wire[0:0] or_624_nl;
  wire[0:0] mux_567_nl;
  wire[0:0] or_619_nl;
  wire[0:0] mux_566_nl;
  wire[0:0] mux_565_nl;
  wire[0:0] or_616_nl;
  wire[0:0] nor_120_nl;
  wire[0:0] mux_600_nl;
  wire[0:0] nor_460_nl;
  wire[0:0] mux_599_nl;
  wire[0:0] nand_30_nl;
  wire[0:0] mux_598_nl;
  wire[0:0] nor_462_nl;
  wire[0:0] or_674_nl;
  wire[0:0] mux_597_nl;
  wire[0:0] or_673_nl;
  wire[0:0] or_672_nl;
  wire[0:0] mux_596_nl;
  wire[0:0] and_408_nl;
  wire[0:0] mux_595_nl;
  wire[0:0] and_498_nl;
  wire[0:0] nor_464_nl;
  wire[0:0] nor_465_nl;
  wire[0:0] mux_594_nl;
  wire[0:0] mux_593_nl;
  wire[0:0] mux_592_nl;
  wire[0:0] nor_466_nl;
  wire[0:0] nor_467_nl;
  wire[0:0] mux_591_nl;
  wire[0:0] or_663_nl;
  wire[0:0] or_661_nl;
  wire[0:0] nor_468_nl;
  wire[0:0] nor_469_nl;
  wire[0:0] mux_590_nl;
  wire[0:0] mux_589_nl;
  wire[0:0] or_656_nl;
  wire[0:0] mux_588_nl;
  wire[0:0] or_655_nl;
  wire[0:0] or_654_nl;
  wire[0:0] nand_28_nl;
  wire[0:0] mux_587_nl;
  wire[0:0] nor_470_nl;
  wire[0:0] or_648_nl;
  wire[0:0] mux_623_nl;
  wire[0:0] mux_622_nl;
  wire[0:0] mux_621_nl;
  wire[0:0] mux_620_nl;
  wire[0:0] or_711_nl;
  wire[0:0] or_709_nl;
  wire[0:0] mux_619_nl;
  wire[0:0] mux_618_nl;
  wire[0:0] mux_617_nl;
  wire[0:0] or_708_nl;
  wire[0:0] or_707_nl;
  wire[0:0] or_705_nl;
  wire[0:0] mux_616_nl;
  wire[0:0] mux_615_nl;
  wire[0:0] mux_614_nl;
  wire[0:0] mux_613_nl;
  wire[0:0] or_704_nl;
  wire[0:0] mux_611_nl;
  wire[0:0] mux_610_nl;
  wire[0:0] or_696_nl;
  wire[0:0] mux_608_nl;
  wire[0:0] mux_607_nl;
  wire[0:0] mux_606_nl;
  wire[0:0] mux_605_nl;
  wire[0:0] or_689_nl;
  wire[0:0] mux_604_nl;
  wire[0:0] or_684_nl;
  wire[0:0] mux_603_nl;
  wire[0:0] mux_602_nl;
  wire[0:0] or_681_nl;
  wire[0:0] nor_126_nl;
  wire[0:0] mux_637_nl;
  wire[0:0] nor_446_nl;
  wire[0:0] mux_636_nl;
  wire[0:0] nand_34_nl;
  wire[0:0] mux_635_nl;
  wire[0:0] nor_448_nl;
  wire[0:0] or_738_nl;
  wire[0:0] mux_634_nl;
  wire[0:0] or_737_nl;
  wire[0:0] or_736_nl;
  wire[0:0] mux_633_nl;
  wire[0:0] and_407_nl;
  wire[0:0] mux_632_nl;
  wire[0:0] and_497_nl;
  wire[0:0] nor_450_nl;
  wire[0:0] nor_451_nl;
  wire[0:0] mux_631_nl;
  wire[0:0] mux_630_nl;
  wire[0:0] mux_629_nl;
  wire[0:0] nor_452_nl;
  wire[0:0] nor_453_nl;
  wire[0:0] mux_628_nl;
  wire[0:0] or_727_nl;
  wire[0:0] or_725_nl;
  wire[0:0] nor_454_nl;
  wire[0:0] nor_455_nl;
  wire[0:0] mux_627_nl;
  wire[0:0] mux_626_nl;
  wire[0:0] or_720_nl;
  wire[0:0] mux_625_nl;
  wire[0:0] or_719_nl;
  wire[0:0] or_718_nl;
  wire[0:0] nand_32_nl;
  wire[0:0] mux_624_nl;
  wire[0:0] nor_456_nl;
  wire[0:0] or_712_nl;
  wire[0:0] mux_660_nl;
  wire[0:0] mux_659_nl;
  wire[0:0] mux_658_nl;
  wire[0:0] mux_657_nl;
  wire[0:0] nand_251_nl;
  wire[0:0] or_773_nl;
  wire[0:0] mux_656_nl;
  wire[0:0] mux_655_nl;
  wire[0:0] mux_654_nl;
  wire[0:0] or_772_nl;
  wire[0:0] nand_252_nl;
  wire[0:0] nand_144_nl;
  wire[0:0] mux_653_nl;
  wire[0:0] mux_652_nl;
  wire[0:0] mux_651_nl;
  wire[0:0] mux_650_nl;
  wire[0:0] nand_250_nl;
  wire[0:0] mux_648_nl;
  wire[0:0] mux_647_nl;
  wire[0:0] or_760_nl;
  wire[0:0] mux_645_nl;
  wire[0:0] mux_644_nl;
  wire[0:0] mux_643_nl;
  wire[0:0] mux_642_nl;
  wire[0:0] nand_147_nl;
  wire[0:0] mux_641_nl;
  wire[0:0] or_748_nl;
  wire[0:0] mux_640_nl;
  wire[0:0] mux_639_nl;
  wire[0:0] nand_149_nl;
  wire[0:0] and_406_nl;
  wire[0:0] mux_674_nl;
  wire[0:0] nor_433_nl;
  wire[0:0] mux_673_nl;
  wire[0:0] nand_38_nl;
  wire[0:0] mux_672_nl;
  wire[0:0] nor_435_nl;
  wire[0:0] or_802_nl;
  wire[0:0] mux_671_nl;
  wire[0:0] nand_134_nl;
  wire[0:0] or_800_nl;
  wire[0:0] mux_670_nl;
  wire[0:0] and_404_nl;
  wire[0:0] mux_669_nl;
  wire[0:0] and_495_nl;
  wire[0:0] nor_437_nl;
  wire[0:0] nor_438_nl;
  wire[0:0] mux_668_nl;
  wire[0:0] mux_667_nl;
  wire[0:0] mux_666_nl;
  wire[0:0] nor_439_nl;
  wire[0:0] nor_440_nl;
  wire[0:0] mux_665_nl;
  wire[0:0] nand_237_nl;
  wire[0:0] or_789_nl;
  wire[0:0] and_405_nl;
  wire[0:0] nor_441_nl;
  wire[0:0] mux_664_nl;
  wire[0:0] mux_663_nl;
  wire[0:0] or_784_nl;
  wire[0:0] mux_662_nl;
  wire[0:0] nand_139_nl;
  wire[0:0] nand_231_nl;
  wire[0:0] nand_36_nl;
  wire[0:0] mux_661_nl;
  wire[0:0] nor_442_nl;
  wire[0:0] or_776_nl;
  wire[0:0] mux_1347_nl;
  wire[0:0] nor_635_nl;
  wire[0:0] nor_636_nl;
  wire[0:0] mux_1346_nl;
  wire[0:0] nor_637_nl;
  wire[0:0] mux_1345_nl;
  wire[0:0] and_nl;
  wire[0:0] mux_1344_nl;
  wire[0:0] or_1438_nl;
  wire[0:0] mux_1372_nl;
  wire[0:0] or_1436_nl;
  wire[10:0] acc_nl;
  wire[11:0] nl_acc_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_7_nl;
  wire[8:0] COMP_LOOP_COMP_LOOP_mux_8_nl;
  wire[0:0] COMP_LOOP_or_44_nl;
  wire[5:0] COMP_LOOP_COMP_LOOP_mux_9_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_8_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_9_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_10_nl;
  wire[2:0] COMP_LOOP_or_45_nl;
  wire[2:0] COMP_LOOP_mux1h_125_nl;
  wire[0:0] and_722_nl;
  wire[0:0] and_723_nl;
  wire[0:0] and_724_nl;
  wire[0:0] and_725_nl;
  wire[0:0] and_726_nl;
  wire[0:0] and_727_nl;
  wire[65:0] acc_2_nl;
  wire[66:0] nl_acc_2_nl;
  wire[63:0] COMP_LOOP_mux1h_126_nl;
  wire[0:0] COMP_LOOP_or_46_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_11_nl;
  wire[2:0] COMP_LOOP_COMP_LOOP_or_12_nl;
  wire[2:0] COMP_LOOP_and_85_nl;
  wire[0:0] COMP_LOOP_nor_107_nl;
  wire[5:0] COMP_LOOP_COMP_LOOP_or_13_nl;
  wire[5:0] COMP_LOOP_mux_41_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_53_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_54_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_55_nl;
  wire[0:0] operator_64_false_1_mux_51_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_56_nl;
  wire[0:0] operator_64_false_1_mux_52_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_57_nl;
  wire[0:0] operator_64_false_1_mux_53_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_58_nl;
  wire[0:0] operator_64_false_1_mux_54_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_59_nl;
  wire[0:0] operator_64_false_1_mux_55_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_60_nl;
  wire[0:0] operator_64_false_1_mux_56_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_61_nl;
  wire[0:0] operator_64_false_1_mux_57_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_62_nl;
  wire[0:0] operator_64_false_1_mux_58_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_63_nl;
  wire[0:0] operator_64_false_1_mux_59_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_64_nl;
  wire[0:0] operator_64_false_1_mux_60_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_65_nl;
  wire[0:0] operator_64_false_1_mux_61_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_66_nl;
  wire[0:0] operator_64_false_1_mux_62_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_67_nl;
  wire[0:0] operator_64_false_1_mux_63_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_68_nl;
  wire[0:0] operator_64_false_1_mux_64_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_69_nl;
  wire[0:0] operator_64_false_1_mux_65_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_70_nl;
  wire[0:0] operator_64_false_1_mux_66_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_71_nl;
  wire[0:0] operator_64_false_1_mux_67_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_72_nl;
  wire[0:0] operator_64_false_1_mux_68_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_73_nl;
  wire[0:0] operator_64_false_1_mux_69_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_74_nl;
  wire[0:0] operator_64_false_1_mux_70_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_75_nl;
  wire[0:0] operator_64_false_1_mux_71_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_76_nl;
  wire[0:0] operator_64_false_1_mux_72_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_77_nl;
  wire[0:0] operator_64_false_1_mux_73_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_78_nl;
  wire[0:0] operator_64_false_1_mux_74_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_79_nl;
  wire[0:0] operator_64_false_1_mux_75_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_80_nl;
  wire[0:0] operator_64_false_1_mux_76_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_81_nl;
  wire[0:0] operator_64_false_1_mux_77_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_82_nl;
  wire[0:0] operator_64_false_1_mux_78_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_83_nl;
  wire[0:0] operator_64_false_1_mux_79_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_84_nl;
  wire[0:0] operator_64_false_1_mux_80_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_85_nl;
  wire[0:0] operator_64_false_1_mux_81_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_86_nl;
  wire[0:0] operator_64_false_1_mux_82_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_87_nl;
  wire[0:0] operator_64_false_1_mux_83_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_88_nl;
  wire[0:0] operator_64_false_1_mux_84_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_89_nl;
  wire[0:0] operator_64_false_1_mux_85_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_90_nl;
  wire[0:0] operator_64_false_1_mux_86_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_91_nl;
  wire[0:0] operator_64_false_1_mux_87_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_92_nl;
  wire[0:0] operator_64_false_1_mux_88_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_93_nl;
  wire[0:0] operator_64_false_1_mux_89_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_94_nl;
  wire[0:0] operator_64_false_1_mux_90_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_95_nl;
  wire[0:0] operator_64_false_1_mux_91_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_96_nl;
  wire[0:0] operator_64_false_1_mux_92_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_97_nl;
  wire[0:0] operator_64_false_1_mux_93_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_98_nl;
  wire[0:0] operator_64_false_1_mux_94_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_99_nl;
  wire[0:0] operator_64_false_1_mux_95_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_100_nl;
  wire[0:0] operator_64_false_1_mux_96_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_101_nl;
  wire[0:0] operator_64_false_1_mux_97_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_102_nl;
  wire[0:0] operator_64_false_1_mux_98_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_103_nl;
  wire[0:0] operator_64_false_1_mux_99_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_104_nl;
  wire[0:0] operator_64_false_1_mux_100_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_105_nl;
  wire[0:0] operator_64_false_1_mux_101_nl;
  wire[3:0] operator_64_false_1_or_7_nl;
  wire[3:0] operator_64_false_1_operator_64_false_1_nor_105_nl;
  wire[3:0] operator_64_false_1_mux1h_4_nl;
  wire[0:0] operator_64_false_1_or_8_nl;
  wire[7:0] operator_64_false_1_mux1h_5_nl;
  wire[6:0] operator_64_false_1_and_53_nl;
  wire[6:0] operator_64_false_1_mux1h_6_nl;
  wire[0:0] operator_64_false_1_not_3_nl;
  wire[2:0] operator_64_false_1_mux1h_7_nl;
  wire[0:0] operator_64_false_1_or_9_nl;
  wire[63:0] modExp_while_if_mux1h_2_nl;
  wire[0:0] and_728_nl;
  wire[0:0] mux_1459_nl;
  wire[0:0] mux_1460_nl;
  wire[0:0] mux_1461_nl;
  wire[0:0] nor_690_nl;
  wire[0:0] nor_691_nl;
  wire[0:0] mux_1462_nl;
  wire[0:0] or_1560_nl;
  wire[0:0] or_1561_nl;
  wire[0:0] mux_1463_nl;
  wire[0:0] nor_692_nl;
  wire[0:0] and_729_nl;
  wire[0:0] mux_1464_nl;
  wire[0:0] nor_693_nl;
  wire[0:0] mux_1465_nl;
  wire[0:0] or_1562_nl;
  wire[0:0] and_730_nl;
  wire[0:0] mux_1466_nl;
  wire[0:0] nor_694_nl;
  wire[0:0] nor_695_nl;
  wire[0:0] mux_1467_nl;
  wire[0:0] mux_1468_nl;
  wire[0:0] nand_279_nl;
  wire[0:0] mux_1469_nl;
  wire[0:0] nor_696_nl;
  wire[0:0] nor_697_nl;
  wire[0:0] mux_1470_nl;
  wire[0:0] mux_1471_nl;
  wire[0:0] mux_1472_nl;
  wire[0:0] or_1564_nl;
  wire[0:0] or_1565_nl;
  wire[0:0] or_1566_nl;
  wire[0:0] mux_1473_nl;
  wire[0:0] or_1567_nl;
  wire[0:0] or_1568_nl;
  wire[0:0] mux_1474_nl;
  wire[0:0] mux_1475_nl;
  wire[0:0] mux_1476_nl;
  wire[0:0] or_1569_nl;
  wire[0:0] mux_1477_nl;
  wire[0:0] or_1570_nl;
  wire[0:0] or_1571_nl;
  wire[0:0] mux_1478_nl;
  wire[0:0] mux_1479_nl;
  wire[0:0] nand_280_nl;
  wire[0:0] mux_1480_nl;
  wire[0:0] nand_281_nl;
  wire[0:0] mux_1481_nl;
  wire[0:0] or_1572_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [10:0] nl_operator_66_true_div_cmp_b;
  assign nl_operator_66_true_div_cmp_b = {1'b0, operator_66_true_div_cmp_b_9_0};
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0 = ~ (z_out_3[64]);
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_62_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_62_tr0 = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_124_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_124_tr0 = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_186_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_186_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_248_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_248_tr0 = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_310_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_310_tr0 = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_372_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_372_tr0 = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_434_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_434_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 = z_out_3[12];
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0 = ~ STAGE_LOOP_acc_itm_2_1;
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd64)) r_rsci (
      .dat(r_rsc_dat),
      .idat(r_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_7_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(vec_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_6_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(vec_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_5_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(vec_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_4_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(vec_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_3_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(vec_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_2_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(vec_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_1_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(vec_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(vec_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd1)) modulo_result_rem_cmp (
      .a(modulo_result_rem_cmp_a),
      .b(modulo_result_rem_cmp_b),
      .z(modulo_result_rem_cmp_z)
    );
  mgc_div #(.width_a(32'sd65),
  .width_b(32'sd11),
  .signd(32'sd1)) operator_66_true_div_cmp (
      .a(operator_66_true_div_cmp_a),
      .b(nl_operator_66_true_div_cmp_b[10:0]),
      .z(operator_66_true_div_cmp_z)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd10)) STAGE_LOOP_lshift_rg (
      .a(1'b1),
      .s(STAGE_LOOP_i_3_0_sva),
      .z(STAGE_LOOP_lshift_psp_sva_mx0w0)
    );
  inPlaceNTT_DIT_core_core_fsm inPlaceNTT_DIT_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .STAGE_LOOP_C_8_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0[0:0]),
      .modExp_while_C_38_tr0(COMP_LOOP_COMP_LOOP_and_11_itm),
      .COMP_LOOP_C_1_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0[0:0]),
      .COMP_LOOP_1_modExp_1_while_C_38_tr0(COMP_LOOP_COMP_LOOP_and_11_itm),
      .COMP_LOOP_C_62_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_62_tr0[0:0]),
      .COMP_LOOP_2_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_124_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_124_tr0[0:0]),
      .COMP_LOOP_3_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_186_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_186_tr0[0:0]),
      .COMP_LOOP_4_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_248_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_248_tr0[0:0]),
      .COMP_LOOP_5_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_310_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_310_tr0[0:0]),
      .COMP_LOOP_6_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_372_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_372_tr0[0:0]),
      .COMP_LOOP_7_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_434_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_434_tr0[0:0]),
      .COMP_LOOP_8_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_496_tr0(COMP_LOOP_COMP_LOOP_and_145_itm),
      .VEC_LOOP_C_0_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0[0:0]),
      .STAGE_LOOP_C_9_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0[0:0])
    );
  assign nand_190_cse = ~((fsm_output[3]) & (fsm_output[2]) & (fsm_output[6]) & (fsm_output[7]));
  assign and_416_cse = (fsm_output[5]) & (fsm_output[4]) & (fsm_output[6]) & (~ (fsm_output[8]));
  assign nand_168_cse = ~((fsm_output[3]) & (fsm_output[6]) & (fsm_output[7]));
  assign and_389_cse = (fsm_output[1:0]==2'b11);
  assign or_838_cse = (fsm_output[1:0]!=2'b00);
  assign or_1391_cse = (fsm_output[2:1]!=2'b00);
  assign nor_425_cse = ~((fsm_output[6:5]!=2'b01));
  assign or_817_cse = (~ (fsm_output[5])) | (fsm_output[3]);
  assign or_816_cse = (fsm_output[5:4]!=2'b01);
  assign or_1392_cse = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[9]);
  assign and_382_cse = or_838_cse & (fsm_output[2]);
  assign or_1394_cse = and_389_cse | (fsm_output[2]);
  assign or_1099_cse = (fsm_output[6]) | (fsm_output[9]);
  assign or_1113_nl = (fsm_output[5]) | (~ (fsm_output[0])) | (fsm_output[9]) | not_tmp_462;
  assign or_1111_nl = (fsm_output[0]) | (~ (fsm_output[9])) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (~ (fsm_output[4]));
  assign or_1109_nl = (~ (fsm_output[0])) | (fsm_output[9]) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[4]));
  assign mux_1119_nl = MUX_s_1_2_2(or_1111_nl, or_1109_nl, fsm_output[5]);
  assign mux_1120_nl = MUX_s_1_2_2(or_1113_nl, mux_1119_nl, fsm_output[1]);
  assign nor_340_nl = ~((fsm_output[6]) | mux_1120_nl);
  assign nor_341_nl = ~((fsm_output[1]) | (~ (fsm_output[5])) | (~ (fsm_output[0]))
      | (~ (fsm_output[9])) | (fsm_output[7]) | (~ (fsm_output[3])) | (fsm_output[4]));
  assign nor_342_nl = ~((fsm_output[9]) | not_tmp_462);
  assign and_492_nl = (fsm_output[9]) & (fsm_output[7]) & (~ (fsm_output[3])) & (fsm_output[4]);
  assign mux_1117_nl = MUX_s_1_2_2(nor_342_nl, and_492_nl, fsm_output[0]);
  assign and_324_nl = (fsm_output[1]) & (fsm_output[5]) & mux_1117_nl;
  assign mux_1118_nl = MUX_s_1_2_2(nor_341_nl, and_324_nl, fsm_output[6]);
  assign mux_1121_nl = MUX_s_1_2_2(nor_340_nl, mux_1118_nl, fsm_output[2]);
  assign nor_344_nl = ~((fsm_output[5]) | (fsm_output[0]) | (fsm_output[9]) | (~
      (fsm_output[7])) | (~ (fsm_output[3])) | (fsm_output[4]));
  assign nor_345_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[0])) | (fsm_output[9])
      | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[4]));
  assign mux_1116_nl = MUX_s_1_2_2(nor_344_nl, nor_345_nl, fsm_output[1]);
  assign and_325_nl = (~((fsm_output[2]) | (~ (fsm_output[6])))) & mux_1116_nl;
  assign mux_1122_nl = MUX_s_1_2_2(mux_1121_nl, and_325_nl, fsm_output[8]);
  assign modExp_while_if_or_nl = and_dcpl_147 | (mux_1122_nl & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign modExp_while_if_and_1_nl = modExp_while_and_3 & not_tmp_414;
  assign modExp_while_if_and_2_nl = modExp_while_and_5 & not_tmp_414;
  assign modExp_while_if_mux1h_nl = MUX1HOT_v_64_5_2(z_out_4, 64'b0000000000000000000000000000000000000000000000000000000000000001,
      modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w1, COMP_LOOP_1_acc_5_mut_mx0w5,
      {modExp_while_if_or_nl , not_tmp_374 , modExp_while_if_and_1_nl , modExp_while_if_and_2_nl
      , not_tmp_312});
  assign and_179_nl = and_dcpl_51 & and_dcpl_58 & and_dcpl_48;
  assign mux_851_nl = MUX_s_1_2_2(or_tmp_113, nor_tmp_23, fsm_output[5]);
  assign mux_852_nl = MUX_s_1_2_2(mux_851_nl, or_247_cse, fsm_output[6]);
  assign mux_849_nl = MUX_s_1_2_2((~ nor_tmp), or_tmp_788, fsm_output[5]);
  assign mux_850_nl = MUX_s_1_2_2(mux_tmp_677, mux_849_nl, fsm_output[6]);
  assign mux_853_nl = MUX_s_1_2_2(mux_852_nl, mux_850_nl, fsm_output[2]);
  assign or_1388_nl = (fsm_output[5]) | mux_tmp_845;
  assign mux_846_nl = MUX_s_1_2_2(mux_tmp_845, (~ or_216_cse), fsm_output[5]);
  assign mux_847_nl = MUX_s_1_2_2(or_1388_nl, mux_846_nl, fsm_output[6]);
  assign or_928_nl = (fsm_output[5]) | and_462_cse;
  assign mux_843_nl = MUX_s_1_2_2((fsm_output[4]), mux_342_cse, fsm_output[5]);
  assign mux_844_nl = MUX_s_1_2_2(or_928_nl, mux_843_nl, fsm_output[6]);
  assign mux_848_nl = MUX_s_1_2_2(mux_847_nl, mux_844_nl, fsm_output[2]);
  assign mux_854_nl = MUX_s_1_2_2(mux_853_nl, mux_848_nl, fsm_output[7]);
  assign and_372_nl = (fsm_output[5]) & (~ mux_tmp_719);
  assign mux_839_nl = MUX_s_1_2_2(or_tmp_788, (~ or_tmp_891), fsm_output[5]);
  assign mux_840_nl = MUX_s_1_2_2(and_372_nl, mux_839_nl, fsm_output[6]);
  assign and_373_nl = (fsm_output[5]) & (~ mux_342_cse);
  assign nor_397_nl = ~((fsm_output[5]) | and_dcpl_50);
  assign mux_838_nl = MUX_s_1_2_2(and_373_nl, nor_397_nl, fsm_output[6]);
  assign mux_841_nl = MUX_s_1_2_2(mux_840_nl, mux_838_nl, fsm_output[2]);
  assign or_925_nl = ((~ (fsm_output[5])) & (fsm_output[0]) & (fsm_output[1]) & (fsm_output[3]))
      | (fsm_output[4]);
  assign mux_835_nl = MUX_s_1_2_2(or_925_nl, mux_tmp_722, fsm_output[6]);
  assign mux_833_nl = MUX_s_1_2_2((~ mux_tmp_688), (fsm_output[4]), fsm_output[5]);
  assign mux_834_nl = MUX_s_1_2_2(mux_833_nl, mux_tmp_718, fsm_output[6]);
  assign mux_836_nl = MUX_s_1_2_2(mux_835_nl, mux_834_nl, fsm_output[2]);
  assign mux_842_nl = MUX_s_1_2_2(mux_841_nl, mux_836_nl, fsm_output[7]);
  assign mux_855_nl = MUX_s_1_2_2((~ mux_854_nl), mux_842_nl, fsm_output[8]);
  assign mux_828_nl = MUX_s_1_2_2(mux_331_cse, (~ or_tmp_788), fsm_output[5]);
  assign mux_826_nl = MUX_s_1_2_2(nor_tmp, mux_tmp_688, fsm_output[5]);
  assign mux_829_nl = MUX_s_1_2_2(mux_828_nl, mux_826_nl, fsm_output[6]);
  assign mux_824_nl = MUX_s_1_2_2(and_705_cse, (~ or_216_cse), fsm_output[5]);
  assign mux_823_nl = MUX_s_1_2_2(and_705_cse, mux_tmp_156, fsm_output[5]);
  assign mux_825_nl = MUX_s_1_2_2(mux_824_nl, mux_823_nl, fsm_output[6]);
  assign mux_830_nl = MUX_s_1_2_2(mux_829_nl, mux_825_nl, fsm_output[2]);
  assign mux_820_nl = MUX_s_1_2_2((~ (fsm_output[4])), and_dcpl_59, fsm_output[5]);
  assign mux_821_nl = MUX_s_1_2_2(mux_820_nl, (~ nor_tmp_146), fsm_output[6]);
  assign mux_818_nl = MUX_s_1_2_2(mux_tmp_689, (~ and_705_cse), fsm_output[5]);
  assign mux_819_nl = MUX_s_1_2_2(mux_tmp_705, mux_818_nl, fsm_output[6]);
  assign mux_822_nl = MUX_s_1_2_2(mux_821_nl, mux_819_nl, fsm_output[2]);
  assign mux_831_nl = MUX_s_1_2_2(mux_830_nl, mux_822_nl, fsm_output[7]);
  assign and_376_nl = (fsm_output[5]) & (~ nor_tmp_23);
  assign mux_816_nl = MUX_s_1_2_2(and_376_nl, or_1202_cse, fsm_output[6]);
  assign mux_815_nl = MUX_s_1_2_2(and_428_cse, (~ (fsm_output[4])), fsm_output[5]);
  assign or_923_nl = (fsm_output[6]) | mux_815_nl;
  assign mux_817_nl = MUX_s_1_2_2(mux_816_nl, or_923_nl, fsm_output[2]);
  assign or_924_nl = (fsm_output[7]) | mux_817_nl;
  assign mux_832_nl = MUX_s_1_2_2(mux_831_nl, or_924_nl, fsm_output[8]);
  assign mux_856_nl = MUX_s_1_2_2(mux_855_nl, mux_832_nl, fsm_output[9]);
  assign operator_64_false_mux1h_2_rgt = MUX1HOT_v_65_3_2(z_out_2, ({2'b00 , operator_64_false_slc_modExp_exp_63_1_3}),
      ({1'b0 , modExp_while_if_mux1h_nl}), {and_179_nl , and_dcpl_156 , (~ mux_856_nl)});
  assign and_705_cse = (fsm_output[4]) & or_136_cse;
  assign or_1385_cse = (fsm_output[2:0]!=3'b000);
  assign nor_393_cse = ~((fsm_output[9:8]!=2'b00));
  assign and_369_cse = (fsm_output[9:8]==2'b11);
  assign and_187_m1c = and_dcpl_137 & and_dcpl_89 & nor_393_cse;
  assign and_491_cse = (fsm_output[6]) & or_tmp;
  assign modExp_result_and_rgt = (~ modExp_while_and_5) & and_187_m1c;
  assign modExp_result_and_1_rgt = modExp_while_and_5 & and_187_m1c;
  assign and_477_cse = (fsm_output[2:0]==3'b111);
  assign and_483_cse = (fsm_output[2:1]==2'b11);
  assign or_1423_cse = and_477_cse | (fsm_output[9]);
  assign or_245_cse = (fsm_output[1]) | (fsm_output[3]);
  assign or_247_cse = (fsm_output[5:4]!=2'b10);
  assign modulo_result_mux_1_cse = MUX_v_64_2_2(modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w1,
      modulo_result_rem_cmp_z[63]);
  assign and_428_cse = (fsm_output[0]) & (fsm_output[1]) & (fsm_output[3]) & (fsm_output[4]);
  assign or_242_cse = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[3]) | (~ (fsm_output[4]));
  assign or_42_nl = (fsm_output[6]) | (fsm_output[2]) | (~ (fsm_output[7])) | (~
      (fsm_output[9])) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign or_41_nl = (~ (fsm_output[6])) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (fsm_output[9]) | (fsm_output[4]) | (~ (fsm_output[8]));
  assign mux_33_nl = MUX_s_1_2_2(or_42_nl, or_41_nl, fsm_output[1]);
  assign or_39_nl = (~ (fsm_output[1])) | (fsm_output[6]) | (~ (fsm_output[2])) |
      (~ (fsm_output[7])) | (fsm_output[9]) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_34_nl = MUX_s_1_2_2(mux_33_nl, or_39_nl, fsm_output[0]);
  assign nor_601_cse = ~((fsm_output[3]) | mux_34_nl);
  assign nor_604_nl = ~((fsm_output[1]) | (~ (fsm_output[6])) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[9]) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_605_nl = ~((~ (fsm_output[1])) | (fsm_output[6]) | (fsm_output[2]) |
      (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[4]) | (fsm_output[8]));
  assign mux_29_cse = MUX_s_1_2_2(nor_604_nl, nor_605_nl, fsm_output[0]);
  assign mux_331_cse = MUX_s_1_2_2(mux_tmp_156, nor_tmp, and_389_cse);
  assign mux_342_cse = MUX_s_1_2_2(mux_tmp_156, nor_tmp, fsm_output[1]);
  assign and_25_cse = (fsm_output[5]) & nor_tmp_23;
  assign nor_386_nl = ~((~ (fsm_output[5])) | (fsm_output[0]) | (fsm_output[3]));
  assign nor_387_nl = ~((fsm_output[5]) | (~((fsm_output[0]) & (fsm_output[3]))));
  assign mux_915_nl = MUX_s_1_2_2(nor_386_nl, nor_387_nl, fsm_output[6]);
  assign and_243_m1c = mux_915_nl & (fsm_output[4]) & (~ (fsm_output[1])) & (~ (fsm_output[2]))
      & (~ (fsm_output[7])) & nor_393_cse;
  assign and_462_cse = (and_389_cse | (fsm_output[3])) & (fsm_output[4]);
  assign or_115_cse = (or_838_cse & (fsm_output[3])) | (fsm_output[4]);
  assign and_502_cse = (fsm_output[6]) & (fsm_output[3]) & (fsm_output[7]) & (fsm_output[2])
      & (fsm_output[8]) & (~ (fsm_output[9])) & (~ (fsm_output[4]));
  assign COMP_LOOP_COMP_LOOP_and_11_cse = (z_out_3[3:1]==3'b101);
  assign modExp_while_or_cse = and_dcpl_84 | and_dcpl_93 | and_dcpl_103 | and_dcpl_112
      | and_dcpl_123 | and_dcpl_130 | and_dcpl_138;
  assign COMP_LOOP_COMP_LOOP_and_37_cse = (z_out_3[3:1]==3'b011);
  assign nand_100_cse = ~((fsm_output[8]) & (fsm_output[4]));
  assign or_1189_cse = (fsm_output[3:2]!=2'b00);
  assign and_316_cse = (fsm_output[3:2]==2'b11);
  assign and_314_cse = (fsm_output[5:4]==2'b11);
  assign and_437_cse = (fsm_output[0]) & (fsm_output[4]);
  assign or_171_cse = (fsm_output[5:4]!=2'b00);
  assign or_210_cse = (fsm_output[4]) | (~ (fsm_output[8]));
  assign or_216_cse = (fsm_output[4:3]!=2'b00);
  assign or_1202_cse = (fsm_output[5:3]!=3'b000);
  assign nand_97_cse = ~((fsm_output[6]) & (fsm_output[8]));
  assign nand_230_cse = ~((fsm_output[9]) & (fsm_output[4]));
  assign nand_89_cse = ~((fsm_output[9]) & (fsm_output[8]) & (fsm_output[4]));
  assign COMP_LOOP_or_2_cse = and_dcpl_69 | and_dcpl_84 | and_dcpl_93 | and_dcpl_103
      | and_dcpl_112 | and_dcpl_123 | and_dcpl_130 | and_dcpl_138;
  assign COMP_LOOP_COMP_LOOP_and_12_cse = (z_out_3[3:1]==3'b110);
  assign COMP_LOOP_COMP_LOOP_and_13_cse = (z_out_3[3:1]==3'b111);
  assign nl_STAGE_LOOP_i_3_0_sva_2 = STAGE_LOOP_i_3_0_sva + 4'b0001;
  assign STAGE_LOOP_i_3_0_sva_2 = nl_STAGE_LOOP_i_3_0_sva_2[3:0];
  assign nl_COMP_LOOP_acc_psp_sva_1 = (VEC_LOOP_j_sva_11_0[11:3]) + conv_u2u_6_9(COMP_LOOP_k_9_3_sva_5_0);
  assign COMP_LOOP_acc_psp_sva_1 = nl_COMP_LOOP_acc_psp_sva_1[8:0];
  assign nl_modulo_qr_sva_1_mx0w1 = modulo_result_rem_cmp_z + p_sva;
  assign modulo_qr_sva_1_mx0w1 = nl_modulo_qr_sva_1_mx0w1[63:0];
  assign nl_COMP_LOOP_1_acc_5_mut_mx0w5 = tmp_10_lpi_4_dfm + modulo_result_mux_1_cse;
  assign COMP_LOOP_1_acc_5_mut_mx0w5 = nl_COMP_LOOP_1_acc_5_mut_mx0w5[63:0];
  assign operator_64_false_slc_modExp_exp_63_1_3 = MUX_v_63_2_2((operator_66_true_div_cmp_z[63:1]),
      (tmp_10_lpi_4_dfm[63:1]), and_dcpl_162);
  assign nl_COMP_LOOP_acc_1_cse_2_sva_mx0w0 = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_3_sva_5_0
      , 3'b001});
  assign COMP_LOOP_acc_1_cse_2_sva_mx0w0 = nl_COMP_LOOP_acc_1_cse_2_sva_mx0w0[11:0];
  assign nl_COMP_LOOP_acc_1_cse_6_sva_1 = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_3_sva_5_0
      , 3'b101});
  assign COMP_LOOP_acc_1_cse_6_sva_1 = nl_COMP_LOOP_acc_1_cse_6_sva_1[11:0];
  assign nl_COMP_LOOP_acc_1_cse_4_sva_1 = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_3_sva_5_0
      , 3'b011});
  assign COMP_LOOP_acc_1_cse_4_sva_1 = nl_COMP_LOOP_acc_1_cse_4_sva_1[11:0];
  assign nl_COMP_LOOP_k_9_3_sva_2 = conv_u2u_6_7(COMP_LOOP_k_9_3_sva_5_0) + 7'b0000001;
  assign COMP_LOOP_k_9_3_sva_2 = nl_COMP_LOOP_k_9_3_sva_2[6:0];
  assign modExp_while_and_3 = (~ (modulo_result_rem_cmp_z[63])) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  assign modExp_while_and_5 = (modulo_result_rem_cmp_z[63]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  assign COMP_LOOP_COMP_LOOP_and_211 = (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]==3'b001);
  assign COMP_LOOP_COMP_LOOP_and_213 = (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]==3'b010);
  assign COMP_LOOP_COMP_LOOP_and_215 = (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]==3'b100);
  assign nor_tmp = (fsm_output[4:3]==2'b11);
  assign or_tmp = (fsm_output[5]) | nor_tmp;
  assign or_81_cse = (fsm_output[9:8]!=2'b01);
  assign or_83_cse = (fsm_output[4]) | (fsm_output[9]);
  assign or_tmp_92 = ~((fsm_output[0]) & (fsm_output[1]) & (~ (fsm_output[3])) &
      (fsm_output[4]));
  assign or_136_cse = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[3]);
  assign nor_tmp_23 = or_245_cse & (fsm_output[4]);
  assign or_tmp_103 = and_389_cse | (fsm_output[4:3]!=2'b00);
  assign nor_tmp_27 = or_838_cse & (fsm_output[4:3]==2'b11);
  assign mux_tmp_156 = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), fsm_output[3]);
  assign or_tmp_113 = ((fsm_output[1]) & (fsm_output[3])) | (fsm_output[4]);
  assign and_dcpl_4 = (fsm_output[0]) & (fsm_output[5]);
  assign or_tmp_154 = (fsm_output[8:7]!=2'b00);
  assign and_dcpl_11 = (fsm_output[9:8]==2'b01);
  assign and_dcpl_14 = ~((fsm_output[0]) | (fsm_output[5]));
  assign and_dcpl_23 = (fsm_output[9:8]==2'b10);
  assign or_1402_nl = (fsm_output[8:0]!=9'b000000000);
  assign and_432_nl = (fsm_output[6:5]==2'b11);
  assign mux_361_nl = MUX_s_1_2_2(and_432_nl, and_491_cse, fsm_output[2]);
  assign nand_199_nl = ~((fsm_output[8]) & ((fsm_output[7]) | mux_361_nl));
  assign not_tmp_131 = MUX_s_1_2_2(or_1402_nl, nand_199_nl, fsm_output[9]);
  assign and_dcpl_46 = ~((fsm_output[6]) | (fsm_output[2]));
  assign and_dcpl_47 = and_dcpl_46 & (~ (fsm_output[7]));
  assign and_dcpl_48 = and_dcpl_47 & nor_393_cse;
  assign and_dcpl_50 = ~((fsm_output[4:3]!=2'b00));
  assign and_dcpl_51 = and_dcpl_50 & (~ (fsm_output[1]));
  assign and_dcpl_56 = (fsm_output[6]) & (~ (fsm_output[2])) & (~ (fsm_output[7]));
  assign and_dcpl_57 = and_dcpl_56 & and_369_cse;
  assign and_dcpl_58 = (fsm_output[0]) & (~ (fsm_output[5]));
  assign and_dcpl_59 = nor_tmp & (fsm_output[1]);
  assign and_dcpl_60 = and_dcpl_59 & and_dcpl_58;
  assign and_dcpl_63 = (fsm_output[4:3]==2'b10);
  assign and_dcpl_64 = and_dcpl_63 & (~ (fsm_output[1]));
  assign and_dcpl_65 = and_dcpl_64 & and_dcpl_4;
  assign and_dcpl_66 = and_dcpl_65 & and_dcpl_48;
  assign and_dcpl_67 = and_dcpl_56 & nor_393_cse;
  assign and_dcpl_68 = and_dcpl_59 & and_dcpl_14;
  assign and_dcpl_69 = and_dcpl_68 & and_dcpl_67;
  assign and_dcpl_70 = and_dcpl_46 & (fsm_output[7]);
  assign and_dcpl_73 = and_dcpl_50 & (fsm_output[1]) & and_dcpl_14;
  assign and_dcpl_80 = (~ (fsm_output[6])) & (fsm_output[2]);
  assign and_dcpl_82 = and_dcpl_80 & (fsm_output[7]) & nor_393_cse;
  assign and_dcpl_84 = and_dcpl_59 & and_dcpl_4 & and_dcpl_82;
  assign and_dcpl_89 = and_dcpl_80 & (~ (fsm_output[7]));
  assign and_dcpl_91 = (~ (fsm_output[0])) & (fsm_output[5]);
  assign and_dcpl_93 = and_dcpl_51 & and_dcpl_91 & and_dcpl_89 & and_dcpl_11;
  assign and_dcpl_100 = (fsm_output[4:3]==2'b01);
  assign and_dcpl_102 = and_dcpl_100 & (~ (fsm_output[1])) & and_dcpl_58;
  assign and_dcpl_103 = and_dcpl_102 & and_dcpl_70 & and_dcpl_11;
  assign and_dcpl_108 = (fsm_output[6]) & (fsm_output[2]) & (fsm_output[7]);
  assign and_dcpl_109 = and_dcpl_108 & and_dcpl_11;
  assign and_dcpl_110 = and_dcpl_100 & (fsm_output[1]);
  assign and_dcpl_112 = and_dcpl_110 & and_dcpl_91 & and_dcpl_109;
  assign and_dcpl_121 = and_dcpl_63 & (fsm_output[1]);
  assign and_dcpl_122 = and_dcpl_121 & and_dcpl_58;
  assign and_dcpl_123 = and_dcpl_122 & and_dcpl_56 & and_dcpl_23;
  assign and_dcpl_127 = and_dcpl_70 & and_dcpl_23;
  assign and_dcpl_128 = nor_tmp & (~ (fsm_output[1]));
  assign and_dcpl_129 = and_dcpl_128 & and_dcpl_91;
  assign and_dcpl_130 = and_dcpl_129 & and_dcpl_127;
  assign and_dcpl_137 = and_dcpl_128 & and_dcpl_58;
  assign and_dcpl_138 = and_dcpl_137 & and_dcpl_89 & and_369_cse;
  assign nand_194_cse = ~((fsm_output[8:7]==2'b11));
  assign or_tmp_268 = (~ (fsm_output[4])) | (fsm_output[9]) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b000) | nand_194_cse;
  assign or_308_nl = (fsm_output[4]) | (VEC_LOOP_j_sva_11_0[0]) | (VEC_LOOP_j_sva_11_0[2])
      | (fsm_output[9:5]!=5'b00100);
  assign or_306_nl = (~ (fsm_output[4])) | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_13_psp_sva[0]) | (fsm_output[8:6]!=3'b000);
  assign mux_381_nl = MUX_s_1_2_2(or_308_nl, or_306_nl, fsm_output[2]);
  assign or_tmp_273 = (VEC_LOOP_j_sva_11_0[1]) | mux_381_nl;
  assign or_329_cse = (fsm_output[9:4]!=6'b011100);
  assign or_327_cse = (fsm_output[9:4]!=6'b110101);
  assign or_325_nl = (fsm_output[9:4]!=6'b001111);
  assign or_323_nl = (fsm_output[9:4]!=6'b101000);
  assign mux_392_cse = MUX_s_1_2_2(or_325_nl, or_323_nl, fsm_output[2]);
  assign or_320_cse = (fsm_output[9:5]!=5'b00100);
  assign nand_246_cse = ~((fsm_output[9:4]==6'b101111));
  assign or_314_cse = (fsm_output[2]) | (fsm_output[4]) | (~ (fsm_output[9])) | (~
      (fsm_output[5])) | (fsm_output[6]) | (fsm_output[8]) | (fsm_output[7]);
  assign or_312_cse = (fsm_output[9:4]!=6'b010101);
  assign not_tmp_165 = ~((fsm_output[7:6]==2'b11));
  assign nand_189_cse = ~((COMP_LOOP_acc_1_cse_4_sva[0]) & (fsm_output[8:7]==2'b11));
  assign or_tmp_335 = (~ (fsm_output[4])) | (fsm_output[9]) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[2:1]!=2'b00) | nand_189_cse;
  assign or_375_nl = (fsm_output[4]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (VEC_LOOP_j_sva_11_0[2])
      | (fsm_output[9:5]!=5'b00100);
  assign or_373_nl = (~ (fsm_output[4])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_13_psp_sva[0]) | (fsm_output[8:6]!=3'b000);
  assign mux_418_nl = MUX_s_1_2_2(or_375_nl, or_373_nl, fsm_output[2]);
  assign or_tmp_340 = (VEC_LOOP_j_sva_11_0[1]) | mux_418_nl;
  assign or_tmp_395 = (~ (fsm_output[4])) | (fsm_output[9]) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b010) | nand_194_cse;
  assign nor_512_nl = ~((fsm_output[4]) | (VEC_LOOP_j_sva_11_0[0]) | (VEC_LOOP_j_sva_11_0[2])
      | (fsm_output[9:5]!=5'b00100));
  assign nor_513_nl = ~((~ (fsm_output[4])) | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_13_psp_sva[0]) | (fsm_output[8:6]!=3'b000));
  assign mux_456_nl = MUX_s_1_2_2(nor_512_nl, nor_513_nl, fsm_output[2]);
  assign nand_tmp_18 = ~((VEC_LOOP_j_sva_11_0[1]) & mux_456_nl);
  assign or_tmp_454 = (~ (fsm_output[4])) | (fsm_output[9]) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[2]) | (~((COMP_LOOP_acc_1_cse_4_sva[1:0]==2'b11)
      & (fsm_output[8:7]==2'b11)));
  assign nor_496_nl = ~((fsm_output[4]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (VEC_LOOP_j_sva_11_0[2])
      | (fsm_output[9:5]!=5'b00100));
  assign nor_497_nl = ~((~ (fsm_output[4])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_13_psp_sva[0]) | (fsm_output[8:6]!=3'b000));
  assign mux_494_nl = MUX_s_1_2_2(nor_496_nl, nor_497_nl, fsm_output[2]);
  assign nand_tmp_21 = ~((VEC_LOOP_j_sva_11_0[1]) & mux_494_nl);
  assign or_tmp_525 = (~ (fsm_output[4])) | (fsm_output[9]) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b100) | nand_194_cse;
  assign or_570_nl = (fsm_output[4]) | (VEC_LOOP_j_sva_11_0[0]) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (fsm_output[9:5]!=5'b00100);
  assign or_568_nl = (~ (fsm_output[4])) | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (~ (COMP_LOOP_acc_13_psp_sva[0])) | (fsm_output[8:6]!=3'b000);
  assign mux_538_nl = MUX_s_1_2_2(or_570_nl, or_568_nl, fsm_output[2]);
  assign or_tmp_535 = (VEC_LOOP_j_sva_11_0[1]) | mux_538_nl;
  assign or_tmp_590 = (~ (fsm_output[4])) | (fsm_output[9]) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[2:1]!=2'b10) | nand_189_cse;
  assign or_635_nl = (fsm_output[4]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (fsm_output[9:5]!=5'b00100);
  assign or_633_nl = (~ (fsm_output[4])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (~ (COMP_LOOP_acc_13_psp_sva[0])) | (fsm_output[8:6]!=3'b000);
  assign mux_575_nl = MUX_s_1_2_2(or_635_nl, or_633_nl, fsm_output[2]);
  assign or_tmp_600 = (VEC_LOOP_j_sva_11_0[1]) | mux_575_nl;
  assign or_tmp_655 = (~ (fsm_output[4])) | (fsm_output[9]) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b110) | nand_194_cse;
  assign nor_458_nl = ~((fsm_output[4]) | (VEC_LOOP_j_sva_11_0[0]) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (fsm_output[9:5]!=5'b00100));
  assign nor_459_nl = ~((~ (fsm_output[4])) | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (~ (COMP_LOOP_acc_13_psp_sva[0])) | (fsm_output[8:6]!=3'b000));
  assign mux_612_nl = MUX_s_1_2_2(nor_458_nl, nor_459_nl, fsm_output[2]);
  assign nand_tmp_31 = ~((VEC_LOOP_j_sva_11_0[1]) & mux_612_nl);
  assign or_tmp_719 = (~ (fsm_output[4])) | (fsm_output[9]) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (~((COMP_LOOP_acc_1_cse_4_sva[2:0]==3'b111) & (fsm_output[8:7]==2'b11)));
  assign nor_444_nl = ~((fsm_output[4]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (fsm_output[9:5]!=5'b00100));
  assign nor_445_nl = ~((~ (fsm_output[4])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (~ (COMP_LOOP_acc_13_psp_sva[0])) | (fsm_output[8:6]!=3'b000));
  assign mux_649_nl = MUX_s_1_2_2(nor_444_nl, nor_445_nl, fsm_output[2]);
  assign nand_tmp_35 = ~((VEC_LOOP_j_sva_11_0[1]) & mux_649_nl);
  assign and_dcpl_140 = ~((fsm_output[2]) | (fsm_output[7]));
  assign and_dcpl_147 = and_dcpl_110 & and_dcpl_14 & and_dcpl_48;
  assign mux_tmp_677 = MUX_s_1_2_2((~ mux_tmp_156), (fsm_output[4]), fsm_output[5]);
  assign mux_tmp_688 = MUX_s_1_2_2(and_dcpl_50, mux_tmp_156, fsm_output[1]);
  assign mux_tmp_689 = MUX_s_1_2_2((~ or_tmp_113), mux_tmp_688, fsm_output[0]);
  assign mux_696_itm = MUX_s_1_2_2(and_dcpl_50, mux_tmp_156, and_389_cse);
  assign nor_tmp_146 = or_817_cse & (fsm_output[4]);
  assign mux_tmp_705 = MUX_s_1_2_2((~ (fsm_output[4])), nor_tmp, fsm_output[5]);
  assign or_tmp_788 = ((fsm_output[0]) & (fsm_output[1]) & (fsm_output[3])) | (fsm_output[4]);
  assign mux_tmp_718 = MUX_s_1_2_2(and_dcpl_51, (fsm_output[4]), fsm_output[5]);
  assign mux_tmp_719 = MUX_s_1_2_2(and_dcpl_50, mux_tmp_156, or_838_cse);
  assign mux_tmp_722 = MUX_s_1_2_2(and_dcpl_50, (fsm_output[4]), fsm_output[5]);
  assign or_tmp_792 = (fsm_output[6]) | (~ or_1385_cse);
  assign nand_tmp_42 = ~((fsm_output[6]) & (~ and_382_cse));
  assign mux_tmp_731 = MUX_s_1_2_2((~ (fsm_output[6])), (fsm_output[6]), fsm_output[5]);
  assign not_tmp_274 = ~((fsm_output[2:0]==3'b111));
  assign not_tmp_280 = ~((fsm_output[6]) | (~((fsm_output[2:1]!=2'b00))));
  assign or_tmp_810 = (fsm_output[6:5]!=2'b10);
  assign or_854_nl = (~ (fsm_output[0])) | (fsm_output[5]) | (fsm_output[2]) | (~
      (fsm_output[7])) | (fsm_output[4]);
  assign or_853_nl = (~ (fsm_output[0])) | (fsm_output[5]) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_tmp_776 = MUX_s_1_2_2(or_854_nl, or_853_nl, fsm_output[9]);
  assign not_tmp_297 = ~((fsm_output[7]) & (fsm_output[4]));
  assign not_tmp_309 = ~((fsm_output[4:3]==2'b11));
  assign or_903_nl = (fsm_output[5]) | (~ (fsm_output[0])) | (~ (fsm_output[1]))
      | (~ (fsm_output[9])) | (fsm_output[3]) | (fsm_output[4]);
  assign or_902_nl = (~ (fsm_output[5])) | (fsm_output[0]) | (fsm_output[1]) | (~
      (fsm_output[9])) | (~ (fsm_output[3])) | (fsm_output[4]);
  assign mux_800_nl = MUX_s_1_2_2(or_903_nl, or_902_nl, fsm_output[6]);
  assign and_489_nl = (fsm_output[1]) & (fsm_output[9]) & (~ (fsm_output[3])) & (fsm_output[4]);
  assign nor_407_nl = ~((fsm_output[1]) | (fsm_output[9]) | not_tmp_309);
  assign mux_799_nl = MUX_s_1_2_2(and_489_nl, nor_407_nl, fsm_output[0]);
  assign nand_49_nl = ~(nor_425_cse & mux_799_nl);
  assign mux_801_nl = MUX_s_1_2_2(mux_800_nl, nand_49_nl, fsm_output[8]);
  assign nor_405_nl = ~((fsm_output[7]) | mux_801_nl);
  assign nor_408_nl = ~((fsm_output[8]) | (~ (fsm_output[6])) | (~ (fsm_output[5]))
      | (~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[9]) | (~ (fsm_output[3]))
      | (fsm_output[4]));
  assign or_895_nl = (fsm_output[1]) | (fsm_output[9]) | (fsm_output[3]) | (~ (fsm_output[4]));
  assign or_893_nl = (fsm_output[1]) | (~ (fsm_output[9])) | (~ (fsm_output[3]))
      | (fsm_output[4]);
  assign mux_796_nl = MUX_s_1_2_2(or_895_nl, or_893_nl, fsm_output[0]);
  assign nor_409_nl = ~((fsm_output[6:5]!=2'b10) | mux_796_nl);
  assign nor_410_nl = ~((fsm_output[6]) | (fsm_output[5]) | (fsm_output[0]) | (~
      (fsm_output[1])) | (fsm_output[9]) | not_tmp_309);
  assign mux_797_nl = MUX_s_1_2_2(nor_409_nl, nor_410_nl, fsm_output[8]);
  assign mux_798_nl = MUX_s_1_2_2(nor_408_nl, mux_797_nl, fsm_output[7]);
  assign not_tmp_312 = MUX_s_1_2_2(nor_405_nl, mux_798_nl, fsm_output[2]);
  assign or_1362_nl = (~ (fsm_output[7])) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign or_913_nl = (~ (fsm_output[7])) | (~ (fsm_output[9])) | (~ (fsm_output[4]))
      | (fsm_output[3]) | (fsm_output[8]);
  assign mux_806_nl = MUX_s_1_2_2(or_1362_nl, or_913_nl, fsm_output[0]);
  assign nor_400_nl = ~((fsm_output[6:5]!=2'b00) | mux_806_nl);
  assign nor_401_nl = ~((~ (fsm_output[5])) | (fsm_output[0]) | (fsm_output[7]) |
      (~ (fsm_output[9])) | (fsm_output[4]) | (~ (fsm_output[3])) | (fsm_output[8]));
  assign and_377_nl = (fsm_output[5]) & (fsm_output[0]) & (fsm_output[7]) & (~ (fsm_output[9]))
      & (fsm_output[4]) & (fsm_output[3]) & (~ (fsm_output[8]));
  assign mux_805_nl = MUX_s_1_2_2(nor_401_nl, and_377_nl, fsm_output[6]);
  assign mux_807_nl = MUX_s_1_2_2(nor_400_nl, mux_805_nl, fsm_output[2]);
  assign nor_402_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[5])) | (fsm_output[0])
      | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[4]) | (fsm_output[3]) | (~
      (fsm_output[8])));
  assign nor_403_nl = ~((~ (fsm_output[0])) | (~ (fsm_output[7])) | (fsm_output[9])
      | (fsm_output[4]) | (fsm_output[3]) | (~ (fsm_output[8])));
  assign nor_404_nl = ~((fsm_output[0]) | (~ (fsm_output[7])) | (~ (fsm_output[9]))
      | (~ (fsm_output[4])) | (fsm_output[3]) | (fsm_output[8]));
  assign mux_803_nl = MUX_s_1_2_2(nor_403_nl, nor_404_nl, fsm_output[5]);
  assign and_378_nl = (fsm_output[6]) & mux_803_nl;
  assign mux_804_nl = MUX_s_1_2_2(nor_402_nl, and_378_nl, fsm_output[2]);
  assign not_tmp_315 = MUX_s_1_2_2(mux_807_nl, mux_804_nl, fsm_output[1]);
  assign mux_809_nl = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), fsm_output[1]);
  assign or_916_nl = (~ (fsm_output[1])) | (fsm_output[3]);
  assign mux_810_nl = MUX_s_1_2_2(mux_809_nl, or_916_nl, fsm_output[0]);
  assign mux_811_nl = MUX_s_1_2_2(mux_810_nl, (fsm_output[3]), fsm_output[2]);
  assign and_dcpl_152 = ~(mux_811_nl | (fsm_output[7:4]!=4'b0000) | (~ nor_393_cse));
  assign nor_398_nl = ~((~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[4]));
  assign nor_399_nl = ~((fsm_output[0]) | (fsm_output[3]) | (~ (fsm_output[4])));
  assign mux_814_nl = MUX_s_1_2_2(nor_398_nl, nor_399_nl, fsm_output[5]);
  assign and_dcpl_156 = mux_814_nl & (~ (fsm_output[1])) & and_dcpl_48;
  assign or_tmp_891 = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[3]) | (fsm_output[4]);
  assign mux_tmp_845 = MUX_s_1_2_2(mux_tmp_156, nor_tmp, or_838_cse);
  assign not_tmp_347 = ~((fsm_output[4]) | (fsm_output[6]) | (fsm_output[8]) | (fsm_output[9]));
  assign and_361_cse = (fsm_output[6]) & (fsm_output[8]) & (fsm_output[9]);
  assign and_dcpl_162 = and_dcpl_64 & and_dcpl_91 & and_dcpl_48;
  assign or_tmp_916 = (fsm_output[6]) | and_314_cse;
  assign or_955_nl = (fsm_output[6]) | and_25_cse;
  assign mux_tmp_886 = MUX_s_1_2_2(or_955_nl, or_tmp_916, fsm_output[2]);
  assign or_tmp_918 = (fsm_output[7]) | mux_tmp_886;
  assign and_tmp_28 = (fsm_output[5]) & or_216_cse;
  assign and_dcpl_164 = ~((fsm_output[9:7]!=3'b000));
  assign and_dcpl_167 = ~((VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (fsm_output[2]) | (~
      and_dcpl_164));
  assign and_dcpl_168 = (fsm_output[6:5]==2'b01);
  assign and_dcpl_171 = and_dcpl_63 & (fsm_output[1:0]==2'b10);
  assign and_dcpl_172 = and_dcpl_171 & and_dcpl_168 & (~ (VEC_LOOP_j_sva_11_0[2]));
  assign and_dcpl_176 = (VEC_LOOP_j_sva_11_0[1:0]==2'b01) & (~ (fsm_output[2])) &
      and_dcpl_164;
  assign and_dcpl_180 = (VEC_LOOP_j_sva_11_0[1:0]==2'b10) & (~ (fsm_output[2])) &
      and_dcpl_164;
  assign and_dcpl_184 = (VEC_LOOP_j_sva_11_0[1:0]==2'b11) & (~ (fsm_output[2])) &
      and_dcpl_164;
  assign and_dcpl_187 = and_dcpl_171 & and_dcpl_168 & (VEC_LOOP_j_sva_11_0[2]);
  assign nor_382_nl = ~((~ (fsm_output[1])) | (fsm_output[6]) | (fsm_output[2]) |
      (fsm_output[7]) | (fsm_output[9]) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign nor_603_nl = ~((fsm_output[7]) | (fsm_output[9]) | (fsm_output[4]) | (~
      (fsm_output[8])));
  assign and_475_nl = (fsm_output[7]) & (fsm_output[9]) & (fsm_output[4]) & (~ (fsm_output[8]));
  assign mux_30_nl = MUX_s_1_2_2(nor_603_nl, and_475_nl, fsm_output[2]);
  assign and_474_nl = (~((fsm_output[1]) | (~ (fsm_output[6])))) & mux_30_nl;
  assign mux_918_nl = MUX_s_1_2_2(nor_382_nl, and_474_nl, fsm_output[0]);
  assign mux_919_nl = MUX_s_1_2_2(mux_918_nl, mux_29_cse, fsm_output[3]);
  assign not_tmp_374 = MUX_s_1_2_2(nor_601_cse, mux_919_nl, fsm_output[5]);
  assign or_1026_nl = (fsm_output[9]) | (fsm_output[2]) | (fsm_output[5]) | nand_100_cse;
  assign or_1024_nl = (~ (fsm_output[9])) | (~ (fsm_output[2])) | (~ (fsm_output[5]))
      | (fsm_output[8]) | (fsm_output[4]);
  assign mux_976_nl = MUX_s_1_2_2(or_1026_nl, or_1024_nl, fsm_output[7]);
  assign nor_366_nl = ~((fsm_output[3]) | (fsm_output[1]) | mux_976_nl);
  assign nor_367_nl = ~((~ (fsm_output[3])) | (~ (fsm_output[1])) | (~ (fsm_output[7]))
      | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[5]) | nand_100_cse);
  assign mux_977_nl = MUX_s_1_2_2(nor_366_nl, nor_367_nl, fsm_output[6]);
  assign nor_368_nl = ~((fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[2]) |
      (fsm_output[5]) | (~ (fsm_output[8])) | (fsm_output[4]));
  assign and_351_nl = (fsm_output[9]) & (fsm_output[2]) & (fsm_output[5]) & (~ (fsm_output[8]))
      & (fsm_output[4]);
  assign nor_369_nl = ~((fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[5])) |
      (fsm_output[8]) | (fsm_output[4]));
  assign mux_973_nl = MUX_s_1_2_2(and_351_nl, nor_369_nl, fsm_output[7]);
  assign mux_974_nl = MUX_s_1_2_2(nor_368_nl, mux_973_nl, fsm_output[1]);
  assign and_350_nl = (fsm_output[3]) & mux_974_nl;
  assign nor_370_nl = ~((fsm_output[3]) | (fsm_output[1]) | (fsm_output[7]) | (fsm_output[9])
      | (~((fsm_output[2]) & (fsm_output[5]) & (fsm_output[8]) & (fsm_output[4]))));
  assign mux_975_nl = MUX_s_1_2_2(and_350_nl, nor_370_nl, fsm_output[6]);
  assign not_tmp_399 = MUX_s_1_2_2(mux_977_nl, mux_975_nl, fsm_output[0]);
  assign not_tmp_400 = ~((fsm_output[0]) & (fsm_output[5]));
  assign not_tmp_406 = ~((fsm_output[7]) & (fsm_output[2]) & (fsm_output[6]));
  assign nor_357_cse = ~((~ (fsm_output[1])) | (~ (fsm_output[3])) | (fsm_output[6])
      | (fsm_output[8]) | (~ (fsm_output[7])) | (~ (fsm_output[2])) | (fsm_output[9])
      | (~ (fsm_output[4])));
  assign and_345_nl = (fsm_output[2]) & (fsm_output[9]) & (fsm_output[4]);
  assign nor_355_nl = ~((fsm_output[2]) | (fsm_output[9]) | (fsm_output[4]));
  assign mux_991_nl = MUX_s_1_2_2(and_345_nl, nor_355_nl, fsm_output[7]);
  assign and_344_nl = (~((~ (fsm_output[3])) | (fsm_output[6]) | (~ (fsm_output[8]))))
      & mux_991_nl;
  assign mux_990_nl = MUX_s_1_2_2(nand_230_cse, or_83_cse, fsm_output[2]);
  assign nor_356_nl = ~((fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[8]) |
      (fsm_output[7]) | mux_990_nl);
  assign mux_992_nl = MUX_s_1_2_2(and_344_nl, nor_356_nl, fsm_output[1]);
  assign mux_993_nl = MUX_s_1_2_2(mux_992_nl, nor_357_cse, fsm_output[5]);
  assign nand_111_nl = ~((fsm_output[7]) & (fsm_output[2]) & (fsm_output[9]) & (fsm_output[4]));
  assign or_1045_nl = (fsm_output[7]) | (fsm_output[2]) | (fsm_output[9]) | (fsm_output[4]);
  assign mux_988_nl = MUX_s_1_2_2(nand_111_nl, or_1045_nl, fsm_output[8]);
  assign nor_358_nl = ~((fsm_output[3]) | (fsm_output[6]) | mux_988_nl);
  assign mux_989_nl = MUX_s_1_2_2(and_502_cse, nor_358_nl, fsm_output[1]);
  assign and_346_nl = (fsm_output[5]) & mux_989_nl;
  assign not_tmp_414 = MUX_s_1_2_2(mux_993_nl, and_346_nl, fsm_output[0]);
  assign mux_tmp_997 = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), fsm_output[5]);
  assign mux_tmp_1006 = MUX_s_1_2_2((fsm_output[5]), or_171_cse, or_1391_cse);
  assign not_tmp_436 = ~((fsm_output[6:5]==2'b11));
  assign not_tmp_462 = ~((fsm_output[7]) & (fsm_output[3]) & (fsm_output[4]));
  assign and_dcpl_219 = and_dcpl_121 & and_dcpl_4 & and_dcpl_48;
  assign not_tmp_480 = ~((fsm_output[8:7]!=2'b00) | mux_tmp_886);
  assign and_320_nl = (fsm_output[6:3]==4'b1111);
  assign and_263_nl = (fsm_output[6:5]==2'b11) & and_705_cse;
  assign mux_1157_nl = MUX_s_1_2_2(and_320_nl, and_263_nl, fsm_output[2]);
  assign or_1183_nl = (fsm_output[8]) | ((fsm_output[7]) & mux_1157_nl);
  assign mux_1158_itm = MUX_s_1_2_2(not_tmp_480, or_1183_nl, fsm_output[9]);
  assign nor_tmp_240 = (fsm_output[5]) & (fsm_output[7]) & (fsm_output[9]);
  assign mux_tmp_1159 = MUX_s_1_2_2(nor_tmp_240, (fsm_output[9]), fsm_output[8]);
  assign nor_tmp_241 = ((fsm_output[5]) | (fsm_output[7])) & (fsm_output[9]);
  assign mux_tmp_1160 = MUX_s_1_2_2(nor_tmp_240, nor_tmp_241, fsm_output[8]);
  assign and_tmp_44 = (fsm_output[8]) & nor_tmp_241;
  assign mux_1161_nl = MUX_s_1_2_2(and_tmp_44, mux_tmp_1160, fsm_output[2]);
  assign mux_tmp_1162 = MUX_s_1_2_2(mux_1161_nl, mux_tmp_1159, fsm_output[3]);
  assign not_tmp_482 = ~((fsm_output[5]) | (fsm_output[7]) | (fsm_output[9]));
  assign nor_tmp_244 = ((~ (fsm_output[5])) | (fsm_output[7])) & (fsm_output[9]);
  assign mux_tmp_1164 = MUX_s_1_2_2(not_tmp_482, nor_tmp_244, fsm_output[8]);
  assign nor_329_nl = ~((fsm_output[7]) | (fsm_output[9]));
  assign mux_tmp_1170 = MUX_s_1_2_2(nor_329_nl, nor_tmp_244, fsm_output[8]);
  assign or_tmp_1144 = (fsm_output[8:6]!=3'b000);
  assign and_tmp_45 = (fsm_output[9]) & or_tmp_1144;
  assign and_tmp_46 = (fsm_output[9]) & or_tmp_154;
  assign mux_tmp_1178 = MUX_s_1_2_2((~ or_tmp_1144), or_tmp_154, fsm_output[9]);
  assign or_tmp_1159 = (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[4])) |
      (fsm_output[6]) | (fsm_output[8]);
  assign or_tmp_1165 = (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_tmp_1202 = MUX_s_1_2_2(or_210_cse, or_tmp_1165, fsm_output[9]);
  assign or_tmp_1174 = (fsm_output[9]) | nand_100_cse;
  assign or_tmp_1176 = (fsm_output[9]) | (fsm_output[4]) | (~ (fsm_output[8]));
  assign and_dcpl_226 = and_dcpl_121 & and_dcpl_91 & and_dcpl_48;
  assign or_1268_nl = (~ (fsm_output[9])) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_1268_nl = MUX_s_1_2_2(mux_tmp_1202, or_1268_nl, and_389_cse);
  assign mux_1269_nl = MUX_s_1_2_2(mux_1268_nl, or_tmp_1165, fsm_output[2]);
  assign mux_1270_nl = MUX_s_1_2_2((~ (fsm_output[8])), mux_1269_nl, fsm_output[5]);
  assign or_1267_nl = (or_1391_cse & (fsm_output[9]) & (fsm_output[4])) | (fsm_output[8]);
  assign mux_1266_nl = MUX_s_1_2_2(or_tmp_1174, or_81_cse, or_1391_cse);
  assign mux_1267_nl = MUX_s_1_2_2(or_1267_nl, mux_1266_nl, fsm_output[5]);
  assign mux_1271_nl = MUX_s_1_2_2(mux_1270_nl, mux_1267_nl, fsm_output[6]);
  assign mux_1263_nl = MUX_s_1_2_2(or_tmp_1176, mux_tmp_1202, or_1385_cse);
  assign or_1263_nl = ((fsm_output[2]) & (fsm_output[0]) & (fsm_output[1]) & (fsm_output[9])
      & (fsm_output[4])) | (fsm_output[8]);
  assign mux_1264_nl = MUX_s_1_2_2(mux_1263_nl, or_1263_nl, fsm_output[5]);
  assign mux_1261_nl = MUX_s_1_2_2(or_tmp_1174, or_81_cse, and_477_cse);
  assign mux_1260_nl = MUX_s_1_2_2(or_tmp_1176, mux_tmp_1202, and_483_cse);
  assign mux_1262_nl = MUX_s_1_2_2(mux_1261_nl, mux_1260_nl, fsm_output[5]);
  assign mux_1265_nl = MUX_s_1_2_2(mux_1264_nl, mux_1262_nl, fsm_output[6]);
  assign mux_1272_nl = MUX_s_1_2_2(mux_1271_nl, mux_1265_nl, fsm_output[7]);
  assign nand_227_nl = ~((~((fsm_output[2]) & (fsm_output[9]) & (fsm_output[4])))
      & (fsm_output[8]));
  assign or_1258_nl = (~(((fsm_output[2]) & (fsm_output[9])) | (fsm_output[4])))
      | (fsm_output[8]);
  assign mux_1257_nl = MUX_s_1_2_2(nand_227_nl, or_1258_nl, fsm_output[5]);
  assign or_1256_nl = (or_1392_cse & (fsm_output[4])) | (fsm_output[8]);
  assign mux_1256_nl = MUX_s_1_2_2(or_1256_nl, or_81_cse, fsm_output[5]);
  assign mux_1258_nl = MUX_s_1_2_2(mux_1257_nl, mux_1256_nl, fsm_output[6]);
  assign or_1254_nl = ((and_483_cse | (fsm_output[9])) & (fsm_output[4])) | (fsm_output[8]);
  assign mux_1254_nl = MUX_s_1_2_2(or_tmp_1165, or_1254_nl, fsm_output[5]);
  assign or_1249_nl = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[9]);
  assign mux_1250_nl = MUX_s_1_2_2(or_210_cse, or_tmp_1165, or_1249_nl);
  assign mux_1252_nl = MUX_s_1_2_2(mux_tmp_1202, mux_1250_nl, fsm_output[2]);
  assign mux_1253_nl = MUX_s_1_2_2(or_81_cse, mux_1252_nl, fsm_output[5]);
  assign mux_1255_nl = MUX_s_1_2_2(mux_1254_nl, mux_1253_nl, fsm_output[6]);
  assign mux_1259_nl = MUX_s_1_2_2(mux_1258_nl, mux_1255_nl, fsm_output[7]);
  assign mux_1273_itm = MUX_s_1_2_2(mux_1272_nl, mux_1259_nl, fsm_output[3]);
  assign nor_310_nl = ~((fsm_output[2]) | (fsm_output[7]) | (fsm_output[4]) | (~
      (fsm_output[8])));
  assign and_295_nl = (fsm_output[2]) & (fsm_output[7]) & (fsm_output[4]) & (~ (fsm_output[8]));
  assign mux_1275_nl = MUX_s_1_2_2(nor_310_nl, and_295_nl, fsm_output[9]);
  assign and_294_nl = (~((~ (fsm_output[0])) | (fsm_output[1]) | (~ (fsm_output[6]))))
      & mux_1275_nl;
  assign mux_1276_nl = MUX_s_1_2_2(and_294_nl, mux_29_cse, fsm_output[3]);
  assign not_tmp_513 = MUX_s_1_2_2(nor_601_cse, mux_1276_nl, fsm_output[5]);
  assign or_1304_nl = (~ (fsm_output[7])) | (~ (fsm_output[8])) | (fsm_output[9])
      | (fsm_output[4]);
  assign or_1303_nl = (fsm_output[7]) | nand_89_cse;
  assign mux_1289_nl = MUX_s_1_2_2(or_1304_nl, or_1303_nl, fsm_output[2]);
  assign nor_300_nl = ~((~ (fsm_output[3])) | (fsm_output[6]) | mux_1289_nl);
  assign nor_628_nl = ~((~ (fsm_output[6])) | (fsm_output[3]) | (fsm_output[7]) |
      (fsm_output[2]) | (fsm_output[8]) | nand_230_cse);
  assign mux_1290_nl = MUX_s_1_2_2(nor_300_nl, nor_628_nl, fsm_output[1]);
  assign mux_1291_nl = MUX_s_1_2_2(mux_1290_nl, nor_357_cse, fsm_output[5]);
  assign or_1093_nl = (fsm_output[9]) | (~ (fsm_output[4]));
  assign mux_1286_nl = MUX_s_1_2_2(or_1093_nl, or_83_cse, fsm_output[8]);
  assign or_1295_nl = (fsm_output[7]) | mux_1286_nl;
  assign or_1292_nl = (fsm_output[8:7]!=2'b01) | nand_230_cse;
  assign mux_1287_nl = MUX_s_1_2_2(or_1295_nl, or_1292_nl, fsm_output[2]);
  assign nor_303_nl = ~((fsm_output[3]) | (fsm_output[6]) | mux_1287_nl);
  assign mux_1288_nl = MUX_s_1_2_2(and_502_cse, nor_303_nl, fsm_output[1]);
  assign and_289_nl = (fsm_output[5]) & mux_1288_nl;
  assign not_tmp_523 = MUX_s_1_2_2(mux_1291_nl, and_289_nl, fsm_output[0]);
  assign or_tmp_1261 = (fsm_output[9]) | (~ (fsm_output[6]));
  assign mux_tmp_1305 = MUX_s_1_2_2((~ (fsm_output[6])), (fsm_output[6]), fsm_output[9]);
  assign STAGE_LOOP_i_3_0_sva_mx0c1 = and_dcpl_60 & and_dcpl_57;
  assign VEC_LOOP_j_sva_11_0_mx0c1 = and_dcpl_68 & and_dcpl_57;
  assign and_363_nl = (fsm_output[0]) & (fsm_output[4]) & (fsm_output[6]) & (fsm_output[8])
      & (fsm_output[9]);
  assign mux_874_nl = MUX_s_1_2_2(not_tmp_347, and_363_nl, fsm_output[1]);
  assign and_364_nl = (fsm_output[4]) & (fsm_output[6]) & (fsm_output[8]) & (fsm_output[9]);
  assign mux_875_nl = MUX_s_1_2_2(mux_874_nl, and_364_nl, fsm_output[2]);
  assign mux_876_nl = MUX_s_1_2_2(not_tmp_347, mux_875_nl, fsm_output[3]);
  assign mux_877_nl = MUX_s_1_2_2(mux_876_nl, and_361_cse, fsm_output[5]);
  assign modExp_result_sva_mx0c0 = MUX_s_1_2_2(mux_877_nl, and_369_cse, fsm_output[7]);
  assign nl_STAGE_LOOP_acc_nl = (STAGE_LOOP_i_3_0_sva_2[3:1]) + 3'b011;
  assign STAGE_LOOP_acc_nl = nl_STAGE_LOOP_acc_nl[2:0];
  assign STAGE_LOOP_acc_itm_2_1 = readslicef_3_1_2(STAGE_LOOP_acc_nl);
  assign and_224_m1c = and_dcpl_122 & and_dcpl_82;
  assign and_226_m1c = and_dcpl_129 & and_dcpl_108 & nor_393_cse;
  assign and_229_m1c = and_dcpl_51 & and_dcpl_4 & and_dcpl_56 & and_dcpl_11;
  assign and_230_m1c = and_dcpl_73 & and_dcpl_109;
  assign and_233_m1c = and_dcpl_110 & and_dcpl_4 & and_dcpl_47 & and_dcpl_23;
  assign and_235_m1c = and_dcpl_64 & and_dcpl_14 & and_dcpl_127;
  assign and_237_m1c = and_dcpl_65 & and_dcpl_108 & and_dcpl_23;
  assign and_244_m1c = and_dcpl_60 & and_dcpl_67;
  assign or_1381_nl = (~ (fsm_output[2])) | (~ (fsm_output[8])) | (fsm_output[1])
      | (fsm_output[6]) | not_tmp_400;
  assign or_1382_nl = (fsm_output[2]) | (fsm_output[8]) | (fsm_output[1]) | (~ (fsm_output[6]))
      | (fsm_output[0]) | (fsm_output[5]);
  assign mux_982_nl = MUX_s_1_2_2(or_1381_nl, or_1382_nl, fsm_output[7]);
  assign nor_362_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[1])) | (fsm_output[6])
      | (fsm_output[0]) | (fsm_output[5]));
  assign and_348_nl = (fsm_output[8]) & (fsm_output[1]) & (fsm_output[6]) & (fsm_output[0])
      & (fsm_output[5]);
  assign mux_981_nl = MUX_s_1_2_2(nor_362_nl, and_348_nl, fsm_output[2]);
  assign nand_113_nl = ~((fsm_output[7]) & mux_981_nl);
  assign mux_983_nl = MUX_s_1_2_2(mux_982_nl, nand_113_nl, fsm_output[3]);
  assign nor_361_nl = ~((fsm_output[9]) | mux_983_nl);
  assign nor_363_nl = ~((fsm_output[7]) | (~ (fsm_output[2])) | (fsm_output[8]) |
      (fsm_output[1]) | (~ (fsm_output[6])) | (fsm_output[0]) | (fsm_output[5]));
  assign nor_364_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[8])) | (~ (fsm_output[1]))
      | (fsm_output[6]) | (fsm_output[0]) | (fsm_output[5]));
  assign nor_365_nl = ~((fsm_output[2]) | (fsm_output[8]) | (fsm_output[1]) | (fsm_output[6])
      | not_tmp_400);
  assign mux_979_nl = MUX_s_1_2_2(nor_364_nl, nor_365_nl, fsm_output[7]);
  assign mux_980_nl = MUX_s_1_2_2(nor_363_nl, mux_979_nl, fsm_output[3]);
  assign and_349_nl = (fsm_output[9]) & mux_980_nl;
  assign mux_984_m1c = MUX_s_1_2_2(nor_361_nl, and_349_nl, fsm_output[4]);
  assign and_91_nl = and_dcpl_73 & and_dcpl_70 & nor_393_cse;
  assign nor_553_nl = ~((fsm_output[1]) | (~ (fsm_output[9])) | (~ (fsm_output[0]))
      | (~ (fsm_output[5])) | (fsm_output[2]));
  assign nor_554_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[9])) | (fsm_output[0])
      | (fsm_output[5]) | (~ (fsm_output[2])));
  assign mux_367_nl = MUX_s_1_2_2(nor_553_nl, nor_554_nl, fsm_output[7]);
  assign and_419_nl = (fsm_output[3]) & mux_367_nl;
  assign nor_555_nl = ~((fsm_output[3]) | (~ (fsm_output[7])) | (fsm_output[1]) |
      (fsm_output[9]) | (~ (fsm_output[0])) | (fsm_output[5]) | (~ (fsm_output[2])));
  assign mux_368_nl = MUX_s_1_2_2(and_419_nl, nor_555_nl, fsm_output[4]);
  assign and_421_nl = (fsm_output[7]) & (fsm_output[1]) & (fsm_output[9]) & (fsm_output[0])
      & (fsm_output[5]) & (~ (fsm_output[2]));
  assign nor_556_nl = ~((~ (fsm_output[7])) | (~ (fsm_output[1])) | (fsm_output[9])
      | (fsm_output[0]) | (~ (fsm_output[5])) | (fsm_output[2]));
  assign mux_366_nl = MUX_s_1_2_2(and_421_nl, nor_556_nl, fsm_output[3]);
  assign and_420_nl = (fsm_output[4]) & mux_366_nl;
  assign mux_369_nl = MUX_s_1_2_2(mux_368_nl, and_420_nl, fsm_output[6]);
  assign nor_557_nl = ~((fsm_output[3]) | (~ (fsm_output[7])) | (fsm_output[1]) |
      (fsm_output[9]) | (fsm_output[0]) | (fsm_output[5]) | (~ (fsm_output[2])));
  assign or_269_nl = (~ (fsm_output[9])) | (fsm_output[0]) | (fsm_output[5]) | (fsm_output[2]);
  assign or_268_nl = (fsm_output[9]) | (~ (fsm_output[0])) | (fsm_output[5]) | (~
      (fsm_output[2]));
  assign mux_364_nl = MUX_s_1_2_2(or_269_nl, or_268_nl, fsm_output[1]);
  assign nor_558_nl = ~((~ (fsm_output[3])) | (fsm_output[7]) | mux_364_nl);
  assign mux_365_nl = MUX_s_1_2_2(nor_557_nl, nor_558_nl, fsm_output[4]);
  assign and_422_nl = (fsm_output[6]) & mux_365_nl;
  assign mux_370_nl = MUX_s_1_2_2(mux_369_nl, and_422_nl, fsm_output[8]);
  assign nor_551_nl = ~((fsm_output[5]) | (fsm_output[0]) | (~ (fsm_output[4])));
  assign nor_552_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[0])) | (fsm_output[4]));
  assign mux_371_nl = MUX_s_1_2_2(nor_551_nl, nor_552_nl, fsm_output[6]);
  assign and_96_nl = mux_371_nl & (~ (fsm_output[3])) & (fsm_output[1]) & (fsm_output[2])
      & (fsm_output[7]) & nor_393_cse;
  assign nor_549_nl = ~((~ (fsm_output[7])) | (fsm_output[2]) | (~((fsm_output[5])
      & (fsm_output[0]) & (fsm_output[1]) & (fsm_output[4]))));
  assign nor_550_nl = ~((fsm_output[7]) | (~ (fsm_output[2])) | (fsm_output[5]) |
      (fsm_output[0]) | (fsm_output[1]) | (fsm_output[4]));
  assign mux_372_nl = MUX_s_1_2_2(nor_549_nl, nor_550_nl, fsm_output[8]);
  assign and_104_nl = mux_372_nl & (fsm_output[3]) & (fsm_output[6]) & (~ (fsm_output[9]));
  assign nor_547_nl = ~((~ (fsm_output[6])) | (fsm_output[0]) | (fsm_output[4]));
  assign nor_548_nl = ~((fsm_output[6]) | (~ and_437_cse));
  assign mux_373_nl = MUX_s_1_2_2(nor_547_nl, nor_548_nl, fsm_output[7]);
  assign and_115_nl = mux_373_nl & (~ (fsm_output[3])) & (~ (fsm_output[1])) & (fsm_output[5])
      & (~ (fsm_output[2])) & and_dcpl_11;
  assign nor_545_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[7])) | (~ (fsm_output[6]))
      | (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[4]));
  assign nor_546_nl = ~((fsm_output[8]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[0])
      | (~((fsm_output[1]) & (fsm_output[4]))));
  assign mux_374_nl = MUX_s_1_2_2(nor_545_nl, nor_546_nl, fsm_output[9]);
  assign and_123_nl = mux_374_nl & (~ (fsm_output[3])) & (~ (fsm_output[5])) & (fsm_output[2]);
  assign nor_544_nl = ~((fsm_output[0]) | (fsm_output[4]));
  assign mux_375_nl = MUX_s_1_2_2(nor_544_nl, and_437_cse, fsm_output[6]);
  assign and_136_nl = mux_375_nl & (fsm_output[3]) & (fsm_output[1]) & (fsm_output[5])
      & (~ (fsm_output[2])) & (~ (fsm_output[7])) & and_dcpl_23;
  assign nor_542_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[5])) | (fsm_output[0])
      | (fsm_output[1]) | (fsm_output[3]));
  assign nor_543_nl = ~((fsm_output[6]) | (fsm_output[5]) | (~((fsm_output[0]) &
      (fsm_output[1]) & (fsm_output[3]))));
  assign mux_376_nl = MUX_s_1_2_2(nor_542_nl, nor_543_nl, fsm_output[2]);
  assign and_143_nl = mux_376_nl & (~ (fsm_output[4])) & (fsm_output[7]) & and_dcpl_23;
  assign and_500_nl = (fsm_output[7]) & (fsm_output[5]) & (~ (fsm_output[0])) & (fsm_output[4]);
  assign nor_541_nl = ~((fsm_output[7]) | (fsm_output[5]) | (~ (fsm_output[0])) |
      (fsm_output[4]));
  assign mux_377_nl = MUX_s_1_2_2(and_500_nl, nor_541_nl, fsm_output[8]);
  assign and_152_nl = mux_377_nl & (~ (fsm_output[3])) & (~ (fsm_output[1])) & (fsm_output[6])
      & (fsm_output[2]) & (fsm_output[9]);
  assign vec_rsc_0_0_i_adra_d_pff = MUX1HOT_v_9_11_2(COMP_LOOP_acc_psp_sva_1, (z_out_3[12:4]),
      COMP_LOOP_acc_psp_sva, (COMP_LOOP_acc_10_cse_12_1_1_sva[11:3]), (COMP_LOOP_acc_1_cse_2_sva[11:3]),
      (COMP_LOOP_acc_11_psp_sva[10:2]), (COMP_LOOP_acc_1_cse_4_sva[11:3]), (COMP_LOOP_acc_13_psp_sva[9:1]),
      (COMP_LOOP_acc_1_cse_6_sva[11:3]), (COMP_LOOP_acc_14_psp_sva[10:2]), (COMP_LOOP_acc_1_cse_sva[11:3]),
      {and_dcpl_66 , COMP_LOOP_or_2_cse , and_91_nl , mux_370_nl , and_96_nl , and_104_nl
      , and_115_nl , and_123_nl , and_136_nl , and_143_nl , and_152_nl});
  assign vec_rsc_0_0_i_da_d_pff = modulo_result_mux_1_cse;
  assign or_331_nl = (fsm_output[4]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[0])
      | (fsm_output[9:5]!=5'b10111);
  assign mux_395_nl = MUX_s_1_2_2(or_331_nl, or_329_cse, fsm_output[2]);
  assign mux_396_nl = MUX_s_1_2_2(mux_395_nl, or_tmp_273, fsm_output[1]);
  assign or_326_nl = (fsm_output[4]) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[0])
      | (fsm_output[9:5]!=5'b01010);
  assign mux_393_nl = MUX_s_1_2_2(or_327_cse, or_326_nl, fsm_output[2]);
  assign mux_394_nl = MUX_s_1_2_2(mux_393_nl, mux_392_cse, fsm_output[1]);
  assign mux_397_nl = MUX_s_1_2_2(mux_396_nl, mux_394_nl, fsm_output[3]);
  assign or_321_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b000) | (fsm_output[9:5]!=5'b11010);
  assign mux_388_nl = MUX_s_1_2_2(or_321_nl, or_320_cse, fsm_output[4]);
  assign mux_389_nl = MUX_s_1_2_2(or_tmp_268, mux_388_nl, fsm_output[2]);
  assign or_316_nl = (fsm_output[4]) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b000) |
      (fsm_output[9:5]!=5'b00111);
  assign mux_387_nl = MUX_s_1_2_2(nand_246_cse, or_316_nl, fsm_output[2]);
  assign mux_390_nl = MUX_s_1_2_2(mux_389_nl, mux_387_nl, fsm_output[1]);
  assign or_313_nl = (~ (fsm_output[4])) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b000) | (fsm_output[8:7]!=2'b00);
  assign mux_385_nl = MUX_s_1_2_2(or_313_nl, or_312_cse, fsm_output[2]);
  assign mux_386_nl = MUX_s_1_2_2(or_314_cse, mux_385_nl, fsm_output[1]);
  assign mux_391_nl = MUX_s_1_2_2(mux_390_nl, mux_386_nl, fsm_output[3]);
  assign mux_398_nl = MUX_s_1_2_2(mux_397_nl, mux_391_nl, fsm_output[0]);
  assign or_311_nl = (fsm_output[2]) | (fsm_output[4]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b00)
      | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[9:5]!=5'b10111);
  assign mux_382_nl = MUX_s_1_2_2(or_311_nl, or_tmp_273, fsm_output[1]);
  assign or_305_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[4]) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b00)
      | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[9:5]!=5'b01010);
  assign mux_383_nl = MUX_s_1_2_2(mux_382_nl, or_305_nl, fsm_output[3]);
  assign or_302_nl = (fsm_output[4]) | (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b000) | (fsm_output[9:5]!=5'b11010);
  assign mux_378_nl = MUX_s_1_2_2(or_tmp_268, or_302_nl, fsm_output[2]);
  assign or_301_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b000)
      | (fsm_output[9:5]!=5'b00111);
  assign mux_379_nl = MUX_s_1_2_2(mux_378_nl, or_301_nl, fsm_output[1]);
  assign or_299_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (~ (fsm_output[4]))
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b000)
      | (fsm_output[8:7]!=2'b00);
  assign mux_380_nl = MUX_s_1_2_2(mux_379_nl, or_299_nl, fsm_output[3]);
  assign mux_384_nl = MUX_s_1_2_2(mux_383_nl, mux_380_nl, fsm_output[0]);
  assign or_298_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b000);
  assign mux_399_nl = MUX_s_1_2_2(mux_398_nl, mux_384_nl, or_298_nl);
  assign vec_rsc_0_0_i_wea_d_pff = ~ mux_399_nl;
  assign nor_529_nl = ~((COMP_LOOP_acc_13_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[1])
      | (~ (fsm_output[2])) | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | not_tmp_165);
  assign nor_530_nl = ~((z_out_3[3:1]!=3'b000) | (fsm_output[2]) | (fsm_output[6])
      | (~ (fsm_output[7])));
  assign mux_411_nl = MUX_s_1_2_2(nor_529_nl, nor_530_nl, fsm_output[3]);
  assign nand_15_nl = ~((fsm_output[0]) & mux_411_nl);
  assign or_358_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[7:6]!=2'b01);
  assign or_357_nl = (z_out_3[3:1]!=3'b000) | (fsm_output[7:6]!=2'b00);
  assign mux_410_nl = MUX_s_1_2_2(or_358_nl, or_357_nl, fsm_output[2]);
  assign or_359_nl = (fsm_output[0]) | (fsm_output[3]) | mux_410_nl;
  assign mux_412_nl = MUX_s_1_2_2(nand_15_nl, or_359_nl, fsm_output[5]);
  assign nor_528_nl = ~((fsm_output[9:8]!=2'b01) | mux_412_nl);
  assign nor_531_nl = ~((~ (fsm_output[0])) | (~ (fsm_output[3])) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b00)
      | (~ (fsm_output[2])) | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[7:6]!=2'b10));
  assign nor_532_nl = ~((fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[2]) |
      (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b000)
      | (fsm_output[7:6]!=2'b00));
  assign mux_408_nl = MUX_s_1_2_2(nor_531_nl, nor_532_nl, fsm_output[5]);
  assign and_417_nl = (fsm_output[9]) & mux_408_nl;
  assign nor_533_nl = ~((fsm_output[9]) | (z_out_3[3:1]!=3'b000) | (~ (fsm_output[5]))
      | (fsm_output[0]) | nand_190_cse);
  assign mux_409_nl = MUX_s_1_2_2(and_417_nl, nor_533_nl, fsm_output[8]);
  assign mux_413_nl = MUX_s_1_2_2(nor_528_nl, mux_409_nl, fsm_output[1]);
  assign nor_534_nl = ~((VEC_LOOP_j_sva_11_0[2]) | (~ (fsm_output[5])) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (VEC_LOOP_j_sva_11_0[1]) | (fsm_output[2]) | (VEC_LOOP_j_sva_11_0[0])
      | (fsm_output[7:6]!=2'b00));
  assign or_347_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b000) | (~ (fsm_output[2]))
      | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | not_tmp_165;
  assign or_345_nl = (z_out_3[3:1]!=3'b000) | (fsm_output[2]) | (fsm_output[6]) |
      (~ (fsm_output[7]));
  assign mux_404_nl = MUX_s_1_2_2(or_347_nl, or_345_nl, fsm_output[3]);
  assign nor_535_nl = ~((~ (fsm_output[5])) | (fsm_output[0]) | mux_404_nl);
  assign mux_405_nl = MUX_s_1_2_2(nor_534_nl, nor_535_nl, fsm_output[9]);
  assign nor_536_nl = ~((~ (fsm_output[9])) | (z_out_3[3:1]!=3'b000) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (~ (fsm_output[2])) | (fsm_output[6])
      | (fsm_output[7]));
  assign mux_406_nl = MUX_s_1_2_2(mux_405_nl, nor_536_nl, fsm_output[8]);
  assign or_339_nl = (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b000) | (~ (fsm_output[2]))
      | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (fsm_output[7:6]!=2'b10);
  assign or_337_nl = (z_out_3[3:1]!=3'b000) | (fsm_output[2]) | (~ (fsm_output[6]))
      | (fsm_output[7]);
  assign mux_401_nl = MUX_s_1_2_2(or_339_nl, or_337_nl, fsm_output[3]);
  assign or_340_nl = (fsm_output[0]) | mux_401_nl;
  assign nor_538_nl = ~((COMP_LOOP_acc_11_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | not_tmp_165);
  assign nor_539_nl = ~((z_out_3[3:1]!=3'b000) | (fsm_output[7:6]!=2'b10));
  assign mux_400_nl = MUX_s_1_2_2(nor_538_nl, nor_539_nl, fsm_output[2]);
  assign nand_13_nl = ~((fsm_output[0]) & (fsm_output[3]) & mux_400_nl);
  assign mux_402_nl = MUX_s_1_2_2(or_340_nl, nand_13_nl, fsm_output[5]);
  assign or_332_nl = (fsm_output[5]) | (~ (fsm_output[0])) | (fsm_output[3]) | (z_out_3[3:1]!=3'b000)
      | (fsm_output[2]) | (~ (fsm_output[6])) | (fsm_output[7]);
  assign mux_403_nl = MUX_s_1_2_2(mux_402_nl, or_332_nl, fsm_output[9]);
  assign nor_537_nl = ~((fsm_output[8]) | mux_403_nl);
  assign mux_407_nl = MUX_s_1_2_2(mux_406_nl, nor_537_nl, fsm_output[1]);
  assign vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_413_nl,
      mux_407_nl, fsm_output[4]);
  assign or_398_nl = (fsm_output[4]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b00) | (~
      (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9:5]!=5'b10111);
  assign mux_432_nl = MUX_s_1_2_2(or_398_nl, or_329_cse, fsm_output[2]);
  assign mux_433_nl = MUX_s_1_2_2(mux_432_nl, or_tmp_340, fsm_output[1]);
  assign or_393_nl = (fsm_output[4]) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b00) | (~
      (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9:5]!=5'b01010);
  assign mux_430_nl = MUX_s_1_2_2(or_327_cse, or_393_nl, fsm_output[2]);
  assign mux_431_nl = MUX_s_1_2_2(mux_430_nl, mux_392_cse, fsm_output[1]);
  assign mux_434_nl = MUX_s_1_2_2(mux_433_nl, mux_431_nl, fsm_output[3]);
  assign or_388_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b001) | (fsm_output[9:5]!=5'b11010);
  assign mux_425_nl = MUX_s_1_2_2(or_388_nl, or_320_cse, fsm_output[4]);
  assign mux_426_nl = MUX_s_1_2_2(or_tmp_335, mux_425_nl, fsm_output[2]);
  assign or_383_nl = (fsm_output[4]) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b001) |
      (fsm_output[9:5]!=5'b00111);
  assign mux_424_nl = MUX_s_1_2_2(nand_246_cse, or_383_nl, fsm_output[2]);
  assign mux_427_nl = MUX_s_1_2_2(mux_426_nl, mux_424_nl, fsm_output[1]);
  assign or_380_nl = (~ (fsm_output[4])) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b001) | (fsm_output[8:7]!=2'b00);
  assign mux_422_nl = MUX_s_1_2_2(or_380_nl, or_312_cse, fsm_output[2]);
  assign mux_423_nl = MUX_s_1_2_2(or_314_cse, mux_422_nl, fsm_output[1]);
  assign mux_428_nl = MUX_s_1_2_2(mux_427_nl, mux_423_nl, fsm_output[3]);
  assign mux_435_nl = MUX_s_1_2_2(mux_434_nl, mux_428_nl, fsm_output[0]);
  assign or_378_nl = (fsm_output[2]) | (fsm_output[4]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b00)
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9:5]!=5'b10111);
  assign mux_419_nl = MUX_s_1_2_2(or_378_nl, or_tmp_340, fsm_output[1]);
  assign or_372_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[4]) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b00)
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9:5]!=5'b01010);
  assign mux_420_nl = MUX_s_1_2_2(mux_419_nl, or_372_nl, fsm_output[3]);
  assign or_369_nl = (fsm_output[4]) | (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b001) | (fsm_output[9:5]!=5'b11010);
  assign mux_415_nl = MUX_s_1_2_2(or_tmp_335, or_369_nl, fsm_output[2]);
  assign or_368_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b001)
      | (fsm_output[9:5]!=5'b00111);
  assign mux_416_nl = MUX_s_1_2_2(mux_415_nl, or_368_nl, fsm_output[1]);
  assign or_366_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (~ (fsm_output[4]))
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b001)
      | (fsm_output[8:7]!=2'b00);
  assign mux_417_nl = MUX_s_1_2_2(mux_416_nl, or_366_nl, fsm_output[3]);
  assign mux_421_nl = MUX_s_1_2_2(mux_420_nl, mux_417_nl, fsm_output[0]);
  assign or_365_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b001);
  assign mux_436_nl = MUX_s_1_2_2(mux_435_nl, mux_421_nl, or_365_nl);
  assign vec_rsc_0_1_i_wea_d_pff = ~ mux_436_nl;
  assign or_423_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5:4]!=2'b10) | nand_97_cse;
  assign or_421_nl = (z_out_3[3:1]!=3'b001) | (~ (fsm_output[5])) | (fsm_output[4])
      | (fsm_output[6]) | (~ (fsm_output[8]));
  assign mux_448_nl = MUX_s_1_2_2(or_423_nl, or_421_nl, fsm_output[2]);
  assign nor_514_nl = ~((fsm_output[3]) | mux_448_nl);
  assign nor_515_nl = ~((VEC_LOOP_j_sva_11_0[2]) | (fsm_output[3]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (fsm_output[2]) | (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[6])
      | (fsm_output[8]));
  assign mux_449_nl = MUX_s_1_2_2(nor_514_nl, nor_515_nl, fsm_output[0]);
  assign nor_516_nl = ~((z_out_3[3:1]!=3'b001) | (~ (fsm_output[0])) | (~ (fsm_output[3]))
      | (~ (fsm_output[2])) | (fsm_output[5]) | (~ (fsm_output[4])) | (fsm_output[6])
      | (~ (fsm_output[8])));
  assign mux_450_nl = MUX_s_1_2_2(mux_449_nl, nor_516_nl, fsm_output[9]);
  assign nor_517_nl = ~((COMP_LOOP_acc_13_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[2])) | (fsm_output[5])
      | (fsm_output[4]) | nand_97_cse);
  assign nor_518_nl = ~((z_out_3[3:1]!=3'b001) | (fsm_output[2]) | (fsm_output[5])
      | (fsm_output[4]) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign mux_446_nl = MUX_s_1_2_2(nor_517_nl, nor_518_nl, fsm_output[3]);
  assign and_414_nl = (fsm_output[0]) & mux_446_nl;
  assign or_411_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b001) | (~ (fsm_output[2]))
      | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5])) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[8]);
  assign or_410_nl = (z_out_3[3:1]!=3'b001) | (fsm_output[2]) | (~ (fsm_output[5]))
      | (~ (fsm_output[4])) | (fsm_output[6]) | (fsm_output[8]);
  assign mux_445_nl = MUX_s_1_2_2(or_411_nl, or_410_nl, fsm_output[3]);
  assign nor_519_nl = ~((fsm_output[0]) | mux_445_nl);
  assign mux_447_nl = MUX_s_1_2_2(and_414_nl, nor_519_nl, fsm_output[9]);
  assign mux_451_nl = MUX_s_1_2_2(mux_450_nl, mux_447_nl, fsm_output[7]);
  assign nor_520_nl = ~((z_out_3[3:1]!=3'b001) | (fsm_output[0]) | (~ (fsm_output[3]))
      | (fsm_output[2]) | (fsm_output[5]) | (~ (fsm_output[4])) | (~ (fsm_output[6]))
      | (fsm_output[8]));
  assign nor_521_nl = ~((~ (fsm_output[3])) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[2]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b001)
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[8]));
  assign nor_522_nl = ~((fsm_output[3]) | (z_out_3[3:1]!=3'b001) | (fsm_output[2])
      | (fsm_output[5]) | (~ (fsm_output[4])) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_442_nl = MUX_s_1_2_2(nor_521_nl, nor_522_nl, fsm_output[0]);
  assign mux_443_nl = MUX_s_1_2_2(nor_520_nl, mux_442_nl, fsm_output[9]);
  assign nor_523_nl = ~((COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b001) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[2])) | (fsm_output[5]) | (~ (fsm_output[4])) | (fsm_output[6])
      | (fsm_output[8]));
  assign nor_524_nl = ~((z_out_3[3:1]!=3'b001) | (~ (fsm_output[2])) | (~ (fsm_output[5]))
      | (fsm_output[4]) | nand_97_cse);
  assign mux_439_nl = MUX_s_1_2_2(nor_523_nl, nor_524_nl, fsm_output[3]);
  assign nor_525_nl = ~((z_out_3[3:1]!=3'b001) | (~ (fsm_output[5])) | (~ (fsm_output[4]))
      | (fsm_output[6]) | (fsm_output[8]));
  assign mux_437_nl = MUX_s_1_2_2(and_416_cse, nor_525_nl, fsm_output[2]);
  assign nor_526_nl = ~((~ (fsm_output[2])) | (z_out_3[3:1]!=3'b001) | (~ (fsm_output[5]))
      | (~ (fsm_output[4])) | (fsm_output[6]) | (fsm_output[8]));
  assign or_400_nl = (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b00) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm);
  assign mux_438_nl = MUX_s_1_2_2(mux_437_nl, nor_526_nl, or_400_nl);
  assign and_415_nl = (fsm_output[3]) & mux_438_nl;
  assign mux_440_nl = MUX_s_1_2_2(mux_439_nl, and_415_nl, fsm_output[0]);
  assign nor_527_nl = ~((COMP_LOOP_acc_14_psp_sva[1:0]!=2'b00) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[2])) | (fsm_output[5]) | (fsm_output[4]) | (fsm_output[6])
      | (fsm_output[8]));
  assign mux_441_nl = MUX_s_1_2_2(mux_440_nl, nor_527_nl, fsm_output[9]);
  assign mux_444_nl = MUX_s_1_2_2(mux_443_nl, mux_441_nl, fsm_output[7]);
  assign vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_451_nl,
      mux_444_nl, fsm_output[1]);
  assign or_457_nl = (fsm_output[4]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_11_0[0])
      | (fsm_output[9:5]!=5'b10111);
  assign mux_470_nl = MUX_s_1_2_2(or_457_nl, or_329_cse, fsm_output[2]);
  assign mux_471_nl = MUX_s_1_2_2(mux_470_nl, nand_tmp_18, fsm_output[1]);
  assign or_452_nl = (fsm_output[4]) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_11_0[0])
      | (fsm_output[9:5]!=5'b01010);
  assign mux_468_nl = MUX_s_1_2_2(or_327_cse, or_452_nl, fsm_output[2]);
  assign mux_469_nl = MUX_s_1_2_2(mux_468_nl, mux_392_cse, fsm_output[1]);
  assign mux_472_nl = MUX_s_1_2_2(mux_471_nl, mux_469_nl, fsm_output[3]);
  assign or_447_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b010) | (fsm_output[9:5]!=5'b11010);
  assign mux_463_nl = MUX_s_1_2_2(or_447_nl, or_320_cse, fsm_output[4]);
  assign mux_464_nl = MUX_s_1_2_2(or_tmp_395, mux_463_nl, fsm_output[2]);
  assign or_442_nl = (fsm_output[4]) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b010) |
      (fsm_output[9:5]!=5'b00111);
  assign mux_462_nl = MUX_s_1_2_2(nand_246_cse, or_442_nl, fsm_output[2]);
  assign mux_465_nl = MUX_s_1_2_2(mux_464_nl, mux_462_nl, fsm_output[1]);
  assign or_439_nl = (~ (fsm_output[4])) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b010) | (fsm_output[8:7]!=2'b00);
  assign mux_460_nl = MUX_s_1_2_2(or_439_nl, or_312_cse, fsm_output[2]);
  assign mux_461_nl = MUX_s_1_2_2(or_314_cse, mux_460_nl, fsm_output[1]);
  assign mux_466_nl = MUX_s_1_2_2(mux_465_nl, mux_461_nl, fsm_output[3]);
  assign mux_473_nl = MUX_s_1_2_2(mux_472_nl, mux_466_nl, fsm_output[0]);
  assign or_437_nl = (fsm_output[2]) | (fsm_output[4]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b01)
      | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[9:5]!=5'b10111);
  assign mux_457_nl = MUX_s_1_2_2(or_437_nl, nand_tmp_18, fsm_output[1]);
  assign or_432_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[4]) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b01)
      | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[9:5]!=5'b01010);
  assign mux_458_nl = MUX_s_1_2_2(mux_457_nl, or_432_nl, fsm_output[3]);
  assign or_429_nl = (fsm_output[4]) | (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b010) | (fsm_output[9:5]!=5'b11010);
  assign mux_453_nl = MUX_s_1_2_2(or_tmp_395, or_429_nl, fsm_output[2]);
  assign or_428_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b010)
      | (fsm_output[9:5]!=5'b00111);
  assign mux_454_nl = MUX_s_1_2_2(mux_453_nl, or_428_nl, fsm_output[1]);
  assign or_426_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (~ (fsm_output[4]))
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b010)
      | (fsm_output[8:7]!=2'b00);
  assign mux_455_nl = MUX_s_1_2_2(mux_454_nl, or_426_nl, fsm_output[3]);
  assign mux_459_nl = MUX_s_1_2_2(mux_458_nl, mux_455_nl, fsm_output[0]);
  assign or_425_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b010);
  assign mux_474_nl = MUX_s_1_2_2(mux_473_nl, mux_459_nl, or_425_nl);
  assign vec_rsc_0_2_i_wea_d_pff = ~ mux_474_nl;
  assign or_482_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[5:4]!=2'b10) | nand_97_cse;
  assign or_480_nl = (z_out_3[3:1]!=3'b010) | (~ (fsm_output[5])) | (fsm_output[4])
      | (fsm_output[6]) | (~ (fsm_output[8]));
  assign mux_486_nl = MUX_s_1_2_2(or_482_nl, or_480_nl, fsm_output[2]);
  assign nor_498_nl = ~((fsm_output[3]) | mux_486_nl);
  assign nor_499_nl = ~((VEC_LOOP_j_sva_11_0[2]) | (fsm_output[3]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10)
      | (fsm_output[2]) | (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[6])
      | (fsm_output[8]));
  assign mux_487_nl = MUX_s_1_2_2(nor_498_nl, nor_499_nl, fsm_output[0]);
  assign nor_500_nl = ~((z_out_3[3:1]!=3'b010) | (~ (fsm_output[0])) | (~ (fsm_output[3]))
      | (~ (fsm_output[2])) | (fsm_output[5]) | (~ (fsm_output[4])) | (fsm_output[6])
      | (~ (fsm_output[8])));
  assign mux_488_nl = MUX_s_1_2_2(mux_487_nl, nor_500_nl, fsm_output[9]);
  assign nor_501_nl = ~((COMP_LOOP_acc_13_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10)
      | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[2])) | (fsm_output[5])
      | (fsm_output[4]) | nand_97_cse);
  assign nor_502_nl = ~((z_out_3[3:1]!=3'b010) | (fsm_output[2]) | (fsm_output[5])
      | (fsm_output[4]) | (fsm_output[6]) | (~ (fsm_output[8])));
  assign mux_484_nl = MUX_s_1_2_2(nor_501_nl, nor_502_nl, fsm_output[3]);
  assign and_411_nl = (fsm_output[0]) & mux_484_nl;
  assign or_470_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b010) | (~ (fsm_output[2]))
      | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5])) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[8]);
  assign or_469_nl = (z_out_3[3:1]!=3'b010) | (fsm_output[2]) | (~ (fsm_output[5]))
      | (~ (fsm_output[4])) | (fsm_output[6]) | (fsm_output[8]);
  assign mux_483_nl = MUX_s_1_2_2(or_470_nl, or_469_nl, fsm_output[3]);
  assign nor_503_nl = ~((fsm_output[0]) | mux_483_nl);
  assign mux_485_nl = MUX_s_1_2_2(and_411_nl, nor_503_nl, fsm_output[9]);
  assign mux_489_nl = MUX_s_1_2_2(mux_488_nl, mux_485_nl, fsm_output[7]);
  assign nor_504_nl = ~((z_out_3[3:1]!=3'b010) | (fsm_output[0]) | (~ (fsm_output[3]))
      | (fsm_output[2]) | (fsm_output[5]) | (~ (fsm_output[4])) | (~ (fsm_output[6]))
      | (fsm_output[8]));
  assign nor_505_nl = ~((~ (fsm_output[3])) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[2]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b010)
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[8]));
  assign nor_506_nl = ~((fsm_output[3]) | (z_out_3[3:1]!=3'b010) | (fsm_output[2])
      | (fsm_output[5]) | (~ (fsm_output[4])) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_480_nl = MUX_s_1_2_2(nor_505_nl, nor_506_nl, fsm_output[0]);
  assign mux_481_nl = MUX_s_1_2_2(nor_504_nl, mux_480_nl, fsm_output[9]);
  assign nor_507_nl = ~((COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b010) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[2])) | (fsm_output[5]) | (~ (fsm_output[4])) | (fsm_output[6])
      | (fsm_output[8]));
  assign nor_508_nl = ~((z_out_3[3:1]!=3'b010) | (~ (fsm_output[2])) | (~ (fsm_output[5]))
      | (fsm_output[4]) | nand_97_cse);
  assign mux_477_nl = MUX_s_1_2_2(nor_507_nl, nor_508_nl, fsm_output[3]);
  assign nor_509_nl = ~((z_out_3[3:1]!=3'b010) | (~ (fsm_output[5])) | (~ (fsm_output[4]))
      | (fsm_output[6]) | (fsm_output[8]));
  assign mux_475_nl = MUX_s_1_2_2(and_416_cse, nor_509_nl, fsm_output[2]);
  assign nor_510_nl = ~((~ (fsm_output[2])) | (z_out_3[3:1]!=3'b010) | (~ (fsm_output[5]))
      | (~ (fsm_output[4])) | (fsm_output[6]) | (fsm_output[8]));
  assign or_459_nl = (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm);
  assign mux_476_nl = MUX_s_1_2_2(mux_475_nl, nor_510_nl, or_459_nl);
  assign and_412_nl = (fsm_output[3]) & mux_476_nl;
  assign mux_478_nl = MUX_s_1_2_2(mux_477_nl, and_412_nl, fsm_output[0]);
  assign nor_511_nl = ~((COMP_LOOP_acc_14_psp_sva[1:0]!=2'b01) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[2])) | (fsm_output[5]) | (fsm_output[4]) | (fsm_output[6])
      | (fsm_output[8]));
  assign mux_479_nl = MUX_s_1_2_2(mux_478_nl, nor_511_nl, fsm_output[9]);
  assign mux_482_nl = MUX_s_1_2_2(mux_481_nl, mux_479_nl, fsm_output[7]);
  assign vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_489_nl,
      mux_482_nl, fsm_output[1]);
  assign or_516_nl = (fsm_output[4]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b01) | (~
      (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9:5]!=5'b10111);
  assign mux_508_nl = MUX_s_1_2_2(or_516_nl, or_329_cse, fsm_output[2]);
  assign mux_509_nl = MUX_s_1_2_2(mux_508_nl, nand_tmp_21, fsm_output[1]);
  assign or_511_nl = (fsm_output[4]) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b01) | (~
      (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9:5]!=5'b01010);
  assign mux_506_nl = MUX_s_1_2_2(or_327_cse, or_511_nl, fsm_output[2]);
  assign mux_507_nl = MUX_s_1_2_2(mux_506_nl, mux_392_cse, fsm_output[1]);
  assign mux_510_nl = MUX_s_1_2_2(mux_509_nl, mux_507_nl, fsm_output[3]);
  assign or_506_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b011) | (fsm_output[9:5]!=5'b11010);
  assign mux_501_nl = MUX_s_1_2_2(or_506_nl, or_320_cse, fsm_output[4]);
  assign mux_502_nl = MUX_s_1_2_2(or_tmp_454, mux_501_nl, fsm_output[2]);
  assign or_501_nl = (fsm_output[4]) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b011) |
      (fsm_output[9:5]!=5'b00111);
  assign mux_500_nl = MUX_s_1_2_2(nand_246_cse, or_501_nl, fsm_output[2]);
  assign mux_503_nl = MUX_s_1_2_2(mux_502_nl, mux_500_nl, fsm_output[1]);
  assign or_498_nl = (~ (fsm_output[4])) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b011) | (fsm_output[8:7]!=2'b00);
  assign mux_498_nl = MUX_s_1_2_2(or_498_nl, or_312_cse, fsm_output[2]);
  assign mux_499_nl = MUX_s_1_2_2(or_314_cse, mux_498_nl, fsm_output[1]);
  assign mux_504_nl = MUX_s_1_2_2(mux_503_nl, mux_499_nl, fsm_output[3]);
  assign mux_511_nl = MUX_s_1_2_2(mux_510_nl, mux_504_nl, fsm_output[0]);
  assign or_496_nl = (fsm_output[2]) | (fsm_output[4]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b01)
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9:5]!=5'b10111);
  assign mux_495_nl = MUX_s_1_2_2(or_496_nl, nand_tmp_21, fsm_output[1]);
  assign or_491_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[4]) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b01)
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9:5]!=5'b01010);
  assign mux_496_nl = MUX_s_1_2_2(mux_495_nl, or_491_nl, fsm_output[3]);
  assign or_488_nl = (fsm_output[4]) | (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b011) | (fsm_output[9:5]!=5'b11010);
  assign mux_491_nl = MUX_s_1_2_2(or_tmp_454, or_488_nl, fsm_output[2]);
  assign or_487_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b011)
      | (fsm_output[9:5]!=5'b00111);
  assign mux_492_nl = MUX_s_1_2_2(mux_491_nl, or_487_nl, fsm_output[1]);
  assign or_485_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (~ (fsm_output[4]))
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b011)
      | (fsm_output[8:7]!=2'b00);
  assign mux_493_nl = MUX_s_1_2_2(mux_492_nl, or_485_nl, fsm_output[3]);
  assign mux_497_nl = MUX_s_1_2_2(mux_496_nl, mux_493_nl, fsm_output[0]);
  assign or_484_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b011);
  assign mux_512_nl = MUX_s_1_2_2(mux_511_nl, mux_497_nl, or_484_nl);
  assign vec_rsc_0_3_i_wea_d_pff = ~ mux_512_nl;
  assign nor_485_nl = ~((~((~ (COMP_LOOP_acc_13_psp_sva[0])) & (VEC_LOOP_j_sva_11_0[1])
      & (fsm_output[2]) & (VEC_LOOP_j_sva_11_0[0]) & COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm))
      | not_tmp_165);
  assign nor_486_nl = ~((z_out_3[3:1]!=3'b011) | (fsm_output[2]) | (fsm_output[6])
      | (~ (fsm_output[7])));
  assign mux_524_nl = MUX_s_1_2_2(nor_485_nl, nor_486_nl, fsm_output[3]);
  assign nand_24_nl = ~((fsm_output[0]) & mux_524_nl);
  assign or_543_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[7:6]!=2'b01);
  assign or_542_nl = (z_out_3[3:1]!=3'b011) | (fsm_output[7:6]!=2'b00);
  assign mux_523_nl = MUX_s_1_2_2(or_543_nl, or_542_nl, fsm_output[2]);
  assign or_544_nl = (fsm_output[0]) | (fsm_output[3]) | mux_523_nl;
  assign mux_525_nl = MUX_s_1_2_2(nand_24_nl, or_544_nl, fsm_output[5]);
  assign nor_484_nl = ~((fsm_output[9:8]!=2'b01) | mux_525_nl);
  assign and_499_nl = (fsm_output[0]) & (fsm_output[3]) & (COMP_LOOP_acc_14_psp_sva[1:0]==2'b01)
      & (fsm_output[2]) & (VEC_LOOP_j_sva_11_0[0]) & COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[7:6]==2'b10);
  assign nor_488_nl = ~((fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[2]) |
      (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b011)
      | (fsm_output[7:6]!=2'b00));
  assign mux_521_nl = MUX_s_1_2_2(and_499_nl, nor_488_nl, fsm_output[5]);
  assign and_410_nl = (fsm_output[9]) & mux_521_nl;
  assign nor_489_nl = ~((fsm_output[9]) | (z_out_3[3:1]!=3'b011) | (~ (fsm_output[5]))
      | (fsm_output[0]) | nand_190_cse);
  assign mux_522_nl = MUX_s_1_2_2(and_410_nl, nor_489_nl, fsm_output[8]);
  assign mux_526_nl = MUX_s_1_2_2(nor_484_nl, mux_522_nl, fsm_output[1]);
  assign nor_490_nl = ~((VEC_LOOP_j_sva_11_0[2]) | (~ (fsm_output[5])) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[2]) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (fsm_output[7:6]!=2'b00));
  assign or_532_nl = (~((COMP_LOOP_acc_1_cse_sva[2:0]==3'b011) & (fsm_output[2])
      & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)) | not_tmp_165;
  assign or_530_nl = (z_out_3[3:1]!=3'b011) | (fsm_output[2]) | (fsm_output[6]) |
      (~ (fsm_output[7]));
  assign mux_517_nl = MUX_s_1_2_2(or_532_nl, or_530_nl, fsm_output[3]);
  assign nor_491_nl = ~((~ (fsm_output[5])) | (fsm_output[0]) | mux_517_nl);
  assign mux_518_nl = MUX_s_1_2_2(nor_490_nl, nor_491_nl, fsm_output[9]);
  assign nor_492_nl = ~((~ (fsm_output[9])) | (z_out_3[3:1]!=3'b011) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[3])) | (~ (fsm_output[2])) | (fsm_output[6])
      | (fsm_output[7]));
  assign mux_519_nl = MUX_s_1_2_2(mux_518_nl, nor_492_nl, fsm_output[8]);
  assign nand_232_nl = ~((COMP_LOOP_acc_1_cse_2_sva[2:0]==3'b011) & (fsm_output[2])
      & COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm & (fsm_output[7:6]==2'b10));
  assign or_522_nl = (z_out_3[3:1]!=3'b011) | (fsm_output[2]) | (~ (fsm_output[6]))
      | (fsm_output[7]);
  assign mux_514_nl = MUX_s_1_2_2(nand_232_nl, or_522_nl, fsm_output[3]);
  assign or_525_nl = (fsm_output[0]) | mux_514_nl;
  assign nor_494_nl = ~((~((COMP_LOOP_acc_11_psp_sva[1:0]==2'b01) & (VEC_LOOP_j_sva_11_0[0])
      & COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)) | not_tmp_165);
  assign nor_495_nl = ~((z_out_3[3:1]!=3'b011) | (fsm_output[7:6]!=2'b10));
  assign mux_513_nl = MUX_s_1_2_2(nor_494_nl, nor_495_nl, fsm_output[2]);
  assign nand_22_nl = ~((fsm_output[0]) & (fsm_output[3]) & mux_513_nl);
  assign mux_515_nl = MUX_s_1_2_2(or_525_nl, nand_22_nl, fsm_output[5]);
  assign or_517_nl = (fsm_output[5]) | (~ (fsm_output[0])) | (fsm_output[3]) | (z_out_3[3:1]!=3'b011)
      | (fsm_output[2]) | (~ (fsm_output[6])) | (fsm_output[7]);
  assign mux_516_nl = MUX_s_1_2_2(mux_515_nl, or_517_nl, fsm_output[9]);
  assign nor_493_nl = ~((fsm_output[8]) | mux_516_nl);
  assign mux_520_nl = MUX_s_1_2_2(mux_519_nl, nor_493_nl, fsm_output[1]);
  assign vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_526_nl,
      mux_520_nl, fsm_output[4]);
  assign or_582_nl = (fsm_output[2]) | (fsm_output[4]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b10)
      | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[9:5]!=5'b10111);
  assign mux_546_nl = MUX_s_1_2_2(or_582_nl, or_tmp_535, fsm_output[1]);
  assign or_580_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[4]) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b10)
      | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[9:5]!=5'b01010);
  assign mux_547_nl = MUX_s_1_2_2(mux_546_nl, or_580_nl, fsm_output[3]);
  assign or_579_nl = (fsm_output[4]) | (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b100) | (fsm_output[9:5]!=5'b11010);
  assign mux_543_nl = MUX_s_1_2_2(or_tmp_525, or_579_nl, fsm_output[2]);
  assign or_578_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b100)
      | (fsm_output[9:5]!=5'b00111);
  assign mux_544_nl = MUX_s_1_2_2(mux_543_nl, or_578_nl, fsm_output[1]);
  assign or_576_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (~ (fsm_output[4]))
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b100)
      | (fsm_output[8:7]!=2'b00);
  assign mux_545_nl = MUX_s_1_2_2(mux_544_nl, or_576_nl, fsm_output[3]);
  assign mux_548_nl = MUX_s_1_2_2(mux_547_nl, mux_545_nl, fsm_output[0]);
  assign or_575_nl = (fsm_output[4]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_11_0[0])
      | (fsm_output[9:5]!=5'b10111);
  assign mux_539_nl = MUX_s_1_2_2(or_575_nl, or_329_cse, fsm_output[2]);
  assign mux_540_nl = MUX_s_1_2_2(mux_539_nl, or_tmp_535, fsm_output[1]);
  assign or_566_nl = (fsm_output[4]) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_11_0[0])
      | (fsm_output[9:5]!=5'b01010);
  assign mux_536_nl = MUX_s_1_2_2(or_327_cse, or_566_nl, fsm_output[2]);
  assign mux_537_nl = MUX_s_1_2_2(mux_536_nl, mux_392_cse, fsm_output[1]);
  assign mux_541_nl = MUX_s_1_2_2(mux_540_nl, mux_537_nl, fsm_output[3]);
  assign or_559_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b100) | (fsm_output[9:5]!=5'b11010);
  assign mux_531_nl = MUX_s_1_2_2(or_559_nl, or_320_cse, fsm_output[4]);
  assign mux_532_nl = MUX_s_1_2_2(or_tmp_525, mux_531_nl, fsm_output[2]);
  assign or_554_nl = (fsm_output[4]) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b100) |
      (fsm_output[9:5]!=5'b00111);
  assign mux_530_nl = MUX_s_1_2_2(nand_246_cse, or_554_nl, fsm_output[2]);
  assign mux_533_nl = MUX_s_1_2_2(mux_532_nl, mux_530_nl, fsm_output[1]);
  assign or_551_nl = (~ (fsm_output[4])) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b100) | (fsm_output[8:7]!=2'b00);
  assign mux_528_nl = MUX_s_1_2_2(or_551_nl, or_312_cse, fsm_output[2]);
  assign mux_529_nl = MUX_s_1_2_2(or_314_cse, mux_528_nl, fsm_output[1]);
  assign mux_534_nl = MUX_s_1_2_2(mux_533_nl, mux_529_nl, fsm_output[3]);
  assign mux_542_nl = MUX_s_1_2_2(mux_541_nl, mux_534_nl, fsm_output[0]);
  assign nor_114_nl = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b100));
  assign mux_549_nl = MUX_s_1_2_2(mux_548_nl, mux_542_nl, nor_114_nl);
  assign vec_rsc_0_4_i_wea_d_pff = ~ mux_549_nl;
  assign nor_473_cse = ~((z_out_3[3:1]!=3'b100) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[7])));
  assign nor_474_nl = ~((~ (COMP_LOOP_acc_13_psp_sva[0])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | not_tmp_165);
  assign mux_561_nl = MUX_s_1_2_2(nor_473_cse, nor_474_nl, fsm_output[2]);
  assign nand_27_nl = ~((fsm_output[0]) & mux_561_nl);
  assign or_608_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[7]);
  assign or_607_nl = (z_out_3[3:1]!=3'b100) | (fsm_output[3]) | (fsm_output[6]) |
      (fsm_output[7]);
  assign mux_560_nl = MUX_s_1_2_2(or_608_nl, or_607_nl, fsm_output[2]);
  assign or_609_nl = (fsm_output[0]) | mux_560_nl;
  assign mux_562_nl = MUX_s_1_2_2(nand_27_nl, or_609_nl, fsm_output[5]);
  assign nor_472_nl = ~((fsm_output[9:8]!=2'b01) | mux_562_nl);
  assign nor_475_nl = ~((~ (fsm_output[0])) | (~ (fsm_output[2])) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b10)
      | (VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[3]))
      | (fsm_output[6]) | (~ (fsm_output[7])));
  assign nor_476_nl = ~((fsm_output[0]) | (fsm_output[2]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b100) | (fsm_output[7:6]!=2'b00));
  assign mux_558_nl = MUX_s_1_2_2(nor_475_nl, nor_476_nl, fsm_output[5]);
  assign and_409_nl = (fsm_output[9]) & mux_558_nl;
  assign nor_477_nl = ~((fsm_output[9]) | (z_out_3[3:1]!=3'b100) | (~ (fsm_output[5]))
      | (fsm_output[0]) | nand_190_cse);
  assign mux_559_nl = MUX_s_1_2_2(and_409_nl, nor_477_nl, fsm_output[8]);
  assign mux_563_nl = MUX_s_1_2_2(nor_472_nl, mux_559_nl, fsm_output[1]);
  assign nor_478_nl = ~((~ (VEC_LOOP_j_sva_11_0[2])) | (~ (fsm_output[5])) | (~ (fsm_output[0]))
      | (fsm_output[2]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[6])
      | (fsm_output[7]));
  assign or_598_nl = (z_out_3[3:1]!=3'b100) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[7]));
  assign or_596_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[3]) | not_tmp_165;
  assign mux_554_nl = MUX_s_1_2_2(or_598_nl, or_596_nl, fsm_output[2]);
  assign nor_479_nl = ~((~ (fsm_output[5])) | (fsm_output[0]) | mux_554_nl);
  assign mux_555_nl = MUX_s_1_2_2(nor_478_nl, nor_479_nl, fsm_output[9]);
  assign nor_480_nl = ~((~ (fsm_output[9])) | (z_out_3[3:1]!=3'b100) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[6])
      | (fsm_output[7]));
  assign mux_556_nl = MUX_s_1_2_2(mux_555_nl, nor_480_nl, fsm_output[8]);
  assign or_590_nl = (z_out_3[3:1]!=3'b100) | (~ (fsm_output[3])) | (~ (fsm_output[6]))
      | (fsm_output[7]);
  assign or_589_nl = (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b100) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[7]));
  assign mux_551_nl = MUX_s_1_2_2(or_590_nl, or_589_nl, fsm_output[2]);
  assign or_591_nl = (fsm_output[0]) | mux_551_nl;
  assign nor_482_nl = ~((COMP_LOOP_acc_11_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | nand_168_cse);
  assign mux_550_nl = MUX_s_1_2_2(nor_482_nl, nor_473_cse, fsm_output[2]);
  assign nand_25_nl = ~((fsm_output[0]) & mux_550_nl);
  assign mux_552_nl = MUX_s_1_2_2(or_591_nl, nand_25_nl, fsm_output[5]);
  assign or_583_nl = (fsm_output[5]) | (~ (fsm_output[0])) | (fsm_output[2]) | (fsm_output[3])
      | (z_out_3[3:1]!=3'b100) | (fsm_output[7:6]!=2'b01);
  assign mux_553_nl = MUX_s_1_2_2(mux_552_nl, or_583_nl, fsm_output[9]);
  assign nor_481_nl = ~((fsm_output[8]) | mux_553_nl);
  assign mux_557_nl = MUX_s_1_2_2(mux_556_nl, nor_481_nl, fsm_output[1]);
  assign vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_563_nl,
      mux_557_nl, fsm_output[4]);
  assign or_647_nl = (fsm_output[2]) | (fsm_output[4]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b10)
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9:5]!=5'b10111);
  assign mux_583_nl = MUX_s_1_2_2(or_647_nl, or_tmp_600, fsm_output[1]);
  assign or_645_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[4]) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b10)
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9:5]!=5'b01010);
  assign mux_584_nl = MUX_s_1_2_2(mux_583_nl, or_645_nl, fsm_output[3]);
  assign or_644_nl = (fsm_output[4]) | (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b101) | (fsm_output[9:5]!=5'b11010);
  assign mux_580_nl = MUX_s_1_2_2(or_tmp_590, or_644_nl, fsm_output[2]);
  assign or_643_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b101)
      | (fsm_output[9:5]!=5'b00111);
  assign mux_581_nl = MUX_s_1_2_2(mux_580_nl, or_643_nl, fsm_output[1]);
  assign or_641_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (~ (fsm_output[4]))
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b101)
      | (fsm_output[8:7]!=2'b00);
  assign mux_582_nl = MUX_s_1_2_2(mux_581_nl, or_641_nl, fsm_output[3]);
  assign mux_585_nl = MUX_s_1_2_2(mux_584_nl, mux_582_nl, fsm_output[0]);
  assign or_640_nl = (fsm_output[4]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b10) | (~
      (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9:5]!=5'b10111);
  assign mux_576_nl = MUX_s_1_2_2(or_640_nl, or_329_cse, fsm_output[2]);
  assign mux_577_nl = MUX_s_1_2_2(mux_576_nl, or_tmp_600, fsm_output[1]);
  assign or_631_nl = (fsm_output[4]) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b10) | (~
      (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9:5]!=5'b01010);
  assign mux_573_nl = MUX_s_1_2_2(or_327_cse, or_631_nl, fsm_output[2]);
  assign mux_574_nl = MUX_s_1_2_2(mux_573_nl, mux_392_cse, fsm_output[1]);
  assign mux_578_nl = MUX_s_1_2_2(mux_577_nl, mux_574_nl, fsm_output[3]);
  assign or_624_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b101) | (fsm_output[9:5]!=5'b11010);
  assign mux_568_nl = MUX_s_1_2_2(or_624_nl, or_320_cse, fsm_output[4]);
  assign mux_569_nl = MUX_s_1_2_2(or_tmp_590, mux_568_nl, fsm_output[2]);
  assign or_619_nl = (fsm_output[4]) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b101) |
      (fsm_output[9:5]!=5'b00111);
  assign mux_567_nl = MUX_s_1_2_2(nand_246_cse, or_619_nl, fsm_output[2]);
  assign mux_570_nl = MUX_s_1_2_2(mux_569_nl, mux_567_nl, fsm_output[1]);
  assign or_616_nl = (~ (fsm_output[4])) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b101) | (fsm_output[8:7]!=2'b00);
  assign mux_565_nl = MUX_s_1_2_2(or_616_nl, or_312_cse, fsm_output[2]);
  assign mux_566_nl = MUX_s_1_2_2(or_314_cse, mux_565_nl, fsm_output[1]);
  assign mux_571_nl = MUX_s_1_2_2(mux_570_nl, mux_566_nl, fsm_output[3]);
  assign mux_579_nl = MUX_s_1_2_2(mux_578_nl, mux_571_nl, fsm_output[0]);
  assign nor_120_nl = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b101));
  assign mux_586_nl = MUX_s_1_2_2(mux_585_nl, mux_579_nl, nor_120_nl);
  assign vec_rsc_0_5_i_wea_d_pff = ~ mux_586_nl;
  assign nor_461_cse = ~((z_out_3[3:1]!=3'b101) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[7])));
  assign nor_462_nl = ~((~ (COMP_LOOP_acc_13_psp_sva[0])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | not_tmp_165);
  assign mux_598_nl = MUX_s_1_2_2(nor_461_cse, nor_462_nl, fsm_output[2]);
  assign nand_30_nl = ~((fsm_output[0]) & mux_598_nl);
  assign or_673_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[7]);
  assign or_672_nl = (z_out_3[3:1]!=3'b101) | (fsm_output[3]) | (fsm_output[6]) |
      (fsm_output[7]);
  assign mux_597_nl = MUX_s_1_2_2(or_673_nl, or_672_nl, fsm_output[2]);
  assign or_674_nl = (fsm_output[0]) | mux_597_nl;
  assign mux_599_nl = MUX_s_1_2_2(nand_30_nl, or_674_nl, fsm_output[5]);
  assign nor_460_nl = ~((fsm_output[9:8]!=2'b01) | mux_599_nl);
  assign and_498_nl = (fsm_output[0]) & (fsm_output[2]) & (COMP_LOOP_acc_14_psp_sva[1:0]==2'b10)
      & (VEC_LOOP_j_sva_11_0[0]) & COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm & (fsm_output[3])
      & (~ (fsm_output[6])) & (fsm_output[7]);
  assign nor_464_nl = ~((fsm_output[0]) | (fsm_output[2]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b101) | (fsm_output[7:6]!=2'b00));
  assign mux_595_nl = MUX_s_1_2_2(and_498_nl, nor_464_nl, fsm_output[5]);
  assign and_408_nl = (fsm_output[9]) & mux_595_nl;
  assign nor_465_nl = ~((fsm_output[9]) | (z_out_3[3:1]!=3'b101) | (~ (fsm_output[5]))
      | (fsm_output[0]) | nand_190_cse);
  assign mux_596_nl = MUX_s_1_2_2(and_408_nl, nor_465_nl, fsm_output[8]);
  assign mux_600_nl = MUX_s_1_2_2(nor_460_nl, mux_596_nl, fsm_output[1]);
  assign nor_466_nl = ~((~ (VEC_LOOP_j_sva_11_0[2])) | (~ (fsm_output[5])) | (~ (fsm_output[0]))
      | (fsm_output[2]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[6])
      | (fsm_output[7]));
  assign or_663_nl = (z_out_3[3:1]!=3'b101) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[7]));
  assign or_661_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[3]) | not_tmp_165;
  assign mux_591_nl = MUX_s_1_2_2(or_663_nl, or_661_nl, fsm_output[2]);
  assign nor_467_nl = ~((~ (fsm_output[5])) | (fsm_output[0]) | mux_591_nl);
  assign mux_592_nl = MUX_s_1_2_2(nor_466_nl, nor_467_nl, fsm_output[9]);
  assign nor_468_nl = ~((~ (fsm_output[9])) | (z_out_3[3:1]!=3'b101) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[6])
      | (fsm_output[7]));
  assign mux_593_nl = MUX_s_1_2_2(mux_592_nl, nor_468_nl, fsm_output[8]);
  assign or_655_nl = (z_out_3[3:1]!=3'b101) | (~ (fsm_output[3])) | (~ (fsm_output[6]))
      | (fsm_output[7]);
  assign or_654_nl = (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b101) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[7]));
  assign mux_588_nl = MUX_s_1_2_2(or_655_nl, or_654_nl, fsm_output[2]);
  assign or_656_nl = (fsm_output[0]) | mux_588_nl;
  assign nor_470_nl = ~((~((COMP_LOOP_acc_11_psp_sva[1:0]==2'b10) & (VEC_LOOP_j_sva_11_0[0])
      & COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)) | nand_168_cse);
  assign mux_587_nl = MUX_s_1_2_2(nor_470_nl, nor_461_cse, fsm_output[2]);
  assign nand_28_nl = ~((fsm_output[0]) & mux_587_nl);
  assign mux_589_nl = MUX_s_1_2_2(or_656_nl, nand_28_nl, fsm_output[5]);
  assign or_648_nl = (fsm_output[5]) | (~ (fsm_output[0])) | (fsm_output[2]) | (fsm_output[3])
      | (z_out_3[3:1]!=3'b101) | (fsm_output[7:6]!=2'b01);
  assign mux_590_nl = MUX_s_1_2_2(mux_589_nl, or_648_nl, fsm_output[9]);
  assign nor_469_nl = ~((fsm_output[8]) | mux_590_nl);
  assign mux_594_nl = MUX_s_1_2_2(mux_593_nl, nor_469_nl, fsm_output[1]);
  assign vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_600_nl,
      mux_594_nl, fsm_output[4]);
  assign or_711_nl = (fsm_output[2]) | (fsm_output[4]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b11)
      | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[9:5]!=5'b10111);
  assign mux_620_nl = MUX_s_1_2_2(or_711_nl, nand_tmp_31, fsm_output[1]);
  assign or_709_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[4]) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b11)
      | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[9:5]!=5'b01010);
  assign mux_621_nl = MUX_s_1_2_2(mux_620_nl, or_709_nl, fsm_output[3]);
  assign or_708_nl = (fsm_output[4]) | (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b110) | (fsm_output[9:5]!=5'b11010);
  assign mux_617_nl = MUX_s_1_2_2(or_tmp_655, or_708_nl, fsm_output[2]);
  assign or_707_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b110)
      | (fsm_output[9:5]!=5'b00111);
  assign mux_618_nl = MUX_s_1_2_2(mux_617_nl, or_707_nl, fsm_output[1]);
  assign or_705_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (~ (fsm_output[4]))
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b110)
      | (fsm_output[8:7]!=2'b00);
  assign mux_619_nl = MUX_s_1_2_2(mux_618_nl, or_705_nl, fsm_output[3]);
  assign mux_622_nl = MUX_s_1_2_2(mux_621_nl, mux_619_nl, fsm_output[0]);
  assign or_704_nl = (fsm_output[4]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_11_0[0])
      | (fsm_output[9:5]!=5'b10111);
  assign mux_613_nl = MUX_s_1_2_2(or_704_nl, or_329_cse, fsm_output[2]);
  assign mux_614_nl = MUX_s_1_2_2(mux_613_nl, nand_tmp_31, fsm_output[1]);
  assign or_696_nl = (fsm_output[4]) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_11_0[0])
      | (fsm_output[9:5]!=5'b01010);
  assign mux_610_nl = MUX_s_1_2_2(or_327_cse, or_696_nl, fsm_output[2]);
  assign mux_611_nl = MUX_s_1_2_2(mux_610_nl, mux_392_cse, fsm_output[1]);
  assign mux_615_nl = MUX_s_1_2_2(mux_614_nl, mux_611_nl, fsm_output[3]);
  assign or_689_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b110) | (fsm_output[9:5]!=5'b11010);
  assign mux_605_nl = MUX_s_1_2_2(or_689_nl, or_320_cse, fsm_output[4]);
  assign mux_606_nl = MUX_s_1_2_2(or_tmp_655, mux_605_nl, fsm_output[2]);
  assign or_684_nl = (fsm_output[4]) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b110) |
      (fsm_output[9:5]!=5'b00111);
  assign mux_604_nl = MUX_s_1_2_2(nand_246_cse, or_684_nl, fsm_output[2]);
  assign mux_607_nl = MUX_s_1_2_2(mux_606_nl, mux_604_nl, fsm_output[1]);
  assign or_681_nl = (~ (fsm_output[4])) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (~ (fsm_output[6])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b110) | (fsm_output[8:7]!=2'b00);
  assign mux_602_nl = MUX_s_1_2_2(or_681_nl, or_312_cse, fsm_output[2]);
  assign mux_603_nl = MUX_s_1_2_2(or_314_cse, mux_602_nl, fsm_output[1]);
  assign mux_608_nl = MUX_s_1_2_2(mux_607_nl, mux_603_nl, fsm_output[3]);
  assign mux_616_nl = MUX_s_1_2_2(mux_615_nl, mux_608_nl, fsm_output[0]);
  assign nor_126_nl = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b110));
  assign mux_623_nl = MUX_s_1_2_2(mux_622_nl, mux_616_nl, nor_126_nl);
  assign vec_rsc_0_6_i_wea_d_pff = ~ mux_623_nl;
  assign nor_447_cse = ~((z_out_3[3:1]!=3'b110) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[7])));
  assign nor_448_nl = ~((~ (COMP_LOOP_acc_13_psp_sva[0])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10)
      | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (fsm_output[3]) | not_tmp_165);
  assign mux_635_nl = MUX_s_1_2_2(nor_447_cse, nor_448_nl, fsm_output[2]);
  assign nand_34_nl = ~((fsm_output[0]) & mux_635_nl);
  assign or_737_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[3]) | (~ (fsm_output[6])) | (fsm_output[7]);
  assign or_736_nl = (z_out_3[3:1]!=3'b110) | (fsm_output[3]) | (fsm_output[6]) |
      (fsm_output[7]);
  assign mux_634_nl = MUX_s_1_2_2(or_737_nl, or_736_nl, fsm_output[2]);
  assign or_738_nl = (fsm_output[0]) | mux_634_nl;
  assign mux_636_nl = MUX_s_1_2_2(nand_34_nl, or_738_nl, fsm_output[5]);
  assign nor_446_nl = ~((fsm_output[9:8]!=2'b01) | mux_636_nl);
  assign and_497_nl = (fsm_output[0]) & (fsm_output[2]) & (COMP_LOOP_acc_14_psp_sva[1:0]==2'b11)
      & (~ (VEC_LOOP_j_sva_11_0[0])) & COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm & (fsm_output[3])
      & (~ (fsm_output[6])) & (fsm_output[7]);
  assign nor_450_nl = ~((fsm_output[0]) | (fsm_output[2]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b110) | (fsm_output[7:6]!=2'b00));
  assign mux_632_nl = MUX_s_1_2_2(and_497_nl, nor_450_nl, fsm_output[5]);
  assign and_407_nl = (fsm_output[9]) & mux_632_nl;
  assign nor_451_nl = ~((fsm_output[9]) | (z_out_3[3:1]!=3'b110) | (~ (fsm_output[5]))
      | (fsm_output[0]) | nand_190_cse);
  assign mux_633_nl = MUX_s_1_2_2(and_407_nl, nor_451_nl, fsm_output[8]);
  assign mux_637_nl = MUX_s_1_2_2(nor_446_nl, mux_633_nl, fsm_output[1]);
  assign nor_452_nl = ~((~ (VEC_LOOP_j_sva_11_0[2])) | (~ (fsm_output[5])) | (~ (fsm_output[0]))
      | (fsm_output[2]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[6])
      | (fsm_output[7]));
  assign or_727_nl = (z_out_3[3:1]!=3'b110) | (~ (fsm_output[3])) | (fsm_output[6])
      | (~ (fsm_output[7]));
  assign or_725_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[3]) | not_tmp_165;
  assign mux_628_nl = MUX_s_1_2_2(or_727_nl, or_725_nl, fsm_output[2]);
  assign nor_453_nl = ~((~ (fsm_output[5])) | (fsm_output[0]) | mux_628_nl);
  assign mux_629_nl = MUX_s_1_2_2(nor_452_nl, nor_453_nl, fsm_output[9]);
  assign nor_454_nl = ~((~ (fsm_output[9])) | (z_out_3[3:1]!=3'b110) | (fsm_output[5])
      | (~ (fsm_output[0])) | (~ (fsm_output[2])) | (~ (fsm_output[3])) | (fsm_output[6])
      | (fsm_output[7]));
  assign mux_630_nl = MUX_s_1_2_2(mux_629_nl, nor_454_nl, fsm_output[8]);
  assign or_719_nl = (z_out_3[3:1]!=3'b110) | (~ (fsm_output[3])) | (~ (fsm_output[6]))
      | (fsm_output[7]);
  assign or_718_nl = (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b110) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[7]));
  assign mux_625_nl = MUX_s_1_2_2(or_719_nl, or_718_nl, fsm_output[2]);
  assign or_720_nl = (fsm_output[0]) | mux_625_nl;
  assign nor_456_nl = ~((~((COMP_LOOP_acc_11_psp_sva[1:0]==2'b11) & (~ (VEC_LOOP_j_sva_11_0[0]))
      & COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)) | nand_168_cse);
  assign mux_624_nl = MUX_s_1_2_2(nor_456_nl, nor_447_cse, fsm_output[2]);
  assign nand_32_nl = ~((fsm_output[0]) & mux_624_nl);
  assign mux_626_nl = MUX_s_1_2_2(or_720_nl, nand_32_nl, fsm_output[5]);
  assign or_712_nl = (fsm_output[5]) | (~ (fsm_output[0])) | (fsm_output[2]) | (fsm_output[3])
      | (z_out_3[3:1]!=3'b110) | (fsm_output[7:6]!=2'b01);
  assign mux_627_nl = MUX_s_1_2_2(mux_626_nl, or_712_nl, fsm_output[9]);
  assign nor_455_nl = ~((fsm_output[8]) | mux_627_nl);
  assign mux_631_nl = MUX_s_1_2_2(mux_630_nl, nor_455_nl, fsm_output[1]);
  assign vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_637_nl,
      mux_631_nl, fsm_output[4]);
  assign nand_251_nl = ~((~ (fsm_output[2])) & (~ (fsm_output[4])) & (COMP_LOOP_acc_14_psp_sva[1:0]==2'b11)
      & (VEC_LOOP_j_sva_11_0[0]) & (fsm_output[9:5]==5'b10111));
  assign mux_657_nl = MUX_s_1_2_2(nand_251_nl, nand_tmp_35, fsm_output[1]);
  assign or_773_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[4]) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b11)
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9:5]!=5'b01010);
  assign mux_658_nl = MUX_s_1_2_2(mux_657_nl, or_773_nl, fsm_output[3]);
  assign or_772_nl = (fsm_output[4]) | (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b111) | (fsm_output[9:5]!=5'b11010);
  assign mux_654_nl = MUX_s_1_2_2(or_tmp_719, or_772_nl, fsm_output[2]);
  assign nand_252_nl = ~((fsm_output[2]) & (~ (fsm_output[4])) & (COMP_LOOP_acc_1_cse_2_sva[2:0]==3'b111)
      & (fsm_output[9:5]==5'b00111));
  assign mux_655_nl = MUX_s_1_2_2(mux_654_nl, nand_252_nl, fsm_output[1]);
  assign nand_144_nl = ~((fsm_output[1]) & (~ (fsm_output[2])) & (fsm_output[4])
      & (fsm_output[9]) & (fsm_output[5]) & (fsm_output[6]) & (COMP_LOOP_acc_1_cse_6_sva[2:0]==3'b111)
      & (fsm_output[8:7]==2'b00));
  assign mux_656_nl = MUX_s_1_2_2(mux_655_nl, nand_144_nl, fsm_output[3]);
  assign mux_659_nl = MUX_s_1_2_2(mux_658_nl, mux_656_nl, fsm_output[0]);
  assign nand_250_nl = ~((~ (fsm_output[4])) & (COMP_LOOP_acc_14_psp_sva[1:0]==2'b11)
      & (VEC_LOOP_j_sva_11_0[0]) & (fsm_output[9:5]==5'b10111));
  assign mux_650_nl = MUX_s_1_2_2(nand_250_nl, or_329_cse, fsm_output[2]);
  assign mux_651_nl = MUX_s_1_2_2(mux_650_nl, nand_tmp_35, fsm_output[1]);
  assign or_760_nl = (fsm_output[4]) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b11) | (~
      (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9:5]!=5'b01010);
  assign mux_647_nl = MUX_s_1_2_2(or_327_cse, or_760_nl, fsm_output[2]);
  assign mux_648_nl = MUX_s_1_2_2(mux_647_nl, mux_392_cse, fsm_output[1]);
  assign mux_652_nl = MUX_s_1_2_2(mux_651_nl, mux_648_nl, fsm_output[3]);
  assign nand_147_nl = ~((COMP_LOOP_acc_1_cse_sva[2:0]==3'b111) & (fsm_output[9:5]==5'b11010));
  assign mux_642_nl = MUX_s_1_2_2(nand_147_nl, or_320_cse, fsm_output[4]);
  assign mux_643_nl = MUX_s_1_2_2(or_tmp_719, mux_642_nl, fsm_output[2]);
  assign or_748_nl = (fsm_output[4]) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b111) |
      (fsm_output[9:5]!=5'b00111);
  assign mux_641_nl = MUX_s_1_2_2(nand_246_cse, or_748_nl, fsm_output[2]);
  assign mux_644_nl = MUX_s_1_2_2(mux_643_nl, mux_641_nl, fsm_output[1]);
  assign nand_149_nl = ~((fsm_output[4]) & (fsm_output[9]) & (fsm_output[5]) & (fsm_output[6])
      & (COMP_LOOP_acc_1_cse_6_sva[2:0]==3'b111) & (fsm_output[8:7]==2'b00));
  assign mux_639_nl = MUX_s_1_2_2(nand_149_nl, or_312_cse, fsm_output[2]);
  assign mux_640_nl = MUX_s_1_2_2(or_314_cse, mux_639_nl, fsm_output[1]);
  assign mux_645_nl = MUX_s_1_2_2(mux_644_nl, mux_640_nl, fsm_output[3]);
  assign mux_653_nl = MUX_s_1_2_2(mux_652_nl, mux_645_nl, fsm_output[0]);
  assign and_406_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]==3'b111);
  assign mux_660_nl = MUX_s_1_2_2(mux_659_nl, mux_653_nl, and_406_nl);
  assign vec_rsc_0_7_i_wea_d_pff = ~ mux_660_nl;
  assign and_494_cse = (z_out_3[3:1]==3'b111) & (fsm_output[3]) & (~ (fsm_output[6]))
      & (fsm_output[7]);
  assign nor_435_nl = ~((~((COMP_LOOP_acc_13_psp_sva[0]) & (VEC_LOOP_j_sva_11_0[1:0]==2'b11)
      & COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm & (~ (fsm_output[3])))) | not_tmp_165);
  assign mux_672_nl = MUX_s_1_2_2(and_494_cse, nor_435_nl, fsm_output[2]);
  assign nand_38_nl = ~((fsm_output[0]) & mux_672_nl);
  assign nand_134_nl = ~((COMP_LOOP_acc_1_cse_4_sva[2:0]==3'b111) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      & (~ (fsm_output[3])) & (fsm_output[6]) & (~ (fsm_output[7])));
  assign or_800_nl = (z_out_3[3:1]!=3'b111) | (fsm_output[3]) | (fsm_output[6]) |
      (fsm_output[7]);
  assign mux_671_nl = MUX_s_1_2_2(nand_134_nl, or_800_nl, fsm_output[2]);
  assign or_802_nl = (fsm_output[0]) | mux_671_nl;
  assign mux_673_nl = MUX_s_1_2_2(nand_38_nl, or_802_nl, fsm_output[5]);
  assign nor_433_nl = ~((fsm_output[9:8]!=2'b01) | mux_673_nl);
  assign and_495_nl = (fsm_output[0]) & (fsm_output[2]) & (COMP_LOOP_acc_14_psp_sva[1:0]==2'b11)
      & (VEC_LOOP_j_sva_11_0[0]) & COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm & (fsm_output[3])
      & (~ (fsm_output[6])) & (fsm_output[7]);
  assign nor_437_nl = ~((fsm_output[0]) | (fsm_output[2]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[3])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b111) | (fsm_output[7:6]!=2'b00));
  assign mux_669_nl = MUX_s_1_2_2(and_495_nl, nor_437_nl, fsm_output[5]);
  assign and_404_nl = (fsm_output[9]) & mux_669_nl;
  assign nor_438_nl = ~((fsm_output[9]) | (z_out_3[3:1]!=3'b111) | (~ (fsm_output[5]))
      | (fsm_output[0]) | nand_190_cse);
  assign mux_670_nl = MUX_s_1_2_2(and_404_nl, nor_438_nl, fsm_output[8]);
  assign mux_674_nl = MUX_s_1_2_2(nor_433_nl, mux_670_nl, fsm_output[1]);
  assign nor_439_nl = ~((~ (VEC_LOOP_j_sva_11_0[2])) | (~ (fsm_output[5])) | (~ (fsm_output[0]))
      | (fsm_output[2]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[6])
      | (fsm_output[7]));
  assign nand_237_nl = ~((z_out_3[3:1]==3'b111) & (fsm_output[3]) & (~ (fsm_output[6]))
      & (fsm_output[7]));
  assign or_789_nl = (~((COMP_LOOP_acc_1_cse_sva[2:0]==3'b111) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      & (~ (fsm_output[3])))) | not_tmp_165;
  assign mux_665_nl = MUX_s_1_2_2(nand_237_nl, or_789_nl, fsm_output[2]);
  assign nor_440_nl = ~((~ (fsm_output[5])) | (fsm_output[0]) | mux_665_nl);
  assign mux_666_nl = MUX_s_1_2_2(nor_439_nl, nor_440_nl, fsm_output[9]);
  assign and_405_nl = (fsm_output[9]) & (z_out_3[3:1]==3'b111) & (~ (fsm_output[5]))
      & (fsm_output[0]) & (fsm_output[2]) & (fsm_output[3]) & (~ (fsm_output[6]))
      & (~ (fsm_output[7]));
  assign mux_667_nl = MUX_s_1_2_2(mux_666_nl, and_405_nl, fsm_output[8]);
  assign nand_139_nl = ~((z_out_3[3:1]==3'b111) & (fsm_output[3]) & (fsm_output[6])
      & (~ (fsm_output[7])));
  assign nand_231_nl = ~((COMP_LOOP_acc_1_cse_2_sva[2:0]==3'b111) & COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm
      & (~ (fsm_output[3])) & (~ (fsm_output[6])) & (fsm_output[7]));
  assign mux_662_nl = MUX_s_1_2_2(nand_139_nl, nand_231_nl, fsm_output[2]);
  assign or_784_nl = (fsm_output[0]) | mux_662_nl;
  assign nor_442_nl = ~((~((COMP_LOOP_acc_11_psp_sva[1:0]==2'b11) & (VEC_LOOP_j_sva_11_0[0])
      & COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)) | nand_168_cse);
  assign mux_661_nl = MUX_s_1_2_2(nor_442_nl, and_494_cse, fsm_output[2]);
  assign nand_36_nl = ~((fsm_output[0]) & mux_661_nl);
  assign mux_663_nl = MUX_s_1_2_2(or_784_nl, nand_36_nl, fsm_output[5]);
  assign or_776_nl = (fsm_output[5]) | (~ (fsm_output[0])) | (fsm_output[2]) | (fsm_output[3])
      | (z_out_3[3:1]!=3'b111) | (fsm_output[7:6]!=2'b01);
  assign mux_664_nl = MUX_s_1_2_2(mux_663_nl, or_776_nl, fsm_output[9]);
  assign nor_441_nl = ~((fsm_output[8]) | mux_664_nl);
  assign mux_668_nl = MUX_s_1_2_2(mux_667_nl, nor_441_nl, fsm_output[1]);
  assign vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_674_nl,
      mux_668_nl, fsm_output[4]);
  assign and_dcpl = (~ (fsm_output[6])) & (fsm_output[0]);
  assign and_511_cse = (fsm_output[4]) & (~ (fsm_output[1])) & (~ (fsm_output[3]))
      & nor_393_cse & (~ (fsm_output[7])) & (fsm_output[5]) & (~ (fsm_output[2]))
      & and_dcpl;
  assign and_dcpl_236 = (fsm_output[6]) & (~ (fsm_output[0]));
  assign and_dcpl_238 = ~((fsm_output[7]) | (fsm_output[5]) | (fsm_output[2]));
  assign and_dcpl_240 = (fsm_output[4]) & (fsm_output[1]);
  assign and_dcpl_242 = and_dcpl_240 & (fsm_output[3]) & nor_393_cse;
  assign and_dcpl_243 = and_dcpl_242 & and_dcpl_238 & and_dcpl_236;
  assign and_dcpl_245 = (fsm_output[7]) & (fsm_output[5]) & (fsm_output[2]);
  assign and_dcpl_247 = and_dcpl_242 & and_dcpl_245 & and_dcpl;
  assign and_dcpl_255 = (~ (fsm_output[4])) & (~ (fsm_output[1])) & (fsm_output[3])
      & and_dcpl_11 & (fsm_output[7]) & (~ (fsm_output[5])) & (~ (fsm_output[2]))
      & and_dcpl;
  assign and_dcpl_260 = (~ (fsm_output[4])) & (fsm_output[1]) & (fsm_output[3]) &
      and_dcpl_11 & and_dcpl_245 & and_dcpl_236;
  assign and_dcpl_266 = and_dcpl_240 & (~ (fsm_output[3])) & (fsm_output[9]) & (~
      (fsm_output[8])) & and_dcpl_238 & (fsm_output[6]) & (fsm_output[0]);
  assign and_dcpl_268 = (fsm_output[7]) & (fsm_output[5]);
  assign and_dcpl_269 = and_dcpl_268 & (fsm_output[2]);
  assign and_dcpl_276 = ~((fsm_output[6]) | (fsm_output[0]));
  assign and_dcpl_298 = ~((fsm_output[7]) | (fsm_output[5]));
  assign and_dcpl_324 = nor_tmp & (~ (fsm_output[1])) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (fsm_output[7]) & (fsm_output[5]) & (~ (fsm_output[2])) & (~ (fsm_output[6]))
      & (~ (fsm_output[0]));
  assign and_dcpl_340 = (~ (fsm_output[4])) & (~ (fsm_output[3])) & (~ (fsm_output[1]))
      & nor_393_cse & and_dcpl_238 & and_dcpl;
  assign and_dcpl_345 = nor_tmp & (fsm_output[1]) & nor_393_cse & and_dcpl_238 &
      (fsm_output[6]) & (~ (fsm_output[0]));
  assign and_dcpl_347 = (~ (fsm_output[7])) & (fsm_output[5]);
  assign and_dcpl_349 = and_dcpl_347 & (~ (fsm_output[2])) & and_dcpl;
  assign and_dcpl_354 = and_dcpl_63 & (~ (fsm_output[1])) & nor_393_cse & and_dcpl_349;
  assign or_tmp_1317 = (fsm_output[1]) | (fsm_output[9]) | (~ (fsm_output[4])) |
      (~ (fsm_output[3])) | (fsm_output[8]);
  assign or_1440_cse = (fsm_output[1]) | (~ (fsm_output[9])) | (~ (fsm_output[4]))
      | (fsm_output[3]) | (fsm_output[8]);
  assign nor_635_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[5])) | (fsm_output[0])
      | (~ (fsm_output[1])) | (fsm_output[9]) | (fsm_output[4]) | (fsm_output[3])
      | (~ (fsm_output[8])));
  assign nor_636_nl = ~((fsm_output[6]) | (~ (fsm_output[5])) | (fsm_output[0]) |
      (fsm_output[1]) | (~ (fsm_output[9])) | (fsm_output[4]) | (~ (fsm_output[3]))
      | (fsm_output[8]));
  assign mux_1347_nl = MUX_s_1_2_2(nor_635_nl, nor_636_nl, fsm_output[2]);
  assign mux_1345_nl = MUX_s_1_2_2(or_tmp_1317, or_1440_cse, fsm_output[0]);
  assign nor_637_nl = ~((fsm_output[6:5]!=2'b00) | mux_1345_nl);
  assign or_1438_nl = (~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[9])
      | (fsm_output[4]) | (fsm_output[3]) | (~ (fsm_output[8]));
  assign or_1436_nl = (~ (fsm_output[1])) | (~ (fsm_output[9])) | (~ (fsm_output[4]))
      | (fsm_output[3]) | (fsm_output[8]);
  assign mux_1372_nl = MUX_s_1_2_2(or_1436_nl, or_tmp_1317, fsm_output[0]);
  assign mux_1344_nl = MUX_s_1_2_2(or_1438_nl, mux_1372_nl, fsm_output[5]);
  assign and_nl = (fsm_output[6]) & (~ mux_1344_nl);
  assign mux_1346_nl = MUX_s_1_2_2(nor_637_nl, and_nl, fsm_output[2]);
  assign not_tmp_581 = MUX_s_1_2_2(mux_1347_nl, mux_1346_nl, fsm_output[7]);
  assign and_dcpl_357 = and_dcpl_298 & (~ (fsm_output[2]));
  assign and_dcpl_362 = and_dcpl_110 & nor_393_cse & and_dcpl_357 & and_dcpl_276;
  assign and_dcpl_364 = and_dcpl_357 & and_dcpl_236;
  assign and_dcpl_367 = and_dcpl_59 & nor_393_cse;
  assign and_dcpl_368 = and_dcpl_367 & and_dcpl_364;
  assign and_dcpl_372 = and_dcpl_367 & and_dcpl_269 & and_dcpl;
  assign and_dcpl_379 = (~ (fsm_output[3])) & (~ (fsm_output[4])) & (~ (fsm_output[1]))
      & and_dcpl_11 & and_dcpl_347 & (fsm_output[2]) & and_dcpl_276;
  assign and_dcpl_383 = and_dcpl_100 & (~ (fsm_output[1]));
  assign and_dcpl_385 = and_dcpl_383 & and_dcpl_11 & (fsm_output[7]) & (~ (fsm_output[5]))
      & (~ (fsm_output[2])) & and_dcpl;
  assign and_dcpl_388 = and_dcpl_110 & and_dcpl_11 & and_dcpl_269 & and_dcpl_236;
  assign and_dcpl_394 = and_dcpl_121 & and_dcpl_23 & and_dcpl_357 & (fsm_output[6])
      & (fsm_output[0]);
  assign and_dcpl_399 = and_dcpl_128 & and_dcpl_23 & and_dcpl_268 & (~ (fsm_output[2]))
      & and_dcpl_276;
  assign and_dcpl_404 = and_dcpl_128 & and_369_cse & and_dcpl_298 & (fsm_output[2])
      & and_dcpl;
  assign and_dcpl_406 = and_dcpl_59 & and_369_cse & and_dcpl_364;
  assign and_dcpl_409 = and_dcpl_383 & nor_393_cse & and_dcpl_357 & and_dcpl;
  assign and_dcpl_411 = and_dcpl_121 & nor_393_cse & and_dcpl_349;
  assign or_tmp_1346 = (fsm_output[8]) | (~((fsm_output[2]) & (fsm_output[9]) & (fsm_output[4])
      & (fsm_output[0])));
  assign or_tmp_1348 = (~ (fsm_output[8])) | (fsm_output[2]) | (fsm_output[9]) |
      (fsm_output[4]) | (~ (fsm_output[0]));
  assign or_tmp_1349 = (~ (fsm_output[7])) | (fsm_output[8]) | (fsm_output[2]) |
      (~ (fsm_output[9])) | (~ (fsm_output[4])) | (fsm_output[0]);
  assign not_tmp_600 = ~((fsm_output[4]) & (fsm_output[0]));
  assign operator_64_false_1_or_4_ssc = and_dcpl_354 | not_tmp_581 | and_dcpl_362
      | and_dcpl_409 | and_dcpl_411;
  assign operator_64_false_1_or_5_ssc = and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404;
  assign or_tmp_1365 = (fsm_output[6]) | (~ (fsm_output[3]));
  assign mux_tmp = MUX_s_1_2_2(or_tmp_1365, (fsm_output[6]), fsm_output[1]);
  assign or_tmp_1367 = (fsm_output[6]) | (fsm_output[3]);
  assign nor_tmp_292 = (fsm_output[6]) & (fsm_output[3]);
  assign mux_tmp_1374 = MUX_s_1_2_2(nor_tmp_292, (fsm_output[6]), fsm_output[4]);
  assign mux_tmp_1377 = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), fsm_output[6]);
  assign mux_tmp_1378 = MUX_s_1_2_2(mux_tmp_1377, or_tmp_1365, or_838_cse);
  assign or_tmp_1370 = (~ (fsm_output[6])) | (fsm_output[3]);
  assign nor_tmp_296 = (fsm_output[0]) & (fsm_output[1]) & (fsm_output[6]) & (fsm_output[3]);
  assign or_tmp_1374 = and_389_cse | (fsm_output[6]) | (fsm_output[3]);
  assign mux_tmp_1399 = MUX_s_1_2_2((fsm_output[6]), or_tmp_1367, fsm_output[1]);
  assign or_tmp_1389 = ~((fsm_output[8:5]==4'b0111));
  assign or_tmp_1394 = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[8:7]!=2'b01);
  assign nor_tmp_301 = (fsm_output[8:7]==2'b11);
  assign or_tmp_1401 = (fsm_output[8:6]!=3'b100);
  assign COMP_LOOP_or_40_itm = and_dcpl_243 | and_dcpl_247 | and_dcpl_255 | and_dcpl_260
      | and_dcpl_266;
  assign operator_64_false_1_or_1_itm = and_dcpl_368 | and_dcpl_372 | and_dcpl_379
      | and_dcpl_385 | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404
      | and_dcpl_406;
  always @(posedge clk) begin
    if ( ~ not_tmp_131 ) begin
      p_sva <= p_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( (and_dcpl_51 & and_dcpl_14 & and_dcpl_48) | STAGE_LOOP_i_3_0_sva_mx0c1 )
        begin
      STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(4'b0001, STAGE_LOOP_i_3_0_sva_2, STAGE_LOOP_i_3_0_sva_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ not_tmp_131 ) begin
      r_sva <= r_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_vec_rsc_triosy_0_7_obj_ld_cse <= 1'b0;
      COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= 1'b0;
      modExp_exp_1_0_1_sva_1 <= 1'b0;
      modExp_exp_1_7_1_sva <= 1'b0;
      modExp_exp_1_2_1_sva <= 1'b0;
      modExp_exp_1_1_1_sva <= 1'b0;
      COMP_LOOP_COMP_LOOP_nor_1_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_12_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_124_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_125_itm <= 1'b0;
    end
    else begin
      reg_vec_rsc_triosy_0_7_obj_ld_cse <= and_dcpl_59 & and_dcpl_58 & (fsm_output[6])
          & and_dcpl_140 & (fsm_output[9:8]==2'b11) & (~ STAGE_LOOP_acc_itm_2_1);
      COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= (COMP_LOOP_mux1h_31_nl & (mux_987_nl
          | (fsm_output[0]))) | (mux_1035_nl & (fsm_output[0]));
      modExp_exp_1_0_1_sva_1 <= (COMP_LOOP_mux_nl & (~(mux_1196_nl & (fsm_output[1]))))
          | (~(mux_1249_nl | (fsm_output[1])));
      modExp_exp_1_7_1_sva <= COMP_LOOP_mux1h_52_nl & mux_1285_nl;
      modExp_exp_1_2_1_sva <= COMP_LOOP_mux1h_66_nl & (~ and_dcpl_226);
      modExp_exp_1_1_1_sva <= (COMP_LOOP_mux1h_68_nl & (mux_1323_nl | (fsm_output[9])))
          | mux_1326_nl;
      COMP_LOOP_COMP_LOOP_nor_1_itm <= ~((z_out_3[3:1]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_12_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_12_cse,
          COMP_LOOP_COMP_LOOP_and_11_cse, modExp_while_or_cse);
      COMP_LOOP_COMP_LOOP_and_124_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_13_cse,
          COMP_LOOP_COMP_LOOP_and_12_cse, modExp_while_or_cse);
      COMP_LOOP_COMP_LOOP_and_125_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_37_cse,
          COMP_LOOP_COMP_LOOP_and_13_cse, modExp_while_or_cse);
    end
  end
  always @(posedge clk) begin
    modulo_result_rem_cmp_a <= MUX1HOT_v_64_5_2(z_out_4, operator_64_false_acc_mut_63_0,
        COMP_LOOP_1_acc_8_itm, COMP_LOOP_1_mul_mut, COMP_LOOP_1_acc_5_mut_mx0w5,
        {modulo_result_or_nl , (~ mux_728_nl) , mux_775_nl , mux_795_nl , not_tmp_312});
    modulo_result_rem_cmp_b <= p_sva;
    operator_66_true_div_cmp_a <= MUX_v_65_2_2(z_out_2, ({operator_64_false_acc_mut_64
        , operator_64_false_acc_mut_63_0}), and_dcpl_152);
    operator_66_true_div_cmp_b_9_0 <= MUX_v_10_2_2(STAGE_LOOP_lshift_psp_sva_mx0w0,
        STAGE_LOOP_lshift_psp_sva, and_dcpl_152);
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(nor_659_nl, and_704_nl, fsm_output[9]) ) begin
      STAGE_LOOP_lshift_psp_sva <= STAGE_LOOP_lshift_psp_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ mux_1423_nl ) begin
      operator_64_false_acc_mut_64 <= operator_64_false_mux1h_2_rgt[64];
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_1453_nl, mux_1437_nl, fsm_output[2]) ) begin
      operator_64_false_acc_mut_63_0 <= operator_64_false_mux1h_2_rgt[63:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      VEC_LOOP_j_sva_11_0 <= 12'b000000000000;
    end
    else if ( and_dcpl_156 | VEC_LOOP_j_sva_11_0_mx0c1 ) begin
      VEC_LOOP_j_sva_11_0 <= MUX_v_12_2_2(12'b000000000000, (z_out_3[11:0]), VEC_LOOP_j_sva_11_0_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_k_9_3_sva_5_0 <= 6'b000000;
    end
    else if ( ~(mux_1457_nl | (fsm_output[7])) ) begin
      COMP_LOOP_k_9_3_sva_5_0 <= MUX_v_6_2_2(6'b000000, (COMP_LOOP_k_9_3_sva_2[5:0]),
          nand_263_nl);
    end
  end
  always @(posedge clk) begin
    if ( (modExp_while_and_3 | modExp_while_and_5 | modExp_result_sva_mx0c0 | (~
        mux_885_nl)) & (modExp_result_sva_mx0c0 | modExp_result_and_rgt | modExp_result_and_1_rgt)
        ) begin
      modExp_result_sva <= MUX1HOT_v_64_3_2(64'b0000000000000000000000000000000000000000000000000000000000000001,
          modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w1, {modExp_result_sva_mx0c0
          , modExp_result_and_rgt , modExp_result_and_1_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_10_lpi_4_dfm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( MUX_s_1_2_2((~ mux_913_nl), mux_896_nl, fsm_output[9]) ) begin
      tmp_10_lpi_4_dfm <= MUX1HOT_v_64_9_2(({1'b0 , operator_64_false_slc_modExp_exp_63_1_3}),
          vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d,
          vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_6_i_qa_d, vec_rsc_0_7_i_qa_d,
          {and_dcpl_156 , COMP_LOOP_or_15_nl , COMP_LOOP_or_16_nl , COMP_LOOP_or_17_nl
          , COMP_LOOP_or_18_nl , COMP_LOOP_or_19_nl , COMP_LOOP_or_20_nl , COMP_LOOP_or_21_nl
          , COMP_LOOP_or_22_nl});
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_971_nl, mux_945_nl, fsm_output[9]) ) begin
      COMP_LOOP_1_mul_mut <= MUX1HOT_v_64_13_2(r_sva, modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w1,
          modExp_result_sva, vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d,
          vec_rsc_0_3_i_qa_d, vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_6_i_qa_d,
          vec_rsc_0_7_i_qa_d, z_out_4, {and_238_nl , COMP_LOOP_or_26_nl , COMP_LOOP_or_27_nl
          , not_tmp_374 , COMP_LOOP_or_7_nl , COMP_LOOP_or_8_nl , COMP_LOOP_or_9_nl
          , COMP_LOOP_or_10_nl , COMP_LOOP_or_11_nl , COMP_LOOP_or_12_nl , COMP_LOOP_or_13_nl
          , COMP_LOOP_or_14_nl , mux_48_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_11_itm <= 1'b0;
    end
    else if ( and_dcpl_147 | and_dcpl_219 | and_dcpl_69 | and_dcpl_84 | and_dcpl_93
        | and_dcpl_103 | and_dcpl_112 | and_dcpl_123 | and_dcpl_130 | and_dcpl_138
        ) begin
      COMP_LOOP_COMP_LOOP_and_11_itm <= MUX1HOT_s_1_4_2((~ (z_out_3[63])), (~ (z_out_3[8])),
          COMP_LOOP_COMP_LOOP_and_11_cse, COMP_LOOP_COMP_LOOP_and_37_cse, {and_dcpl_147
          , and_dcpl_219 , and_dcpl_69 , modExp_while_or_cse});
    end
  end
  always @(posedge clk) begin
    if ( mux_1139_nl | not_tmp_312 ) begin
      COMP_LOOP_1_acc_8_itm <= MUX_v_64_2_2(z_out_4, COMP_LOOP_1_acc_8_nl, not_tmp_312);
    end
  end
  always @(posedge clk) begin
    if ( ~((fsm_output!=10'b0000110001)) ) begin
      COMP_LOOP_acc_psp_sva <= COMP_LOOP_acc_psp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_2_sva <= 12'b000000000000;
    end
    else if ( ~(mux_1156_nl & nor_393_cse) ) begin
      COMP_LOOP_acc_1_cse_2_sva <= COMP_LOOP_acc_1_cse_2_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_4_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_86_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_30_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_89_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_32_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_33_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_34_itm <= 1'b0;
    end
    else if ( mux_1158_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_4_itm <= ~((COMP_LOOP_acc_1_cse_2_sva_mx0w0[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_86_itm <= (COMP_LOOP_acc_1_cse_4_sva_1[2:0]==3'b011);
      COMP_LOOP_COMP_LOOP_and_30_itm <= (COMP_LOOP_acc_1_cse_2_sva_mx0w0[2:0]==3'b011);
      COMP_LOOP_COMP_LOOP_and_89_itm <= (COMP_LOOP_acc_1_cse_4_sva_1[2:0]==3'b110);
      COMP_LOOP_COMP_LOOP_and_32_itm <= (COMP_LOOP_acc_1_cse_2_sva_mx0w0[2:0]==3'b101);
      COMP_LOOP_COMP_LOOP_and_33_itm <= (COMP_LOOP_acc_1_cse_2_sva_mx0w0[2:0]==3'b110);
      COMP_LOOP_COMP_LOOP_and_34_itm <= (COMP_LOOP_acc_1_cse_2_sva_mx0w0[2:0]==3'b111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_145_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_1174_nl, mux_1173_nl, fsm_output[4]) ) begin
      COMP_LOOP_COMP_LOOP_and_145_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_145_nl,
          (~ (readslicef_10_1_9(COMP_LOOP_1_acc_nl))), and_dcpl_138);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_6_sva <= 12'b000000000000;
    end
    else if ( MUX_s_1_2_2(mux_tmp_1178, mux_1181_nl, and_314_cse) ) begin
      COMP_LOOP_acc_1_cse_6_sva <= COMP_LOOP_acc_1_cse_6_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_4_sva <= 12'b000000000000;
    end
    else if ( ~(mux_1184_nl & (~ (fsm_output[9]))) ) begin
      COMP_LOOP_acc_1_cse_4_sva <= COMP_LOOP_acc_1_cse_4_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_11_psp_sva <= 11'b00000000000;
    end
    else if ( ~(mux_1186_nl & (~ (fsm_output[9]))) ) begin
      COMP_LOOP_acc_11_psp_sva <= nl_COMP_LOOP_acc_11_psp_sva[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_13_psp_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_480, or_1200_nl, fsm_output[9]) ) begin
      COMP_LOOP_acc_13_psp_sva <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_14_psp_sva <= 11'b00000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_480, or_1201_nl, fsm_output[9]) ) begin
      COMP_LOOP_acc_14_psp_sva <= nl_COMP_LOOP_acc_14_psp_sva[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_sva <= 12'b000000000000;
    end
    else if ( MUX_s_1_2_2(mux_1192_nl, and_369_cse, fsm_output[7]) ) begin
      COMP_LOOP_acc_1_cse_sva <= z_out_2[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_6_1_sva <= 1'b0;
      modExp_exp_1_5_1_sva <= 1'b0;
      modExp_exp_1_4_1_sva <= 1'b0;
      modExp_exp_1_3_1_sva <= 1'b0;
    end
    else if ( mux_1273_itm ) begin
      modExp_exp_1_6_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_3_sva_5_0[3]), modExp_exp_1_7_1_sva,
          (COMP_LOOP_k_9_3_sva_5_0[4]), {and_dcpl_226 , not_tmp_523 , not_tmp_513});
      modExp_exp_1_5_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_3_sva_5_0[2]), modExp_exp_1_6_1_sva,
          (COMP_LOOP_k_9_3_sva_5_0[3]), {and_dcpl_226 , not_tmp_523 , not_tmp_513});
      modExp_exp_1_4_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_3_sva_5_0[1]), modExp_exp_1_5_1_sva,
          (COMP_LOOP_k_9_3_sva_5_0[2]), {and_dcpl_226 , not_tmp_523 , not_tmp_513});
      modExp_exp_1_3_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_3_sva_5_0[0]), modExp_exp_1_4_1_sva,
          (COMP_LOOP_k_9_3_sva_5_0[1]), {and_dcpl_226 , not_tmp_523 , not_tmp_513});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_12_1_1_sva <= 12'b000000000000;
    end
    else if ( COMP_LOOP_or_2_cse ) begin
      COMP_LOOP_acc_10_cse_12_1_1_sva <= z_out_3[12:1];
    end
  end
  always @(posedge clk) begin
    if ( and_dcpl_69 | not_tmp_315 | and_dcpl_84 | and_dcpl_103 | and_dcpl_112 |
        and_dcpl_123 ) begin
      COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm <= MUX_s_1_2_2((z_out[9]), (z_out_3[8]),
          not_tmp_315);
    end
  end
  assign or_864_nl = (fsm_output[9]) | (fsm_output[0]) | (fsm_output[5]) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[4]));
  assign mux_780_nl = MUX_s_1_2_2(mux_tmp_776, or_864_nl, fsm_output[3]);
  assign or_862_nl = (fsm_output[3]) | (fsm_output[9]) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[2]) | not_tmp_297;
  assign mux_781_nl = MUX_s_1_2_2(mux_780_nl, or_862_nl, fsm_output[8]);
  assign and_388_nl = (fsm_output[6]) & (~ mux_781_nl);
  assign or_859_nl = (fsm_output[9]) | (~ (fsm_output[0])) | (~ (fsm_output[5]))
      | (fsm_output[2]) | (fsm_output[7]) | (~ (fsm_output[4]));
  assign or_857_nl = (~ (fsm_output[9])) | (fsm_output[0]) | (~ (fsm_output[5]))
      | (fsm_output[2]) | not_tmp_297;
  assign mux_778_nl = MUX_s_1_2_2(or_859_nl, or_857_nl, fsm_output[3]);
  assign or_855_nl = (fsm_output[9]) | (fsm_output[0]) | (~ (fsm_output[5])) | (~
      (fsm_output[2])) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_777_nl = MUX_s_1_2_2(or_855_nl, mux_tmp_776, fsm_output[3]);
  assign mux_779_nl = MUX_s_1_2_2(mux_778_nl, mux_777_nl, fsm_output[8]);
  assign nor_422_nl = ~((fsm_output[6]) | mux_779_nl);
  assign mux_782_nl = MUX_s_1_2_2(and_388_nl, nor_422_nl, fsm_output[1]);
  assign modulo_result_or_nl = and_dcpl_147 | not_tmp_315 | mux_782_nl;
  assign mux_723_nl = MUX_s_1_2_2(or_tmp_788, nor_tmp, fsm_output[5]);
  assign mux_724_nl = MUX_s_1_2_2(mux_723_nl, mux_tmp_722, fsm_output[6]);
  assign mux_720_nl = MUX_s_1_2_2((~ mux_tmp_719), (fsm_output[4]), fsm_output[5]);
  assign mux_721_nl = MUX_s_1_2_2(mux_720_nl, mux_tmp_718, fsm_output[6]);
  assign mux_725_nl = MUX_s_1_2_2(mux_724_nl, mux_721_nl, fsm_output[2]);
  assign mux_715_nl = MUX_s_1_2_2(and_dcpl_51, or_tmp_788, fsm_output[5]);
  assign mux_714_nl = MUX_s_1_2_2((~ nor_tmp), or_216_cse, fsm_output[5]);
  assign mux_716_nl = MUX_s_1_2_2((~ mux_715_nl), mux_714_nl, fsm_output[6]);
  assign nand_41_nl = ~((fsm_output[5]) & (~ mux_tmp_688));
  assign mux_712_nl = MUX_s_1_2_2((~ and_705_cse), or_tmp_103, fsm_output[5]);
  assign mux_713_nl = MUX_s_1_2_2(nand_41_nl, mux_712_nl, fsm_output[6]);
  assign mux_717_nl = MUX_s_1_2_2(mux_716_nl, mux_713_nl, fsm_output[2]);
  assign mux_726_nl = MUX_s_1_2_2((~ mux_725_nl), mux_717_nl, fsm_output[7]);
  assign mux_706_nl = MUX_s_1_2_2(and_dcpl_50, nor_tmp, fsm_output[1]);
  assign mux_707_nl = MUX_s_1_2_2(mux_tmp_688, mux_706_nl, fsm_output[0]);
  assign mux_708_nl = MUX_s_1_2_2((fsm_output[4]), mux_707_nl, fsm_output[5]);
  assign mux_709_nl = MUX_s_1_2_2(mux_708_nl, mux_tmp_705, fsm_output[6]);
  assign mux_703_nl = MUX_s_1_2_2(and_dcpl_50, and_705_cse, fsm_output[5]);
  assign mux_704_nl = MUX_s_1_2_2(nor_tmp_146, mux_703_nl, fsm_output[6]);
  assign mux_710_nl = MUX_s_1_2_2(mux_709_nl, mux_704_nl, fsm_output[2]);
  assign mux_700_nl = MUX_s_1_2_2(or_216_cse, and_705_cse, fsm_output[5]);
  assign mux_699_nl = MUX_s_1_2_2((~ and_dcpl_59), (fsm_output[4]), fsm_output[5]);
  assign mux_701_nl = MUX_s_1_2_2(mux_700_nl, mux_699_nl, fsm_output[6]);
  assign mux_697_nl = MUX_s_1_2_2((~ mux_696_itm), (fsm_output[4]), fsm_output[5]);
  assign mux_695_nl = MUX_s_1_2_2((~ nor_tmp), or_115_cse, fsm_output[5]);
  assign mux_698_nl = MUX_s_1_2_2(mux_697_nl, mux_695_nl, fsm_output[6]);
  assign mux_702_nl = MUX_s_1_2_2(mux_701_nl, mux_698_nl, fsm_output[2]);
  assign mux_711_nl = MUX_s_1_2_2((~ mux_710_nl), mux_702_nl, fsm_output[7]);
  assign mux_727_nl = MUX_s_1_2_2(mux_726_nl, mux_711_nl, fsm_output[8]);
  assign or_819_nl = (fsm_output[5]) | mux_tmp_156;
  assign mux_690_nl = MUX_s_1_2_2(nor_tmp_23, mux_tmp_689, fsm_output[5]);
  assign mux_691_nl = MUX_s_1_2_2(or_819_nl, mux_690_nl, fsm_output[6]);
  assign mux_686_nl = MUX_s_1_2_2(nor_tmp_23, (~ and_428_cse), fsm_output[5]);
  assign mux_685_nl = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), or_817_cse);
  assign mux_687_nl = MUX_s_1_2_2(mux_686_nl, mux_685_nl, fsm_output[6]);
  assign mux_692_nl = MUX_s_1_2_2(mux_691_nl, mux_687_nl, fsm_output[2]);
  assign nand_40_nl = ~((fsm_output[5]) & (~ mux_tmp_156));
  assign mux_683_nl = MUX_s_1_2_2(nand_40_nl, or_816_cse, fsm_output[6]);
  assign nand_39_nl = ~((fsm_output[5]) & (~ and_462_cse));
  assign or_815_nl = (fsm_output[5]) | (~ or_tmp_113);
  assign mux_682_nl = MUX_s_1_2_2(nand_39_nl, or_815_nl, fsm_output[6]);
  assign mux_684_nl = MUX_s_1_2_2(mux_683_nl, mux_682_nl, fsm_output[2]);
  assign mux_693_nl = MUX_s_1_2_2(mux_692_nl, mux_684_nl, fsm_output[7]);
  assign mux_679_nl = MUX_s_1_2_2(or_115_cse, and_462_cse, fsm_output[5]);
  assign mux_680_nl = MUX_s_1_2_2((~ mux_679_nl), or_1202_cse, fsm_output[6]);
  assign or_808_nl = (fsm_output[5]) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[3])
      | (fsm_output[4]);
  assign mux_678_nl = MUX_s_1_2_2((~ mux_tmp_677), or_808_nl, fsm_output[6]);
  assign mux_681_nl = MUX_s_1_2_2(mux_680_nl, mux_678_nl, fsm_output[2]);
  assign or_813_nl = (fsm_output[7]) | mux_681_nl;
  assign mux_694_nl = MUX_s_1_2_2(mux_693_nl, or_813_nl, fsm_output[8]);
  assign mux_728_nl = MUX_s_1_2_2(mux_727_nl, mux_694_nl, fsm_output[9]);
  assign nand_130_nl = ~((fsm_output[6]) & (fsm_output[1]) & (fsm_output[2]));
  assign mux_770_nl = MUX_s_1_2_2(nand_130_nl, (fsm_output[6]), fsm_output[5]);
  assign nand_44_nl = ~((fsm_output[6]) & not_tmp_274);
  assign mux_769_nl = MUX_s_1_2_2(not_tmp_280, nand_44_nl, fsm_output[5]);
  assign mux_771_nl = MUX_s_1_2_2((~ mux_770_nl), mux_769_nl, fsm_output[7]);
  assign nor_423_nl = ~((fsm_output[6]) | and_382_cse);
  assign mux_767_nl = MUX_s_1_2_2(nor_423_nl, (fsm_output[6]), fsm_output[5]);
  assign mux_768_nl = MUX_s_1_2_2((~ or_tmp_810), mux_767_nl, fsm_output[7]);
  assign mux_772_nl = MUX_s_1_2_2(mux_771_nl, mux_768_nl, fsm_output[4]);
  assign or_850_nl = (fsm_output[6]) | (~ or_1394_cse);
  assign mux_764_nl = MUX_s_1_2_2((~ (fsm_output[6])), or_850_nl, fsm_output[5]);
  assign mux_765_nl = MUX_s_1_2_2((~ mux_tmp_731), mux_764_nl, fsm_output[7]);
  assign mux_762_nl = MUX_s_1_2_2((~ and_382_cse), or_1385_cse, fsm_output[6]);
  assign nor_424_nl = ~((fsm_output[5]) | mux_762_nl);
  assign mux_760_nl = MUX_s_1_2_2((~ (fsm_output[2])), (fsm_output[2]), fsm_output[1]);
  assign and_167_nl = (fsm_output[6]) & mux_760_nl;
  assign mux_761_nl = MUX_s_1_2_2((~ or_tmp_792), and_167_nl, fsm_output[5]);
  assign mux_763_nl = MUX_s_1_2_2(nor_424_nl, mux_761_nl, fsm_output[7]);
  assign mux_766_nl = MUX_s_1_2_2(mux_765_nl, mux_763_nl, fsm_output[4]);
  assign mux_773_nl = MUX_s_1_2_2(mux_772_nl, mux_766_nl, fsm_output[3]);
  assign nand_249_nl = ~((fsm_output[6]) & or_1394_cse);
  assign mux_756_nl = MUX_s_1_2_2((fsm_output[6]), nand_249_nl, fsm_output[5]);
  assign or_848_nl = (fsm_output[5]) | (~ (fsm_output[6])) | (fsm_output[2]);
  assign mux_757_nl = MUX_s_1_2_2(mux_756_nl, or_848_nl, fsm_output[7]);
  assign mux_754_nl = MUX_s_1_2_2((~ (fsm_output[6])), nand_tmp_42, fsm_output[5]);
  assign mux_753_nl = MUX_s_1_2_2((~ (fsm_output[6])), or_tmp_792, fsm_output[5]);
  assign mux_755_nl = MUX_s_1_2_2(mux_754_nl, mux_753_nl, fsm_output[7]);
  assign mux_758_nl = MUX_s_1_2_2(mux_757_nl, mux_755_nl, fsm_output[4]);
  assign or_847_nl = (~ (fsm_output[6])) | (fsm_output[2]);
  assign mux_750_nl = MUX_s_1_2_2(or_847_nl, (fsm_output[6]), fsm_output[5]);
  assign mux_751_nl = MUX_s_1_2_2((~ mux_750_nl), or_tmp_810, fsm_output[7]);
  assign nand_43_nl = ~((~((fsm_output[6:5]!=2'b10))) & not_tmp_274);
  assign or_845_nl = (~ (fsm_output[6])) | (fsm_output[1]) | (fsm_output[2]);
  assign mux_748_nl = MUX_s_1_2_2(or_845_nl, (fsm_output[6]), fsm_output[5]);
  assign mux_749_nl = MUX_s_1_2_2(nand_43_nl, mux_748_nl, fsm_output[7]);
  assign mux_752_nl = MUX_s_1_2_2(mux_751_nl, mux_749_nl, fsm_output[4]);
  assign mux_759_nl = MUX_s_1_2_2(mux_758_nl, mux_752_nl, fsm_output[3]);
  assign mux_774_nl = MUX_s_1_2_2(mux_773_nl, (~ mux_759_nl), fsm_output[8]);
  assign or_843_nl = (fsm_output[6]) | (~ (fsm_output[2]));
  assign mux_743_nl = MUX_s_1_2_2((~ (fsm_output[6])), or_843_nl, fsm_output[5]);
  assign mux_744_nl = MUX_s_1_2_2(nor_425_cse, mux_743_nl, fsm_output[7]);
  assign or_842_nl = (fsm_output[6]) | (~ and_483_cse);
  assign mux_741_nl = MUX_s_1_2_2(or_842_nl, (fsm_output[6]), fsm_output[5]);
  assign mux_739_nl = MUX_s_1_2_2((~ (fsm_output[2])), (fsm_output[2]), and_389_cse);
  assign and_165_nl = (fsm_output[6]) & mux_739_nl;
  assign mux_740_nl = MUX_s_1_2_2(not_tmp_280, and_165_nl, fsm_output[5]);
  assign mux_742_nl = MUX_s_1_2_2((~ mux_741_nl), mux_740_nl, fsm_output[7]);
  assign mux_745_nl = MUX_s_1_2_2(mux_744_nl, mux_742_nl, fsm_output[4]);
  assign mux_736_nl = MUX_s_1_2_2((fsm_output[2]), (~ (fsm_output[2])), or_838_cse);
  assign nor_426_nl = ~((fsm_output[6:5]!=2'b01) | mux_736_nl);
  assign nor_427_nl = ~((fsm_output[6]) | and_483_cse);
  assign mux_735_nl = MUX_s_1_2_2(nor_427_nl, (fsm_output[6]), fsm_output[5]);
  assign mux_737_nl = MUX_s_1_2_2(nor_426_nl, mux_735_nl, fsm_output[7]);
  assign mux_732_nl = MUX_s_1_2_2(not_tmp_274, or_1394_cse, fsm_output[6]);
  assign mux_733_nl = MUX_s_1_2_2((~ (fsm_output[6])), mux_732_nl, fsm_output[5]);
  assign mux_734_nl = MUX_s_1_2_2(mux_733_nl, mux_tmp_731, fsm_output[7]);
  assign mux_738_nl = MUX_s_1_2_2(mux_737_nl, mux_734_nl, fsm_output[4]);
  assign mux_746_nl = MUX_s_1_2_2(mux_745_nl, mux_738_nl, fsm_output[3]);
  assign nor_428_nl = ~((fsm_output[7]) | (fsm_output[5]) | (~ nand_tmp_42));
  assign nor_429_nl = ~((fsm_output[7:5]!=3'b010));
  assign mux_729_nl = MUX_s_1_2_2(nor_428_nl, nor_429_nl, fsm_output[4]);
  assign nor_430_nl = ~((fsm_output[4]) | (fsm_output[7]) | (fsm_output[5]) | (~
      or_tmp_792));
  assign mux_730_nl = MUX_s_1_2_2(mux_729_nl, nor_430_nl, fsm_output[3]);
  assign mux_747_nl = MUX_s_1_2_2(mux_746_nl, mux_730_nl, fsm_output[8]);
  assign mux_775_nl = MUX_s_1_2_2(mux_774_nl, mux_747_nl, fsm_output[9]);
  assign nor_411_nl = ~((fsm_output[8]) | (fsm_output[6]) | (fsm_output[3]) | and_389_cse
      | (fsm_output[2]) | (~ (fsm_output[9])));
  assign and_380_nl = (fsm_output[6]) & (~((fsm_output[3]) & or_1423_cse));
  assign nor_412_nl = ~((fsm_output[6]) | (~((fsm_output[3]) | or_1423_cse)));
  assign mux_792_nl = MUX_s_1_2_2(and_380_nl, nor_412_nl, fsm_output[8]);
  assign mux_793_nl = MUX_s_1_2_2(nor_411_nl, mux_792_nl, fsm_output[5]);
  assign and_381_nl = (fsm_output[1]) & (fsm_output[2]) & (fsm_output[9]);
  assign or_881_nl = and_382_cse | (fsm_output[9]);
  assign mux_790_nl = MUX_s_1_2_2(and_381_nl, or_881_nl, fsm_output[3]);
  assign nor_414_nl = ~((fsm_output[8]) | (~((fsm_output[6]) & mux_790_nl)));
  assign and_383_nl = or_1391_cse & (fsm_output[9]);
  assign or_877_nl = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[2]) | (fsm_output[9]);
  assign mux_789_nl = MUX_s_1_2_2(and_383_nl, or_877_nl, fsm_output[3]);
  assign nor_415_nl = ~((~ (fsm_output[8])) | (fsm_output[6]) | mux_789_nl);
  assign mux_791_nl = MUX_s_1_2_2(nor_414_nl, nor_415_nl, fsm_output[5]);
  assign mux_794_nl = MUX_s_1_2_2(mux_793_nl, mux_791_nl, fsm_output[4]);
  assign nand_127_nl = ~(or_838_cse & (fsm_output[2]) & (fsm_output[9]));
  assign mux_786_nl = MUX_s_1_2_2(or_1392_cse, nand_127_nl, fsm_output[3]);
  assign nand_47_nl = ~((fsm_output[6]) & mux_786_nl);
  assign or_872_nl = (fsm_output[6]) | (~ (fsm_output[3])) | (~ (fsm_output[2]))
      | (fsm_output[9]);
  assign mux_787_nl = MUX_s_1_2_2(nand_47_nl, or_872_nl, fsm_output[8]);
  assign nor_416_nl = ~((fsm_output[5]) | mux_787_nl);
  assign nor_417_nl = ~((~ (fsm_output[6])) | (fsm_output[3]) | (fsm_output[2]) |
      (fsm_output[9]));
  assign nor_418_nl = ~((fsm_output[6]) | ((fsm_output[3:1]==3'b111)) | (fsm_output[9]));
  assign mux_784_nl = MUX_s_1_2_2(nor_417_nl, nor_418_nl, fsm_output[8]);
  assign nor_419_nl = ~((fsm_output[6]) | (~((fsm_output[3]) & or_1394_cse & (fsm_output[9]))));
  assign and_386_nl = (fsm_output[6]) & (~((~((fsm_output[3:0]!=4'b0000))) | (fsm_output[9])));
  assign mux_783_nl = MUX_s_1_2_2(nor_419_nl, and_386_nl, fsm_output[8]);
  assign mux_785_nl = MUX_s_1_2_2(mux_784_nl, mux_783_nl, fsm_output[5]);
  assign mux_788_nl = MUX_s_1_2_2(nor_416_nl, mux_785_nl, fsm_output[4]);
  assign mux_795_nl = MUX_s_1_2_2(mux_794_nl, mux_788_nl, fsm_output[7]);
  assign nl_COMP_LOOP_acc_12_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[9:3]))})
      + conv_u2u_7_8({COMP_LOOP_k_9_3_sva_5_0 , 1'b0}) + 8'b00000001;
  assign COMP_LOOP_acc_12_nl = nl_COMP_LOOP_acc_12_nl[7:0];
  assign COMP_LOOP_and_76_nl = (~ and_dcpl_162) & and_dcpl_156;
  assign mux_1026_nl = MUX_s_1_2_2((~ or_816_cse), (fsm_output[4]), and_389_cse);
  assign mux_1027_nl = MUX_s_1_2_2(mux_1026_nl, (fsm_output[4]), fsm_output[2]);
  assign nor_205_nl = ~((fsm_output[2:0]!=3'b110));
  assign mux_1025_nl = MUX_s_1_2_2((fsm_output[5]), or_816_cse, nor_205_nl);
  assign mux_1028_nl = MUX_s_1_2_2(mux_1027_nl, (~ mux_1025_nl), fsm_output[6]);
  assign mux_1029_nl = MUX_s_1_2_2(mux_1028_nl, nor_425_cse, fsm_output[7]);
  assign or_1072_nl = (~((~ (fsm_output[1])) | (fsm_output[5]))) | (fsm_output[4]);
  assign mux_1021_nl = MUX_s_1_2_2(or_247_cse, mux_tmp_997, or_838_cse);
  assign mux_1022_nl = MUX_s_1_2_2(or_1072_nl, mux_1021_nl, fsm_output[2]);
  assign mux_1023_nl = MUX_s_1_2_2(mux_1022_nl, (~ mux_tmp_1006), fsm_output[6]);
  assign mux_1019_nl = MUX_s_1_2_2(or_171_cse, (~ mux_tmp_997), and_483_cse);
  assign and_252_nl = (fsm_output[2]) & or_838_cse & (fsm_output[5:4]==2'b11);
  assign mux_1020_nl = MUX_s_1_2_2(mux_1019_nl, and_252_nl, fsm_output[6]);
  assign mux_1024_nl = MUX_s_1_2_2(mux_1023_nl, mux_1020_nl, fsm_output[7]);
  assign mux_1030_nl = MUX_s_1_2_2(mux_1029_nl, mux_1024_nl, fsm_output[3]);
  assign and_340_nl = (fsm_output[0]) & (fsm_output[1]) & (fsm_output[5]) & (~ (fsm_output[4]));
  assign nor_351_nl = ~((fsm_output[0]) | (fsm_output[1]) | (~ (fsm_output[5])) |
      (fsm_output[4]));
  assign mux_1015_nl = MUX_s_1_2_2(and_340_nl, nor_351_nl, fsm_output[2]);
  assign nor_352_nl = ~((fsm_output[2]) | (fsm_output[1]) | (~ (fsm_output[5])) |
      (fsm_output[4]));
  assign mux_1016_nl = MUX_s_1_2_2(mux_1015_nl, nor_352_nl, fsm_output[6]);
  assign mux_1013_nl = MUX_s_1_2_2(mux_tmp_997, and_314_cse, and_477_cse);
  assign mux_1014_nl = MUX_s_1_2_2(or_171_cse, mux_1013_nl, fsm_output[6]);
  assign mux_1017_nl = MUX_s_1_2_2(mux_1016_nl, mux_1014_nl, fsm_output[7]);
  assign mux_1011_nl = MUX_s_1_2_2(and_314_cse, (fsm_output[5]), or_838_cse);
  assign mux_1012_nl = MUX_s_1_2_2(and_314_cse, mux_1011_nl, fsm_output[2]);
  assign and_251_nl = (fsm_output[7]) & (~((fsm_output[6]) & (~ mux_1012_nl)));
  assign mux_1018_nl = MUX_s_1_2_2(mux_1017_nl, and_251_nl, fsm_output[3]);
  assign mux_1031_nl = MUX_s_1_2_2(mux_1030_nl, (~ mux_1018_nl), fsm_output[8]);
  assign mux_1007_nl = MUX_s_1_2_2(and_314_cse, (~ mux_tmp_1006), fsm_output[6]);
  assign mux_1003_nl = MUX_s_1_2_2((fsm_output[5]), or_171_cse, or_838_cse);
  assign mux_1002_nl = MUX_s_1_2_2(or_171_cse, (~ mux_tmp_997), and_389_cse);
  assign mux_1004_nl = MUX_s_1_2_2(mux_1003_nl, mux_1002_nl, fsm_output[2]);
  assign or_1061_nl = (fsm_output[2:1]!=2'b10) | (~ and_314_cse);
  assign mux_1005_nl = MUX_s_1_2_2(mux_1004_nl, or_1061_nl, fsm_output[6]);
  assign mux_1008_nl = MUX_s_1_2_2(mux_1007_nl, mux_1005_nl, fsm_output[7]);
  assign mux_999_nl = MUX_s_1_2_2(and_314_cse, (fsm_output[5]), fsm_output[2]);
  assign mux_1000_nl = MUX_s_1_2_2(mux_999_nl, (~ or_171_cse), fsm_output[6]);
  assign mux_998_nl = MUX_s_1_2_2((~ mux_tmp_997), or_171_cse, or_1385_cse);
  assign or_1059_nl = (fsm_output[6]) | mux_998_nl;
  assign mux_1001_nl = MUX_s_1_2_2(mux_1000_nl, or_1059_nl, fsm_output[7]);
  assign mux_1009_nl = MUX_s_1_2_2(mux_1008_nl, mux_1001_nl, fsm_output[3]);
  assign nor_353_nl = ~((fsm_output[7:5]!=3'b000));
  assign mux_995_nl = MUX_s_1_2_2((fsm_output[5]), or_171_cse, fsm_output[2]);
  assign nor_354_nl = ~((fsm_output[7:6]!=2'b00) | mux_995_nl);
  assign mux_996_nl = MUX_s_1_2_2(nor_353_nl, nor_354_nl, fsm_output[3]);
  assign mux_1010_nl = MUX_s_1_2_2(mux_1009_nl, mux_996_nl, fsm_output[8]);
  assign mux_1032_nl = MUX_s_1_2_2(mux_1031_nl, mux_1010_nl, fsm_output[9]);
  assign COMP_LOOP_mux1h_31_nl = MUX1HOT_s_1_7_2((operator_66_true_div_cmp_z[0]),
      (tmp_10_lpi_4_dfm[0]), (z_out_3[6]), modExp_exp_1_0_1_sva_1, COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm,
      (readslicef_8_1_7(COMP_LOOP_acc_12_nl)), (z_out_2[6]), {COMP_LOOP_and_76_nl
      , and_dcpl_162 , and_dcpl_66 , not_tmp_414 , mux_1032_nl , and_dcpl_93 , and_dcpl_130});
  assign or_1432_nl = (~ (fsm_output[8])) | (~ (fsm_output[1])) | (fsm_output[5])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_406;
  assign or_1040_nl = (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[7]))
      | (fsm_output[2]) | (fsm_output[6]);
  assign or_1039_nl = (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_406;
  assign mux_985_nl = MUX_s_1_2_2(or_1040_nl, or_1039_nl, fsm_output[5]);
  assign or_1037_nl = (~ (fsm_output[5])) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[7])
      | (fsm_output[2]) | (fsm_output[6]);
  assign mux_986_nl = MUX_s_1_2_2(mux_985_nl, or_1037_nl, fsm_output[1]);
  assign or_1433_nl = (fsm_output[8]) | mux_986_nl;
  assign mux_987_nl = MUX_s_1_2_2(or_1432_nl, or_1433_nl, fsm_output[4]);
  assign nand_108_nl = ~((fsm_output[9]) & (fsm_output[3]) & (fsm_output[1]) & (~
      (fsm_output[6])) & (fsm_output[5]));
  assign or_1082_nl = (fsm_output[9]) | (fsm_output[3]) | (fsm_output[1]) | not_tmp_436;
  assign mux_1034_nl = MUX_s_1_2_2(nand_108_nl, or_1082_nl, fsm_output[8]);
  assign nor_347_nl = ~((fsm_output[4]) | (fsm_output[7]) | mux_1034_nl);
  assign or_1078_nl = (fsm_output[3]) | (~ (fsm_output[1])) | (fsm_output[6]) | (fsm_output[5]);
  assign or_1077_nl = (fsm_output[3]) | (fsm_output[1]) | not_tmp_436;
  assign mux_1033_nl = MUX_s_1_2_2(or_1078_nl, or_1077_nl, fsm_output[9]);
  assign nor_348_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[7])) | (fsm_output[8])
      | mux_1033_nl);
  assign mux_1035_nl = MUX_s_1_2_2(nor_347_nl, nor_348_nl, fsm_output[2]);
  assign nor_316_nl = ~((fsm_output[5]) | (fsm_output[2]) | (~ (fsm_output[7])) |
      (~ (fsm_output[8])) | (fsm_output[4]));
  assign nor_317_nl = ~((fsm_output[5]) | (~ (fsm_output[2])) | (fsm_output[7]) |
      nand_100_cse);
  assign mux_1243_nl = MUX_s_1_2_2(nor_316_nl, nor_317_nl, fsm_output[9]);
  assign nor_318_nl = ~((fsm_output[9]) | (~ (fsm_output[5])) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[4])));
  assign mux_1244_nl = MUX_s_1_2_2(mux_1243_nl, nor_318_nl, fsm_output[1]);
  assign and_306_nl = (fsm_output[3]) & mux_1244_nl;
  assign nor_319_nl = ~((fsm_output[3]) | (~ (fsm_output[1])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[8]) | (~
      (fsm_output[4])));
  assign mux_1245_nl = MUX_s_1_2_2(and_306_nl, nor_319_nl, fsm_output[6]);
  assign nor_320_nl = ~((~ (fsm_output[5])) | (fsm_output[2]) | (fsm_output[7]) |
      (~ (fsm_output[8])) | (fsm_output[4]));
  assign and_493_nl = (fsm_output[5]) & (fsm_output[2]) & (fsm_output[7]) & (~ (fsm_output[8]))
      & (fsm_output[4]);
  assign mux_1241_nl = MUX_s_1_2_2(nor_320_nl, and_493_nl, fsm_output[9]);
  assign and_307_nl = (~((fsm_output[3]) | (~ (fsm_output[1])))) & mux_1241_nl;
  assign or_1229_nl = (fsm_output[2]) | (fsm_output[7]) | (fsm_output[8]) | (~ (fsm_output[4]));
  assign nand_95_nl = ~((fsm_output[2]) & (fsm_output[7]) & (fsm_output[8]) & (~
      (fsm_output[4])));
  assign mux_1240_nl = MUX_s_1_2_2(or_1229_nl, nand_95_nl, fsm_output[5]);
  assign nor_322_nl = ~((~ (fsm_output[3])) | (fsm_output[1]) | (fsm_output[9]) |
      mux_1240_nl);
  assign mux_1242_nl = MUX_s_1_2_2(and_307_nl, nor_322_nl, fsm_output[6]);
  assign mux_1246_nl = MUX_s_1_2_2(mux_1245_nl, mux_1242_nl, fsm_output[0]);
  assign COMP_LOOP_mux_nl = MUX_s_1_2_2(modExp_exp_1_0_1_sva_1, modExp_exp_1_1_1_sva,
      mux_1246_nl);
  assign or_1210_nl = (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[4])
      | (fsm_output[6]) | (fsm_output[8]);
  assign mux_1195_nl = MUX_s_1_2_2(or_tmp_1159, or_1210_nl, fsm_output[0]);
  assign nor_324_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | mux_1195_nl);
  assign or_1208_nl = (fsm_output[3]) | (fsm_output[9]) | (fsm_output[4]) | nand_97_cse;
  assign mux_1194_nl = MUX_s_1_2_2(or_1208_nl, or_tmp_1159, fsm_output[0]);
  assign nor_325_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | mux_1194_nl);
  assign mux_1196_nl = MUX_s_1_2_2(nor_324_nl, nor_325_nl, fsm_output[2]);
  assign or_1430_nl = (fsm_output[7]) | (~ (fsm_output[8])) | (fsm_output[9]) | (~
      (fsm_output[0])) | (fsm_output[2]) | (fsm_output[3]) | not_tmp_436;
  assign or_1245_nl = (fsm_output[0]) | (~((fsm_output[2]) & (fsm_output[3]) & (fsm_output[5])
      & (fsm_output[6])));
  assign or_1244_nl = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[5]) | (fsm_output[6]);
  assign or_1243_nl = (fsm_output[3:2]!=2'b01) | not_tmp_436;
  assign mux_1247_nl = MUX_s_1_2_2(or_1244_nl, or_1243_nl, fsm_output[0]);
  assign mux_1248_nl = MUX_s_1_2_2(or_1245_nl, mux_1247_nl, fsm_output[9]);
  assign or_1431_nl = (fsm_output[8:7]!=2'b01) | mux_1248_nl;
  assign mux_1249_nl = MUX_s_1_2_2(or_1430_nl, or_1431_nl, fsm_output[4]);
  assign COMP_LOOP_mux1h_52_nl = MUX1HOT_s_1_4_2((COMP_LOOP_k_9_3_sva_5_0[4]), modExp_exp_1_1_1_sva,
      modExp_exp_1_7_1_sva, (COMP_LOOP_k_9_3_sva_5_0[5]), {and_dcpl_226 , and_dcpl_219
      , (~ mux_1273_itm) , not_tmp_513});
  assign nor_304_nl = ~((~ (fsm_output[7])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[4]));
  assign nor_305_nl = ~((fsm_output[7]) | nand_89_cse);
  assign mux_1283_nl = MUX_s_1_2_2(nor_304_nl, nor_305_nl, fsm_output[2]);
  assign nand_259_nl = ~((~((fsm_output[5]) | (fsm_output[0]) | (~ (fsm_output[3]))))
      & mux_1283_nl);
  assign nand_260_nl = ~((fsm_output[5]) & (fsm_output[0]) & (fsm_output[3]) & (fsm_output[2])
      & (fsm_output[7]) & (~ (fsm_output[9])) & (fsm_output[8]) & (~ (fsm_output[4])));
  assign mux_1284_nl = MUX_s_1_2_2(nand_259_nl, nand_260_nl, fsm_output[6]);
  assign nor_306_nl = ~((~ (fsm_output[3])) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[4])));
  assign or_1283_nl = (fsm_output[7]) | (fsm_output[9]) | (~ (fsm_output[8])) | (fsm_output[4]);
  assign nand_226_nl = ~((fsm_output[7]) & (fsm_output[9]) & (~ (fsm_output[8]))
      & (fsm_output[4]));
  assign mux_1280_nl = MUX_s_1_2_2(or_1283_nl, nand_226_nl, fsm_output[2]);
  assign nor_307_nl = ~((fsm_output[3]) | mux_1280_nl);
  assign mux_1281_nl = MUX_s_1_2_2(nor_306_nl, nor_307_nl, fsm_output[0]);
  assign nand_261_nl = ~((fsm_output[5]) & mux_1281_nl);
  assign or_1483_nl = (fsm_output[5]) | (fsm_output[0]) | (fsm_output[3]) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[4]));
  assign mux_1282_nl = MUX_s_1_2_2(nand_261_nl, or_1483_nl, fsm_output[6]);
  assign mux_1285_nl = MUX_s_1_2_2(mux_1284_nl, mux_1282_nl, fsm_output[1]);
  assign COMP_LOOP_mux1h_66_nl = MUX1HOT_s_1_3_2(modExp_exp_1_3_1_sva, modExp_exp_1_2_1_sva,
      (COMP_LOOP_k_9_3_sva_5_0[0]), {not_tmp_523 , (~ mux_1273_itm) , not_tmp_513});
  assign nand_86_nl = ~((fsm_output[3]) & (fsm_output[2]) & (fsm_output[9]) & (~
      (fsm_output[6])));
  assign mux_1317_nl = MUX_s_1_2_2((~ (fsm_output[6])), nand_86_nl, fsm_output[5]);
  assign or_1323_nl = (fsm_output[6:5]!=2'b01);
  assign mux_1318_nl = MUX_s_1_2_2(mux_1317_nl, or_1323_nl, fsm_output[7]);
  assign nand_247_nl = ~((~(or_1391_cse & (fsm_output[9]))) & (fsm_output[6]));
  assign or_1366_nl = (fsm_output[2]) | (fsm_output[1]) | (fsm_output[0]) | (fsm_output[9])
      | (~ (fsm_output[6]));
  assign mux_1314_nl = MUX_s_1_2_2(nand_247_nl, or_1366_nl, fsm_output[3]);
  assign or_1367_nl = (~((fsm_output[3]) | (fsm_output[2]) | (fsm_output[9]))) |
      (fsm_output[6]);
  assign mux_1315_nl = MUX_s_1_2_2(mux_1314_nl, or_1367_nl, fsm_output[5]);
  assign or_1316_nl = (~((fsm_output[2:0]!=3'b000))) | (~ (fsm_output[9])) | (fsm_output[6]);
  assign mux_1312_nl = MUX_s_1_2_2(or_1316_nl, (fsm_output[6]), fsm_output[3]);
  assign mux_1309_nl = MUX_s_1_2_2(or_tmp_1261, mux_tmp_1305, fsm_output[0]);
  assign mux_1310_nl = MUX_s_1_2_2((~ (fsm_output[6])), mux_1309_nl, and_483_cse);
  assign or_1314_nl = (~ (fsm_output[9])) | (fsm_output[6]);
  assign mux_1306_nl = MUX_s_1_2_2(mux_tmp_1305, or_1314_nl, fsm_output[0]);
  assign mux_1307_nl = MUX_s_1_2_2(mux_1306_nl, (fsm_output[6]), fsm_output[1]);
  assign mux_1308_nl = MUX_s_1_2_2(mux_tmp_1305, mux_1307_nl, fsm_output[2]);
  assign mux_1311_nl = MUX_s_1_2_2(mux_1310_nl, mux_1308_nl, fsm_output[3]);
  assign mux_1313_nl = MUX_s_1_2_2(mux_1312_nl, (~ mux_1311_nl), fsm_output[5]);
  assign mux_1316_nl = MUX_s_1_2_2(mux_1315_nl, mux_1313_nl, fsm_output[7]);
  assign mux_1319_nl = MUX_s_1_2_2(mux_1318_nl, mux_1316_nl, fsm_output[4]);
  assign mux_1299_nl = MUX_s_1_2_2((fsm_output[9]), or_tmp_1261, fsm_output[0]);
  assign mux_1300_nl = MUX_s_1_2_2(or_1099_cse, mux_1299_nl, fsm_output[1]);
  assign mux_1301_nl = MUX_s_1_2_2(mux_1300_nl, or_tmp_1261, or_1189_cse);
  assign mux_1302_nl = MUX_s_1_2_2((fsm_output[6]), mux_1301_nl, fsm_output[5]);
  assign mux_1296_nl = MUX_s_1_2_2(or_1099_cse, (fsm_output[9]), and_477_cse);
  assign mux_1297_nl = MUX_s_1_2_2(mux_1296_nl, or_tmp_1261, fsm_output[3]);
  assign or_1311_nl = (fsm_output[1]) | (fsm_output[0]) | (fsm_output[9]) | (~ (fsm_output[6]));
  assign mux_1295_nl = MUX_s_1_2_2(or_tmp_1261, or_1311_nl, and_316_cse);
  assign mux_1298_nl = MUX_s_1_2_2(mux_1297_nl, mux_1295_nl, fsm_output[5]);
  assign mux_1303_nl = MUX_s_1_2_2(mux_1302_nl, mux_1298_nl, fsm_output[7]);
  assign or_1309_nl = ((fsm_output[3]) & (fsm_output[2]) & (fsm_output[9])) | (fsm_output[6]);
  assign mux_1293_nl = MUX_s_1_2_2(or_1309_nl, or_tmp_1261, fsm_output[5]);
  assign or_1307_nl = (fsm_output[5]) | (fsm_output[9]) | (~ (fsm_output[6]));
  assign mux_1294_nl = MUX_s_1_2_2(mux_1293_nl, or_1307_nl, fsm_output[7]);
  assign mux_1304_nl = MUX_s_1_2_2(mux_1303_nl, mux_1294_nl, fsm_output[4]);
  assign mux_1320_nl = MUX_s_1_2_2(mux_1319_nl, mux_1304_nl, fsm_output[8]);
  assign COMP_LOOP_mux1h_68_nl = MUX1HOT_s_1_3_2((COMP_LOOP_k_9_3_sva_5_0[5]), modExp_exp_1_2_1_sva,
      modExp_exp_1_1_1_sva, {and_dcpl_226 , not_tmp_523 , (~ mux_1320_nl)});
  assign or_1434_nl = (~ (fsm_output[8])) | (fsm_output[3]) | (~ (fsm_output[5]))
      | (~ (fsm_output[0])) | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[1])
      | (~ (fsm_output[6]));
  assign or_1329_nl = (fsm_output[5]) | (~ (fsm_output[0])) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (fsm_output[1])) | (fsm_output[6]);
  assign or_1328_nl = (~ (fsm_output[0])) | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[1])
      | (~ (fsm_output[6]));
  assign or_1326_nl = (fsm_output[0]) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (fsm_output[1]) | (~ (fsm_output[6]));
  assign mux_1321_nl = MUX_s_1_2_2(or_1328_nl, or_1326_nl, fsm_output[5]);
  assign mux_1322_nl = MUX_s_1_2_2(or_1329_nl, mux_1321_nl, fsm_output[3]);
  assign or_1435_nl = (fsm_output[8]) | mux_1322_nl;
  assign mux_1323_nl = MUX_s_1_2_2(or_1434_nl, or_1435_nl, fsm_output[4]);
  assign nor_293_nl = ~((fsm_output[5]) | (fsm_output[2]) | (fsm_output[6]));
  assign and_283_nl = (fsm_output[5]) & (fsm_output[2]) & (fsm_output[6]);
  assign mux_1324_nl = MUX_s_1_2_2(nor_293_nl, and_283_nl, fsm_output[0]);
  assign nor_292_nl = ~((fsm_output[4:3]!=2'b10) | (~((fsm_output[7]) & mux_1324_nl)));
  assign nor_294_nl = ~((fsm_output[4]) | (~ (fsm_output[3])) | (fsm_output[7]) |
      (~ (fsm_output[0])) | (~ (fsm_output[5])) | (fsm_output[2]) | (fsm_output[6]));
  assign mux_1325_nl = MUX_s_1_2_2(nor_292_nl, nor_294_nl, fsm_output[1]);
  assign and_282_nl = (fsm_output[9]) & mux_1325_nl;
  assign nor_295_nl = ~((fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[4]) |
      (fsm_output[3]) | (~ (fsm_output[7])) | (fsm_output[0]) | (fsm_output[5]) |
      (~((fsm_output[2]) & (fsm_output[6]))));
  assign mux_1326_nl = MUX_s_1_2_2(and_282_nl, nor_295_nl, fsm_output[8]);
  assign nor_659_nl = ~((fsm_output[8:1]!=8'b00000000));
  assign and_176_nl = (fsm_output[6]) & ((fsm_output[5]) | and_428_cse);
  assign mux_812_nl = MUX_s_1_2_2(and_176_nl, and_491_cse, fsm_output[2]);
  assign and_704_nl = (fsm_output[8]) & ((fsm_output[7]) | mux_812_nl);
  assign or_1499_nl = (~ (fsm_output[1])) | (fsm_output[6]) | (fsm_output[3]);
  assign mux_1418_nl = MUX_s_1_2_2(mux_tmp_1399, or_1499_nl, fsm_output[0]);
  assign or_1550_nl = (fsm_output[4]) | mux_1418_nl;
  assign mux_1417_nl = MUX_s_1_2_2(or_tmp_1367, (~ (fsm_output[3])), fsm_output[4]);
  assign mux_1419_nl = MUX_s_1_2_2(or_1550_nl, mux_1417_nl, fsm_output[2]);
  assign mux_1415_nl = MUX_s_1_2_2((~ or_136_cse), (fsm_output[3]), fsm_output[4]);
  assign and_707_nl = (fsm_output[4]) & or_tmp_1374;
  assign mux_1416_nl = MUX_s_1_2_2(mux_1415_nl, and_707_nl, fsm_output[2]);
  assign mux_1420_nl = MUX_s_1_2_2(mux_1419_nl, mux_1416_nl, fsm_output[7]);
  assign and_706_nl = (fsm_output[4]) & ((~ (fsm_output[0])) | (fsm_output[1]) |
      (fsm_output[6]) | (fsm_output[3]));
  assign or_1497_nl = (fsm_output[4]) | nor_tmp_296;
  assign mux_1413_nl = MUX_s_1_2_2(and_706_nl, or_1497_nl, fsm_output[2]);
  assign mux_1410_nl = MUX_s_1_2_2(nor_tmp_292, (fsm_output[6]), fsm_output[1]);
  assign mux_1411_nl = MUX_s_1_2_2((~ mux_1410_nl), or_tmp_1370, fsm_output[4]);
  assign mux_1412_nl = MUX_s_1_2_2((~ mux_tmp_1374), mux_1411_nl, fsm_output[2]);
  assign mux_1414_nl = MUX_s_1_2_2(mux_1413_nl, mux_1412_nl, fsm_output[7]);
  assign mux_1421_nl = MUX_s_1_2_2(mux_1420_nl, mux_1414_nl, fsm_output[5]);
  assign mux_1406_nl = MUX_s_1_2_2(nor_tmp_296, (fsm_output[6]), fsm_output[4]);
  assign mux_1407_nl = MUX_s_1_2_2(mux_1406_nl, mux_tmp_1374, fsm_output[2]);
  assign mux_1403_nl = MUX_s_1_2_2(or_tmp_1370, mux_tmp_1377, and_389_cse);
  assign mux_1404_nl = MUX_s_1_2_2(mux_1403_nl, (fsm_output[6]), fsm_output[4]);
  assign mux_1401_nl = MUX_s_1_2_2(mux_tmp_1377, or_tmp_1365, fsm_output[1]);
  assign mux_1402_nl = MUX_s_1_2_2(mux_1401_nl, mux_tmp_1399, fsm_output[4]);
  assign mux_1405_nl = MUX_s_1_2_2(mux_1404_nl, mux_1402_nl, fsm_output[2]);
  assign mux_1408_nl = MUX_s_1_2_2(mux_1407_nl, (~ mux_1405_nl), fsm_output[7]);
  assign mux_1396_nl = MUX_s_1_2_2((fsm_output[6]), or_tmp_1367, or_838_cse);
  assign mux_1397_nl = MUX_s_1_2_2(mux_tmp_1378, mux_1396_nl, fsm_output[4]);
  assign mux_1395_nl = MUX_s_1_2_2(mux_tmp, or_tmp_1367, fsm_output[4]);
  assign mux_1398_nl = MUX_s_1_2_2(mux_1397_nl, mux_1395_nl, fsm_output[2]);
  assign mux_1399_nl = MUX_s_1_2_2((~ mux_1398_nl), (fsm_output[4]), fsm_output[7]);
  assign mux_1409_nl = MUX_s_1_2_2(mux_1408_nl, mux_1399_nl, fsm_output[5]);
  assign mux_1422_nl = MUX_s_1_2_2((~ mux_1421_nl), mux_1409_nl, fsm_output[8]);
  assign mux_1390_nl = MUX_s_1_2_2((~ or_tmp_1374), (fsm_output[3]), fsm_output[4]);
  assign mux_1391_nl = MUX_s_1_2_2(mux_1390_nl, and_705_cse, fsm_output[2]);
  assign nand_275_nl = ~(or_838_cse & (fsm_output[6]) & (fsm_output[3]));
  assign mux_1388_nl = MUX_s_1_2_2(nand_275_nl, nor_tmp_296, fsm_output[4]);
  assign mux_1389_nl = MUX_s_1_2_2((~ (fsm_output[4])), mux_1388_nl, fsm_output[2]);
  assign mux_1392_nl = MUX_s_1_2_2(mux_1391_nl, mux_1389_nl, fsm_output[7]);
  assign nand_276_nl = ~((and_389_cse | (fsm_output[6])) & (fsm_output[3]));
  assign and_717_nl = (fsm_output[1]) & (fsm_output[6]) & (fsm_output[3]);
  assign mux_1385_nl = MUX_s_1_2_2(nand_276_nl, and_717_nl, fsm_output[4]);
  assign mux_1384_nl = MUX_s_1_2_2((~ (fsm_output[3])), nor_tmp_292, fsm_output[4]);
  assign mux_1386_nl = MUX_s_1_2_2(mux_1385_nl, mux_1384_nl, fsm_output[2]);
  assign mux_1381_nl = MUX_s_1_2_2(or_tmp_1370, mux_tmp_1377, fsm_output[1]);
  assign mux_1382_nl = MUX_s_1_2_2((~ (fsm_output[6])), mux_1381_nl, fsm_output[4]);
  assign mux_1380_nl = MUX_s_1_2_2((~ (fsm_output[6])), mux_tmp_1378, fsm_output[4]);
  assign mux_1383_nl = MUX_s_1_2_2(mux_1382_nl, mux_1380_nl, fsm_output[2]);
  assign mux_1387_nl = MUX_s_1_2_2(mux_1386_nl, (~ mux_1383_nl), fsm_output[7]);
  assign mux_1393_nl = MUX_s_1_2_2(mux_1392_nl, mux_1387_nl, fsm_output[5]);
  assign and_718_nl = (fsm_output[4]) & (fsm_output[0]) & (fsm_output[1]);
  assign mux_1374_nl = MUX_s_1_2_2((fsm_output[6]), or_tmp_1367, and_718_nl);
  assign mux_1376_nl = MUX_s_1_2_2(mux_tmp_1374, mux_1374_nl, fsm_output[2]);
  assign or_1489_nl = (fsm_output[7]) | mux_1376_nl;
  assign nand_266_nl = ~((fsm_output[4]) & (~ mux_tmp));
  assign or_1485_nl = (~ (fsm_output[4])) | (fsm_output[6]);
  assign mux_1373_nl = MUX_s_1_2_2(nand_266_nl, or_1485_nl, fsm_output[2]);
  assign or_1487_nl = (fsm_output[7]) | mux_1373_nl;
  assign mux_1377_nl = MUX_s_1_2_2(or_1489_nl, or_1487_nl, fsm_output[5]);
  assign mux_1394_nl = MUX_s_1_2_2(mux_1393_nl, mux_1377_nl, fsm_output[8]);
  assign mux_1423_nl = MUX_s_1_2_2(mux_1422_nl, mux_1394_nl, fsm_output[9]);
  assign or_1540_nl = (fsm_output[8:5]!=4'b0001);
  assign or_1539_nl = (fsm_output[8:5]!=4'b0100);
  assign or_1537_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[8:7]!=2'b00);
  assign mux_1448_nl = MUX_s_1_2_2(or_tmp_1394, or_1537_nl, fsm_output[6]);
  assign mux_1449_nl = MUX_s_1_2_2(mux_1448_nl, or_tmp_1401, fsm_output[5]);
  assign mux_1450_nl = MUX_s_1_2_2(or_1539_nl, mux_1449_nl, fsm_output[1]);
  assign mux_1451_nl = MUX_s_1_2_2(or_1540_nl, mux_1450_nl, fsm_output[9]);
  assign and_710_nl = (fsm_output[4]) & (~ mux_1451_nl);
  assign or_1535_nl = (fsm_output[5]) | (~(COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm &
      (fsm_output[8:7]==2'b11)));
  assign or_1534_nl = (fsm_output[8:5]!=4'b0000);
  assign mux_1446_nl = MUX_s_1_2_2(or_1535_nl, or_1534_nl, fsm_output[1]);
  assign or_1533_nl = (fsm_output[1]) | (~ (fsm_output[5])) | (~ (fsm_output[6]))
      | (fsm_output[8]) | (fsm_output[7]);
  assign mux_1447_nl = MUX_s_1_2_2(mux_1446_nl, or_1533_nl, fsm_output[9]);
  assign nor_676_nl = ~((fsm_output[4]) | mux_1447_nl);
  assign mux_1452_nl = MUX_s_1_2_2(and_710_nl, nor_676_nl, fsm_output[3]);
  assign nor_677_nl = ~((fsm_output[8:6]!=3'b000));
  assign nor_678_nl = ~((fsm_output[8:6]!=3'b101));
  assign mux_1441_nl = MUX_s_1_2_2(nor_677_nl, nor_678_nl, fsm_output[5]);
  assign and_711_nl = (fsm_output[5]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & (fsm_output[8:7]==2'b10);
  assign mux_1442_nl = MUX_s_1_2_2(mux_1441_nl, and_711_nl, fsm_output[1]);
  assign nor_679_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[6]) |
      (fsm_output[8]) | (fsm_output[7]));
  assign mux_1443_nl = MUX_s_1_2_2(mux_1442_nl, nor_679_nl, fsm_output[9]);
  assign nor_680_nl = ~((fsm_output[9]) | (~ (fsm_output[1])) | (~ (fsm_output[5]))
      | (fsm_output[6]) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[8:7]!=2'b00));
  assign mux_1444_nl = MUX_s_1_2_2(mux_1443_nl, nor_680_nl, fsm_output[4]);
  assign nor_681_nl = ~((fsm_output[1]) | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[8])
      | (fsm_output[7]));
  assign nor_682_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[5])) | (fsm_output[6])
      | (fsm_output[8]) | (fsm_output[7]));
  assign mux_1439_nl = MUX_s_1_2_2(nor_681_nl, nor_682_nl, fsm_output[9]);
  assign or_1524_nl = (fsm_output[6]) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[8:7]!=2'b01);
  assign mux_1438_nl = MUX_s_1_2_2(or_1524_nl, or_tmp_1401, fsm_output[5]);
  assign nor_683_nl = ~((fsm_output[9]) | (fsm_output[1]) | mux_1438_nl);
  assign mux_1440_nl = MUX_s_1_2_2(mux_1439_nl, nor_683_nl, fsm_output[4]);
  assign mux_1445_nl = MUX_s_1_2_2(mux_1444_nl, mux_1440_nl, fsm_output[3]);
  assign mux_1453_nl = MUX_s_1_2_2(mux_1452_nl, mux_1445_nl, fsm_output[0]);
  assign mux_1433_nl = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[8]);
  assign mux_1434_nl = MUX_s_1_2_2(nor_tmp_301, mux_1433_nl, COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign nor_684_nl = ~((fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[5]) |
      (~((fsm_output[6]) & mux_1434_nl)));
  assign nor_685_nl = ~((fsm_output[9]) | (fsm_output[1]) | (fsm_output[5]) | (~
      (fsm_output[6])) | (fsm_output[8]) | (~ (fsm_output[7])));
  assign mux_1435_nl = MUX_s_1_2_2(nor_684_nl, nor_685_nl, fsm_output[4]);
  assign or_1516_nl = (fsm_output[6]) | (~ nor_tmp_301);
  assign mux_1430_nl = MUX_s_1_2_2(or_1516_nl, or_tmp_1394, fsm_output[5]);
  assign mux_1431_nl = MUX_s_1_2_2(or_tmp_1389, mux_1430_nl, fsm_output[1]);
  assign or_1513_nl = (fsm_output[1]) | (fsm_output[5]) | (fsm_output[6]) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[8:7]!=2'b10);
  assign mux_1432_nl = MUX_s_1_2_2(mux_1431_nl, or_1513_nl, fsm_output[9]);
  assign and_712_nl = (fsm_output[4]) & (~ mux_1432_nl);
  assign mux_1436_nl = MUX_s_1_2_2(mux_1435_nl, and_712_nl, fsm_output[3]);
  assign or_1512_nl = (~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[8])
      | (~ (fsm_output[7]));
  assign nand_278_nl = ~((fsm_output[5]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm &
      (fsm_output[8:7]==2'b01));
  assign mux_1427_nl = MUX_s_1_2_2(or_tmp_1389, nand_278_nl, fsm_output[1]);
  assign mux_1428_nl = MUX_s_1_2_2(or_1512_nl, mux_1427_nl, fsm_output[9]);
  assign and_713_nl = (fsm_output[4]) & (~ mux_1428_nl);
  assign nand_274_nl = ~((fsm_output[6:5]==2'b11) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      & (fsm_output[8:7]==2'b11));
  assign or_1505_nl = (fsm_output[8:5]!=4'b0011);
  assign mux_1425_nl = MUX_s_1_2_2(nand_274_nl, or_1505_nl, fsm_output[1]);
  assign or_1503_nl = (fsm_output[8:6]!=3'b011);
  assign or_1501_nl = (fsm_output[6]) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[8:7]!=2'b00);
  assign mux_1424_nl = MUX_s_1_2_2(or_1503_nl, or_1501_nl, fsm_output[5]);
  assign or_1504_nl = (fsm_output[1]) | mux_1424_nl;
  assign mux_1426_nl = MUX_s_1_2_2(mux_1425_nl, or_1504_nl, fsm_output[9]);
  assign nor_686_nl = ~((fsm_output[4]) | mux_1426_nl);
  assign mux_1429_nl = MUX_s_1_2_2(and_713_nl, nor_686_nl, fsm_output[3]);
  assign mux_1437_nl = MUX_s_1_2_2(mux_1436_nl, mux_1429_nl, fsm_output[0]);
  assign or_940_nl = (~ (fsm_output[0])) | (fsm_output[1]) | (~ (fsm_output[3]))
      | (fsm_output[4]);
  assign mux_864_nl = MUX_s_1_2_2(or_940_nl, or_242_cse, fsm_output[5]);
  assign nor_630_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_864_nl);
  assign nor_631_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[6])) | (fsm_output[5])
      | (fsm_output[0]) | (~ and_dcpl_59));
  assign mux_865_nl = MUX_s_1_2_2(nor_630_nl, nor_631_nl, fsm_output[9]);
  assign nand_263_nl = ~(mux_865_nl & and_dcpl_140);
  assign or_1547_nl = (fsm_output[2]) | (~ (fsm_output[0])) | (fsm_output[6]) | (fsm_output[1])
      | (fsm_output[5]) | (~ (fsm_output[3]));
  assign or_1545_nl = (fsm_output[2]) | (fsm_output[0]) | (fsm_output[6]) | (fsm_output[1])
      | (~ (fsm_output[5])) | (fsm_output[3]);
  assign mux_1456_nl = MUX_s_1_2_2(or_1547_nl, or_1545_nl, fsm_output[4]);
  assign or_1549_nl = (fsm_output[8]) | mux_1456_nl;
  assign nor_674_nl = ~((fsm_output[0]) | (~ (fsm_output[6])) | (~ (fsm_output[1]))
      | (fsm_output[5]) | (~ (fsm_output[3])));
  assign nor_675_nl = ~((~ (fsm_output[0])) | (fsm_output[6]) | (fsm_output[1]) |
      (fsm_output[5]) | (~ (fsm_output[3])));
  assign mux_1455_nl = MUX_s_1_2_2(nor_674_nl, nor_675_nl, fsm_output[2]);
  assign nand_271_nl = ~((fsm_output[8]) & (fsm_output[4]) & mux_1455_nl);
  assign mux_1457_nl = MUX_s_1_2_2(or_1549_nl, nand_271_nl, fsm_output[9]);
  assign nor_389_nl = ~((fsm_output[6]) | (fsm_output[8]) | (fsm_output[9]));
  assign nor_390_nl = ~((fsm_output[1]) | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[8])
      | (fsm_output[9]));
  assign mux_882_nl = MUX_s_1_2_2(nor_389_nl, nor_390_nl, fsm_output[3]);
  assign and_360_nl = (fsm_output[2]) & (fsm_output[6]) & (fsm_output[8]) & (fsm_output[9]);
  assign mux_879_nl = MUX_s_1_2_2(nor_393_cse, and_369_cse, fsm_output[6]);
  assign and_184_nl = (fsm_output[2]) & mux_879_nl;
  assign mux_880_nl = MUX_s_1_2_2(and_184_nl, and_361_cse, fsm_output[1]);
  assign mux_881_nl = MUX_s_1_2_2(and_360_nl, mux_880_nl, fsm_output[0]);
  assign and_185_nl = (fsm_output[3]) & mux_881_nl;
  assign mux_883_nl = MUX_s_1_2_2(mux_882_nl, and_185_nl, fsm_output[4]);
  assign mux_884_nl = MUX_s_1_2_2(mux_883_nl, and_361_cse, fsm_output[5]);
  assign mux_885_nl = MUX_s_1_2_2(mux_884_nl, and_369_cse, fsm_output[7]);
  assign COMP_LOOP_or_15_nl = (and_dcpl_172 & and_dcpl_167) | (COMP_LOOP_COMP_LOOP_nor_4_itm
      & and_224_m1c) | (COMP_LOOP_COMP_LOOP_and_34_itm & and_226_m1c) | (COMP_LOOP_COMP_LOOP_and_33_itm
      & and_229_m1c) | (COMP_LOOP_COMP_LOOP_and_32_itm & and_230_m1c) | (COMP_LOOP_COMP_LOOP_and_89_itm
      & and_233_m1c) | (COMP_LOOP_COMP_LOOP_and_30_itm & and_235_m1c) | (COMP_LOOP_COMP_LOOP_and_145_itm
      & and_237_m1c);
  assign COMP_LOOP_or_16_nl = (and_dcpl_172 & and_dcpl_176) | (COMP_LOOP_COMP_LOOP_and_86_itm
      & and_224_m1c) | (COMP_LOOP_COMP_LOOP_nor_4_itm & and_226_m1c) | (COMP_LOOP_COMP_LOOP_and_34_itm
      & and_229_m1c) | (COMP_LOOP_COMP_LOOP_and_33_itm & and_230_m1c) | (COMP_LOOP_COMP_LOOP_and_32_itm
      & and_233_m1c) | (COMP_LOOP_COMP_LOOP_and_89_itm & and_235_m1c) | (COMP_LOOP_COMP_LOOP_and_30_itm
      & and_237_m1c);
  assign COMP_LOOP_or_17_nl = (and_dcpl_172 & and_dcpl_180) | (COMP_LOOP_COMP_LOOP_and_145_itm
      & and_224_m1c) | (COMP_LOOP_COMP_LOOP_and_86_itm & and_226_m1c) | (COMP_LOOP_COMP_LOOP_nor_4_itm
      & and_229_m1c) | (COMP_LOOP_COMP_LOOP_and_34_itm & and_230_m1c) | (COMP_LOOP_COMP_LOOP_and_33_itm
      & and_233_m1c) | (COMP_LOOP_COMP_LOOP_and_32_itm & and_235_m1c) | (COMP_LOOP_COMP_LOOP_and_89_itm
      & and_237_m1c);
  assign COMP_LOOP_or_18_nl = (and_dcpl_172 & and_dcpl_184) | (COMP_LOOP_COMP_LOOP_and_30_itm
      & and_224_m1c) | (COMP_LOOP_COMP_LOOP_and_145_itm & and_226_m1c) | (COMP_LOOP_COMP_LOOP_and_86_itm
      & and_229_m1c) | (COMP_LOOP_COMP_LOOP_nor_4_itm & and_230_m1c) | (COMP_LOOP_COMP_LOOP_and_34_itm
      & and_233_m1c) | (COMP_LOOP_COMP_LOOP_and_33_itm & and_235_m1c) | (COMP_LOOP_COMP_LOOP_and_32_itm
      & and_237_m1c);
  assign COMP_LOOP_or_19_nl = (and_dcpl_187 & and_dcpl_167) | (COMP_LOOP_COMP_LOOP_and_89_itm
      & and_224_m1c) | (COMP_LOOP_COMP_LOOP_and_30_itm & and_226_m1c) | (COMP_LOOP_COMP_LOOP_and_145_itm
      & and_229_m1c) | (COMP_LOOP_COMP_LOOP_and_86_itm & and_230_m1c) | (COMP_LOOP_COMP_LOOP_nor_4_itm
      & and_233_m1c) | (COMP_LOOP_COMP_LOOP_and_34_itm & and_235_m1c) | (COMP_LOOP_COMP_LOOP_and_33_itm
      & and_237_m1c);
  assign COMP_LOOP_or_20_nl = (and_dcpl_187 & and_dcpl_176) | (COMP_LOOP_COMP_LOOP_and_32_itm
      & and_224_m1c) | (COMP_LOOP_COMP_LOOP_and_89_itm & and_226_m1c) | (COMP_LOOP_COMP_LOOP_and_30_itm
      & and_229_m1c) | (COMP_LOOP_COMP_LOOP_and_145_itm & and_230_m1c) | (COMP_LOOP_COMP_LOOP_and_86_itm
      & and_233_m1c) | (COMP_LOOP_COMP_LOOP_nor_4_itm & and_235_m1c) | (COMP_LOOP_COMP_LOOP_and_34_itm
      & and_237_m1c);
  assign COMP_LOOP_or_21_nl = (and_dcpl_187 & and_dcpl_180) | (COMP_LOOP_COMP_LOOP_and_33_itm
      & and_224_m1c) | (COMP_LOOP_COMP_LOOP_and_32_itm & and_226_m1c) | (COMP_LOOP_COMP_LOOP_and_89_itm
      & and_229_m1c) | (COMP_LOOP_COMP_LOOP_and_30_itm & and_230_m1c) | (COMP_LOOP_COMP_LOOP_and_145_itm
      & and_233_m1c) | (COMP_LOOP_COMP_LOOP_and_86_itm & and_235_m1c) | (COMP_LOOP_COMP_LOOP_nor_4_itm
      & and_237_m1c);
  assign COMP_LOOP_or_22_nl = (and_dcpl_187 & and_dcpl_184) | (COMP_LOOP_COMP_LOOP_and_34_itm
      & and_224_m1c) | (COMP_LOOP_COMP_LOOP_and_33_itm & and_226_m1c) | (COMP_LOOP_COMP_LOOP_and_32_itm
      & and_229_m1c) | (COMP_LOOP_COMP_LOOP_and_89_itm & and_230_m1c) | (COMP_LOOP_COMP_LOOP_and_30_itm
      & and_233_m1c) | (COMP_LOOP_COMP_LOOP_and_145_itm & and_235_m1c) | (COMP_LOOP_COMP_LOOP_and_86_itm
      & and_237_m1c);
  assign or_964_nl = and_389_cse | (fsm_output[4:3]!=2'b10);
  assign mux_909_nl = MUX_s_1_2_2(or_tmp_113, or_964_nl, fsm_output[5]);
  assign mux_910_nl = MUX_s_1_2_2(mux_909_nl, (~ and_314_cse), fsm_output[6]);
  assign nand_120_nl = ~((fsm_output[5]) & or_tmp_788);
  assign mux_908_nl = MUX_s_1_2_2(or_1202_cse, nand_120_nl, fsm_output[6]);
  assign mux_911_nl = MUX_s_1_2_2(mux_910_nl, mux_908_nl, fsm_output[2]);
  assign mux_906_nl = MUX_s_1_2_2(or_tmp, (~ or_tmp), fsm_output[6]);
  assign mux_904_nl = MUX_s_1_2_2((~ (fsm_output[4])), nor_tmp_27, fsm_output[5]);
  assign mux_905_nl = MUX_s_1_2_2(or_tmp, mux_904_nl, fsm_output[6]);
  assign mux_907_nl = MUX_s_1_2_2(mux_906_nl, mux_905_nl, fsm_output[2]);
  assign mux_912_nl = MUX_s_1_2_2(mux_911_nl, mux_907_nl, fsm_output[7]);
  assign nand_121_nl = ~((fsm_output[5]) & nor_tmp_27);
  assign and_192_nl = (fsm_output[5]) & ((fsm_output[1]) | (fsm_output[3]) | (fsm_output[4]));
  assign mux_901_nl = MUX_s_1_2_2(nand_121_nl, and_192_nl, fsm_output[6]);
  assign nand_122_nl = ~((fsm_output[5:3]==3'b111));
  assign mux_900_nl = MUX_s_1_2_2(nand_122_nl, (fsm_output[5]), fsm_output[6]);
  assign mux_902_nl = MUX_s_1_2_2(mux_901_nl, mux_900_nl, fsm_output[2]);
  assign mux_898_nl = MUX_s_1_2_2((~ (fsm_output[5])), or_1202_cse, fsm_output[6]);
  assign nor_388_nl = ~((fsm_output[5]) | and_dcpl_59);
  assign or_959_nl = (fsm_output[5]) | or_tmp_103;
  assign mux_897_nl = MUX_s_1_2_2(nor_388_nl, or_959_nl, fsm_output[6]);
  assign mux_899_nl = MUX_s_1_2_2(mux_898_nl, mux_897_nl, fsm_output[2]);
  assign mux_903_nl = MUX_s_1_2_2(mux_902_nl, mux_899_nl, fsm_output[7]);
  assign mux_913_nl = MUX_s_1_2_2(mux_912_nl, mux_903_nl, fsm_output[8]);
  assign mux_892_nl = MUX_s_1_2_2(or_tmp_103, (~ (fsm_output[4])), fsm_output[5]);
  assign mux_893_nl = MUX_s_1_2_2(mux_892_nl, and_tmp_28, fsm_output[6]);
  assign mux_891_nl = MUX_s_1_2_2((~ and_tmp_28), and_tmp_28, fsm_output[6]);
  assign mux_894_nl = MUX_s_1_2_2(mux_893_nl, mux_891_nl, fsm_output[2]);
  assign or_958_nl = (fsm_output[5]) | and_705_cse;
  assign mux_889_nl = MUX_s_1_2_2(or_958_nl, mux_tmp_705, fsm_output[6]);
  assign mux_887_nl = MUX_s_1_2_2((~ or_115_cse), nor_tmp_23, fsm_output[5]);
  assign mux_888_nl = MUX_s_1_2_2(or_171_cse, mux_887_nl, fsm_output[6]);
  assign mux_890_nl = MUX_s_1_2_2(mux_889_nl, mux_888_nl, fsm_output[2]);
  assign mux_895_nl = MUX_s_1_2_2(mux_894_nl, (~ mux_890_nl), fsm_output[7]);
  assign mux_896_nl = MUX_s_1_2_2(mux_895_nl, or_tmp_918, fsm_output[8]);
  assign and_238_nl = and_dcpl_102 & and_dcpl_48;
  assign COMP_LOOP_or_26_nl = ((~ (modulo_result_rem_cmp_z[63])) & and_243_m1c) |
      (not_tmp_399 & (~ (modulo_result_rem_cmp_z[63])));
  assign COMP_LOOP_or_27_nl = ((modulo_result_rem_cmp_z[63]) & and_243_m1c) | (not_tmp_399
      & (modulo_result_rem_cmp_z[63]));
  assign COMP_LOOP_or_7_nl = (COMP_LOOP_COMP_LOOP_nor_1_itm & and_244_m1c) | (COMP_LOOP_COMP_LOOP_nor_1_itm
      & mux_984_m1c);
  assign COMP_LOOP_or_8_nl = (COMP_LOOP_COMP_LOOP_and_211 & and_244_m1c) | (COMP_LOOP_COMP_LOOP_and_211
      & mux_984_m1c);
  assign COMP_LOOP_or_9_nl = (COMP_LOOP_COMP_LOOP_and_213 & and_244_m1c) | (COMP_LOOP_COMP_LOOP_and_213
      & mux_984_m1c);
  assign COMP_LOOP_or_10_nl = (COMP_LOOP_COMP_LOOP_and_125_itm & and_244_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & mux_984_m1c);
  assign COMP_LOOP_or_11_nl = (COMP_LOOP_COMP_LOOP_and_215 & and_244_m1c) | (COMP_LOOP_COMP_LOOP_and_215
      & mux_984_m1c);
  assign COMP_LOOP_or_12_nl = (COMP_LOOP_COMP_LOOP_and_11_itm & and_244_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & mux_984_m1c);
  assign COMP_LOOP_or_13_nl = (COMP_LOOP_COMP_LOOP_and_12_itm & and_244_m1c) | (COMP_LOOP_COMP_LOOP_and_124_itm
      & mux_984_m1c);
  assign COMP_LOOP_or_14_nl = (COMP_LOOP_COMP_LOOP_and_124_itm & and_244_m1c) | (COMP_LOOP_COMP_LOOP_and_125_itm
      & mux_984_m1c);
  assign nor_591_nl = ~((~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[9]) |
      (fsm_output[4]) | (fsm_output[1]) | (~ (fsm_output[6])));
  assign nor_592_nl = ~((fsm_output[0]) | (~ (fsm_output[3])) | (~ (fsm_output[9]))
      | (~ (fsm_output[4])) | (~ (fsm_output[1])) | (fsm_output[6]));
  assign mux_46_nl = MUX_s_1_2_2(nor_591_nl, nor_592_nl, fsm_output[5]);
  assign nor_593_nl = ~((~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[9])
      | (fsm_output[4]) | (~ (fsm_output[1])) | (fsm_output[6]));
  assign nor_594_nl = ~((fsm_output[0]) | (fsm_output[3]) | (fsm_output[9]) | (~
      (fsm_output[4])) | (fsm_output[1]) | (~ (fsm_output[6])));
  assign mux_45_nl = MUX_s_1_2_2(nor_593_nl, nor_594_nl, fsm_output[5]);
  assign mux_47_nl = MUX_s_1_2_2(mux_46_nl, mux_45_nl, fsm_output[8]);
  assign and_470_nl = (fsm_output[7]) & mux_47_nl;
  assign or_61_nl = (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[4])) |
      (fsm_output[1]) | (~ (fsm_output[6]));
  assign or_59_nl = (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[4])) |
      (fsm_output[1]) | (~ (fsm_output[6]));
  assign mux_43_nl = MUX_s_1_2_2(or_61_nl, or_59_nl, fsm_output[0]);
  assign or_62_nl = (fsm_output[5]) | mux_43_nl;
  assign nand_224_nl = ~((fsm_output[0]) & (fsm_output[3]) & (fsm_output[9]) & (fsm_output[4])
      & (fsm_output[1]) & (~ (fsm_output[6])));
  assign or_56_nl = (fsm_output[0]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[4])
      | (~ (fsm_output[1])) | (fsm_output[6]);
  assign mux_42_nl = MUX_s_1_2_2(nand_224_nl, or_56_nl, fsm_output[5]);
  assign mux_44_nl = MUX_s_1_2_2(or_62_nl, mux_42_nl, fsm_output[8]);
  assign nor_595_nl = ~((fsm_output[7]) | mux_44_nl);
  assign mux_48_nl = MUX_s_1_2_2(and_470_nl, nor_595_nl, fsm_output[2]);
  assign or_248_nl = (fsm_output[0]) | (~ (fsm_output[1])) | (~ (fsm_output[3]))
      | (fsm_output[4]);
  assign mux_347_nl = MUX_s_1_2_2(or_248_nl, or_tmp_92, fsm_output[5]);
  assign mux_348_nl = MUX_s_1_2_2(mux_347_nl, or_247_cse, fsm_output[6]);
  assign mux_346_nl = MUX_s_1_2_2(nor_tmp_27, (~ or_tmp_113), fsm_output[5]);
  assign nand_9_nl = ~((fsm_output[6]) & mux_346_nl);
  assign mux_349_nl = MUX_s_1_2_2(mux_348_nl, nand_9_nl, fsm_output[2]);
  assign nor_371_nl = ~((fsm_output[1:0]!=2'b00) | (~ nor_tmp));
  assign mux_963_nl = MUX_s_1_2_2(nor_371_nl, (fsm_output[4]), fsm_output[5]);
  assign mux_341_nl = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), or_245_cse);
  assign mux_343_nl = MUX_s_1_2_2(mux_342_cse, mux_341_nl, fsm_output[0]);
  assign or_246_nl = (fsm_output[5]) | mux_343_nl;
  assign mux_964_nl = MUX_s_1_2_2((~ mux_963_nl), or_246_nl, fsm_output[6]);
  assign nand_56_nl = ~((fsm_output[5]) & (~ mux_696_itm));
  assign or_1009_nl = (fsm_output[1:0]!=2'b01) | (~ nor_tmp);
  assign mux_959_nl = MUX_s_1_2_2((fsm_output[4]), or_1009_nl, fsm_output[5]);
  assign mux_960_nl = MUX_s_1_2_2(nand_56_nl, mux_959_nl, fsm_output[6]);
  assign mux_965_nl = MUX_s_1_2_2(mux_964_nl, mux_960_nl, fsm_output[2]);
  assign mux_970_nl = MUX_s_1_2_2(mux_349_nl, mux_965_nl, fsm_output[7]);
  assign mux_955_nl = MUX_s_1_2_2(and_705_cse, (~ nor_tmp), fsm_output[5]);
  assign nor_190_nl = ~((fsm_output[1:0]!=2'b10));
  assign mux_954_nl = MUX_s_1_2_2(nor_tmp, mux_tmp_156, nor_190_nl);
  assign and_246_nl = (fsm_output[5]) & mux_954_nl;
  assign mux_956_nl = MUX_s_1_2_2(mux_955_nl, and_246_nl, fsm_output[6]);
  assign mux_332_nl = MUX_s_1_2_2((fsm_output[4]), (~ mux_331_cse), fsm_output[5]);
  assign mux_333_nl = MUX_s_1_2_2(mux_332_nl, and_25_cse, fsm_output[6]);
  assign mux_957_nl = MUX_s_1_2_2(mux_956_nl, mux_333_nl, fsm_output[2]);
  assign nor_372_nl = ~((fsm_output[5]) | (~((~((fsm_output[1:0]!=2'b00))) | (fsm_output[4:3]!=2'b01))));
  assign mux_328_nl = MUX_s_1_2_2(and_428_cse, or_242_cse, fsm_output[5]);
  assign mux_950_nl = MUX_s_1_2_2(nor_372_nl, mux_328_nl, fsm_output[6]);
  assign nor_560_nl = ~((fsm_output[5]) | nor_tmp_27);
  assign mux_334_nl = MUX_s_1_2_2(nor_tmp, mux_tmp_156, and_389_cse);
  assign or_1003_nl = (~ (fsm_output[1])) | (~ (fsm_output[3])) | (fsm_output[4]);
  assign mux_947_nl = MUX_s_1_2_2(mux_334_nl, or_1003_nl, fsm_output[5]);
  assign mux_948_nl = MUX_s_1_2_2(nor_560_nl, mux_947_nl, fsm_output[6]);
  assign mux_951_nl = MUX_s_1_2_2(mux_950_nl, mux_948_nl, fsm_output[2]);
  assign mux_958_nl = MUX_s_1_2_2(mux_957_nl, mux_951_nl, fsm_output[7]);
  assign mux_971_nl = MUX_s_1_2_2(mux_970_nl, (~ mux_958_nl), fsm_output[8]);
  assign or_1002_nl = (fsm_output[5]) | (fsm_output[1]) | (fsm_output[3]) | (fsm_output[4]);
  assign mux_941_nl = MUX_s_1_2_2((~ or_tmp_92), or_216_cse, fsm_output[5]);
  assign mux_942_nl = MUX_s_1_2_2(or_1002_nl, mux_941_nl, fsm_output[6]);
  assign or_999_nl = (~ (fsm_output[5])) | (fsm_output[0]) | (fsm_output[1]) | (~
      (fsm_output[3])) | (fsm_output[4]);
  assign mux_939_nl = MUX_s_1_2_2(and_dcpl_64, or_tmp_103, fsm_output[5]);
  assign mux_940_nl = MUX_s_1_2_2(or_999_nl, mux_939_nl, fsm_output[6]);
  assign mux_943_nl = MUX_s_1_2_2(mux_942_nl, mux_940_nl, fsm_output[2]);
  assign or_1383_nl = (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[3]) | (~
      (fsm_output[4]));
  assign mux_935_nl = MUX_s_1_2_2(mux_tmp_156, (~ or_216_cse), and_389_cse);
  assign mux_936_nl = MUX_s_1_2_2(or_1383_nl, mux_935_nl, fsm_output[5]);
  assign mux_937_nl = MUX_s_1_2_2(mux_936_nl, or_171_cse, fsm_output[6]);
  assign nand_117_nl = ~((fsm_output[5]) & or_tmp_891);
  assign or_996_nl = (fsm_output[0]) | (~ (fsm_output[1])) | (fsm_output[3]) | (~
      (fsm_output[4]));
  assign mux_933_nl = MUX_s_1_2_2(or_216_cse, or_996_nl, fsm_output[5]);
  assign mux_934_nl = MUX_s_1_2_2(nand_117_nl, mux_933_nl, fsm_output[6]);
  assign mux_938_nl = MUX_s_1_2_2(mux_937_nl, mux_934_nl, fsm_output[2]);
  assign mux_944_nl = MUX_s_1_2_2(mux_943_nl, mux_938_nl, fsm_output[7]);
  assign mux_313_nl = MUX_s_1_2_2((~ or_tmp_113), and_705_cse, fsm_output[5]);
  assign or_231_nl = (fsm_output[6]) | mux_313_nl;
  assign mux_930_nl = MUX_s_1_2_2(mux_tmp_719, (fsm_output[4]), fsm_output[5]);
  assign or_992_nl = (fsm_output[6]) | mux_930_nl;
  assign mux_932_nl = MUX_s_1_2_2(or_231_nl, or_992_nl, fsm_output[2]);
  assign or_994_nl = (fsm_output[7]) | mux_932_nl;
  assign mux_945_nl = MUX_s_1_2_2(mux_944_nl, or_994_nl, fsm_output[8]);
  assign nl_COMP_LOOP_1_acc_8_nl = tmp_10_lpi_4_dfm - modulo_result_mux_1_cse;
  assign COMP_LOOP_1_acc_8_nl = nl_COMP_LOOP_1_acc_8_nl[63:0];
  assign or_1146_nl = (fsm_output[9]) | (~ (fsm_output[4])) | (fsm_output[6]) | (~
      (fsm_output[3])) | (fsm_output[8]);
  assign or_1145_nl = (~ (fsm_output[9])) | (~ (fsm_output[4])) | (fsm_output[6])
      | (fsm_output[3]) | (fsm_output[8]);
  assign mux_1137_nl = MUX_s_1_2_2(or_1146_nl, or_1145_nl, fsm_output[0]);
  assign nor_334_nl = ~((~ (fsm_output[7])) | (fsm_output[5]) | mux_1137_nl);
  assign or_1142_nl = (~ (fsm_output[4])) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[8]);
  assign or_1141_nl = (fsm_output[4]) | (fsm_output[6]) | (~ (fsm_output[3])) | (fsm_output[8]);
  assign mux_1135_nl = MUX_s_1_2_2(or_1142_nl, or_1141_nl, fsm_output[9]);
  assign nor_335_nl = ~((~ (fsm_output[5])) | (fsm_output[0]) | mux_1135_nl);
  assign and_321_nl = (fsm_output[5]) & (fsm_output[0]) & (~ (fsm_output[9])) & (fsm_output[4])
      & (fsm_output[6]) & (fsm_output[3]) & (~ (fsm_output[8]));
  assign mux_1136_nl = MUX_s_1_2_2(nor_335_nl, and_321_nl, fsm_output[7]);
  assign mux_1138_nl = MUX_s_1_2_2(nor_334_nl, mux_1136_nl, fsm_output[2]);
  assign or_1137_nl = (~ (fsm_output[0])) | (fsm_output[9]) | (fsm_output[4]) | (fsm_output[6])
      | (~ (fsm_output[3])) | (fsm_output[8]);
  assign or_1136_nl = (fsm_output[0]) | (fsm_output[9]) | (fsm_output[4]) | (~ (fsm_output[6]))
      | (fsm_output[3]) | (~ (fsm_output[8]));
  assign mux_1133_nl = MUX_s_1_2_2(or_1137_nl, or_1136_nl, fsm_output[5]);
  assign nor_336_nl = ~((fsm_output[7]) | mux_1133_nl);
  assign nor_337_nl = ~((~ (fsm_output[0])) | (fsm_output[9]) | (fsm_output[4]) |
      (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[8])));
  assign nor_338_nl = ~((fsm_output[0]) | (~ (fsm_output[9])) | (~ (fsm_output[4]))
      | (~ (fsm_output[6])) | (fsm_output[3]) | (fsm_output[8]));
  assign mux_1132_nl = MUX_s_1_2_2(nor_337_nl, nor_338_nl, fsm_output[5]);
  assign and_322_nl = (fsm_output[7]) & mux_1132_nl;
  assign mux_1134_nl = MUX_s_1_2_2(nor_336_nl, and_322_nl, fsm_output[2]);
  assign mux_1139_nl = MUX_s_1_2_2(mux_1138_nl, mux_1134_nl, fsm_output[1]);
  assign nand_98_nl = ~((fsm_output[6:5]==2'b11) & or_216_cse);
  assign nand_99_nl = ~((fsm_output[6:5]==2'b11) & or_tmp_103);
  assign mux_1155_nl = MUX_s_1_2_2(nand_98_nl, nand_99_nl, fsm_output[2]);
  assign mux_1156_nl = MUX_s_1_2_2(mux_tmp_886, mux_1155_nl, fsm_output[7]);
  assign COMP_LOOP_COMP_LOOP_and_145_nl = (COMP_LOOP_acc_1_cse_6_sva_1[2:0]==3'b110);
  assign nl_COMP_LOOP_1_acc_nl = ({COMP_LOOP_k_9_3_sva_2 , 3'b000}) + ({1'b1 , (~
      (STAGE_LOOP_lshift_psp_sva[9:1]))}) + 10'b0000000001;
  assign COMP_LOOP_1_acc_nl = nl_COMP_LOOP_1_acc_nl[9:0];
  assign mux_1174_nl = MUX_s_1_2_2(mux_tmp_1170, and_tmp_44, fsm_output[6]);
  assign mux_1171_nl = MUX_s_1_2_2(mux_tmp_1170, mux_tmp_1164, or_1189_cse);
  assign mux_1167_nl = MUX_s_1_2_2(mux_tmp_1160, mux_tmp_1159, fsm_output[2]);
  assign mux_1168_nl = MUX_s_1_2_2(and_tmp_44, mux_1167_nl, fsm_output[3]);
  assign mux_1169_nl = MUX_s_1_2_2(mux_1168_nl, mux_tmp_1162, fsm_output[0]);
  assign mux_1172_nl = MUX_s_1_2_2(mux_1171_nl, mux_1169_nl, fsm_output[6]);
  assign and_315_nl = (fsm_output[7]) & (fsm_output[9]);
  assign mux_1163_nl = MUX_s_1_2_2(not_tmp_482, and_315_nl, fsm_output[8]);
  assign mux_1165_nl = MUX_s_1_2_2(mux_tmp_1164, mux_1163_nl, and_316_cse);
  assign mux_1166_nl = MUX_s_1_2_2(mux_1165_nl, mux_tmp_1162, fsm_output[6]);
  assign mux_1173_nl = MUX_s_1_2_2(mux_1172_nl, mux_1166_nl, fsm_output[1]);
  assign mux_1179_nl = MUX_s_1_2_2(mux_tmp_1178, and_tmp_46, fsm_output[3]);
  assign and_313_nl = (fsm_output[0]) & (fsm_output[3]);
  assign mux_1177_nl = MUX_s_1_2_2(and_tmp_46, and_tmp_45, and_313_nl);
  assign mux_1180_nl = MUX_s_1_2_2(mux_1179_nl, mux_1177_nl, fsm_output[1]);
  assign mux_1176_nl = MUX_s_1_2_2(and_tmp_46, and_tmp_45, fsm_output[3]);
  assign mux_1181_nl = MUX_s_1_2_2(mux_1180_nl, mux_1176_nl, fsm_output[2]);
  assign or_1193_nl = (fsm_output[6]) | ((fsm_output[5]) & and_705_cse);
  assign mux_1183_nl = MUX_s_1_2_2(or_1193_nl, or_tmp_916, fsm_output[2]);
  assign nand_234_nl = ~((fsm_output[7]) & mux_1183_nl);
  assign mux_1184_nl = MUX_s_1_2_2(or_tmp_918, nand_234_nl, fsm_output[8]);
  assign nl_COMP_LOOP_acc_11_psp_sva  = (VEC_LOOP_j_sva_11_0[11:1]) + conv_u2u_8_11({COMP_LOOP_k_9_3_sva_5_0
      , 2'b01});
  assign and_272_nl = (fsm_output[6]) & or_171_cse;
  assign and_271_nl = (fsm_output[6]) & or_1202_cse;
  assign mux_1185_nl = MUX_s_1_2_2(and_272_nl, and_271_nl, fsm_output[2]);
  assign nor_328_nl = ~((fsm_output[7]) | mux_1185_nl);
  assign mux_1186_nl = MUX_s_1_2_2(or_tmp_918, nor_328_nl, fsm_output[8]);
  assign or_100_nl = (fsm_output[6:5]!=2'b00) | nor_tmp;
  assign or_1197_nl = (fsm_output[6:5]!=2'b00) | nor_tmp_23;
  assign mux_1187_nl = MUX_s_1_2_2(or_100_nl, or_1197_nl, fsm_output[2]);
  assign or_1200_nl = (fsm_output[8:7]!=2'b00) | mux_1187_nl;
  assign nl_COMP_LOOP_acc_14_psp_sva  = (VEC_LOOP_j_sva_11_0[11:1]) + conv_u2u_8_11({COMP_LOOP_k_9_3_sva_5_0
      , 2'b11});
  assign or_1201_nl = (fsm_output[8]) | ((fsm_output[7:5]==3'b111));
  assign nor_327_nl = ~((fsm_output[3]) | (fsm_output[2]) | (fsm_output[1]) | (fsm_output[8])
      | (fsm_output[9]));
  assign mux_1191_nl = MUX_s_1_2_2(nor_393_cse, nor_327_nl, and_314_cse);
  assign and_274_nl = (fsm_output[2]) & or_838_cse & (fsm_output[9:8]==2'b11);
  assign mux_1190_nl = MUX_s_1_2_2(and_274_nl, and_369_cse, or_1202_cse);
  assign mux_1192_nl = MUX_s_1_2_2(mux_1191_nl, mux_1190_nl, fsm_output[6]);
  assign COMP_LOOP_COMP_LOOP_or_7_nl = (VEC_LOOP_j_sva_11_0[11]) | and_dcpl_243 |
      and_dcpl_247 | and_dcpl_255 | and_dcpl_260 | and_dcpl_266;
  assign COMP_LOOP_COMP_LOOP_mux_8_nl = MUX_v_9_2_2((VEC_LOOP_j_sva_11_0[10:2]),
      (~ (STAGE_LOOP_lshift_psp_sva[9:1])), COMP_LOOP_or_40_itm);
  assign COMP_LOOP_or_44_nl = (~ and_511_cse) | and_dcpl_243 | and_dcpl_247 | and_dcpl_255
      | and_dcpl_260 | and_dcpl_266;
  assign COMP_LOOP_COMP_LOOP_mux_9_nl = MUX_v_6_2_2(({2'b00 , (COMP_LOOP_k_9_3_sva_5_0[5:2])}),
      COMP_LOOP_k_9_3_sva_5_0, COMP_LOOP_or_40_itm);
  assign COMP_LOOP_COMP_LOOP_or_8_nl = ((COMP_LOOP_k_9_3_sva_5_0[1]) & (~(and_dcpl_243
      | and_dcpl_247))) | and_dcpl_255 | and_dcpl_260 | and_dcpl_266;
  assign COMP_LOOP_COMP_LOOP_or_9_nl = ((COMP_LOOP_k_9_3_sva_5_0[0]) & (~(and_dcpl_243
      | and_dcpl_255 | and_dcpl_260))) | and_dcpl_247 | and_dcpl_266;
  assign COMP_LOOP_COMP_LOOP_or_10_nl = (~(and_dcpl_247 | and_dcpl_255 | and_dcpl_266))
      | and_511_cse | and_dcpl_243 | and_dcpl_260;
  assign nl_acc_nl = ({COMP_LOOP_COMP_LOOP_or_7_nl , COMP_LOOP_COMP_LOOP_mux_8_nl
      , COMP_LOOP_or_44_nl}) + conv_u2u_10_11({COMP_LOOP_COMP_LOOP_mux_9_nl , COMP_LOOP_COMP_LOOP_or_8_nl
      , COMP_LOOP_COMP_LOOP_or_9_nl , COMP_LOOP_COMP_LOOP_or_10_nl , 1'b1});
  assign acc_nl = nl_acc_nl[10:0];
  assign z_out = readslicef_11_10_1(acc_nl);
  assign and_722_nl = nor_tmp & (fsm_output[1]) & (~ (fsm_output[9])) & (~ (fsm_output[8]))
      & and_dcpl_269 & and_dcpl;
  assign and_723_nl = (~ (fsm_output[3])) & (~ (fsm_output[4])) & (~ (fsm_output[1]))
      & and_dcpl_11 & (~ (fsm_output[7])) & (fsm_output[5]) & (fsm_output[2]) & and_dcpl_276;
  assign and_724_nl = and_dcpl_100 & (~ (fsm_output[1])) & and_dcpl_11 & (fsm_output[7])
      & (~ (fsm_output[5])) & (~ (fsm_output[2])) & and_dcpl;
  assign and_725_nl = and_dcpl_100 & (fsm_output[1]) & and_dcpl_11 & and_dcpl_269
      & (fsm_output[6]) & (~ (fsm_output[0]));
  assign and_726_nl = (~ (fsm_output[3])) & (fsm_output[4]) & (fsm_output[1]) & and_dcpl_23
      & and_dcpl_298 & (~ (fsm_output[2])) & (fsm_output[6]) & (fsm_output[0]);
  assign COMP_LOOP_mux1h_125_nl = MUX1HOT_v_3_6_2(3'b001, 3'b010, 3'b011, 3'b100,
      3'b101, 3'b110, {and_722_nl , and_723_nl , and_724_nl , and_725_nl , and_726_nl
      , and_dcpl_399});
  assign and_727_nl = and_dcpl_128 & (fsm_output[9:8]==2'b11) & and_dcpl_298 & (fsm_output[2])
      & and_dcpl;
  assign COMP_LOOP_or_45_nl = MUX_v_3_2_2(COMP_LOOP_mux1h_125_nl, 3'b111, and_727_nl);
  assign nl_z_out_1 = STAGE_LOOP_lshift_psp_sva + conv_u2u_9_10({COMP_LOOP_k_9_3_sva_5_0
      , COMP_LOOP_or_45_nl});
  assign z_out_1 = nl_z_out_1[9:0];
  assign COMP_LOOP_mux1h_126_nl = MUX1HOT_v_64_4_2(({58'b0000000000000000000000000000000000000000000000000000000001
      , (~ (STAGE_LOOP_lshift_psp_sva[9:4]))}), ({52'b0000000000000000000000000000000000000000000000000000
      , VEC_LOOP_j_sva_11_0}), p_sva, ({57'b000000000000000000000000000000000000000000000000000000000
      , (STAGE_LOOP_lshift_psp_sva[9:3])}), {and_dcpl_324 , and_511_cse , and_dcpl_340
      , and_dcpl_345});
  assign COMP_LOOP_or_46_nl = (~(and_511_cse | and_dcpl_340 | and_dcpl_345)) | and_dcpl_324;
  assign COMP_LOOP_COMP_LOOP_or_11_nl = (~(and_dcpl_324 | and_511_cse | and_dcpl_345))
      | and_dcpl_340;
  assign COMP_LOOP_nor_107_nl = ~(and_dcpl_324 | and_dcpl_345);
  assign COMP_LOOP_and_85_nl = MUX_v_3_2_2(3'b000, (COMP_LOOP_k_9_3_sva_5_0[5:3]),
      COMP_LOOP_nor_107_nl);
  assign COMP_LOOP_COMP_LOOP_or_12_nl = MUX_v_3_2_2(COMP_LOOP_and_85_nl, 3'b111,
      and_dcpl_340);
  assign COMP_LOOP_mux_41_nl = MUX_v_6_2_2(COMP_LOOP_k_9_3_sva_5_0, ({(COMP_LOOP_k_9_3_sva_5_0[2:0])
      , 3'b111}), and_511_cse);
  assign COMP_LOOP_COMP_LOOP_or_13_nl = MUX_v_6_2_2(COMP_LOOP_mux_41_nl, 6'b111111,
      and_dcpl_340);
  assign nl_acc_2_nl = conv_u2u_65_66({COMP_LOOP_mux1h_126_nl , COMP_LOOP_or_46_nl})
      + conv_s2u_11_66({COMP_LOOP_COMP_LOOP_or_11_nl , COMP_LOOP_COMP_LOOP_or_12_nl
      , COMP_LOOP_COMP_LOOP_or_13_nl , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[65:0];
  assign z_out_2 = readslicef_66_65_1(acc_2_nl);
  assign operator_64_false_1_operator_64_false_1_or_53_nl = (~(and_dcpl_354 | and_dcpl_368
      | and_dcpl_372 | and_dcpl_379 | and_dcpl_385 | and_dcpl_388 | and_dcpl_394
      | and_dcpl_399 | and_dcpl_404 | and_dcpl_406)) | not_tmp_581 | and_dcpl_362
      | and_dcpl_411 | and_dcpl_409;
  assign operator_64_false_1_operator_64_false_1_or_54_nl = (~((operator_66_true_div_cmp_z[63])
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_362 | and_dcpl_411;
  assign operator_64_false_1_mux_51_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[62]),
      (operator_66_true_div_cmp_z[62]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_55_nl = (~(operator_64_false_1_mux_51_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_52_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[61]),
      (operator_66_true_div_cmp_z[61]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_56_nl = (~(operator_64_false_1_mux_52_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_53_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[60]),
      (operator_66_true_div_cmp_z[60]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_57_nl = (~(operator_64_false_1_mux_53_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_54_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[59]),
      (operator_66_true_div_cmp_z[59]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_58_nl = (~(operator_64_false_1_mux_54_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_55_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[58]),
      (operator_66_true_div_cmp_z[58]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_59_nl = (~(operator_64_false_1_mux_55_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_56_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[57]),
      (operator_66_true_div_cmp_z[57]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_60_nl = (~(operator_64_false_1_mux_56_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_57_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[56]),
      (operator_66_true_div_cmp_z[56]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_61_nl = (~(operator_64_false_1_mux_57_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_58_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[55]),
      (operator_66_true_div_cmp_z[55]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_62_nl = (~(operator_64_false_1_mux_58_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_59_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[54]),
      (operator_66_true_div_cmp_z[54]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_63_nl = (~(operator_64_false_1_mux_59_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_60_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[53]),
      (operator_66_true_div_cmp_z[53]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_64_nl = (~(operator_64_false_1_mux_60_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_61_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[52]),
      (operator_66_true_div_cmp_z[52]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_65_nl = (~(operator_64_false_1_mux_61_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_62_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[51]),
      (operator_66_true_div_cmp_z[51]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_66_nl = (~(operator_64_false_1_mux_62_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_63_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[50]),
      (operator_66_true_div_cmp_z[50]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_67_nl = (~(operator_64_false_1_mux_63_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_64_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[49]),
      (operator_66_true_div_cmp_z[49]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_68_nl = (~(operator_64_false_1_mux_64_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_65_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[48]),
      (operator_66_true_div_cmp_z[48]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_69_nl = (~(operator_64_false_1_mux_65_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_66_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[47]),
      (operator_66_true_div_cmp_z[47]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_70_nl = (~(operator_64_false_1_mux_66_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_67_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[46]),
      (operator_66_true_div_cmp_z[46]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_71_nl = (~(operator_64_false_1_mux_67_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_68_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[45]),
      (operator_66_true_div_cmp_z[45]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_72_nl = (~(operator_64_false_1_mux_68_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_69_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[44]),
      (operator_66_true_div_cmp_z[44]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_73_nl = (~(operator_64_false_1_mux_69_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_70_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[43]),
      (operator_66_true_div_cmp_z[43]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_74_nl = (~(operator_64_false_1_mux_70_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_71_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[42]),
      (operator_66_true_div_cmp_z[42]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_75_nl = (~(operator_64_false_1_mux_71_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_72_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[41]),
      (operator_66_true_div_cmp_z[41]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_76_nl = (~(operator_64_false_1_mux_72_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_73_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[40]),
      (operator_66_true_div_cmp_z[40]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_77_nl = (~(operator_64_false_1_mux_73_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_74_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[39]),
      (operator_66_true_div_cmp_z[39]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_78_nl = (~(operator_64_false_1_mux_74_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_75_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[38]),
      (operator_66_true_div_cmp_z[38]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_79_nl = (~(operator_64_false_1_mux_75_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_76_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[37]),
      (operator_66_true_div_cmp_z[37]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_80_nl = (~(operator_64_false_1_mux_76_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_77_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[36]),
      (operator_66_true_div_cmp_z[36]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_81_nl = (~(operator_64_false_1_mux_77_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_78_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[35]),
      (operator_66_true_div_cmp_z[35]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_82_nl = (~(operator_64_false_1_mux_78_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_79_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[34]),
      (operator_66_true_div_cmp_z[34]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_83_nl = (~(operator_64_false_1_mux_79_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_80_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[33]),
      (operator_66_true_div_cmp_z[33]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_84_nl = (~(operator_64_false_1_mux_80_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_81_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[32]),
      (operator_66_true_div_cmp_z[32]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_85_nl = (~(operator_64_false_1_mux_81_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_82_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[31]),
      (operator_66_true_div_cmp_z[31]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_86_nl = (~(operator_64_false_1_mux_82_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_83_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[30]),
      (operator_66_true_div_cmp_z[30]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_87_nl = (~(operator_64_false_1_mux_83_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_84_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[29]),
      (operator_66_true_div_cmp_z[29]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_88_nl = (~(operator_64_false_1_mux_84_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_85_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[28]),
      (operator_66_true_div_cmp_z[28]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_89_nl = (~(operator_64_false_1_mux_85_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_86_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[27]),
      (operator_66_true_div_cmp_z[27]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_90_nl = (~(operator_64_false_1_mux_86_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_87_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[26]),
      (operator_66_true_div_cmp_z[26]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_91_nl = (~(operator_64_false_1_mux_87_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_88_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[25]),
      (operator_66_true_div_cmp_z[25]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_92_nl = (~(operator_64_false_1_mux_88_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_89_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[24]),
      (operator_66_true_div_cmp_z[24]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_93_nl = (~(operator_64_false_1_mux_89_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_90_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[23]),
      (operator_66_true_div_cmp_z[23]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_94_nl = (~(operator_64_false_1_mux_90_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_91_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[22]),
      (operator_66_true_div_cmp_z[22]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_95_nl = (~(operator_64_false_1_mux_91_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_92_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[21]),
      (operator_66_true_div_cmp_z[21]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_96_nl = (~(operator_64_false_1_mux_92_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_93_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[20]),
      (operator_66_true_div_cmp_z[20]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_97_nl = (~(operator_64_false_1_mux_93_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_94_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[19]),
      (operator_66_true_div_cmp_z[19]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_98_nl = (~(operator_64_false_1_mux_94_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_95_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[18]),
      (operator_66_true_div_cmp_z[18]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_99_nl = (~(operator_64_false_1_mux_95_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_96_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[17]),
      (operator_66_true_div_cmp_z[17]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_100_nl = (~(operator_64_false_1_mux_96_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_97_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[16]),
      (operator_66_true_div_cmp_z[16]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_101_nl = (~(operator_64_false_1_mux_97_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_98_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[15]),
      (operator_66_true_div_cmp_z[15]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_102_nl = (~(operator_64_false_1_mux_98_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_99_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[14]),
      (operator_66_true_div_cmp_z[14]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_103_nl = (~(operator_64_false_1_mux_99_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_100_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[13]),
      (operator_66_true_div_cmp_z[13]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_104_nl = (~(operator_64_false_1_mux_100_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux_101_nl = MUX_s_1_2_2((operator_64_false_acc_mut_63_0[12]),
      (operator_66_true_div_cmp_z[12]), and_dcpl_409);
  assign operator_64_false_1_operator_64_false_1_or_105_nl = (~(operator_64_false_1_mux_101_nl
      | and_dcpl_354 | and_dcpl_368 | and_dcpl_372 | and_dcpl_379 | and_dcpl_385
      | and_dcpl_388 | and_dcpl_394 | and_dcpl_399 | and_dcpl_404 | and_dcpl_406))
      | not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_mux1h_4_nl = MUX1HOT_v_4_3_2((operator_64_false_acc_mut_63_0[11:8]),
      (~ (VEC_LOOP_j_sva_11_0[11:8])), (operator_66_true_div_cmp_z[11:8]), {and_dcpl_362
      , operator_64_false_1_or_1_itm , and_dcpl_409});
  assign operator_64_false_1_operator_64_false_1_nor_105_nl = ~(MUX_v_4_2_2(operator_64_false_1_mux1h_4_nl,
      4'b1111, and_dcpl_354));
  assign operator_64_false_1_or_8_nl = not_tmp_581 | and_dcpl_411;
  assign operator_64_false_1_or_7_nl = MUX_v_4_2_2(operator_64_false_1_operator_64_false_1_nor_105_nl,
      4'b1111, operator_64_false_1_or_8_nl);
  assign operator_64_false_1_mux1h_5_nl = MUX1HOT_v_8_6_2(({2'b01 , (~ COMP_LOOP_k_9_3_sva_5_0)}),
      ({(~ modExp_exp_1_7_1_sva) , (~ modExp_exp_1_6_1_sva) , (~ modExp_exp_1_5_1_sva)
      , (~ modExp_exp_1_4_1_sva) , (~ modExp_exp_1_3_1_sva) , (~ modExp_exp_1_2_1_sva)
      , (~ modExp_exp_1_1_1_sva) , (~ modExp_exp_1_0_1_sva_1)}), (~ (operator_64_false_acc_mut_63_0[7:0])),
      (VEC_LOOP_j_sva_11_0[7:0]), (~ (operator_66_true_div_cmp_z[7:0])), ({(~ modExp_exp_1_1_1_sva)
      , (~ modExp_exp_1_7_1_sva) , (~ modExp_exp_1_6_1_sva) , (~ modExp_exp_1_5_1_sva)
      , (~ modExp_exp_1_4_1_sva) , (~ modExp_exp_1_3_1_sva) , (~ modExp_exp_1_2_1_sva)
      , (~ modExp_exp_1_0_1_sva_1)}), {and_dcpl_354 , not_tmp_581 , and_dcpl_362
      , operator_64_false_1_or_1_itm , and_dcpl_409 , and_dcpl_411});
  assign operator_64_false_1_mux1h_6_nl = MUX1HOT_v_7_3_2((z_out_2[6:0]), (z_out_1[9:3]),
      (STAGE_LOOP_lshift_psp_sva[9:3]), {and_dcpl_368 , operator_64_false_1_or_5_ssc
      , and_dcpl_406});
  assign operator_64_false_1_not_3_nl = ~ operator_64_false_1_or_4_ssc;
  assign operator_64_false_1_and_53_nl = MUX_v_7_2_2(7'b0000000, operator_64_false_1_mux1h_6_nl,
      operator_64_false_1_not_3_nl);
  assign operator_64_false_1_or_9_nl = and_dcpl_368 | and_dcpl_406;
  assign operator_64_false_1_mux1h_7_nl = MUX1HOT_v_3_3_2(3'b001, (STAGE_LOOP_lshift_psp_sva[2:0]),
      (z_out_1[2:0]), {operator_64_false_1_or_4_ssc , operator_64_false_1_or_9_nl
      , operator_64_false_1_or_5_ssc});
  assign nl_z_out_3 = ({operator_64_false_1_operator_64_false_1_or_53_nl , operator_64_false_1_operator_64_false_1_or_54_nl
      , operator_64_false_1_operator_64_false_1_or_55_nl , operator_64_false_1_operator_64_false_1_or_56_nl
      , operator_64_false_1_operator_64_false_1_or_57_nl , operator_64_false_1_operator_64_false_1_or_58_nl
      , operator_64_false_1_operator_64_false_1_or_59_nl , operator_64_false_1_operator_64_false_1_or_60_nl
      , operator_64_false_1_operator_64_false_1_or_61_nl , operator_64_false_1_operator_64_false_1_or_62_nl
      , operator_64_false_1_operator_64_false_1_or_63_nl , operator_64_false_1_operator_64_false_1_or_64_nl
      , operator_64_false_1_operator_64_false_1_or_65_nl , operator_64_false_1_operator_64_false_1_or_66_nl
      , operator_64_false_1_operator_64_false_1_or_67_nl , operator_64_false_1_operator_64_false_1_or_68_nl
      , operator_64_false_1_operator_64_false_1_or_69_nl , operator_64_false_1_operator_64_false_1_or_70_nl
      , operator_64_false_1_operator_64_false_1_or_71_nl , operator_64_false_1_operator_64_false_1_or_72_nl
      , operator_64_false_1_operator_64_false_1_or_73_nl , operator_64_false_1_operator_64_false_1_or_74_nl
      , operator_64_false_1_operator_64_false_1_or_75_nl , operator_64_false_1_operator_64_false_1_or_76_nl
      , operator_64_false_1_operator_64_false_1_or_77_nl , operator_64_false_1_operator_64_false_1_or_78_nl
      , operator_64_false_1_operator_64_false_1_or_79_nl , operator_64_false_1_operator_64_false_1_or_80_nl
      , operator_64_false_1_operator_64_false_1_or_81_nl , operator_64_false_1_operator_64_false_1_or_82_nl
      , operator_64_false_1_operator_64_false_1_or_83_nl , operator_64_false_1_operator_64_false_1_or_84_nl
      , operator_64_false_1_operator_64_false_1_or_85_nl , operator_64_false_1_operator_64_false_1_or_86_nl
      , operator_64_false_1_operator_64_false_1_or_87_nl , operator_64_false_1_operator_64_false_1_or_88_nl
      , operator_64_false_1_operator_64_false_1_or_89_nl , operator_64_false_1_operator_64_false_1_or_90_nl
      , operator_64_false_1_operator_64_false_1_or_91_nl , operator_64_false_1_operator_64_false_1_or_92_nl
      , operator_64_false_1_operator_64_false_1_or_93_nl , operator_64_false_1_operator_64_false_1_or_94_nl
      , operator_64_false_1_operator_64_false_1_or_95_nl , operator_64_false_1_operator_64_false_1_or_96_nl
      , operator_64_false_1_operator_64_false_1_or_97_nl , operator_64_false_1_operator_64_false_1_or_98_nl
      , operator_64_false_1_operator_64_false_1_or_99_nl , operator_64_false_1_operator_64_false_1_or_100_nl
      , operator_64_false_1_operator_64_false_1_or_101_nl , operator_64_false_1_operator_64_false_1_or_102_nl
      , operator_64_false_1_operator_64_false_1_or_103_nl , operator_64_false_1_operator_64_false_1_or_104_nl
      , operator_64_false_1_operator_64_false_1_or_105_nl , operator_64_false_1_or_7_nl
      , operator_64_false_1_mux1h_5_nl}) + conv_u2u_10_65({operator_64_false_1_and_53_nl
      , operator_64_false_1_mux1h_7_nl});
  assign z_out_3 = nl_z_out_3[64:0];
  assign and_728_nl = (~ (fsm_output[4])) & (fsm_output[3]) & (fsm_output[1]) & nor_393_cse
      & and_dcpl_238 & and_dcpl_276;
  assign nor_690_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (fsm_output[8]) |
      (fsm_output[9]) | (fsm_output[1]) | not_tmp_309);
  assign or_1560_nl = (fsm_output[1]) | (fsm_output[3]) | (~ (fsm_output[4]));
  assign or_1561_nl = (fsm_output[1]) | (~ (fsm_output[3])) | (fsm_output[4]);
  assign mux_1462_nl = MUX_s_1_2_2(or_1560_nl, or_1561_nl, fsm_output[9]);
  assign nor_691_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[8]) |
      mux_1462_nl);
  assign mux_1461_nl = MUX_s_1_2_2(nor_690_nl, nor_691_nl, fsm_output[2]);
  assign nor_692_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (~ (fsm_output[8]))
      | (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[3]) | (fsm_output[4]));
  assign and_729_nl = (fsm_output[5]) & (fsm_output[7]) & (~ (fsm_output[8])) & (fsm_output[9])
      & (fsm_output[1]) & (~ (fsm_output[3])) & (fsm_output[4]);
  assign mux_1463_nl = MUX_s_1_2_2(nor_692_nl, and_729_nl, fsm_output[2]);
  assign mux_1460_nl = MUX_s_1_2_2(mux_1461_nl, mux_1463_nl, fsm_output[6]);
  assign or_1562_nl = (fsm_output[8]) | (fsm_output[9]) | (~ (fsm_output[1])) | (~
      (fsm_output[3])) | (fsm_output[4]);
  assign mux_1465_nl = MUX_s_1_2_2(or_1562_nl, or_1440_cse, fsm_output[7]);
  assign nor_693_nl = ~((fsm_output[2]) | (fsm_output[5]) | mux_1465_nl);
  assign nor_694_nl = ~((~ (fsm_output[7])) | (~ (fsm_output[8])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (fsm_output[3]) | (fsm_output[4]));
  assign nor_695_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (fsm_output[9]) |
      (fsm_output[1]) | not_tmp_309);
  assign mux_1466_nl = MUX_s_1_2_2(nor_694_nl, nor_695_nl, fsm_output[5]);
  assign and_730_nl = (fsm_output[2]) & mux_1466_nl;
  assign mux_1464_nl = MUX_s_1_2_2(nor_693_nl, and_730_nl, fsm_output[6]);
  assign mux_1459_nl = MUX_s_1_2_2(mux_1460_nl, mux_1464_nl, fsm_output[0]);
  assign nor_696_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (fsm_output[2]) |
      (fsm_output[9]) | not_tmp_600);
  assign nor_697_nl = ~((fsm_output[7]) | (fsm_output[8]) | (~ (fsm_output[2])) |
      (~ (fsm_output[9])) | (fsm_output[4]) | (~ (fsm_output[0])));
  assign mux_1469_nl = MUX_s_1_2_2(nor_696_nl, nor_697_nl, fsm_output[5]);
  assign nand_279_nl = ~((fsm_output[3]) & mux_1469_nl);
  assign or_1564_nl = (fsm_output[8]) | (fsm_output[2]) | (fsm_output[9]) | (fsm_output[4])
      | (~ (fsm_output[0]));
  assign mux_1472_nl = MUX_s_1_2_2(or_tmp_1346, or_1564_nl, fsm_output[7]);
  assign or_1565_nl = (~ (fsm_output[7])) | (~ (fsm_output[8])) | (fsm_output[2])
      | (fsm_output[9]) | (~ (fsm_output[4])) | (fsm_output[0]);
  assign mux_1471_nl = MUX_s_1_2_2(mux_1472_nl, or_1565_nl, fsm_output[5]);
  assign or_1567_nl = (fsm_output[8]) | (~ (fsm_output[2])) | (fsm_output[9]) | (~
      (fsm_output[4])) | (fsm_output[0]);
  assign or_1568_nl = (~ (fsm_output[8])) | (fsm_output[2]) | (fsm_output[9]) | (fsm_output[4])
      | (fsm_output[0]);
  assign mux_1473_nl = MUX_s_1_2_2(or_1567_nl, or_1568_nl, fsm_output[7]);
  assign or_1566_nl = (fsm_output[5]) | mux_1473_nl;
  assign mux_1470_nl = MUX_s_1_2_2(mux_1471_nl, or_1566_nl, fsm_output[3]);
  assign mux_1468_nl = MUX_s_1_2_2(nand_279_nl, mux_1470_nl, fsm_output[6]);
  assign or_1570_nl = (fsm_output[2]) | (fsm_output[9]) | not_tmp_600;
  assign or_1571_nl = (~ (fsm_output[2])) | (fsm_output[9]) | (fsm_output[4]) | (fsm_output[0]);
  assign mux_1477_nl = MUX_s_1_2_2(or_1570_nl, or_1571_nl, fsm_output[8]);
  assign or_1569_nl = (fsm_output[7]) | mux_1477_nl;
  assign mux_1476_nl = MUX_s_1_2_2(or_tmp_1349, or_1569_nl, fsm_output[5]);
  assign nand_280_nl = ~((fsm_output[8]) & (fsm_output[2]) & (fsm_output[9]) & (fsm_output[4])
      & (fsm_output[0]));
  assign mux_1479_nl = MUX_s_1_2_2(nand_280_nl, or_tmp_1348, fsm_output[7]);
  assign mux_1478_nl = MUX_s_1_2_2(mux_1479_nl, or_tmp_1349, fsm_output[5]);
  assign mux_1475_nl = MUX_s_1_2_2(mux_1476_nl, mux_1478_nl, fsm_output[3]);
  assign mux_1481_nl = MUX_s_1_2_2(or_tmp_1348, or_tmp_1346, fsm_output[7]);
  assign nand_281_nl = ~((fsm_output[5]) & (~ mux_1481_nl));
  assign or_1572_nl = (~ (fsm_output[5])) | (~ (fsm_output[7])) | (fsm_output[8])
      | (~ (fsm_output[2])) | (fsm_output[9]) | (~ (fsm_output[4])) | (fsm_output[0]);
  assign mux_1480_nl = MUX_s_1_2_2(nand_281_nl, or_1572_nl, fsm_output[3]);
  assign mux_1474_nl = MUX_s_1_2_2(mux_1475_nl, mux_1480_nl, fsm_output[6]);
  assign mux_1467_nl = MUX_s_1_2_2(mux_1468_nl, mux_1474_nl, fsm_output[1]);
  assign modExp_while_if_mux1h_2_nl = MUX1HOT_v_64_3_2(modExp_result_sva, COMP_LOOP_1_mul_mut,
      operator_64_false_acc_mut_63_0, {and_728_nl , mux_1459_nl , (~ mux_1467_nl)});
  assign nl_z_out_4 = $signed(conv_u2s_64_65(modExp_while_if_mux1h_2_nl)) * $signed(COMP_LOOP_1_mul_mut);
  assign z_out_4 = nl_z_out_4[63:0];

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_7_2;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [6:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_6_2;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [5:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    result = result | ( input_4 & {3{sel[4]}});
    result = result | ( input_5 & {3{sel[5]}});
    MUX1HOT_v_3_6_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_13_2;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [12:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    MUX1HOT_v_64_13_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_4_2;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [3:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    MUX1HOT_v_64_4_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_5_2;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [4:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    MUX1HOT_v_64_5_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_9_2;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [8:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    MUX1HOT_v_64_9_2 = result;
  end
  endfunction


  function automatic [64:0] MUX1HOT_v_65_3_2;
    input [64:0] input_2;
    input [64:0] input_1;
    input [64:0] input_0;
    input [2:0] sel;
    reg [64:0] result;
  begin
    result = input_0 & {65{sel[0]}};
    result = result | ( input_1 & {65{sel[1]}});
    result = result | ( input_2 & {65{sel[2]}});
    MUX1HOT_v_65_3_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_6_2;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [5:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    result = result | ( input_5 & {8{sel[5]}});
    MUX1HOT_v_8_6_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_11_2;
    input [8:0] input_10;
    input [8:0] input_9;
    input [8:0] input_8;
    input [8:0] input_7;
    input [8:0] input_6;
    input [8:0] input_5;
    input [8:0] input_4;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [10:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    result = result | ( input_3 & {9{sel[3]}});
    result = result | ( input_4 & {9{sel[4]}});
    result = result | ( input_5 & {9{sel[5]}});
    result = result | ( input_6 & {9{sel[6]}});
    result = result | ( input_7 & {9{sel[7]}});
    result = result | ( input_8 & {9{sel[8]}});
    result = result | ( input_9 & {9{sel[9]}});
    result = result | ( input_10 & {9{sel[10]}});
    MUX1HOT_v_9_11_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [0:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [62:0] MUX_v_63_2_2;
    input [62:0] input_0;
    input [62:0] input_1;
    input [0:0] sel;
    reg [62:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_63_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [64:0] MUX_v_65_2_2;
    input [64:0] input_0;
    input [64:0] input_1;
    input [0:0] sel;
    reg [64:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_65_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [9:0] readslicef_11_10_1;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_11_10_1 = tmp[9:0];
  end
  endfunction


  function automatic [0:0] readslicef_3_1_2;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_3_1_2 = tmp[0:0];
  end
  endfunction


  function automatic [64:0] readslicef_66_65_1;
    input [65:0] vector;
    reg [65:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_66_65_1 = tmp[64:0];
  end
  endfunction


  function automatic [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function automatic [65:0] conv_s2u_11_66 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_66 = {{55{vector[10]}}, vector};
  end
  endfunction


  function automatic [64:0] conv_u2s_64_65 ;
    input [63:0]  vector ;
  begin
    conv_u2s_64_65 =  {1'b0, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_6_9 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_9 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_8_11 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_11 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_9_12 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_12 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [64:0] conv_u2u_10_65 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_65 = {{55{1'b0}}, vector};
  end
  endfunction


  function automatic [65:0] conv_u2u_65_66 ;
    input [64:0]  vector ;
  begin
    conv_u2u_65_66 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT
// ------------------------------------------------------------------


module inPlaceNTT_DIT (
  clk, rst, vec_rsc_0_0_adra, vec_rsc_0_0_da, vec_rsc_0_0_wea, vec_rsc_0_0_qa, vec_rsc_triosy_0_0_lz,
      vec_rsc_0_1_adra, vec_rsc_0_1_da, vec_rsc_0_1_wea, vec_rsc_0_1_qa, vec_rsc_triosy_0_1_lz,
      vec_rsc_0_2_adra, vec_rsc_0_2_da, vec_rsc_0_2_wea, vec_rsc_0_2_qa, vec_rsc_triosy_0_2_lz,
      vec_rsc_0_3_adra, vec_rsc_0_3_da, vec_rsc_0_3_wea, vec_rsc_0_3_qa, vec_rsc_triosy_0_3_lz,
      vec_rsc_0_4_adra, vec_rsc_0_4_da, vec_rsc_0_4_wea, vec_rsc_0_4_qa, vec_rsc_triosy_0_4_lz,
      vec_rsc_0_5_adra, vec_rsc_0_5_da, vec_rsc_0_5_wea, vec_rsc_0_5_qa, vec_rsc_triosy_0_5_lz,
      vec_rsc_0_6_adra, vec_rsc_0_6_da, vec_rsc_0_6_wea, vec_rsc_0_6_qa, vec_rsc_triosy_0_6_lz,
      vec_rsc_0_7_adra, vec_rsc_0_7_da, vec_rsc_0_7_wea, vec_rsc_0_7_qa, vec_rsc_triosy_0_7_lz,
      p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz
);
  input clk;
  input rst;
  output [8:0] vec_rsc_0_0_adra;
  output [63:0] vec_rsc_0_0_da;
  output vec_rsc_0_0_wea;
  input [63:0] vec_rsc_0_0_qa;
  output vec_rsc_triosy_0_0_lz;
  output [8:0] vec_rsc_0_1_adra;
  output [63:0] vec_rsc_0_1_da;
  output vec_rsc_0_1_wea;
  input [63:0] vec_rsc_0_1_qa;
  output vec_rsc_triosy_0_1_lz;
  output [8:0] vec_rsc_0_2_adra;
  output [63:0] vec_rsc_0_2_da;
  output vec_rsc_0_2_wea;
  input [63:0] vec_rsc_0_2_qa;
  output vec_rsc_triosy_0_2_lz;
  output [8:0] vec_rsc_0_3_adra;
  output [63:0] vec_rsc_0_3_da;
  output vec_rsc_0_3_wea;
  input [63:0] vec_rsc_0_3_qa;
  output vec_rsc_triosy_0_3_lz;
  output [8:0] vec_rsc_0_4_adra;
  output [63:0] vec_rsc_0_4_da;
  output vec_rsc_0_4_wea;
  input [63:0] vec_rsc_0_4_qa;
  output vec_rsc_triosy_0_4_lz;
  output [8:0] vec_rsc_0_5_adra;
  output [63:0] vec_rsc_0_5_da;
  output vec_rsc_0_5_wea;
  input [63:0] vec_rsc_0_5_qa;
  output vec_rsc_triosy_0_5_lz;
  output [8:0] vec_rsc_0_6_adra;
  output [63:0] vec_rsc_0_6_da;
  output vec_rsc_0_6_wea;
  input [63:0] vec_rsc_0_6_qa;
  output vec_rsc_triosy_0_6_lz;
  output [8:0] vec_rsc_0_7_adra;
  output [63:0] vec_rsc_0_7_da;
  output vec_rsc_0_7_wea;
  input [63:0] vec_rsc_0_7_qa;
  output vec_rsc_triosy_0_7_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;


  // Interconnect Declarations
  wire [63:0] vec_rsc_0_0_i_qa_d;
  wire vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_1_i_qa_d;
  wire vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_2_i_qa_d;
  wire vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_3_i_qa_d;
  wire vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_4_i_qa_d;
  wire vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_5_i_qa_d;
  wire vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_6_i_qa_d;
  wire vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_7_i_qa_d;
  wire vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [8:0] vec_rsc_0_0_i_adra_d_iff;
  wire [63:0] vec_rsc_0_0_i_da_d_iff;
  wire vec_rsc_0_0_i_wea_d_iff;
  wire vec_rsc_0_1_i_wea_d_iff;
  wire vec_rsc_0_2_i_wea_d_iff;
  wire vec_rsc_0_3_i_wea_d_iff;
  wire vec_rsc_0_4_i_wea_d_iff;
  wire vec_rsc_0_5_i_wea_d_iff;
  wire vec_rsc_0_6_i_wea_d_iff;
  wire vec_rsc_0_7_i_wea_d_iff;


  // Interconnect Declarations for Component Instantiations 
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_9_64_512_512_64_1_gen vec_rsc_0_0_i
      (
      .qa(vec_rsc_0_0_qa),
      .wea(vec_rsc_0_0_wea),
      .da(vec_rsc_0_0_da),
      .adra(vec_rsc_0_0_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_0_i_qa_d),
      .wea_d(vec_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_0_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_9_64_512_512_64_1_gen vec_rsc_0_1_i
      (
      .qa(vec_rsc_0_1_qa),
      .wea(vec_rsc_0_1_wea),
      .da(vec_rsc_0_1_da),
      .adra(vec_rsc_0_1_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_1_i_qa_d),
      .wea_d(vec_rsc_0_1_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_1_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_9_64_512_512_64_1_gen vec_rsc_0_2_i
      (
      .qa(vec_rsc_0_2_qa),
      .wea(vec_rsc_0_2_wea),
      .da(vec_rsc_0_2_da),
      .adra(vec_rsc_0_2_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_2_i_qa_d),
      .wea_d(vec_rsc_0_2_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_2_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_9_64_512_512_64_1_gen vec_rsc_0_3_i
      (
      .qa(vec_rsc_0_3_qa),
      .wea(vec_rsc_0_3_wea),
      .da(vec_rsc_0_3_da),
      .adra(vec_rsc_0_3_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_3_i_qa_d),
      .wea_d(vec_rsc_0_3_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_3_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_9_64_512_512_64_1_gen vec_rsc_0_4_i
      (
      .qa(vec_rsc_0_4_qa),
      .wea(vec_rsc_0_4_wea),
      .da(vec_rsc_0_4_da),
      .adra(vec_rsc_0_4_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_4_i_qa_d),
      .wea_d(vec_rsc_0_4_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_4_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_9_64_512_512_64_1_gen vec_rsc_0_5_i
      (
      .qa(vec_rsc_0_5_qa),
      .wea(vec_rsc_0_5_wea),
      .da(vec_rsc_0_5_da),
      .adra(vec_rsc_0_5_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_5_i_qa_d),
      .wea_d(vec_rsc_0_5_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_5_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_9_64_512_512_64_1_gen
      vec_rsc_0_6_i (
      .qa(vec_rsc_0_6_qa),
      .wea(vec_rsc_0_6_wea),
      .da(vec_rsc_0_6_da),
      .adra(vec_rsc_0_6_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_6_i_qa_d),
      .wea_d(vec_rsc_0_6_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_6_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_9_64_512_512_64_1_gen
      vec_rsc_0_7_i (
      .qa(vec_rsc_0_7_qa),
      .wea(vec_rsc_0_7_wea),
      .da(vec_rsc_0_7_da),
      .adra(vec_rsc_0_7_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_7_i_qa_d),
      .wea_d(vec_rsc_0_7_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_7_i_wea_d_iff)
    );
  inPlaceNTT_DIT_core inPlaceNTT_DIT_core_inst (
      .clk(clk),
      .rst(rst),
      .vec_rsc_triosy_0_0_lz(vec_rsc_triosy_0_0_lz),
      .vec_rsc_triosy_0_1_lz(vec_rsc_triosy_0_1_lz),
      .vec_rsc_triosy_0_2_lz(vec_rsc_triosy_0_2_lz),
      .vec_rsc_triosy_0_3_lz(vec_rsc_triosy_0_3_lz),
      .vec_rsc_triosy_0_4_lz(vec_rsc_triosy_0_4_lz),
      .vec_rsc_triosy_0_5_lz(vec_rsc_triosy_0_5_lz),
      .vec_rsc_triosy_0_6_lz(vec_rsc_triosy_0_6_lz),
      .vec_rsc_triosy_0_7_lz(vec_rsc_triosy_0_7_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_dat(r_rsc_dat),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .vec_rsc_0_0_i_qa_d(vec_rsc_0_0_i_qa_d),
      .vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_1_i_qa_d(vec_rsc_0_1_i_qa_d),
      .vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_2_i_qa_d(vec_rsc_0_2_i_qa_d),
      .vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_3_i_qa_d(vec_rsc_0_3_i_qa_d),
      .vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_4_i_qa_d(vec_rsc_0_4_i_qa_d),
      .vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_5_i_qa_d(vec_rsc_0_5_i_qa_d),
      .vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_6_i_qa_d(vec_rsc_0_6_i_qa_d),
      .vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_7_i_qa_d(vec_rsc_0_7_i_qa_d),
      .vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_0_i_adra_d_pff(vec_rsc_0_0_i_adra_d_iff),
      .vec_rsc_0_0_i_da_d_pff(vec_rsc_0_0_i_da_d_iff),
      .vec_rsc_0_0_i_wea_d_pff(vec_rsc_0_0_i_wea_d_iff),
      .vec_rsc_0_1_i_wea_d_pff(vec_rsc_0_1_i_wea_d_iff),
      .vec_rsc_0_2_i_wea_d_pff(vec_rsc_0_2_i_wea_d_iff),
      .vec_rsc_0_3_i_wea_d_pff(vec_rsc_0_3_i_wea_d_iff),
      .vec_rsc_0_4_i_wea_d_pff(vec_rsc_0_4_i_wea_d_iff),
      .vec_rsc_0_5_i_wea_d_pff(vec_rsc_0_5_i_wea_d_iff),
      .vec_rsc_0_6_i_wea_d_pff(vec_rsc_0_6_i_wea_d_iff),
      .vec_rsc_0_7_i_wea_d_pff(vec_rsc_0_7_i_wea_d_iff)
    );
endmodule



